VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO caravel_motto
  CLASS BLOCK ;
  FOREIGN caravel_motto ;
  ORIGIN 0 0 ;
  SIZE 95.050 BY 17.000 ;
  OBS
      LAYER Metal5 ;
        RECT 9337.650 385.490 9338.730 389.810 ;
        RECT 9339.810 385.490 9340.890 389.810 ;
        RECT 9344.420 385.850 9346.940 386.210 ;
        RECT 9344.060 385.490 9346.940 385.850 ;
        RECT 9343.700 384.770 9346.940 385.490 ;
        RECT 9343.700 383.330 9344.780 384.770 ;
        RECT 9354.400 384.000 9356.560 386.160 ;
        RECT 9349.100 383.640 9351.980 384.000 ;
        RECT 9343.700 382.970 9346.220 383.330 ;
        RECT 9343.700 382.610 9346.580 382.970 ;
        RECT 9349.100 382.920 9352.340 383.640 ;
        RECT 9344.060 382.250 9346.940 382.610 ;
        RECT 9344.420 381.890 9346.940 382.250 ;
        RECT 9345.860 380.090 9346.940 381.890 ;
        RECT 9351.260 381.840 9352.340 382.920 ;
        RECT 9354.400 381.840 9356.560 382.920 ;
        RECT 9349.460 381.480 9352.340 381.840 ;
        RECT 9343.700 379.370 9346.940 380.090 ;
        RECT 9349.100 380.760 9352.340 381.480 ;
        RECT 9349.100 379.680 9350.180 380.760 ;
        RECT 9351.260 379.680 9352.340 380.760 ;
        RECT 9355.480 379.680 9356.560 381.840 ;
        RECT 9343.700 379.010 9346.580 379.370 ;
        RECT 9343.700 378.650 9346.220 379.010 ;
        RECT 9349.100 378.960 9352.340 379.680 ;
        RECT 9349.460 378.600 9352.340 378.960 ;
        RECT 9354.400 378.600 9356.560 379.680 ;
        RECT 9358.550 378.550 9359.630 386.110 ;
        RECT 9361.900 383.950 9364.060 386.110 ;
        RECT 9383.400 385.030 9386.640 386.110 ;
        RECT 9365.850 383.590 9368.370 383.950 ;
        RECT 9371.570 383.590 9373.370 383.950 ;
        RECT 9365.850 383.230 9368.730 383.590 ;
        RECT 9371.210 383.230 9373.730 383.590 ;
        RECT 9361.900 381.790 9364.060 382.870 ;
        RECT 9362.980 379.630 9364.060 381.790 ;
        RECT 9361.900 378.550 9364.060 379.630 ;
        RECT 9365.850 382.510 9369.090 383.230 ;
        RECT 9365.850 378.550 9366.930 382.510 ;
        RECT 9368.010 378.550 9369.090 382.510 ;
        RECT 9370.850 382.510 9374.090 383.230 ;
        RECT 9370.850 379.990 9371.930 382.510 ;
        RECT 9373.010 379.990 9374.090 382.510 ;
        RECT 9370.850 379.270 9374.090 379.990 ;
        RECT 9371.210 378.910 9374.090 379.270 ;
        RECT 9371.570 378.550 9374.090 378.910 ;
        RECT 9384.480 378.550 9385.560 385.030 ;
        RECT 9388.650 383.950 9389.730 386.110 ;
        RECT 9406.800 385.080 9410.040 386.160 ;
        RECT 9413.470 385.700 9415.990 386.060 ;
        RECT 9413.110 385.340 9415.990 385.700 ;
        RECT 9424.250 385.490 9425.330 389.810 ;
        RECT 9426.410 385.490 9427.490 389.810 ;
        RECT 9388.650 383.590 9391.170 383.950 ;
        RECT 9394.310 383.590 9396.830 383.950 ;
        RECT 9388.650 383.230 9391.530 383.590 ;
        RECT 9388.650 382.510 9391.890 383.230 ;
        RECT 9388.650 378.550 9389.730 382.510 ;
        RECT 9390.810 378.550 9391.890 382.510 ;
        RECT 9393.950 382.870 9397.190 383.590 ;
        RECT 9393.950 381.790 9395.030 382.870 ;
        RECT 9396.110 381.790 9397.190 382.870 ;
        RECT 9393.950 381.070 9397.190 381.790 ;
        RECT 9393.950 380.710 9396.830 381.070 ;
        RECT 9393.950 379.630 9395.030 380.710 ;
        RECT 9407.880 379.680 9408.960 385.080 ;
        RECT 9412.750 384.620 9415.990 385.340 ;
        RECT 9412.750 379.940 9413.830 384.620 ;
        RECT 9419.370 383.590 9421.890 383.950 ;
        RECT 9419.010 383.230 9421.890 383.590 ;
        RECT 9418.650 382.870 9421.890 383.230 ;
        RECT 9418.650 381.790 9420.090 382.870 ;
        RECT 9418.650 381.430 9421.170 381.790 ;
        RECT 9419.010 381.070 9421.530 381.430 ;
        RECT 9419.370 380.710 9421.890 381.070 ;
        RECT 9393.950 378.910 9397.190 379.630 ;
        RECT 9394.310 378.550 9397.190 378.910 ;
        RECT 9406.800 378.600 9410.040 379.680 ;
        RECT 9412.750 379.220 9415.990 379.940 ;
        RECT 9420.450 379.630 9421.890 380.710 ;
        RECT 9413.110 378.860 9415.990 379.220 ;
        RECT 9372.650 377.470 9374.090 378.550 ;
        RECT 9413.470 378.500 9415.990 378.860 ;
        RECT 9418.650 379.270 9421.890 379.630 ;
        RECT 9418.650 378.910 9421.530 379.270 ;
        RECT 9418.650 378.550 9421.170 378.910 ;
        RECT 9370.850 377.110 9374.090 377.470 ;
        RECT 9370.850 376.750 9373.730 377.110 ;
        RECT 9370.850 376.390 9373.370 376.750 ;
  END
END caravel_motto
END LIBRARY

