magic
tech gf180mcuC
magscale 1 5
timestamp 1655473382
<< checkpaint >>
rect -1530 -1200 236506 101200
<< obsm1 >>
rect 560 1051 234416 99917
<< metal2 >>
rect 252 99600 308 100200
rect 868 99600 924 100200
rect 1484 99600 1540 100200
rect 2156 99600 2212 100200
rect 2772 99600 2828 100200
rect 3444 99600 3500 100200
rect 4060 99600 4116 100200
rect 4732 99600 4788 100200
rect 5348 99600 5404 100200
rect 5964 99600 6020 100200
rect 6636 99600 6692 100200
rect 7252 99600 7308 100200
rect 7924 99600 7980 100200
rect 8540 99600 8596 100200
rect 9212 99600 9268 100200
rect 9828 99600 9884 100200
rect 10444 99600 10500 100200
rect 11116 99600 11172 100200
rect 11732 99600 11788 100200
rect 12404 99600 12460 100200
rect 13020 99600 13076 100200
rect 13692 99600 13748 100200
rect 14308 99600 14364 100200
rect 14980 99600 15036 100200
rect 15596 99600 15652 100200
rect 16212 99600 16268 100200
rect 16884 99600 16940 100200
rect 17500 99600 17556 100200
rect 18172 99600 18228 100200
rect 18788 99600 18844 100200
rect 19460 99600 19516 100200
rect 20076 99600 20132 100200
rect 20692 99600 20748 100200
rect 21364 99600 21420 100200
rect 21980 99600 22036 100200
rect 22652 99600 22708 100200
rect 23268 99600 23324 100200
rect 23940 99600 23996 100200
rect 24556 99600 24612 100200
rect 25228 99600 25284 100200
rect 25844 99600 25900 100200
rect 26460 99600 26516 100200
rect 27132 99600 27188 100200
rect 27748 99600 27804 100200
rect 28420 99600 28476 100200
rect 29036 99600 29092 100200
rect 29708 99600 29764 100200
rect 30324 99600 30380 100200
rect 30940 99600 30996 100200
rect 31612 99600 31668 100200
rect 32228 99600 32284 100200
rect 32900 99600 32956 100200
rect 33516 99600 33572 100200
rect 34188 99600 34244 100200
rect 34804 99600 34860 100200
rect 35420 99600 35476 100200
rect 36092 99600 36148 100200
rect 36708 99600 36764 100200
rect 37380 99600 37436 100200
rect 37996 99600 38052 100200
rect 38668 99600 38724 100200
rect 39284 99600 39340 100200
rect 39956 99600 40012 100200
rect 40572 99600 40628 100200
rect 41188 99600 41244 100200
rect 41860 99600 41916 100200
rect 42476 99600 42532 100200
rect 43148 99600 43204 100200
rect 43764 99600 43820 100200
rect 44436 99600 44492 100200
rect 45052 99600 45108 100200
rect 45668 99600 45724 100200
rect 46340 99600 46396 100200
rect 46956 99600 47012 100200
rect 47628 99600 47684 100200
rect 48244 99600 48300 100200
rect 48916 99600 48972 100200
rect 49532 99600 49588 100200
rect 50204 99600 50260 100200
rect 50820 99600 50876 100200
rect 51436 99600 51492 100200
rect 52108 99600 52164 100200
rect 52724 99600 52780 100200
rect 53396 99600 53452 100200
rect 54012 99600 54068 100200
rect 54684 99600 54740 100200
rect 55300 99600 55356 100200
rect 55916 99600 55972 100200
rect 56588 99600 56644 100200
rect 57204 99600 57260 100200
rect 57876 99600 57932 100200
rect 58492 99600 58548 100200
rect 59164 99600 59220 100200
rect 59780 99600 59836 100200
rect 60396 99600 60452 100200
rect 61068 99600 61124 100200
rect 61684 99600 61740 100200
rect 62356 99600 62412 100200
rect 62972 99600 63028 100200
rect 63644 99600 63700 100200
rect 64260 99600 64316 100200
rect 64932 99600 64988 100200
rect 65548 99600 65604 100200
rect 66164 99600 66220 100200
rect 66836 99600 66892 100200
rect 67452 99600 67508 100200
rect 68124 99600 68180 100200
rect 68740 99600 68796 100200
rect 69412 99600 69468 100200
rect 70028 99600 70084 100200
rect 70644 99600 70700 100200
rect 71316 99600 71372 100200
rect 71932 99600 71988 100200
rect 72604 99600 72660 100200
rect 73220 99600 73276 100200
rect 73892 99600 73948 100200
rect 74508 99600 74564 100200
rect 75180 99600 75236 100200
rect 75796 99600 75852 100200
rect 76412 99600 76468 100200
rect 77084 99600 77140 100200
rect 77700 99600 77756 100200
rect 78372 99600 78428 100200
rect 78988 99600 79044 100200
rect 79660 99600 79716 100200
rect 80276 99600 80332 100200
rect 80892 99600 80948 100200
rect 81564 99600 81620 100200
rect 82180 99600 82236 100200
rect 82852 99600 82908 100200
rect 83468 99600 83524 100200
rect 84140 99600 84196 100200
rect 84756 99600 84812 100200
rect 85372 99600 85428 100200
rect 86044 99600 86100 100200
rect 86660 99600 86716 100200
rect 87332 99600 87388 100200
rect 87948 99600 88004 100200
rect 88620 99600 88676 100200
rect 89236 99600 89292 100200
rect 89908 99600 89964 100200
rect 90524 99600 90580 100200
rect 91140 99600 91196 100200
rect 91812 99600 91868 100200
rect 92428 99600 92484 100200
rect 93100 99600 93156 100200
rect 93716 99600 93772 100200
rect 94388 99600 94444 100200
rect 95004 99600 95060 100200
rect 95620 99600 95676 100200
rect 96292 99600 96348 100200
rect 96908 99600 96964 100200
rect 97580 99600 97636 100200
rect 98196 99600 98252 100200
rect 98868 99600 98924 100200
rect 99484 99600 99540 100200
rect 100156 99600 100212 100200
rect 100772 99600 100828 100200
rect 101388 99600 101444 100200
rect 102060 99600 102116 100200
rect 102676 99600 102732 100200
rect 103348 99600 103404 100200
rect 103964 99600 104020 100200
rect 104636 99600 104692 100200
rect 105252 99600 105308 100200
rect 105868 99600 105924 100200
rect 106540 99600 106596 100200
rect 107156 99600 107212 100200
rect 107828 99600 107884 100200
rect 108444 99600 108500 100200
rect 109116 99600 109172 100200
rect 109732 99600 109788 100200
rect 110348 99600 110404 100200
rect 111020 99600 111076 100200
rect 111636 99600 111692 100200
rect 112308 99600 112364 100200
rect 112924 99600 112980 100200
rect 113596 99600 113652 100200
rect 114212 99600 114268 100200
rect 114884 99600 114940 100200
rect 115500 99600 115556 100200
rect 116116 99600 116172 100200
rect 116788 99600 116844 100200
rect 117404 99600 117460 100200
rect 118076 99600 118132 100200
rect 118692 99600 118748 100200
rect 119364 99600 119420 100200
rect 119980 99600 120036 100200
rect 120596 99600 120652 100200
rect 121268 99600 121324 100200
rect 121884 99600 121940 100200
rect 122556 99600 122612 100200
rect 123172 99600 123228 100200
rect 123844 99600 123900 100200
rect 124460 99600 124516 100200
rect 125132 99600 125188 100200
rect 125748 99600 125804 100200
rect 126364 99600 126420 100200
rect 127036 99600 127092 100200
rect 127652 99600 127708 100200
rect 128324 99600 128380 100200
rect 128940 99600 128996 100200
rect 129612 99600 129668 100200
rect 130228 99600 130284 100200
rect 130844 99600 130900 100200
rect 131516 99600 131572 100200
rect 132132 99600 132188 100200
rect 132804 99600 132860 100200
rect 133420 99600 133476 100200
rect 134092 99600 134148 100200
rect 134708 99600 134764 100200
rect 135324 99600 135380 100200
rect 135996 99600 136052 100200
rect 136612 99600 136668 100200
rect 137284 99600 137340 100200
rect 137900 99600 137956 100200
rect 138572 99600 138628 100200
rect 139188 99600 139244 100200
rect 139860 99600 139916 100200
rect 140476 99600 140532 100200
rect 141092 99600 141148 100200
rect 141764 99600 141820 100200
rect 142380 99600 142436 100200
rect 143052 99600 143108 100200
rect 143668 99600 143724 100200
rect 144340 99600 144396 100200
rect 144956 99600 145012 100200
rect 145572 99600 145628 100200
rect 146244 99600 146300 100200
rect 146860 99600 146916 100200
rect 147532 99600 147588 100200
rect 148148 99600 148204 100200
rect 148820 99600 148876 100200
rect 149436 99600 149492 100200
rect 150108 99600 150164 100200
rect 150724 99600 150780 100200
rect 151340 99600 151396 100200
rect 152012 99600 152068 100200
rect 152628 99600 152684 100200
rect 153300 99600 153356 100200
rect 153916 99600 153972 100200
rect 154588 99600 154644 100200
rect 155204 99600 155260 100200
rect 155820 99600 155876 100200
rect 156492 99600 156548 100200
rect 157108 99600 157164 100200
rect 157780 99600 157836 100200
rect 158396 99600 158452 100200
rect 159068 99600 159124 100200
rect 159684 99600 159740 100200
rect 160300 99600 160356 100200
rect 160972 99600 161028 100200
rect 161588 99600 161644 100200
rect 162260 99600 162316 100200
rect 162876 99600 162932 100200
rect 163548 99600 163604 100200
rect 164164 99600 164220 100200
rect 164836 99600 164892 100200
rect 165452 99600 165508 100200
rect 166068 99600 166124 100200
rect 166740 99600 166796 100200
rect 167356 99600 167412 100200
rect 168028 99600 168084 100200
rect 168644 99600 168700 100200
rect 169316 99600 169372 100200
rect 169932 99600 169988 100200
rect 170548 99600 170604 100200
rect 171220 99600 171276 100200
rect 171836 99600 171892 100200
rect 172508 99600 172564 100200
rect 173124 99600 173180 100200
rect 173796 99600 173852 100200
rect 174412 99600 174468 100200
rect 175084 99600 175140 100200
rect 175700 99600 175756 100200
rect 176316 99600 176372 100200
rect 176988 99600 177044 100200
rect 177604 99600 177660 100200
rect 178276 99600 178332 100200
rect 178892 99600 178948 100200
rect 179564 99600 179620 100200
rect 180180 99600 180236 100200
rect 180796 99600 180852 100200
rect 181468 99600 181524 100200
rect 182084 99600 182140 100200
rect 182756 99600 182812 100200
rect 183372 99600 183428 100200
rect 184044 99600 184100 100200
rect 184660 99600 184716 100200
rect 185276 99600 185332 100200
rect 185948 99600 186004 100200
rect 186564 99600 186620 100200
rect 187236 99600 187292 100200
rect 187852 99600 187908 100200
rect 188524 99600 188580 100200
rect 189140 99600 189196 100200
rect 189812 99600 189868 100200
rect 190428 99600 190484 100200
rect 191044 99600 191100 100200
rect 191716 99600 191772 100200
rect 192332 99600 192388 100200
rect 193004 99600 193060 100200
rect 193620 99600 193676 100200
rect 194292 99600 194348 100200
rect 194908 99600 194964 100200
rect 195524 99600 195580 100200
rect 196196 99600 196252 100200
rect 196812 99600 196868 100200
rect 197484 99600 197540 100200
rect 198100 99600 198156 100200
rect 198772 99600 198828 100200
rect 199388 99600 199444 100200
rect 200060 99600 200116 100200
rect 200676 99600 200732 100200
rect 201292 99600 201348 100200
rect 201964 99600 202020 100200
rect 202580 99600 202636 100200
rect 203252 99600 203308 100200
rect 203868 99600 203924 100200
rect 204540 99600 204596 100200
rect 205156 99600 205212 100200
rect 205772 99600 205828 100200
rect 206444 99600 206500 100200
rect 207060 99600 207116 100200
rect 207732 99600 207788 100200
rect 208348 99600 208404 100200
rect 209020 99600 209076 100200
rect 209636 99600 209692 100200
rect 210252 99600 210308 100200
rect 210924 99600 210980 100200
rect 211540 99600 211596 100200
rect 212212 99600 212268 100200
rect 212828 99600 212884 100200
rect 213500 99600 213556 100200
rect 214116 99600 214172 100200
rect 214788 99600 214844 100200
rect 215404 99600 215460 100200
rect 216020 99600 216076 100200
rect 216692 99600 216748 100200
rect 217308 99600 217364 100200
rect 217980 99600 218036 100200
rect 218596 99600 218652 100200
rect 219268 99600 219324 100200
rect 219884 99600 219940 100200
rect 220500 99600 220556 100200
rect 221172 99600 221228 100200
rect 221788 99600 221844 100200
rect 222460 99600 222516 100200
rect 223076 99600 223132 100200
rect 223748 99600 223804 100200
rect 224364 99600 224420 100200
rect 225036 99600 225092 100200
rect 225652 99600 225708 100200
rect 226268 99600 226324 100200
rect 226940 99600 226996 100200
rect 227556 99600 227612 100200
rect 228228 99600 228284 100200
rect 228844 99600 228900 100200
rect 229516 99600 229572 100200
rect 230132 99600 230188 100200
rect 230748 99600 230804 100200
rect 231420 99600 231476 100200
rect 232036 99600 232092 100200
rect 232708 99600 232764 100200
rect 233324 99600 233380 100200
rect 233996 99600 234052 100200
rect 234612 99600 234668 100200
rect 16716 -200 16772 400
rect 50260 -200 50316 400
rect 83860 -200 83916 400
rect 117404 -200 117460 400
rect 151004 -200 151060 400
rect 184548 -200 184604 400
rect 218148 -200 218204 400
<< obsm2 >>
rect 338 99570 838 99979
rect 954 99570 1454 99979
rect 1570 99570 2126 99979
rect 2242 99570 2742 99979
rect 2858 99570 3414 99979
rect 3530 99570 4030 99979
rect 4146 99570 4702 99979
rect 4818 99570 5318 99979
rect 5434 99570 5934 99979
rect 6050 99570 6606 99979
rect 6722 99570 7222 99979
rect 7338 99570 7894 99979
rect 8010 99570 8510 99979
rect 8626 99570 9182 99979
rect 9298 99570 9798 99979
rect 9914 99570 10414 99979
rect 10530 99570 11086 99979
rect 11202 99570 11702 99979
rect 11818 99570 12374 99979
rect 12490 99570 12990 99979
rect 13106 99570 13662 99979
rect 13778 99570 14278 99979
rect 14394 99570 14950 99979
rect 15066 99570 15566 99979
rect 15682 99570 16182 99979
rect 16298 99570 16854 99979
rect 16970 99570 17470 99979
rect 17586 99570 18142 99979
rect 18258 99570 18758 99979
rect 18874 99570 19430 99979
rect 19546 99570 20046 99979
rect 20162 99570 20662 99979
rect 20778 99570 21334 99979
rect 21450 99570 21950 99979
rect 22066 99570 22622 99979
rect 22738 99570 23238 99979
rect 23354 99570 23910 99979
rect 24026 99570 24526 99979
rect 24642 99570 25198 99979
rect 25314 99570 25814 99979
rect 25930 99570 26430 99979
rect 26546 99570 27102 99979
rect 27218 99570 27718 99979
rect 27834 99570 28390 99979
rect 28506 99570 29006 99979
rect 29122 99570 29678 99979
rect 29794 99570 30294 99979
rect 30410 99570 30910 99979
rect 31026 99570 31582 99979
rect 31698 99570 32198 99979
rect 32314 99570 32870 99979
rect 32986 99570 33486 99979
rect 33602 99570 34158 99979
rect 34274 99570 34774 99979
rect 34890 99570 35390 99979
rect 35506 99570 36062 99979
rect 36178 99570 36678 99979
rect 36794 99570 37350 99979
rect 37466 99570 37966 99979
rect 38082 99570 38638 99979
rect 38754 99570 39254 99979
rect 39370 99570 39926 99979
rect 40042 99570 40542 99979
rect 40658 99570 41158 99979
rect 41274 99570 41830 99979
rect 41946 99570 42446 99979
rect 42562 99570 43118 99979
rect 43234 99570 43734 99979
rect 43850 99570 44406 99979
rect 44522 99570 45022 99979
rect 45138 99570 45638 99979
rect 45754 99570 46310 99979
rect 46426 99570 46926 99979
rect 47042 99570 47598 99979
rect 47714 99570 48214 99979
rect 48330 99570 48886 99979
rect 49002 99570 49502 99979
rect 49618 99570 50174 99979
rect 50290 99570 50790 99979
rect 50906 99570 51406 99979
rect 51522 99570 52078 99979
rect 52194 99570 52694 99979
rect 52810 99570 53366 99979
rect 53482 99570 53982 99979
rect 54098 99570 54654 99979
rect 54770 99570 55270 99979
rect 55386 99570 55886 99979
rect 56002 99570 56558 99979
rect 56674 99570 57174 99979
rect 57290 99570 57846 99979
rect 57962 99570 58462 99979
rect 58578 99570 59134 99979
rect 59250 99570 59750 99979
rect 59866 99570 60366 99979
rect 60482 99570 61038 99979
rect 61154 99570 61654 99979
rect 61770 99570 62326 99979
rect 62442 99570 62942 99979
rect 63058 99570 63614 99979
rect 63730 99570 64230 99979
rect 64346 99570 64902 99979
rect 65018 99570 65518 99979
rect 65634 99570 66134 99979
rect 66250 99570 66806 99979
rect 66922 99570 67422 99979
rect 67538 99570 68094 99979
rect 68210 99570 68710 99979
rect 68826 99570 69382 99979
rect 69498 99570 69998 99979
rect 70114 99570 70614 99979
rect 70730 99570 71286 99979
rect 71402 99570 71902 99979
rect 72018 99570 72574 99979
rect 72690 99570 73190 99979
rect 73306 99570 73862 99979
rect 73978 99570 74478 99979
rect 74594 99570 75150 99979
rect 75266 99570 75766 99979
rect 75882 99570 76382 99979
rect 76498 99570 77054 99979
rect 77170 99570 77670 99979
rect 77786 99570 78342 99979
rect 78458 99570 78958 99979
rect 79074 99570 79630 99979
rect 79746 99570 80246 99979
rect 80362 99570 80862 99979
rect 80978 99570 81534 99979
rect 81650 99570 82150 99979
rect 82266 99570 82822 99979
rect 82938 99570 83438 99979
rect 83554 99570 84110 99979
rect 84226 99570 84726 99979
rect 84842 99570 85342 99979
rect 85458 99570 86014 99979
rect 86130 99570 86630 99979
rect 86746 99570 87302 99979
rect 87418 99570 87918 99979
rect 88034 99570 88590 99979
rect 88706 99570 89206 99979
rect 89322 99570 89878 99979
rect 89994 99570 90494 99979
rect 90610 99570 91110 99979
rect 91226 99570 91782 99979
rect 91898 99570 92398 99979
rect 92514 99570 93070 99979
rect 93186 99570 93686 99979
rect 93802 99570 94358 99979
rect 94474 99570 94974 99979
rect 95090 99570 95590 99979
rect 95706 99570 96262 99979
rect 96378 99570 96878 99979
rect 96994 99570 97550 99979
rect 97666 99570 98166 99979
rect 98282 99570 98838 99979
rect 98954 99570 99454 99979
rect 99570 99570 100126 99979
rect 100242 99570 100742 99979
rect 100858 99570 101358 99979
rect 101474 99570 102030 99979
rect 102146 99570 102646 99979
rect 102762 99570 103318 99979
rect 103434 99570 103934 99979
rect 104050 99570 104606 99979
rect 104722 99570 105222 99979
rect 105338 99570 105838 99979
rect 105954 99570 106510 99979
rect 106626 99570 107126 99979
rect 107242 99570 107798 99979
rect 107914 99570 108414 99979
rect 108530 99570 109086 99979
rect 109202 99570 109702 99979
rect 109818 99570 110318 99979
rect 110434 99570 110990 99979
rect 111106 99570 111606 99979
rect 111722 99570 112278 99979
rect 112394 99570 112894 99979
rect 113010 99570 113566 99979
rect 113682 99570 114182 99979
rect 114298 99570 114854 99979
rect 114970 99570 115470 99979
rect 115586 99570 116086 99979
rect 116202 99570 116758 99979
rect 116874 99570 117374 99979
rect 117490 99570 118046 99979
rect 118162 99570 118662 99979
rect 118778 99570 119334 99979
rect 119450 99570 119950 99979
rect 120066 99570 120566 99979
rect 120682 99570 121238 99979
rect 121354 99570 121854 99979
rect 121970 99570 122526 99979
rect 122642 99570 123142 99979
rect 123258 99570 123814 99979
rect 123930 99570 124430 99979
rect 124546 99570 125102 99979
rect 125218 99570 125718 99979
rect 125834 99570 126334 99979
rect 126450 99570 127006 99979
rect 127122 99570 127622 99979
rect 127738 99570 128294 99979
rect 128410 99570 128910 99979
rect 129026 99570 129582 99979
rect 129698 99570 130198 99979
rect 130314 99570 130814 99979
rect 130930 99570 131486 99979
rect 131602 99570 132102 99979
rect 132218 99570 132774 99979
rect 132890 99570 133390 99979
rect 133506 99570 134062 99979
rect 134178 99570 134678 99979
rect 134794 99570 135294 99979
rect 135410 99570 135966 99979
rect 136082 99570 136582 99979
rect 136698 99570 137254 99979
rect 137370 99570 137870 99979
rect 137986 99570 138542 99979
rect 138658 99570 139158 99979
rect 139274 99570 139830 99979
rect 139946 99570 140446 99979
rect 140562 99570 141062 99979
rect 141178 99570 141734 99979
rect 141850 99570 142350 99979
rect 142466 99570 143022 99979
rect 143138 99570 143638 99979
rect 143754 99570 144310 99979
rect 144426 99570 144926 99979
rect 145042 99570 145542 99979
rect 145658 99570 146214 99979
rect 146330 99570 146830 99979
rect 146946 99570 147502 99979
rect 147618 99570 148118 99979
rect 148234 99570 148790 99979
rect 148906 99570 149406 99979
rect 149522 99570 150078 99979
rect 150194 99570 150694 99979
rect 150810 99570 151310 99979
rect 151426 99570 151982 99979
rect 152098 99570 152598 99979
rect 152714 99570 153270 99979
rect 153386 99570 153886 99979
rect 154002 99570 154558 99979
rect 154674 99570 155174 99979
rect 155290 99570 155790 99979
rect 155906 99570 156462 99979
rect 156578 99570 157078 99979
rect 157194 99570 157750 99979
rect 157866 99570 158366 99979
rect 158482 99570 159038 99979
rect 159154 99570 159654 99979
rect 159770 99570 160270 99979
rect 160386 99570 160942 99979
rect 161058 99570 161558 99979
rect 161674 99570 162230 99979
rect 162346 99570 162846 99979
rect 162962 99570 163518 99979
rect 163634 99570 164134 99979
rect 164250 99570 164806 99979
rect 164922 99570 165422 99979
rect 165538 99570 166038 99979
rect 166154 99570 166710 99979
rect 166826 99570 167326 99979
rect 167442 99570 167998 99979
rect 168114 99570 168614 99979
rect 168730 99570 169286 99979
rect 169402 99570 169902 99979
rect 170018 99570 170518 99979
rect 170634 99570 171190 99979
rect 171306 99570 171806 99979
rect 171922 99570 172478 99979
rect 172594 99570 173094 99979
rect 173210 99570 173766 99979
rect 173882 99570 174382 99979
rect 174498 99570 175054 99979
rect 175170 99570 175670 99979
rect 175786 99570 176286 99979
rect 176402 99570 176958 99979
rect 177074 99570 177574 99979
rect 177690 99570 178246 99979
rect 178362 99570 178862 99979
rect 178978 99570 179534 99979
rect 179650 99570 180150 99979
rect 180266 99570 180766 99979
rect 180882 99570 181438 99979
rect 181554 99570 182054 99979
rect 182170 99570 182726 99979
rect 182842 99570 183342 99979
rect 183458 99570 184014 99979
rect 184130 99570 184630 99979
rect 184746 99570 185246 99979
rect 185362 99570 185918 99979
rect 186034 99570 186534 99979
rect 186650 99570 187206 99979
rect 187322 99570 187822 99979
rect 187938 99570 188494 99979
rect 188610 99570 189110 99979
rect 189226 99570 189782 99979
rect 189898 99570 190398 99979
rect 190514 99570 191014 99979
rect 191130 99570 191686 99979
rect 191802 99570 192302 99979
rect 192418 99570 192974 99979
rect 193090 99570 193590 99979
rect 193706 99570 194262 99979
rect 194378 99570 194878 99979
rect 194994 99570 195494 99979
rect 195610 99570 196166 99979
rect 196282 99570 196782 99979
rect 196898 99570 197454 99979
rect 197570 99570 198070 99979
rect 198186 99570 198742 99979
rect 198858 99570 199358 99979
rect 199474 99570 200030 99979
rect 200146 99570 200646 99979
rect 200762 99570 201262 99979
rect 201378 99570 201934 99979
rect 202050 99570 202550 99979
rect 202666 99570 203222 99979
rect 203338 99570 203838 99979
rect 203954 99570 204510 99979
rect 204626 99570 205126 99979
rect 205242 99570 205742 99979
rect 205858 99570 206414 99979
rect 206530 99570 207030 99979
rect 207146 99570 207702 99979
rect 207818 99570 208318 99979
rect 208434 99570 208990 99979
rect 209106 99570 209606 99979
rect 209722 99570 210222 99979
rect 210338 99570 210894 99979
rect 211010 99570 211510 99979
rect 211626 99570 212182 99979
rect 212298 99570 212798 99979
rect 212914 99570 213470 99979
rect 213586 99570 214086 99979
rect 214202 99570 214758 99979
rect 214874 99570 215374 99979
rect 215490 99570 215990 99979
rect 216106 99570 216662 99979
rect 216778 99570 217278 99979
rect 217394 99570 217950 99979
rect 218066 99570 218566 99979
rect 218682 99570 219238 99979
rect 219354 99570 219854 99979
rect 219970 99570 220470 99979
rect 220586 99570 221142 99979
rect 221258 99570 221758 99979
rect 221874 99570 222430 99979
rect 222546 99570 223046 99979
rect 223162 99570 223718 99979
rect 223834 99570 224334 99979
rect 224450 99570 225006 99979
rect 225122 99570 225622 99979
rect 225738 99570 226238 99979
rect 226354 99570 226910 99979
rect 227026 99570 227526 99979
rect 227642 99570 228198 99979
rect 228314 99570 228814 99979
rect 228930 99570 229486 99979
rect 229602 99570 230102 99979
rect 230218 99570 230718 99979
rect 230834 99570 231390 99979
rect 231506 99570 232006 99979
rect 232122 99570 232678 99979
rect 232794 99570 233294 99979
rect 233410 99570 233966 99979
rect 234082 99570 234582 99979
rect 266 430 234654 99570
rect 266 400 16686 430
rect 16802 400 50230 430
rect 50346 400 83830 430
rect 83946 400 117374 430
rect 117490 400 150974 430
rect 151090 400 184518 430
rect 184634 400 218118 430
rect 218234 400 234654 430
<< metal3 >>
rect 234600 99204 235200 99260
rect 234600 97748 235200 97804
rect 234600 96292 235200 96348
rect 234600 94836 235200 94892
rect 234600 93324 235200 93380
rect 234600 91868 235200 91924
rect 234600 90412 235200 90468
rect 234600 88956 235200 89012
rect 234600 87444 235200 87500
rect 234600 85988 235200 86044
rect 234600 84532 235200 84588
rect 234600 83076 235200 83132
rect 234600 81564 235200 81620
rect 234600 80108 235200 80164
rect 234600 78652 235200 78708
rect 234600 77196 235200 77252
rect 234600 75684 235200 75740
rect 234600 74228 235200 74284
rect 234600 72772 235200 72828
rect 234600 71316 235200 71372
rect 234600 69804 235200 69860
rect 234600 68348 235200 68404
rect 234600 66892 235200 66948
rect 234600 65436 235200 65492
rect 234600 63924 235200 63980
rect 234600 62468 235200 62524
rect 234600 61012 235200 61068
rect 234600 59556 235200 59612
rect 234600 58044 235200 58100
rect 234600 56588 235200 56644
rect 234600 55132 235200 55188
rect 234600 53676 235200 53732
rect 234600 52164 235200 52220
rect 234600 50708 235200 50764
rect 234600 49252 235200 49308
rect 234600 47796 235200 47852
rect 234600 46284 235200 46340
rect 234600 44828 235200 44884
rect 234600 43372 235200 43428
rect 234600 41916 235200 41972
rect 234600 40404 235200 40460
rect 234600 38948 235200 39004
rect 234600 37492 235200 37548
rect 234600 36036 235200 36092
rect 234600 34524 235200 34580
rect 234600 33068 235200 33124
rect 234600 31612 235200 31668
rect 234600 30156 235200 30212
rect 234600 28644 235200 28700
rect 234600 27188 235200 27244
rect 234600 25732 235200 25788
rect 234600 24276 235200 24332
rect 234600 22764 235200 22820
rect 234600 21308 235200 21364
rect 234600 19852 235200 19908
rect 234600 18396 235200 18452
rect 234600 16884 235200 16940
rect 234600 15428 235200 15484
rect 234600 13972 235200 14028
rect 234600 12516 235200 12572
rect 234600 11004 235200 11060
rect 234600 9548 235200 9604
rect 234600 8092 235200 8148
rect 234600 6636 235200 6692
rect 234600 5124 235200 5180
rect 234600 3668 235200 3724
rect 234600 2212 235200 2268
rect 234600 756 235200 812
<< obsm3 >>
rect 765 99290 234600 99974
rect 765 99174 234570 99290
rect 765 97834 234600 99174
rect 765 97718 234570 97834
rect 765 96378 234600 97718
rect 765 96262 234570 96378
rect 765 94922 234600 96262
rect 765 94806 234570 94922
rect 765 93410 234600 94806
rect 765 93294 234570 93410
rect 765 91954 234600 93294
rect 765 91838 234570 91954
rect 765 90498 234600 91838
rect 765 90382 234570 90498
rect 765 89042 234600 90382
rect 765 88926 234570 89042
rect 765 87530 234600 88926
rect 765 87414 234570 87530
rect 765 86074 234600 87414
rect 765 85958 234570 86074
rect 765 84618 234600 85958
rect 765 84502 234570 84618
rect 765 83162 234600 84502
rect 765 83046 234570 83162
rect 765 81650 234600 83046
rect 765 81534 234570 81650
rect 765 80194 234600 81534
rect 765 80078 234570 80194
rect 765 78738 234600 80078
rect 765 78622 234570 78738
rect 765 77282 234600 78622
rect 765 77166 234570 77282
rect 765 75770 234600 77166
rect 765 75654 234570 75770
rect 765 74314 234600 75654
rect 765 74198 234570 74314
rect 765 72858 234600 74198
rect 765 72742 234570 72858
rect 765 71402 234600 72742
rect 765 71286 234570 71402
rect 765 69890 234600 71286
rect 765 69774 234570 69890
rect 765 68434 234600 69774
rect 765 68318 234570 68434
rect 765 66978 234600 68318
rect 765 66862 234570 66978
rect 765 65522 234600 66862
rect 765 65406 234570 65522
rect 765 64010 234600 65406
rect 765 63894 234570 64010
rect 765 62554 234600 63894
rect 765 62438 234570 62554
rect 765 61098 234600 62438
rect 765 60982 234570 61098
rect 765 59642 234600 60982
rect 765 59526 234570 59642
rect 765 58130 234600 59526
rect 765 58014 234570 58130
rect 765 56674 234600 58014
rect 765 56558 234570 56674
rect 765 55218 234600 56558
rect 765 55102 234570 55218
rect 765 53762 234600 55102
rect 765 53646 234570 53762
rect 765 52250 234600 53646
rect 765 52134 234570 52250
rect 765 50794 234600 52134
rect 765 50678 234570 50794
rect 765 49338 234600 50678
rect 765 49222 234570 49338
rect 765 47882 234600 49222
rect 765 47766 234570 47882
rect 765 46370 234600 47766
rect 765 46254 234570 46370
rect 765 44914 234600 46254
rect 765 44798 234570 44914
rect 765 43458 234600 44798
rect 765 43342 234570 43458
rect 765 42002 234600 43342
rect 765 41886 234570 42002
rect 765 40490 234600 41886
rect 765 40374 234570 40490
rect 765 39034 234600 40374
rect 765 38918 234570 39034
rect 765 37578 234600 38918
rect 765 37462 234570 37578
rect 765 36122 234600 37462
rect 765 36006 234570 36122
rect 765 34610 234600 36006
rect 765 34494 234570 34610
rect 765 33154 234600 34494
rect 765 33038 234570 33154
rect 765 31698 234600 33038
rect 765 31582 234570 31698
rect 765 30242 234600 31582
rect 765 30126 234570 30242
rect 765 28730 234600 30126
rect 765 28614 234570 28730
rect 765 27274 234600 28614
rect 765 27158 234570 27274
rect 765 25818 234600 27158
rect 765 25702 234570 25818
rect 765 24362 234600 25702
rect 765 24246 234570 24362
rect 765 22850 234600 24246
rect 765 22734 234570 22850
rect 765 21394 234600 22734
rect 765 21278 234570 21394
rect 765 19938 234600 21278
rect 765 19822 234570 19938
rect 765 18482 234600 19822
rect 765 18366 234570 18482
rect 765 16970 234600 18366
rect 765 16854 234570 16970
rect 765 15514 234600 16854
rect 765 15398 234570 15514
rect 765 14058 234600 15398
rect 765 13942 234570 14058
rect 765 12602 234600 13942
rect 765 12486 234570 12602
rect 765 11090 234600 12486
rect 765 10974 234570 11090
rect 765 9634 234600 10974
rect 765 9518 234570 9634
rect 765 8178 234600 9518
rect 765 8062 234570 8178
rect 765 6722 234600 8062
rect 765 6606 234570 6722
rect 765 5210 234600 6606
rect 765 5094 234570 5210
rect 765 3754 234600 5094
rect 765 3638 234570 3754
rect 765 2298 234600 3638
rect 765 2182 234570 2298
rect 765 842 234600 2182
rect 765 726 234570 842
rect 765 658 234600 726
<< metal4 >>
rect -530 86 -370 99874
rect -200 416 -40 99544
rect 2112 86 2272 99874
rect 4612 86 4772 99874
rect 7112 86 7272 99874
rect 9612 86 9772 99874
rect 12112 86 12272 99874
rect 14612 86 14772 99874
rect 17112 86 17272 99874
rect 19612 86 19772 99874
rect 22112 86 22272 99874
rect 24612 86 24772 99874
rect 27112 86 27272 99874
rect 29612 86 29772 99874
rect 32112 86 32272 99874
rect 34612 86 34772 99874
rect 37112 86 37272 99874
rect 39612 86 39772 99874
rect 42112 86 42272 99874
rect 44612 86 44772 99874
rect 47112 86 47272 99874
rect 49612 86 49772 99874
rect 52112 86 52272 99874
rect 54612 86 54772 99874
rect 57112 86 57272 99874
rect 59612 86 59772 99874
rect 62112 86 62272 99874
rect 64612 86 64772 99874
rect 67112 86 67272 99874
rect 69612 86 69772 99874
rect 72112 86 72272 99874
rect 74612 86 74772 99874
rect 77112 86 77272 99874
rect 79612 86 79772 99874
rect 82112 86 82272 99874
rect 84612 86 84772 99874
rect 87112 86 87272 99874
rect 89612 86 89772 99874
rect 92112 86 92272 99874
rect 94612 86 94772 99874
rect 97112 86 97272 99874
rect 99612 86 99772 99874
rect 102112 86 102272 99874
rect 104612 86 104772 99874
rect 107112 86 107272 99874
rect 109612 86 109772 99874
rect 112112 86 112272 99874
rect 114612 86 114772 99874
rect 117112 86 117272 99874
rect 119612 86 119772 99874
rect 122112 86 122272 99874
rect 124612 86 124772 99874
rect 127112 86 127272 99874
rect 129612 86 129772 99874
rect 132112 86 132272 99874
rect 134612 86 134772 99874
rect 137112 86 137272 99874
rect 139612 86 139772 99874
rect 142112 86 142272 99874
rect 144612 86 144772 99874
rect 147112 86 147272 99874
rect 149612 86 149772 99874
rect 152112 86 152272 99874
rect 154612 86 154772 99874
rect 157112 86 157272 99874
rect 159612 86 159772 99874
rect 162112 86 162272 99874
rect 164612 86 164772 99874
rect 167112 86 167272 99874
rect 169612 86 169772 99874
rect 172112 86 172272 99874
rect 174612 86 174772 99874
rect 177112 86 177272 99874
rect 179612 86 179772 99874
rect 182112 86 182272 99874
rect 184612 86 184772 99874
rect 187112 86 187272 99874
rect 189612 86 189772 99874
rect 192112 86 192272 99874
rect 194612 86 194772 99874
rect 197112 86 197272 99874
rect 199612 86 199772 99874
rect 202112 86 202272 99874
rect 204612 86 204772 99874
rect 207112 86 207272 99874
rect 209612 86 209772 99874
rect 212112 86 212272 99874
rect 214612 86 214772 99874
rect 217112 86 217272 99874
rect 219612 86 219772 99874
rect 222112 86 222272 99874
rect 224612 86 224772 99874
rect 227112 86 227272 99874
rect 229612 86 229772 99874
rect 232112 86 232272 99874
rect 235016 416 235176 99544
rect 235346 86 235506 99874
<< obsm4 >>
rect 2002 99904 234094 99979
rect 2002 1317 2082 99904
rect 2302 1317 4582 99904
rect 4802 1317 7082 99904
rect 7302 1317 9582 99904
rect 9802 1317 12082 99904
rect 12302 1317 14582 99904
rect 14802 1317 17082 99904
rect 17302 1317 19582 99904
rect 19802 1317 22082 99904
rect 22302 1317 24582 99904
rect 24802 1317 27082 99904
rect 27302 1317 29582 99904
rect 29802 1317 32082 99904
rect 32302 1317 34582 99904
rect 34802 1317 37082 99904
rect 37302 1317 39582 99904
rect 39802 1317 42082 99904
rect 42302 1317 44582 99904
rect 44802 1317 47082 99904
rect 47302 1317 49582 99904
rect 49802 1317 52082 99904
rect 52302 1317 54582 99904
rect 54802 1317 57082 99904
rect 57302 1317 59582 99904
rect 59802 1317 62082 99904
rect 62302 1317 64582 99904
rect 64802 1317 67082 99904
rect 67302 1317 69582 99904
rect 69802 1317 72082 99904
rect 72302 1317 74582 99904
rect 74802 1317 77082 99904
rect 77302 1317 79582 99904
rect 79802 1317 82082 99904
rect 82302 1317 84582 99904
rect 84802 1317 87082 99904
rect 87302 1317 89582 99904
rect 89802 1317 92082 99904
rect 92302 1317 94582 99904
rect 94802 1317 97082 99904
rect 97302 1317 99582 99904
rect 99802 1317 102082 99904
rect 102302 1317 104582 99904
rect 104802 1317 107082 99904
rect 107302 1317 109582 99904
rect 109802 1317 112082 99904
rect 112302 1317 114582 99904
rect 114802 1317 117082 99904
rect 117302 1317 119582 99904
rect 119802 1317 122082 99904
rect 122302 1317 124582 99904
rect 124802 1317 127082 99904
rect 127302 1317 129582 99904
rect 129802 1317 132082 99904
rect 132302 1317 134582 99904
rect 134802 1317 137082 99904
rect 137302 1317 139582 99904
rect 139802 1317 142082 99904
rect 142302 1317 144582 99904
rect 144802 1317 147082 99904
rect 147302 1317 149582 99904
rect 149802 1317 152082 99904
rect 152302 1317 154582 99904
rect 154802 1317 157082 99904
rect 157302 1317 159582 99904
rect 159802 1317 162082 99904
rect 162302 1317 164582 99904
rect 164802 1317 167082 99904
rect 167302 1317 169582 99904
rect 169802 1317 172082 99904
rect 172302 1317 174582 99904
rect 174802 1317 177082 99904
rect 177302 1317 179582 99904
rect 179802 1317 182082 99904
rect 182302 1317 184582 99904
rect 184802 1317 187082 99904
rect 187302 1317 189582 99904
rect 189802 1317 192082 99904
rect 192302 1317 194582 99904
rect 194802 1317 197082 99904
rect 197302 1317 199582 99904
rect 199802 1317 202082 99904
rect 202302 1317 204582 99904
rect 204802 1317 207082 99904
rect 207302 1317 209582 99904
rect 209802 1317 212082 99904
rect 212302 1317 214582 99904
rect 214802 1317 217082 99904
rect 217302 1317 219582 99904
rect 219802 1317 222082 99904
rect 222302 1317 224582 99904
rect 224802 1317 227082 99904
rect 227302 1317 229582 99904
rect 229802 1317 232082 99904
rect 232302 1317 234094 99904
<< metal5 >>
rect -530 99714 235506 99874
rect -200 99384 235176 99544
rect -530 93761 235506 93921
rect -530 87261 235506 87421
rect -530 80761 235506 80921
rect -530 74261 235506 74421
rect -530 67761 235506 67921
rect -530 61261 235506 61421
rect -530 54761 235506 54921
rect -530 48261 235506 48421
rect -530 41761 235506 41921
rect -530 35261 235506 35421
rect -530 28761 235506 28921
rect -530 22261 235506 22421
rect -530 15761 235506 15921
rect -530 9261 235506 9421
rect -530 2761 235506 2921
rect -200 416 235176 576
rect -530 86 235506 246
<< obsm5 >>
rect 2330 99594 234102 99652
rect 2330 93971 234102 99334
rect 2330 87471 234102 93711
rect 2330 80971 234102 87211
rect 2330 74471 234102 80711
rect 2330 67971 234102 74211
rect 2330 61471 234102 67711
rect 2330 54971 234102 61211
rect 2330 48471 234102 54711
rect 2330 41971 234102 48211
rect 2330 35471 234102 41711
rect 2330 28971 234102 35211
rect 2330 22471 234102 28711
rect 2330 15971 234102 22211
rect 2330 9471 234102 15711
rect 2330 2971 234102 9211
rect 2330 1328 234102 2711
<< labels >>
rlabel metal4 s -200 416 -40 99544 4 VDD
port 1 nsew power bidirectional
rlabel metal5 s -200 416 235176 576 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s -200 99384 235176 99544 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 235016 416 235176 99544 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 2112 86 2272 99874 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 7112 86 7272 99874 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 12112 86 12272 99874 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 17112 86 17272 99874 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 22112 86 22272 99874 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 27112 86 27272 99874 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 32112 86 32272 99874 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 37112 86 37272 99874 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 42112 86 42272 99874 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 47112 86 47272 99874 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 52112 86 52272 99874 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 57112 86 57272 99874 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 62112 86 62272 99874 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 67112 86 67272 99874 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 72112 86 72272 99874 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 77112 86 77272 99874 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 82112 86 82272 99874 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 87112 86 87272 99874 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 92112 86 92272 99874 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 97112 86 97272 99874 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 102112 86 102272 99874 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 107112 86 107272 99874 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 112112 86 112272 99874 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 117112 86 117272 99874 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 122112 86 122272 99874 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 127112 86 127272 99874 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 132112 86 132272 99874 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 137112 86 137272 99874 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 142112 86 142272 99874 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 147112 86 147272 99874 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 152112 86 152272 99874 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 157112 86 157272 99874 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 162112 86 162272 99874 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 167112 86 167272 99874 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 172112 86 172272 99874 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 177112 86 177272 99874 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 182112 86 182272 99874 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 187112 86 187272 99874 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 192112 86 192272 99874 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 197112 86 197272 99874 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 202112 86 202272 99874 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 207112 86 207272 99874 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 212112 86 212272 99874 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 217112 86 217272 99874 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 222112 86 222272 99874 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 227112 86 227272 99874 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 232112 86 232272 99874 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s -530 2761 235506 2921 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s -530 15761 235506 15921 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s -530 28761 235506 28921 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s -530 41761 235506 41921 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s -530 54761 235506 54921 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s -530 67761 235506 67921 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s -530 80761 235506 80921 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s -530 93761 235506 93921 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s -530 86 -370 99874 4 VSS
port 2 nsew ground bidirectional
rlabel metal5 s -530 86 235506 246 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s -530 99714 235506 99874 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 235346 86 235506 99874 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 4612 86 4772 99874 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 9612 86 9772 99874 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 14612 86 14772 99874 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 19612 86 19772 99874 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 24612 86 24772 99874 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 29612 86 29772 99874 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 34612 86 34772 99874 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 39612 86 39772 99874 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 44612 86 44772 99874 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 49612 86 49772 99874 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 54612 86 54772 99874 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 59612 86 59772 99874 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 64612 86 64772 99874 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 69612 86 69772 99874 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 74612 86 74772 99874 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 79612 86 79772 99874 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 84612 86 84772 99874 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 89612 86 89772 99874 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 94612 86 94772 99874 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 99612 86 99772 99874 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 104612 86 104772 99874 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 109612 86 109772 99874 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 114612 86 114772 99874 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 119612 86 119772 99874 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 124612 86 124772 99874 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 129612 86 129772 99874 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 134612 86 134772 99874 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 139612 86 139772 99874 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 144612 86 144772 99874 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 149612 86 149772 99874 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 154612 86 154772 99874 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 159612 86 159772 99874 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 164612 86 164772 99874 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 169612 86 169772 99874 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 174612 86 174772 99874 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 179612 86 179772 99874 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 184612 86 184772 99874 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 189612 86 189772 99874 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 194612 86 194772 99874 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 199612 86 199772 99874 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 204612 86 204772 99874 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 209612 86 209772 99874 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 214612 86 214772 99874 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 219612 86 219772 99874 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 224612 86 224772 99874 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 229612 86 229772 99874 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s -530 9261 235506 9421 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s -530 22261 235506 22421 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s -530 35261 235506 35421 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s -530 48261 235506 48421 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s -530 61261 235506 61421 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s -530 74261 235506 74421 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s -530 87261 235506 87421 6 VSS
port 2 nsew ground bidirectional
rlabel metal3 s 234600 27188 235200 27244 6 core_clk
port 3 nsew signal input
rlabel metal2 s 50260 -200 50316 400 6 core_rstn
port 4 nsew signal input
rlabel metal3 s 234600 756 235200 812 6 debug_in
port 5 nsew signal input
rlabel metal3 s 234600 2212 235200 2268 6 debug_mode
port 6 nsew signal output
rlabel metal3 s 234600 3668 235200 3724 6 debug_oeb
port 7 nsew signal output
rlabel metal3 s 234600 5124 235200 5180 6 debug_out
port 8 nsew signal output
rlabel metal3 s 234600 81564 235200 81620 6 flash_clk
port 9 nsew signal output
rlabel metal3 s 234600 80108 235200 80164 6 flash_csb
port 10 nsew signal output
rlabel metal3 s 234600 83076 235200 83132 6 flash_io0_di
port 11 nsew signal input
rlabel metal3 s 234600 84532 235200 84588 6 flash_io0_do
port 12 nsew signal output
rlabel metal3 s 234600 85988 235200 86044 6 flash_io0_oeb
port 13 nsew signal output
rlabel metal3 s 234600 87444 235200 87500 6 flash_io1_di
port 14 nsew signal input
rlabel metal3 s 234600 88956 235200 89012 6 flash_io1_do
port 15 nsew signal output
rlabel metal3 s 234600 90412 235200 90468 6 flash_io1_oeb
port 16 nsew signal output
rlabel metal3 s 234600 91868 235200 91924 6 flash_io2_di
port 17 nsew signal input
rlabel metal3 s 234600 93324 235200 93380 6 flash_io2_do
port 18 nsew signal output
rlabel metal3 s 234600 94836 235200 94892 6 flash_io2_oeb
port 19 nsew signal output
rlabel metal3 s 234600 96292 235200 96348 6 flash_io3_di
port 20 nsew signal input
rlabel metal3 s 234600 97748 235200 97804 6 flash_io3_do
port 21 nsew signal output
rlabel metal3 s 234600 99204 235200 99260 6 flash_io3_oeb
port 22 nsew signal output
rlabel metal2 s 16716 -200 16772 400 6 gpio_in_pad
port 23 nsew signal input
rlabel metal2 s 83860 -200 83916 400 6 gpio_inenb_pad
port 24 nsew signal output
rlabel metal2 s 117404 -200 117460 400 6 gpio_mode0_pad
port 25 nsew signal output
rlabel metal2 s 151004 -200 151060 400 6 gpio_mode1_pad
port 26 nsew signal output
rlabel metal2 s 184548 -200 184604 400 6 gpio_out_pad
port 27 nsew signal output
rlabel metal2 s 218148 -200 218204 400 6 gpio_outenb_pad
port 28 nsew signal output
rlabel metal3 s 234600 28644 235200 28700 6 hk_ack_i
port 29 nsew signal input
rlabel metal3 s 234600 31612 235200 31668 6 hk_cyc_o
port 30 nsew signal output
rlabel metal3 s 234600 33068 235200 33124 6 hk_dat_i[0]
port 31 nsew signal input
rlabel metal3 s 234600 47796 235200 47852 6 hk_dat_i[10]
port 32 nsew signal input
rlabel metal3 s 234600 49252 235200 49308 6 hk_dat_i[11]
port 33 nsew signal input
rlabel metal3 s 234600 50708 235200 50764 6 hk_dat_i[12]
port 34 nsew signal input
rlabel metal3 s 234600 52164 235200 52220 6 hk_dat_i[13]
port 35 nsew signal input
rlabel metal3 s 234600 53676 235200 53732 6 hk_dat_i[14]
port 36 nsew signal input
rlabel metal3 s 234600 55132 235200 55188 6 hk_dat_i[15]
port 37 nsew signal input
rlabel metal3 s 234600 56588 235200 56644 6 hk_dat_i[16]
port 38 nsew signal input
rlabel metal3 s 234600 58044 235200 58100 6 hk_dat_i[17]
port 39 nsew signal input
rlabel metal3 s 234600 59556 235200 59612 6 hk_dat_i[18]
port 40 nsew signal input
rlabel metal3 s 234600 61012 235200 61068 6 hk_dat_i[19]
port 41 nsew signal input
rlabel metal3 s 234600 34524 235200 34580 6 hk_dat_i[1]
port 42 nsew signal input
rlabel metal3 s 234600 62468 235200 62524 6 hk_dat_i[20]
port 43 nsew signal input
rlabel metal3 s 234600 63924 235200 63980 6 hk_dat_i[21]
port 44 nsew signal input
rlabel metal3 s 234600 65436 235200 65492 6 hk_dat_i[22]
port 45 nsew signal input
rlabel metal3 s 234600 66892 235200 66948 6 hk_dat_i[23]
port 46 nsew signal input
rlabel metal3 s 234600 68348 235200 68404 6 hk_dat_i[24]
port 47 nsew signal input
rlabel metal3 s 234600 69804 235200 69860 6 hk_dat_i[25]
port 48 nsew signal input
rlabel metal3 s 234600 71316 235200 71372 6 hk_dat_i[26]
port 49 nsew signal input
rlabel metal3 s 234600 72772 235200 72828 6 hk_dat_i[27]
port 50 nsew signal input
rlabel metal3 s 234600 74228 235200 74284 6 hk_dat_i[28]
port 51 nsew signal input
rlabel metal3 s 234600 75684 235200 75740 6 hk_dat_i[29]
port 52 nsew signal input
rlabel metal3 s 234600 36036 235200 36092 6 hk_dat_i[2]
port 53 nsew signal input
rlabel metal3 s 234600 77196 235200 77252 6 hk_dat_i[30]
port 54 nsew signal input
rlabel metal3 s 234600 78652 235200 78708 6 hk_dat_i[31]
port 55 nsew signal input
rlabel metal3 s 234600 37492 235200 37548 6 hk_dat_i[3]
port 56 nsew signal input
rlabel metal3 s 234600 38948 235200 39004 6 hk_dat_i[4]
port 57 nsew signal input
rlabel metal3 s 234600 40404 235200 40460 6 hk_dat_i[5]
port 58 nsew signal input
rlabel metal3 s 234600 41916 235200 41972 6 hk_dat_i[6]
port 59 nsew signal input
rlabel metal3 s 234600 43372 235200 43428 6 hk_dat_i[7]
port 60 nsew signal input
rlabel metal3 s 234600 44828 235200 44884 6 hk_dat_i[8]
port 61 nsew signal input
rlabel metal3 s 234600 46284 235200 46340 6 hk_dat_i[9]
port 62 nsew signal input
rlabel metal3 s 234600 30156 235200 30212 6 hk_stb_o
port 63 nsew signal output
rlabel metal2 s 233324 99600 233380 100200 6 irq[0]
port 64 nsew signal input
rlabel metal2 s 233996 99600 234052 100200 6 irq[1]
port 65 nsew signal input
rlabel metal2 s 234612 99600 234668 100200 6 irq[2]
port 66 nsew signal input
rlabel metal3 s 234600 11004 235200 11060 6 irq[3]
port 67 nsew signal input
rlabel metal3 s 234600 9548 235200 9604 6 irq[4]
port 68 nsew signal input
rlabel metal3 s 234600 8092 235200 8148 6 irq[5]
port 69 nsew signal input
rlabel metal2 s 123172 99600 123228 100200 6 la_iena[0]
port 70 nsew signal output
rlabel metal2 s 129612 99600 129668 100200 6 la_iena[10]
port 71 nsew signal output
rlabel metal2 s 130228 99600 130284 100200 6 la_iena[11]
port 72 nsew signal output
rlabel metal2 s 130844 99600 130900 100200 6 la_iena[12]
port 73 nsew signal output
rlabel metal2 s 131516 99600 131572 100200 6 la_iena[13]
port 74 nsew signal output
rlabel metal2 s 132132 99600 132188 100200 6 la_iena[14]
port 75 nsew signal output
rlabel metal2 s 132804 99600 132860 100200 6 la_iena[15]
port 76 nsew signal output
rlabel metal2 s 133420 99600 133476 100200 6 la_iena[16]
port 77 nsew signal output
rlabel metal2 s 134092 99600 134148 100200 6 la_iena[17]
port 78 nsew signal output
rlabel metal2 s 134708 99600 134764 100200 6 la_iena[18]
port 79 nsew signal output
rlabel metal2 s 135324 99600 135380 100200 6 la_iena[19]
port 80 nsew signal output
rlabel metal2 s 123844 99600 123900 100200 6 la_iena[1]
port 81 nsew signal output
rlabel metal2 s 135996 99600 136052 100200 6 la_iena[20]
port 82 nsew signal output
rlabel metal2 s 136612 99600 136668 100200 6 la_iena[21]
port 83 nsew signal output
rlabel metal2 s 137284 99600 137340 100200 6 la_iena[22]
port 84 nsew signal output
rlabel metal2 s 137900 99600 137956 100200 6 la_iena[23]
port 85 nsew signal output
rlabel metal2 s 138572 99600 138628 100200 6 la_iena[24]
port 86 nsew signal output
rlabel metal2 s 139188 99600 139244 100200 6 la_iena[25]
port 87 nsew signal output
rlabel metal2 s 139860 99600 139916 100200 6 la_iena[26]
port 88 nsew signal output
rlabel metal2 s 140476 99600 140532 100200 6 la_iena[27]
port 89 nsew signal output
rlabel metal2 s 141092 99600 141148 100200 6 la_iena[28]
port 90 nsew signal output
rlabel metal2 s 141764 99600 141820 100200 6 la_iena[29]
port 91 nsew signal output
rlabel metal2 s 124460 99600 124516 100200 6 la_iena[2]
port 92 nsew signal output
rlabel metal2 s 142380 99600 142436 100200 6 la_iena[30]
port 93 nsew signal output
rlabel metal2 s 143052 99600 143108 100200 6 la_iena[31]
port 94 nsew signal output
rlabel metal2 s 143668 99600 143724 100200 6 la_iena[32]
port 95 nsew signal output
rlabel metal2 s 144340 99600 144396 100200 6 la_iena[33]
port 96 nsew signal output
rlabel metal2 s 144956 99600 145012 100200 6 la_iena[34]
port 97 nsew signal output
rlabel metal2 s 145572 99600 145628 100200 6 la_iena[35]
port 98 nsew signal output
rlabel metal2 s 146244 99600 146300 100200 6 la_iena[36]
port 99 nsew signal output
rlabel metal2 s 146860 99600 146916 100200 6 la_iena[37]
port 100 nsew signal output
rlabel metal2 s 147532 99600 147588 100200 6 la_iena[38]
port 101 nsew signal output
rlabel metal2 s 148148 99600 148204 100200 6 la_iena[39]
port 102 nsew signal output
rlabel metal2 s 125132 99600 125188 100200 6 la_iena[3]
port 103 nsew signal output
rlabel metal2 s 148820 99600 148876 100200 6 la_iena[40]
port 104 nsew signal output
rlabel metal2 s 149436 99600 149492 100200 6 la_iena[41]
port 105 nsew signal output
rlabel metal2 s 150108 99600 150164 100200 6 la_iena[42]
port 106 nsew signal output
rlabel metal2 s 150724 99600 150780 100200 6 la_iena[43]
port 107 nsew signal output
rlabel metal2 s 151340 99600 151396 100200 6 la_iena[44]
port 108 nsew signal output
rlabel metal2 s 152012 99600 152068 100200 6 la_iena[45]
port 109 nsew signal output
rlabel metal2 s 152628 99600 152684 100200 6 la_iena[46]
port 110 nsew signal output
rlabel metal2 s 153300 99600 153356 100200 6 la_iena[47]
port 111 nsew signal output
rlabel metal2 s 153916 99600 153972 100200 6 la_iena[48]
port 112 nsew signal output
rlabel metal2 s 154588 99600 154644 100200 6 la_iena[49]
port 113 nsew signal output
rlabel metal2 s 125748 99600 125804 100200 6 la_iena[4]
port 114 nsew signal output
rlabel metal2 s 155204 99600 155260 100200 6 la_iena[50]
port 115 nsew signal output
rlabel metal2 s 155820 99600 155876 100200 6 la_iena[51]
port 116 nsew signal output
rlabel metal2 s 156492 99600 156548 100200 6 la_iena[52]
port 117 nsew signal output
rlabel metal2 s 157108 99600 157164 100200 6 la_iena[53]
port 118 nsew signal output
rlabel metal2 s 157780 99600 157836 100200 6 la_iena[54]
port 119 nsew signal output
rlabel metal2 s 158396 99600 158452 100200 6 la_iena[55]
port 120 nsew signal output
rlabel metal2 s 159068 99600 159124 100200 6 la_iena[56]
port 121 nsew signal output
rlabel metal2 s 159684 99600 159740 100200 6 la_iena[57]
port 122 nsew signal output
rlabel metal2 s 160300 99600 160356 100200 6 la_iena[58]
port 123 nsew signal output
rlabel metal2 s 160972 99600 161028 100200 6 la_iena[59]
port 124 nsew signal output
rlabel metal2 s 126364 99600 126420 100200 6 la_iena[5]
port 125 nsew signal output
rlabel metal2 s 161588 99600 161644 100200 6 la_iena[60]
port 126 nsew signal output
rlabel metal2 s 162260 99600 162316 100200 6 la_iena[61]
port 127 nsew signal output
rlabel metal2 s 162876 99600 162932 100200 6 la_iena[62]
port 128 nsew signal output
rlabel metal2 s 163548 99600 163604 100200 6 la_iena[63]
port 129 nsew signal output
rlabel metal2 s 127036 99600 127092 100200 6 la_iena[6]
port 130 nsew signal output
rlabel metal2 s 127652 99600 127708 100200 6 la_iena[7]
port 131 nsew signal output
rlabel metal2 s 128324 99600 128380 100200 6 la_iena[8]
port 132 nsew signal output
rlabel metal2 s 128940 99600 128996 100200 6 la_iena[9]
port 133 nsew signal output
rlabel metal2 s 252 99600 308 100200 6 la_input[0]
port 134 nsew signal input
rlabel metal2 s 6636 99600 6692 100200 6 la_input[10]
port 135 nsew signal input
rlabel metal2 s 7252 99600 7308 100200 6 la_input[11]
port 136 nsew signal input
rlabel metal2 s 7924 99600 7980 100200 6 la_input[12]
port 137 nsew signal input
rlabel metal2 s 8540 99600 8596 100200 6 la_input[13]
port 138 nsew signal input
rlabel metal2 s 9212 99600 9268 100200 6 la_input[14]
port 139 nsew signal input
rlabel metal2 s 9828 99600 9884 100200 6 la_input[15]
port 140 nsew signal input
rlabel metal2 s 10444 99600 10500 100200 6 la_input[16]
port 141 nsew signal input
rlabel metal2 s 11116 99600 11172 100200 6 la_input[17]
port 142 nsew signal input
rlabel metal2 s 11732 99600 11788 100200 6 la_input[18]
port 143 nsew signal input
rlabel metal2 s 12404 99600 12460 100200 6 la_input[19]
port 144 nsew signal input
rlabel metal2 s 868 99600 924 100200 6 la_input[1]
port 145 nsew signal input
rlabel metal2 s 13020 99600 13076 100200 6 la_input[20]
port 146 nsew signal input
rlabel metal2 s 13692 99600 13748 100200 6 la_input[21]
port 147 nsew signal input
rlabel metal2 s 14308 99600 14364 100200 6 la_input[22]
port 148 nsew signal input
rlabel metal2 s 14980 99600 15036 100200 6 la_input[23]
port 149 nsew signal input
rlabel metal2 s 15596 99600 15652 100200 6 la_input[24]
port 150 nsew signal input
rlabel metal2 s 16212 99600 16268 100200 6 la_input[25]
port 151 nsew signal input
rlabel metal2 s 16884 99600 16940 100200 6 la_input[26]
port 152 nsew signal input
rlabel metal2 s 17500 99600 17556 100200 6 la_input[27]
port 153 nsew signal input
rlabel metal2 s 18172 99600 18228 100200 6 la_input[28]
port 154 nsew signal input
rlabel metal2 s 18788 99600 18844 100200 6 la_input[29]
port 155 nsew signal input
rlabel metal2 s 1484 99600 1540 100200 6 la_input[2]
port 156 nsew signal input
rlabel metal2 s 19460 99600 19516 100200 6 la_input[30]
port 157 nsew signal input
rlabel metal2 s 20076 99600 20132 100200 6 la_input[31]
port 158 nsew signal input
rlabel metal2 s 20692 99600 20748 100200 6 la_input[32]
port 159 nsew signal input
rlabel metal2 s 21364 99600 21420 100200 6 la_input[33]
port 160 nsew signal input
rlabel metal2 s 21980 99600 22036 100200 6 la_input[34]
port 161 nsew signal input
rlabel metal2 s 22652 99600 22708 100200 6 la_input[35]
port 162 nsew signal input
rlabel metal2 s 23268 99600 23324 100200 6 la_input[36]
port 163 nsew signal input
rlabel metal2 s 23940 99600 23996 100200 6 la_input[37]
port 164 nsew signal input
rlabel metal2 s 24556 99600 24612 100200 6 la_input[38]
port 165 nsew signal input
rlabel metal2 s 25228 99600 25284 100200 6 la_input[39]
port 166 nsew signal input
rlabel metal2 s 2156 99600 2212 100200 6 la_input[3]
port 167 nsew signal input
rlabel metal2 s 25844 99600 25900 100200 6 la_input[40]
port 168 nsew signal input
rlabel metal2 s 26460 99600 26516 100200 6 la_input[41]
port 169 nsew signal input
rlabel metal2 s 27132 99600 27188 100200 6 la_input[42]
port 170 nsew signal input
rlabel metal2 s 27748 99600 27804 100200 6 la_input[43]
port 171 nsew signal input
rlabel metal2 s 28420 99600 28476 100200 6 la_input[44]
port 172 nsew signal input
rlabel metal2 s 29036 99600 29092 100200 6 la_input[45]
port 173 nsew signal input
rlabel metal2 s 29708 99600 29764 100200 6 la_input[46]
port 174 nsew signal input
rlabel metal2 s 30324 99600 30380 100200 6 la_input[47]
port 175 nsew signal input
rlabel metal2 s 30940 99600 30996 100200 6 la_input[48]
port 176 nsew signal input
rlabel metal2 s 31612 99600 31668 100200 6 la_input[49]
port 177 nsew signal input
rlabel metal2 s 2772 99600 2828 100200 6 la_input[4]
port 178 nsew signal input
rlabel metal2 s 32228 99600 32284 100200 6 la_input[50]
port 179 nsew signal input
rlabel metal2 s 32900 99600 32956 100200 6 la_input[51]
port 180 nsew signal input
rlabel metal2 s 33516 99600 33572 100200 6 la_input[52]
port 181 nsew signal input
rlabel metal2 s 34188 99600 34244 100200 6 la_input[53]
port 182 nsew signal input
rlabel metal2 s 34804 99600 34860 100200 6 la_input[54]
port 183 nsew signal input
rlabel metal2 s 35420 99600 35476 100200 6 la_input[55]
port 184 nsew signal input
rlabel metal2 s 36092 99600 36148 100200 6 la_input[56]
port 185 nsew signal input
rlabel metal2 s 36708 99600 36764 100200 6 la_input[57]
port 186 nsew signal input
rlabel metal2 s 37380 99600 37436 100200 6 la_input[58]
port 187 nsew signal input
rlabel metal2 s 37996 99600 38052 100200 6 la_input[59]
port 188 nsew signal input
rlabel metal2 s 3444 99600 3500 100200 6 la_input[5]
port 189 nsew signal input
rlabel metal2 s 38668 99600 38724 100200 6 la_input[60]
port 190 nsew signal input
rlabel metal2 s 39284 99600 39340 100200 6 la_input[61]
port 191 nsew signal input
rlabel metal2 s 39956 99600 40012 100200 6 la_input[62]
port 192 nsew signal input
rlabel metal2 s 40572 99600 40628 100200 6 la_input[63]
port 193 nsew signal input
rlabel metal2 s 4060 99600 4116 100200 6 la_input[6]
port 194 nsew signal input
rlabel metal2 s 4732 99600 4788 100200 6 la_input[7]
port 195 nsew signal input
rlabel metal2 s 5348 99600 5404 100200 6 la_input[8]
port 196 nsew signal input
rlabel metal2 s 5964 99600 6020 100200 6 la_input[9]
port 197 nsew signal input
rlabel metal2 s 82180 99600 82236 100200 6 la_oenb[0]
port 198 nsew signal output
rlabel metal2 s 88620 99600 88676 100200 6 la_oenb[10]
port 199 nsew signal output
rlabel metal2 s 89236 99600 89292 100200 6 la_oenb[11]
port 200 nsew signal output
rlabel metal2 s 89908 99600 89964 100200 6 la_oenb[12]
port 201 nsew signal output
rlabel metal2 s 90524 99600 90580 100200 6 la_oenb[13]
port 202 nsew signal output
rlabel metal2 s 91140 99600 91196 100200 6 la_oenb[14]
port 203 nsew signal output
rlabel metal2 s 91812 99600 91868 100200 6 la_oenb[15]
port 204 nsew signal output
rlabel metal2 s 92428 99600 92484 100200 6 la_oenb[16]
port 205 nsew signal output
rlabel metal2 s 93100 99600 93156 100200 6 la_oenb[17]
port 206 nsew signal output
rlabel metal2 s 93716 99600 93772 100200 6 la_oenb[18]
port 207 nsew signal output
rlabel metal2 s 94388 99600 94444 100200 6 la_oenb[19]
port 208 nsew signal output
rlabel metal2 s 82852 99600 82908 100200 6 la_oenb[1]
port 209 nsew signal output
rlabel metal2 s 95004 99600 95060 100200 6 la_oenb[20]
port 210 nsew signal output
rlabel metal2 s 95620 99600 95676 100200 6 la_oenb[21]
port 211 nsew signal output
rlabel metal2 s 96292 99600 96348 100200 6 la_oenb[22]
port 212 nsew signal output
rlabel metal2 s 96908 99600 96964 100200 6 la_oenb[23]
port 213 nsew signal output
rlabel metal2 s 97580 99600 97636 100200 6 la_oenb[24]
port 214 nsew signal output
rlabel metal2 s 98196 99600 98252 100200 6 la_oenb[25]
port 215 nsew signal output
rlabel metal2 s 98868 99600 98924 100200 6 la_oenb[26]
port 216 nsew signal output
rlabel metal2 s 99484 99600 99540 100200 6 la_oenb[27]
port 217 nsew signal output
rlabel metal2 s 100156 99600 100212 100200 6 la_oenb[28]
port 218 nsew signal output
rlabel metal2 s 100772 99600 100828 100200 6 la_oenb[29]
port 219 nsew signal output
rlabel metal2 s 83468 99600 83524 100200 6 la_oenb[2]
port 220 nsew signal output
rlabel metal2 s 101388 99600 101444 100200 6 la_oenb[30]
port 221 nsew signal output
rlabel metal2 s 102060 99600 102116 100200 6 la_oenb[31]
port 222 nsew signal output
rlabel metal2 s 102676 99600 102732 100200 6 la_oenb[32]
port 223 nsew signal output
rlabel metal2 s 103348 99600 103404 100200 6 la_oenb[33]
port 224 nsew signal output
rlabel metal2 s 103964 99600 104020 100200 6 la_oenb[34]
port 225 nsew signal output
rlabel metal2 s 104636 99600 104692 100200 6 la_oenb[35]
port 226 nsew signal output
rlabel metal2 s 105252 99600 105308 100200 6 la_oenb[36]
port 227 nsew signal output
rlabel metal2 s 105868 99600 105924 100200 6 la_oenb[37]
port 228 nsew signal output
rlabel metal2 s 106540 99600 106596 100200 6 la_oenb[38]
port 229 nsew signal output
rlabel metal2 s 107156 99600 107212 100200 6 la_oenb[39]
port 230 nsew signal output
rlabel metal2 s 84140 99600 84196 100200 6 la_oenb[3]
port 231 nsew signal output
rlabel metal2 s 107828 99600 107884 100200 6 la_oenb[40]
port 232 nsew signal output
rlabel metal2 s 108444 99600 108500 100200 6 la_oenb[41]
port 233 nsew signal output
rlabel metal2 s 109116 99600 109172 100200 6 la_oenb[42]
port 234 nsew signal output
rlabel metal2 s 109732 99600 109788 100200 6 la_oenb[43]
port 235 nsew signal output
rlabel metal2 s 110348 99600 110404 100200 6 la_oenb[44]
port 236 nsew signal output
rlabel metal2 s 111020 99600 111076 100200 6 la_oenb[45]
port 237 nsew signal output
rlabel metal2 s 111636 99600 111692 100200 6 la_oenb[46]
port 238 nsew signal output
rlabel metal2 s 112308 99600 112364 100200 6 la_oenb[47]
port 239 nsew signal output
rlabel metal2 s 112924 99600 112980 100200 6 la_oenb[48]
port 240 nsew signal output
rlabel metal2 s 113596 99600 113652 100200 6 la_oenb[49]
port 241 nsew signal output
rlabel metal2 s 84756 99600 84812 100200 6 la_oenb[4]
port 242 nsew signal output
rlabel metal2 s 114212 99600 114268 100200 6 la_oenb[50]
port 243 nsew signal output
rlabel metal2 s 114884 99600 114940 100200 6 la_oenb[51]
port 244 nsew signal output
rlabel metal2 s 115500 99600 115556 100200 6 la_oenb[52]
port 245 nsew signal output
rlabel metal2 s 116116 99600 116172 100200 6 la_oenb[53]
port 246 nsew signal output
rlabel metal2 s 116788 99600 116844 100200 6 la_oenb[54]
port 247 nsew signal output
rlabel metal2 s 117404 99600 117460 100200 6 la_oenb[55]
port 248 nsew signal output
rlabel metal2 s 118076 99600 118132 100200 6 la_oenb[56]
port 249 nsew signal output
rlabel metal2 s 118692 99600 118748 100200 6 la_oenb[57]
port 250 nsew signal output
rlabel metal2 s 119364 99600 119420 100200 6 la_oenb[58]
port 251 nsew signal output
rlabel metal2 s 119980 99600 120036 100200 6 la_oenb[59]
port 252 nsew signal output
rlabel metal2 s 85372 99600 85428 100200 6 la_oenb[5]
port 253 nsew signal output
rlabel metal2 s 120596 99600 120652 100200 6 la_oenb[60]
port 254 nsew signal output
rlabel metal2 s 121268 99600 121324 100200 6 la_oenb[61]
port 255 nsew signal output
rlabel metal2 s 121884 99600 121940 100200 6 la_oenb[62]
port 256 nsew signal output
rlabel metal2 s 122556 99600 122612 100200 6 la_oenb[63]
port 257 nsew signal output
rlabel metal2 s 86044 99600 86100 100200 6 la_oenb[6]
port 258 nsew signal output
rlabel metal2 s 86660 99600 86716 100200 6 la_oenb[7]
port 259 nsew signal output
rlabel metal2 s 87332 99600 87388 100200 6 la_oenb[8]
port 260 nsew signal output
rlabel metal2 s 87948 99600 88004 100200 6 la_oenb[9]
port 261 nsew signal output
rlabel metal2 s 41188 99600 41244 100200 6 la_output[0]
port 262 nsew signal output
rlabel metal2 s 47628 99600 47684 100200 6 la_output[10]
port 263 nsew signal output
rlabel metal2 s 48244 99600 48300 100200 6 la_output[11]
port 264 nsew signal output
rlabel metal2 s 48916 99600 48972 100200 6 la_output[12]
port 265 nsew signal output
rlabel metal2 s 49532 99600 49588 100200 6 la_output[13]
port 266 nsew signal output
rlabel metal2 s 50204 99600 50260 100200 6 la_output[14]
port 267 nsew signal output
rlabel metal2 s 50820 99600 50876 100200 6 la_output[15]
port 268 nsew signal output
rlabel metal2 s 51436 99600 51492 100200 6 la_output[16]
port 269 nsew signal output
rlabel metal2 s 52108 99600 52164 100200 6 la_output[17]
port 270 nsew signal output
rlabel metal2 s 52724 99600 52780 100200 6 la_output[18]
port 271 nsew signal output
rlabel metal2 s 53396 99600 53452 100200 6 la_output[19]
port 272 nsew signal output
rlabel metal2 s 41860 99600 41916 100200 6 la_output[1]
port 273 nsew signal output
rlabel metal2 s 54012 99600 54068 100200 6 la_output[20]
port 274 nsew signal output
rlabel metal2 s 54684 99600 54740 100200 6 la_output[21]
port 275 nsew signal output
rlabel metal2 s 55300 99600 55356 100200 6 la_output[22]
port 276 nsew signal output
rlabel metal2 s 55916 99600 55972 100200 6 la_output[23]
port 277 nsew signal output
rlabel metal2 s 56588 99600 56644 100200 6 la_output[24]
port 278 nsew signal output
rlabel metal2 s 57204 99600 57260 100200 6 la_output[25]
port 279 nsew signal output
rlabel metal2 s 57876 99600 57932 100200 6 la_output[26]
port 280 nsew signal output
rlabel metal2 s 58492 99600 58548 100200 6 la_output[27]
port 281 nsew signal output
rlabel metal2 s 59164 99600 59220 100200 6 la_output[28]
port 282 nsew signal output
rlabel metal2 s 59780 99600 59836 100200 6 la_output[29]
port 283 nsew signal output
rlabel metal2 s 42476 99600 42532 100200 6 la_output[2]
port 284 nsew signal output
rlabel metal2 s 60396 99600 60452 100200 6 la_output[30]
port 285 nsew signal output
rlabel metal2 s 61068 99600 61124 100200 6 la_output[31]
port 286 nsew signal output
rlabel metal2 s 61684 99600 61740 100200 6 la_output[32]
port 287 nsew signal output
rlabel metal2 s 62356 99600 62412 100200 6 la_output[33]
port 288 nsew signal output
rlabel metal2 s 62972 99600 63028 100200 6 la_output[34]
port 289 nsew signal output
rlabel metal2 s 63644 99600 63700 100200 6 la_output[35]
port 290 nsew signal output
rlabel metal2 s 64260 99600 64316 100200 6 la_output[36]
port 291 nsew signal output
rlabel metal2 s 64932 99600 64988 100200 6 la_output[37]
port 292 nsew signal output
rlabel metal2 s 65548 99600 65604 100200 6 la_output[38]
port 293 nsew signal output
rlabel metal2 s 66164 99600 66220 100200 6 la_output[39]
port 294 nsew signal output
rlabel metal2 s 43148 99600 43204 100200 6 la_output[3]
port 295 nsew signal output
rlabel metal2 s 66836 99600 66892 100200 6 la_output[40]
port 296 nsew signal output
rlabel metal2 s 67452 99600 67508 100200 6 la_output[41]
port 297 nsew signal output
rlabel metal2 s 68124 99600 68180 100200 6 la_output[42]
port 298 nsew signal output
rlabel metal2 s 68740 99600 68796 100200 6 la_output[43]
port 299 nsew signal output
rlabel metal2 s 69412 99600 69468 100200 6 la_output[44]
port 300 nsew signal output
rlabel metal2 s 70028 99600 70084 100200 6 la_output[45]
port 301 nsew signal output
rlabel metal2 s 70644 99600 70700 100200 6 la_output[46]
port 302 nsew signal output
rlabel metal2 s 71316 99600 71372 100200 6 la_output[47]
port 303 nsew signal output
rlabel metal2 s 71932 99600 71988 100200 6 la_output[48]
port 304 nsew signal output
rlabel metal2 s 72604 99600 72660 100200 6 la_output[49]
port 305 nsew signal output
rlabel metal2 s 43764 99600 43820 100200 6 la_output[4]
port 306 nsew signal output
rlabel metal2 s 73220 99600 73276 100200 6 la_output[50]
port 307 nsew signal output
rlabel metal2 s 73892 99600 73948 100200 6 la_output[51]
port 308 nsew signal output
rlabel metal2 s 74508 99600 74564 100200 6 la_output[52]
port 309 nsew signal output
rlabel metal2 s 75180 99600 75236 100200 6 la_output[53]
port 310 nsew signal output
rlabel metal2 s 75796 99600 75852 100200 6 la_output[54]
port 311 nsew signal output
rlabel metal2 s 76412 99600 76468 100200 6 la_output[55]
port 312 nsew signal output
rlabel metal2 s 77084 99600 77140 100200 6 la_output[56]
port 313 nsew signal output
rlabel metal2 s 77700 99600 77756 100200 6 la_output[57]
port 314 nsew signal output
rlabel metal2 s 78372 99600 78428 100200 6 la_output[58]
port 315 nsew signal output
rlabel metal2 s 78988 99600 79044 100200 6 la_output[59]
port 316 nsew signal output
rlabel metal2 s 44436 99600 44492 100200 6 la_output[5]
port 317 nsew signal output
rlabel metal2 s 79660 99600 79716 100200 6 la_output[60]
port 318 nsew signal output
rlabel metal2 s 80276 99600 80332 100200 6 la_output[61]
port 319 nsew signal output
rlabel metal2 s 80892 99600 80948 100200 6 la_output[62]
port 320 nsew signal output
rlabel metal2 s 81564 99600 81620 100200 6 la_output[63]
port 321 nsew signal output
rlabel metal2 s 45052 99600 45108 100200 6 la_output[6]
port 322 nsew signal output
rlabel metal2 s 45668 99600 45724 100200 6 la_output[7]
port 323 nsew signal output
rlabel metal2 s 46340 99600 46396 100200 6 la_output[8]
port 324 nsew signal output
rlabel metal2 s 46956 99600 47012 100200 6 la_output[9]
port 325 nsew signal output
rlabel metal2 s 232036 99600 232092 100200 6 mprj_ack_i
port 326 nsew signal input
rlabel metal2 s 189140 99600 189196 100200 6 mprj_adr_o[0]
port 327 nsew signal output
rlabel metal2 s 195524 99600 195580 100200 6 mprj_adr_o[10]
port 328 nsew signal output
rlabel metal2 s 196196 99600 196252 100200 6 mprj_adr_o[11]
port 329 nsew signal output
rlabel metal2 s 196812 99600 196868 100200 6 mprj_adr_o[12]
port 330 nsew signal output
rlabel metal2 s 197484 99600 197540 100200 6 mprj_adr_o[13]
port 331 nsew signal output
rlabel metal2 s 198100 99600 198156 100200 6 mprj_adr_o[14]
port 332 nsew signal output
rlabel metal2 s 198772 99600 198828 100200 6 mprj_adr_o[15]
port 333 nsew signal output
rlabel metal2 s 199388 99600 199444 100200 6 mprj_adr_o[16]
port 334 nsew signal output
rlabel metal2 s 200060 99600 200116 100200 6 mprj_adr_o[17]
port 335 nsew signal output
rlabel metal2 s 200676 99600 200732 100200 6 mprj_adr_o[18]
port 336 nsew signal output
rlabel metal2 s 201292 99600 201348 100200 6 mprj_adr_o[19]
port 337 nsew signal output
rlabel metal2 s 189812 99600 189868 100200 6 mprj_adr_o[1]
port 338 nsew signal output
rlabel metal2 s 201964 99600 202020 100200 6 mprj_adr_o[20]
port 339 nsew signal output
rlabel metal2 s 202580 99600 202636 100200 6 mprj_adr_o[21]
port 340 nsew signal output
rlabel metal2 s 203252 99600 203308 100200 6 mprj_adr_o[22]
port 341 nsew signal output
rlabel metal2 s 203868 99600 203924 100200 6 mprj_adr_o[23]
port 342 nsew signal output
rlabel metal2 s 204540 99600 204596 100200 6 mprj_adr_o[24]
port 343 nsew signal output
rlabel metal2 s 205156 99600 205212 100200 6 mprj_adr_o[25]
port 344 nsew signal output
rlabel metal2 s 205772 99600 205828 100200 6 mprj_adr_o[26]
port 345 nsew signal output
rlabel metal2 s 206444 99600 206500 100200 6 mprj_adr_o[27]
port 346 nsew signal output
rlabel metal2 s 207060 99600 207116 100200 6 mprj_adr_o[28]
port 347 nsew signal output
rlabel metal2 s 207732 99600 207788 100200 6 mprj_adr_o[29]
port 348 nsew signal output
rlabel metal2 s 190428 99600 190484 100200 6 mprj_adr_o[2]
port 349 nsew signal output
rlabel metal2 s 208348 99600 208404 100200 6 mprj_adr_o[30]
port 350 nsew signal output
rlabel metal2 s 209020 99600 209076 100200 6 mprj_adr_o[31]
port 351 nsew signal output
rlabel metal2 s 191044 99600 191100 100200 6 mprj_adr_o[3]
port 352 nsew signal output
rlabel metal2 s 191716 99600 191772 100200 6 mprj_adr_o[4]
port 353 nsew signal output
rlabel metal2 s 192332 99600 192388 100200 6 mprj_adr_o[5]
port 354 nsew signal output
rlabel metal2 s 193004 99600 193060 100200 6 mprj_adr_o[6]
port 355 nsew signal output
rlabel metal2 s 193620 99600 193676 100200 6 mprj_adr_o[7]
port 356 nsew signal output
rlabel metal2 s 194292 99600 194348 100200 6 mprj_adr_o[8]
port 357 nsew signal output
rlabel metal2 s 194908 99600 194964 100200 6 mprj_adr_o[9]
port 358 nsew signal output
rlabel metal2 s 230748 99600 230804 100200 6 mprj_cyc_o
port 359 nsew signal output
rlabel metal2 s 164164 99600 164220 100200 6 mprj_dat_i[0]
port 360 nsew signal input
rlabel metal2 s 170548 99600 170604 100200 6 mprj_dat_i[10]
port 361 nsew signal input
rlabel metal2 s 171220 99600 171276 100200 6 mprj_dat_i[11]
port 362 nsew signal input
rlabel metal2 s 171836 99600 171892 100200 6 mprj_dat_i[12]
port 363 nsew signal input
rlabel metal2 s 172508 99600 172564 100200 6 mprj_dat_i[13]
port 364 nsew signal input
rlabel metal2 s 173124 99600 173180 100200 6 mprj_dat_i[14]
port 365 nsew signal input
rlabel metal2 s 173796 99600 173852 100200 6 mprj_dat_i[15]
port 366 nsew signal input
rlabel metal2 s 174412 99600 174468 100200 6 mprj_dat_i[16]
port 367 nsew signal input
rlabel metal2 s 175084 99600 175140 100200 6 mprj_dat_i[17]
port 368 nsew signal input
rlabel metal2 s 175700 99600 175756 100200 6 mprj_dat_i[18]
port 369 nsew signal input
rlabel metal2 s 176316 99600 176372 100200 6 mprj_dat_i[19]
port 370 nsew signal input
rlabel metal2 s 164836 99600 164892 100200 6 mprj_dat_i[1]
port 371 nsew signal input
rlabel metal2 s 176988 99600 177044 100200 6 mprj_dat_i[20]
port 372 nsew signal input
rlabel metal2 s 177604 99600 177660 100200 6 mprj_dat_i[21]
port 373 nsew signal input
rlabel metal2 s 178276 99600 178332 100200 6 mprj_dat_i[22]
port 374 nsew signal input
rlabel metal2 s 178892 99600 178948 100200 6 mprj_dat_i[23]
port 375 nsew signal input
rlabel metal2 s 179564 99600 179620 100200 6 mprj_dat_i[24]
port 376 nsew signal input
rlabel metal2 s 180180 99600 180236 100200 6 mprj_dat_i[25]
port 377 nsew signal input
rlabel metal2 s 180796 99600 180852 100200 6 mprj_dat_i[26]
port 378 nsew signal input
rlabel metal2 s 181468 99600 181524 100200 6 mprj_dat_i[27]
port 379 nsew signal input
rlabel metal2 s 182084 99600 182140 100200 6 mprj_dat_i[28]
port 380 nsew signal input
rlabel metal2 s 182756 99600 182812 100200 6 mprj_dat_i[29]
port 381 nsew signal input
rlabel metal2 s 165452 99600 165508 100200 6 mprj_dat_i[2]
port 382 nsew signal input
rlabel metal2 s 183372 99600 183428 100200 6 mprj_dat_i[30]
port 383 nsew signal input
rlabel metal2 s 184044 99600 184100 100200 6 mprj_dat_i[31]
port 384 nsew signal input
rlabel metal2 s 166068 99600 166124 100200 6 mprj_dat_i[3]
port 385 nsew signal input
rlabel metal2 s 166740 99600 166796 100200 6 mprj_dat_i[4]
port 386 nsew signal input
rlabel metal2 s 167356 99600 167412 100200 6 mprj_dat_i[5]
port 387 nsew signal input
rlabel metal2 s 168028 99600 168084 100200 6 mprj_dat_i[6]
port 388 nsew signal input
rlabel metal2 s 168644 99600 168700 100200 6 mprj_dat_i[7]
port 389 nsew signal input
rlabel metal2 s 169316 99600 169372 100200 6 mprj_dat_i[8]
port 390 nsew signal input
rlabel metal2 s 169932 99600 169988 100200 6 mprj_dat_i[9]
port 391 nsew signal input
rlabel metal2 s 209636 99600 209692 100200 6 mprj_dat_o[0]
port 392 nsew signal output
rlabel metal2 s 216020 99600 216076 100200 6 mprj_dat_o[10]
port 393 nsew signal output
rlabel metal2 s 216692 99600 216748 100200 6 mprj_dat_o[11]
port 394 nsew signal output
rlabel metal2 s 217308 99600 217364 100200 6 mprj_dat_o[12]
port 395 nsew signal output
rlabel metal2 s 217980 99600 218036 100200 6 mprj_dat_o[13]
port 396 nsew signal output
rlabel metal2 s 218596 99600 218652 100200 6 mprj_dat_o[14]
port 397 nsew signal output
rlabel metal2 s 219268 99600 219324 100200 6 mprj_dat_o[15]
port 398 nsew signal output
rlabel metal2 s 219884 99600 219940 100200 6 mprj_dat_o[16]
port 399 nsew signal output
rlabel metal2 s 220500 99600 220556 100200 6 mprj_dat_o[17]
port 400 nsew signal output
rlabel metal2 s 221172 99600 221228 100200 6 mprj_dat_o[18]
port 401 nsew signal output
rlabel metal2 s 221788 99600 221844 100200 6 mprj_dat_o[19]
port 402 nsew signal output
rlabel metal2 s 210252 99600 210308 100200 6 mprj_dat_o[1]
port 403 nsew signal output
rlabel metal2 s 222460 99600 222516 100200 6 mprj_dat_o[20]
port 404 nsew signal output
rlabel metal2 s 223076 99600 223132 100200 6 mprj_dat_o[21]
port 405 nsew signal output
rlabel metal2 s 223748 99600 223804 100200 6 mprj_dat_o[22]
port 406 nsew signal output
rlabel metal2 s 224364 99600 224420 100200 6 mprj_dat_o[23]
port 407 nsew signal output
rlabel metal2 s 225036 99600 225092 100200 6 mprj_dat_o[24]
port 408 nsew signal output
rlabel metal2 s 225652 99600 225708 100200 6 mprj_dat_o[25]
port 409 nsew signal output
rlabel metal2 s 226268 99600 226324 100200 6 mprj_dat_o[26]
port 410 nsew signal output
rlabel metal2 s 226940 99600 226996 100200 6 mprj_dat_o[27]
port 411 nsew signal output
rlabel metal2 s 227556 99600 227612 100200 6 mprj_dat_o[28]
port 412 nsew signal output
rlabel metal2 s 228228 99600 228284 100200 6 mprj_dat_o[29]
port 413 nsew signal output
rlabel metal2 s 210924 99600 210980 100200 6 mprj_dat_o[2]
port 414 nsew signal output
rlabel metal2 s 228844 99600 228900 100200 6 mprj_dat_o[30]
port 415 nsew signal output
rlabel metal2 s 229516 99600 229572 100200 6 mprj_dat_o[31]
port 416 nsew signal output
rlabel metal2 s 211540 99600 211596 100200 6 mprj_dat_o[3]
port 417 nsew signal output
rlabel metal2 s 212212 99600 212268 100200 6 mprj_dat_o[4]
port 418 nsew signal output
rlabel metal2 s 212828 99600 212884 100200 6 mprj_dat_o[5]
port 419 nsew signal output
rlabel metal2 s 213500 99600 213556 100200 6 mprj_dat_o[6]
port 420 nsew signal output
rlabel metal2 s 214116 99600 214172 100200 6 mprj_dat_o[7]
port 421 nsew signal output
rlabel metal2 s 214788 99600 214844 100200 6 mprj_dat_o[8]
port 422 nsew signal output
rlabel metal2 s 215404 99600 215460 100200 6 mprj_dat_o[9]
port 423 nsew signal output
rlabel metal2 s 186564 99600 186620 100200 6 mprj_sel_o[0]
port 424 nsew signal output
rlabel metal2 s 187236 99600 187292 100200 6 mprj_sel_o[1]
port 425 nsew signal output
rlabel metal2 s 187852 99600 187908 100200 6 mprj_sel_o[2]
port 426 nsew signal output
rlabel metal2 s 188524 99600 188580 100200 6 mprj_sel_o[3]
port 427 nsew signal output
rlabel metal2 s 231420 99600 231476 100200 6 mprj_stb_o
port 428 nsew signal output
rlabel metal2 s 232708 99600 232764 100200 6 mprj_wb_iena
port 429 nsew signal output
rlabel metal2 s 230132 99600 230188 100200 6 mprj_we_o
port 430 nsew signal output
rlabel metal3 s 234600 25732 235200 25788 6 qspi_enabled
port 431 nsew signal output
rlabel metal3 s 234600 19852 235200 19908 6 ser_rx
port 432 nsew signal input
rlabel metal3 s 234600 21308 235200 21364 6 ser_tx
port 433 nsew signal output
rlabel metal3 s 234600 16884 235200 16940 6 spi_csb
port 434 nsew signal output
rlabel metal3 s 234600 22764 235200 22820 6 spi_enabled
port 435 nsew signal output
rlabel metal3 s 234600 15428 235200 15484 6 spi_sck
port 436 nsew signal output
rlabel metal3 s 234600 18396 235200 18452 6 spi_sdi
port 437 nsew signal input
rlabel metal3 s 234600 13972 235200 14028 6 spi_sdo
port 438 nsew signal output
rlabel metal3 s 234600 12516 235200 12572 6 spi_sdoenb
port 439 nsew signal output
rlabel metal3 s 234600 6636 235200 6692 6 trap
port 440 nsew signal output
rlabel metal3 s 234600 24276 235200 24332 6 uart_enabled
port 441 nsew signal output
rlabel metal2 s 184660 99600 184716 100200 6 user_irq_ena[0]
port 442 nsew signal output
rlabel metal2 s 185276 99600 185332 100200 6 user_irq_ena[1]
port 443 nsew signal output
rlabel metal2 s 185948 99600 186004 100200 6 user_irq_ena[2]
port 444 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 235000 100000
string LEFclass BLOCK
string LEFview TRUE
<< end >>
