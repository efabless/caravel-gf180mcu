magic
tech gf180mcuC
magscale 1 10
timestamp 1670447278
<< metal5 >>
tri 2594 5158 2684 5248 se
rect 2684 5158 3584 5428
tri 3584 5158 3674 5248 sw
tri 2504 4888 2594 4978 se
rect 2594 4888 3674 5158
tri 3674 4888 3764 4978 sw
tri 1064 4709 1243 4888 se
tri 1243 4798 1333 4888 sw
rect 1243 4709 1423 4798
rect 1064 4708 1423 4709
tri 1423 4708 1513 4798 sw
rect 2504 4708 3764 4888
tri 4935 4798 5025 4888 se
tri 4755 4708 4845 4798 se
rect 4845 4709 5025 4798
tri 5025 4709 5204 4888 sw
rect 4845 4708 5204 4709
tri 704 4348 1064 4708 se
rect 1064 4618 1603 4708
tri 1603 4618 1693 4708 sw
tri 2323 4618 2413 4708 se
rect 2413 4618 3855 4708
rect 1064 4438 1783 4618
tri 1783 4438 1963 4618 sw
tri 2233 4528 2323 4618 se
rect 2323 4528 3855 4618
tri 3855 4528 4035 4708 sw
tri 4575 4618 4665 4708 se
rect 4665 4618 5204 4708
tri 4395 4528 4485 4618 se
rect 4485 4528 5204 4618
tri 1963 4438 2053 4528 se
rect 2053 4438 4215 4528
tri 4215 4438 4305 4528 sw
tri 4305 4438 4395 4528 se
rect 4395 4438 5204 4528
rect 1064 4348 5204 4438
tri 5204 4348 5564 4708 sw
tri 704 4168 884 4348 ne
rect 884 4078 5384 4348
tri 5384 4168 5564 4348 nw
tri 884 3808 1154 4078 ne
tri 1064 3448 1154 3538 se
rect 1154 3448 5114 4078
tri 5114 3808 5384 4078 nw
tri 5114 3448 5204 3538 sw
rect 6680 3519 6980 3579
rect 7400 3519 7700 3579
rect 8060 3519 8480 3579
rect 8720 3519 9140 3579
rect 9920 3519 10340 3579
rect 10640 3519 10940 3579
rect 6620 3459 7040 3519
rect 7340 3459 7760 3519
rect 1064 3358 2864 3448
tri 2864 3358 2954 3448 nw
tri 3314 3358 3404 3448 ne
rect 3404 3358 5204 3448
tri 884 3088 1064 3268 se
rect 1064 3088 2324 3358
tri 434 2998 524 3088 se
rect 524 2998 2324 3088
rect 164 2188 2324 2998
tri 2324 2908 2774 3358 nw
tri 3494 2908 3944 3358 ne
rect 3944 3088 5204 3358
rect 6560 3339 7100 3459
tri 5204 3088 5384 3268 sw
rect 3944 2998 5744 3088
tri 5744 2998 5834 3088 sw
rect 3944 2188 6104 2998
rect 6560 2919 6740 3339
rect 6920 2919 7100 3339
rect 6560 2799 7100 2919
rect 7280 3339 7820 3459
rect 7280 2919 7460 3339
rect 7640 2919 7820 3339
rect 7280 2799 7820 2919
rect 8000 3399 8540 3519
rect 8000 3219 8180 3399
rect 8360 3219 8540 3399
rect 8000 3099 8540 3219
rect 8720 3459 9200 3519
rect 9860 3459 10340 3519
rect 10580 3459 11000 3519
rect 8720 3339 9260 3459
rect 8000 3039 8480 3099
rect 8000 2859 8180 3039
rect 6620 2739 7040 2799
rect 7280 2739 7760 2799
rect 8000 2739 8540 2859
rect 6680 2679 6980 2739
rect 7280 2679 7700 2739
rect 8060 2679 8540 2739
rect 8720 2679 8900 3339
rect 9080 2679 9260 3339
rect 9800 3399 10340 3459
rect 9800 3219 10040 3399
rect 10520 3339 11060 3459
rect 9800 3159 10220 3219
rect 9860 3099 10280 3159
rect 9920 3039 10340 3099
rect 10100 2859 10340 3039
rect 9800 2799 10340 2859
rect 10520 2919 10700 3339
rect 10880 2919 11060 3339
rect 10520 2799 11060 2919
rect 11240 2919 11420 3579
rect 11600 2919 11780 3579
rect 11240 2799 11780 2919
rect 11960 3519 12380 3579
rect 12800 3519 13100 3579
rect 13460 3519 13880 3579
rect 11960 3459 12440 3519
rect 12740 3459 13160 3519
rect 11960 3339 12500 3459
rect 9800 2739 10280 2799
rect 10580 2739 11000 2799
rect 11300 2739 11720 2799
rect 9800 2679 10220 2739
rect 10640 2679 10940 2739
rect 11360 2679 11660 2739
rect 11960 2679 12140 3339
rect 12320 3219 12500 3339
rect 12680 3339 13220 3459
rect 12680 2919 12860 3339
rect 13040 3219 13220 3339
rect 13400 3399 13940 3519
rect 13400 3219 13580 3399
rect 13760 3219 13940 3399
rect 13400 3099 13940 3219
rect 13400 3039 13880 3099
rect 13040 2919 13220 3039
rect 12680 2799 13220 2919
rect 13400 2859 13580 3039
rect 12740 2739 13160 2799
rect 13400 2739 13940 2859
rect 12800 2679 13100 2739
rect 13460 2679 13940 2739
rect 7280 2319 7460 2679
rect 9800 2319 9980 2679
rect 7280 2259 7700 2319
rect 8000 2259 8480 2319
rect 8720 2259 9140 2319
rect 9560 2259 9980 2319
rect 7280 2199 7760 2259
tri 434 2098 524 2188 ne
rect 524 2098 2324 2188
tri 794 1918 974 2098 ne
rect 974 1828 2324 2098
tri 2324 1828 2684 2188 sw
rect 974 1738 2684 1828
tri 974 1648 1064 1738 ne
rect 1064 1648 2684 1738
rect 1064 1558 2594 1648
tri 2594 1558 2684 1648 nw
tri 3584 1828 3944 2188 se
rect 3944 2098 5744 2188
tri 5744 2098 5834 2188 nw
rect 3944 1828 5294 2098
tri 5294 1918 5474 2098 nw
rect 7280 2079 7820 2199
rect 8000 2139 8540 2259
rect 3584 1738 5294 1828
rect 3584 1648 5204 1738
tri 5204 1648 5294 1738 nw
tri 3584 1558 3674 1648 ne
rect 3674 1558 5204 1648
tri 1064 1468 1154 1558 ne
tri 1064 1378 1154 1468 se
rect 1154 1378 2594 1558
tri 884 1108 1064 1288 se
rect 1064 1198 2504 1378
tri 2504 1288 2594 1378 nw
rect 3674 1378 5114 1558
tri 5114 1468 5204 1558 nw
tri 5114 1378 5204 1468 sw
rect 7280 1419 7460 2079
rect 7640 1419 7820 2079
rect 8360 1959 8540 2139
rect 8000 1779 8540 1959
rect 8000 1599 8180 1779
rect 8360 1599 8540 1779
rect 8000 1479 8540 1599
rect 8060 1419 8540 1479
rect 8720 2199 9200 2259
rect 9500 2199 9980 2259
rect 8720 2079 9260 2199
rect 8720 1419 8900 2079
rect 9080 1959 9260 2079
rect 9440 2079 9980 2199
rect 9440 1659 9620 2079
rect 9800 1659 9980 2079
rect 9440 1539 9980 1659
rect 10160 1659 10340 2319
rect 10520 1659 10700 2319
rect 10880 1659 11060 2319
rect 11240 2259 11720 2319
rect 11960 2259 12380 2319
rect 12740 2259 13160 2319
rect 11240 2139 11780 2259
rect 11600 1959 11780 2139
rect 11300 1899 11780 1959
rect 10160 1539 11060 1659
rect 11240 1779 11780 1899
rect 11240 1599 11420 1779
rect 11600 1599 11780 1779
rect 9500 1479 9980 1539
rect 10220 1479 11000 1539
rect 11240 1479 11780 1599
rect 9560 1419 9980 1479
rect 10280 1419 10520 1479
rect 10700 1419 10940 1479
rect 11300 1419 11780 1479
rect 11960 2199 12440 2259
rect 11960 2079 12500 2199
rect 11960 1419 12140 2079
rect 12320 1959 12500 2079
rect 12680 2139 13220 2259
rect 12680 1959 12860 2139
rect 13040 1959 13220 2139
rect 12680 1779 13220 1959
rect 12680 1599 12860 1779
rect 12680 1479 13220 1599
rect 12740 1419 13220 1479
tri 3674 1288 3764 1378 ne
rect 1064 1108 2414 1198
tri 2414 1108 2504 1198 nw
rect 3764 1198 5204 1378
tri 3764 1108 3854 1198 ne
rect 3854 1108 5204 1198
tri 5204 1108 5384 1288 sw
tri 704 838 884 1018 se
rect 884 928 2414 1108
rect 884 838 2324 928
tri 2324 838 2414 928 nw
rect 3854 928 5384 1108
tri 3854 838 3944 928 ne
rect 3944 838 5384 928
tri 5384 838 5564 1018 sw
tri 704 298 1244 838 ne
rect 1244 748 2324 838
rect 1244 658 2258 748
tri 2258 682 2324 748 nw
rect 3944 748 5024 838
tri 3944 682 4010 748 ne
rect 1244 568 1784 658
tri 1784 568 1874 658 nw
tri 1939 568 2029 658 ne
rect 2029 592 2258 658
rect 2029 568 2144 592
rect 1244 478 1604 568
tri 1604 478 1694 568 nw
tri 2029 478 2119 568 ne
rect 2119 478 2144 568
tri 2144 478 2258 592 nw
rect 4010 658 5024 748
rect 4010 592 4149 658
tri 4010 478 4124 592 ne
rect 4124 478 4149 592
tri 4149 478 4329 658 nw
tri 4394 568 4484 658 ne
rect 4484 568 5024 658
tri 4574 478 4664 568 ne
rect 4664 478 5024 568
rect 1244 298 1334 478
tri 1334 298 1514 478 nw
tri 4754 298 4934 478 ne
rect 4934 298 5024 478
tri 5024 298 5564 838 nw
<< fillblock >>
rect 0 0 6227 5539
rect 6420 1242 14139 3770
<< end >>
