magic
tech gf180mcuC
magscale 1 5
timestamp 1654634570
<< metal5 >>
rect 0 432 108 756
rect 216 432 324 756
rect 0 324 324 432
rect 0 0 108 324
rect 216 0 324 324
<< properties >>
string FIXED_BBOX 0 -216 432 756
<< end >>
