magic
tech gf180mcuC
magscale 1 5
timestamp 1654634570
<< metal5 >>
rect 144 720 648 756
rect 108 684 684 720
rect 72 648 720 684
rect 36 612 216 648
rect 576 612 756 648
rect 0 576 180 612
rect 612 576 756 612
rect 0 540 144 576
rect 0 0 108 540
rect 288 504 468 540
rect 252 468 504 504
rect 216 396 540 468
rect 216 144 324 396
rect 432 144 540 396
rect 648 144 756 576
rect 216 72 756 144
rect 252 36 720 72
rect 288 0 432 36
rect 540 0 684 36
rect 0 -36 144 0
rect 0 -72 180 -36
rect 36 -108 216 -72
rect 72 -144 648 -108
rect 108 -180 648 -144
rect 144 -216 648 -180
<< properties >>
string FIXED_BBOX 0 -216 864 756
<< end >>
