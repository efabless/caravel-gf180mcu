* NGSPICE file created from housekeeping.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1 D RN CLKN Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 D RN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 D RN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyd_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyd_4 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 D SETN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_4 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_4 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_4 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_4 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_16 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_4 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffsnq_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffsnq_4 D SETN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_20 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_20 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_2 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_20 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_20 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_4 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrnq_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_4 D RN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_4 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffnsnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffnsnq_1 D SETN CLKN Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_12 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_12 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_16 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyd_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyd_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_2 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_4 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_16 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_2 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_2 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffsnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffsnq_2 D SETN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_20 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_20 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tieh abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tieh Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_4 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_4 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_12 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_12 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_4 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_2 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_4 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_2 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyc_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyc_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_4 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_2 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_4 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_8 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_8 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_4 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_3 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_12 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_12 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 I ZN VDD VSS
.ends

.subckt housekeeping VDD VSS debug_in debug_mode debug_oeb debug_out irq[0] irq[1]
+ irq[2] mask_rev_in[0] mask_rev_in[10] mask_rev_in[11] mask_rev_in[12] mask_rev_in[13]
+ mask_rev_in[14] mask_rev_in[15] mask_rev_in[16] mask_rev_in[17] mask_rev_in[18]
+ mask_rev_in[19] mask_rev_in[1] mask_rev_in[20] mask_rev_in[21] mask_rev_in[22] mask_rev_in[23]
+ mask_rev_in[24] mask_rev_in[25] mask_rev_in[26] mask_rev_in[27] mask_rev_in[28]
+ mask_rev_in[29] mask_rev_in[2] mask_rev_in[30] mask_rev_in[31] mask_rev_in[3] mask_rev_in[4]
+ mask_rev_in[5] mask_rev_in[6] mask_rev_in[7] mask_rev_in[8] mask_rev_in[9] mgmt_gpio_in[0]
+ mgmt_gpio_in[10] mgmt_gpio_in[11] mgmt_gpio_in[12] mgmt_gpio_in[13] mgmt_gpio_in[14]
+ mgmt_gpio_in[15] mgmt_gpio_in[16] mgmt_gpio_in[17] mgmt_gpio_in[18] mgmt_gpio_in[19]
+ mgmt_gpio_in[1] mgmt_gpio_in[20] mgmt_gpio_in[21] mgmt_gpio_in[22] mgmt_gpio_in[23]
+ mgmt_gpio_in[24] mgmt_gpio_in[25] mgmt_gpio_in[26] mgmt_gpio_in[27] mgmt_gpio_in[28]
+ mgmt_gpio_in[29] mgmt_gpio_in[2] mgmt_gpio_in[30] mgmt_gpio_in[31] mgmt_gpio_in[32]
+ mgmt_gpio_in[33] mgmt_gpio_in[34] mgmt_gpio_in[35] mgmt_gpio_in[36] mgmt_gpio_in[37]
+ mgmt_gpio_in[3] mgmt_gpio_in[4] mgmt_gpio_in[5] mgmt_gpio_in[6] mgmt_gpio_in[7]
+ mgmt_gpio_in[8] mgmt_gpio_in[9] mgmt_gpio_oeb[0] mgmt_gpio_oeb[10] mgmt_gpio_oeb[11]
+ mgmt_gpio_oeb[12] mgmt_gpio_oeb[13] mgmt_gpio_oeb[14] mgmt_gpio_oeb[15] mgmt_gpio_oeb[16]
+ mgmt_gpio_oeb[17] mgmt_gpio_oeb[18] mgmt_gpio_oeb[19] mgmt_gpio_oeb[1] mgmt_gpio_oeb[20]
+ mgmt_gpio_oeb[21] mgmt_gpio_oeb[22] mgmt_gpio_oeb[23] mgmt_gpio_oeb[24] mgmt_gpio_oeb[25]
+ mgmt_gpio_oeb[26] mgmt_gpio_oeb[27] mgmt_gpio_oeb[28] mgmt_gpio_oeb[29] mgmt_gpio_oeb[2]
+ mgmt_gpio_oeb[30] mgmt_gpio_oeb[31] mgmt_gpio_oeb[32] mgmt_gpio_oeb[33] mgmt_gpio_oeb[34]
+ mgmt_gpio_oeb[35] mgmt_gpio_oeb[36] mgmt_gpio_oeb[37] mgmt_gpio_oeb[3] mgmt_gpio_oeb[4]
+ mgmt_gpio_oeb[5] mgmt_gpio_oeb[6] mgmt_gpio_oeb[7] mgmt_gpio_oeb[8] mgmt_gpio_oeb[9]
+ mgmt_gpio_out[0] mgmt_gpio_out[10] mgmt_gpio_out[11] mgmt_gpio_out[12] mgmt_gpio_out[13]
+ mgmt_gpio_out[14] mgmt_gpio_out[15] mgmt_gpio_out[16] mgmt_gpio_out[17] mgmt_gpio_out[18]
+ mgmt_gpio_out[19] mgmt_gpio_out[1] mgmt_gpio_out[20] mgmt_gpio_out[21] mgmt_gpio_out[22]
+ mgmt_gpio_out[23] mgmt_gpio_out[24] mgmt_gpio_out[25] mgmt_gpio_out[26] mgmt_gpio_out[27]
+ mgmt_gpio_out[28] mgmt_gpio_out[29] mgmt_gpio_out[2] mgmt_gpio_out[30] mgmt_gpio_out[31]
+ mgmt_gpio_out[32] mgmt_gpio_out[33] mgmt_gpio_out[34] mgmt_gpio_out[35] mgmt_gpio_out[36]
+ mgmt_gpio_out[37] mgmt_gpio_out[3] mgmt_gpio_out[4] mgmt_gpio_out[5] mgmt_gpio_out[6]
+ mgmt_gpio_out[7] mgmt_gpio_out[8] mgmt_gpio_out[9] pad_flash_clk pad_flash_clk_oe
+ pad_flash_csb pad_flash_csb_oe pad_flash_io0_di pad_flash_io0_do pad_flash_io0_ie
+ pad_flash_io0_oe pad_flash_io1_di pad_flash_io1_do pad_flash_io1_ie pad_flash_io1_oe
+ pll90_sel[0] pll90_sel[1] pll90_sel[2] pll_bypass pll_dco_ena pll_div[0] pll_div[1]
+ pll_div[2] pll_div[3] pll_div[4] pll_ena pll_sel[0] pll_sel[1] pll_sel[2] pll_trim[0]
+ pll_trim[10] pll_trim[11] pll_trim[12] pll_trim[13] pll_trim[14] pll_trim[15] pll_trim[16]
+ pll_trim[17] pll_trim[18] pll_trim[19] pll_trim[1] pll_trim[20] pll_trim[21] pll_trim[22]
+ pll_trim[23] pll_trim[24] pll_trim[25] pll_trim[2] pll_trim[3] pll_trim[4] pll_trim[5]
+ pll_trim[6] pll_trim[7] pll_trim[8] pll_trim[9] porb pwr_ctrl_out qspi_enabled reset
+ ser_rx ser_tx serial_clock serial_data_1 serial_data_2 serial_load serial_resetn
+ spi_csb spi_enabled spi_sck spi_sdi spi_sdo spi_sdoenb spimemio_flash_clk spimemio_flash_csb
+ spimemio_flash_io0_di spimemio_flash_io0_do spimemio_flash_io0_oeb spimemio_flash_io1_di
+ spimemio_flash_io1_do spimemio_flash_io1_oeb spimemio_flash_io2_di spimemio_flash_io2_do
+ spimemio_flash_io2_oeb spimemio_flash_io3_di spimemio_flash_io3_do spimemio_flash_io3_oeb
+ trap uart_enabled user_clock wb_ack_o wb_adr_i[0] wb_adr_i[10] wb_adr_i[11] wb_adr_i[12]
+ wb_adr_i[13] wb_adr_i[14] wb_adr_i[15] wb_adr_i[16] wb_adr_i[17] wb_adr_i[18] wb_adr_i[19]
+ wb_adr_i[1] wb_adr_i[20] wb_adr_i[21] wb_adr_i[22] wb_adr_i[23] wb_adr_i[24] wb_adr_i[25]
+ wb_adr_i[26] wb_adr_i[27] wb_adr_i[28] wb_adr_i[29] wb_adr_i[2] wb_adr_i[30] wb_adr_i[31]
+ wb_adr_i[3] wb_adr_i[4] wb_adr_i[5] wb_adr_i[6] wb_adr_i[7] wb_adr_i[8] wb_adr_i[9]
+ wb_clk_i wb_cyc_i wb_dat_i[0] wb_dat_i[10] wb_dat_i[11] wb_dat_i[12] wb_dat_i[13]
+ wb_dat_i[14] wb_dat_i[15] wb_dat_i[16] wb_dat_i[17] wb_dat_i[18] wb_dat_i[19] wb_dat_i[1]
+ wb_dat_i[20] wb_dat_i[21] wb_dat_i[22] wb_dat_i[23] wb_dat_i[24] wb_dat_i[25] wb_dat_i[26]
+ wb_dat_i[27] wb_dat_i[28] wb_dat_i[29] wb_dat_i[2] wb_dat_i[30] wb_dat_i[31] wb_dat_i[3]
+ wb_dat_i[4] wb_dat_i[5] wb_dat_i[6] wb_dat_i[7] wb_dat_i[8] wb_dat_i[9] wb_dat_o[0]
+ wb_dat_o[10] wb_dat_o[11] wb_dat_o[12] wb_dat_o[13] wb_dat_o[14] wb_dat_o[15] wb_dat_o[16]
+ wb_dat_o[17] wb_dat_o[18] wb_dat_o[19] wb_dat_o[1] wb_dat_o[20] wb_dat_o[21] wb_dat_o[22]
+ wb_dat_o[23] wb_dat_o[24] wb_dat_o[25] wb_dat_o[26] wb_dat_o[27] wb_dat_o[28] wb_dat_o[29]
+ wb_dat_o[2] wb_dat_o[30] wb_dat_o[31] wb_dat_o[3] wb_dat_o[4] wb_dat_o[5] wb_dat_o[6]
+ wb_dat_o[7] wb_dat_o[8] wb_dat_o[9] wb_rstn_i wb_sel_i[0] wb_sel_i[1] wb_sel_i[2]
+ wb_sel_i[3] wb_stb_i wb_we_i
XFILLER_100_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6914_ _6914_/D _6672_/Z _4111_/I1 _6914_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_54_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6845_ _6845_/D _6862_/CLK _6845_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_168_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3988_ _3991_/A2 _6707_/Q _6708_/Q _3989_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6776_ _6776_/D _6667_/Z _4111_/I1 _6776_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_5727_ _5784_/A2 _5535_/B _5727_/A3 _5802_/A2 _5735_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_182_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5658_ hold25/Z hold527/Z _5663_/S _7042_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4609_ _4443_/Z _5459_/A3 _5404_/B2 _5225_/A2 _4609_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_163_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5589_ hold58/Z hold355/Z _5590_/S _5589_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7328_ _7328_/D _6682_/Z _4089_/I1 _7328_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_117_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold351 _5769_/Z _7140_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold340 _7119_/Q hold340/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold362 _7046_/Q hold362/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold395 _5560_/Z _6956_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold373 _5624_/Z _7013_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7259_ _7259_/D _7341_/RN _7259_/CLK _7259_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_89_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold384 _4167_/Z _6732_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2512 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_165_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1833 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1855 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1844 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1888 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1877 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_876 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4960_ _4958_/B _4777_/C _4960_/B _4960_/C _5104_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_64_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3911_ _6887_/Q _5655_/A4 _4405_/A3 _5546_/A2 _3954_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_4891_ _4891_/A1 _5263_/A3 _4891_/A3 _5469_/A4 _4893_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6630_ _6630_/I0 _7318_/Q _6642_/S _7318_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_177_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3842_ _7065_/Q _3980_/A2 _3842_/B _3845_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_177_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6561_ _6902_/Q _6563_/A3 _6561_/A3 _6563_/A4 _6565_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_164_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3773_ _3773_/A1 _3773_/A2 _3773_/A3 _3773_/A4 _3790_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5512_ _5856_/A1 _5745_/A4 _5552_/A2 _5838_/A4 _5517_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_146_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6492_ hold60/I _6285_/Z _6294_/Z _7038_/Q _6564_/C1 _7086_/Q _6499_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_9_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5443_ _5481_/A1 _5443_/A2 _5504_/A2 _5487_/A2 _5448_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_5374_ _5376_/A1 _5374_/A2 _5498_/A2 _5454_/A2 _5374_/C _5412_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_4325_ _6600_/I0 _6840_/Q _4328_/S _6840_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7113_ _7113_/D _7302_/RN _7113_/CLK _7113_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_87_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4256_ hold313/Z hold164/Z _4262_/S _4256_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xnet483_109 net483_129/I _7160_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7044_ _7044_/D _7302_/RN _7044_/CLK _7044_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4187_ hold5/Z hold235/Z _4189_/S _4187_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_27_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6828_ _6828_/D _7302_/RN _6828_/CLK _6828_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_50_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6759_ _6759_/D _7341_/RN _6759_/CLK _6759_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_152_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold170 _6704_/Q hold170/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_105_731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold192 _7256_/Q hold192/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold181 _7108_/Q hold181/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_59_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2364 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1674 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1652 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_612 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_678 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5090_ _5315_/A4 _5476_/A2 _5301_/A2 _3379_/I _5382_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_96_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4110_ input84/Z input67/Z _7344_/Q _4110_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_111_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4041_ _6532_/C _4041_/A2 _6788_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_110_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5992_ _6211_/B _7274_/Q _6232_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_37_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4943_ _5370_/A1 _5454_/A1 _5003_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6613_ _6613_/A1 _6613_/A2 _6614_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4874_ _4874_/A1 _4874_/A2 _4874_/A3 _5256_/A3 _4877_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_177_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3825_ _6711_/Q _5784_/A3 _5532_/A3 _6653_/A2 _3843_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_177_299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6544_ _7340_/Q _6279_/Z _6299_/Z _6889_/Q _6575_/B1 _6885_/Q _6548_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_3756_ _7026_/Q _5727_/A3 _4378_/A1 _5856_/A2 _3788_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_180_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6475_ _7093_/Q _6578_/A2 _6310_/Z _6981_/Q _6578_/C1 _7175_/Q _6480_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_118_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5426_ _5426_/A1 _5466_/A2 _5327_/B _5426_/B1 _5426_/B2 _5427_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_3687_ _3687_/A1 _3687_/A2 _3687_/A3 _3687_/A4 _3715_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_134_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput242 _7353_/Z mgmt_gpio_out[5] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput253 _4115_/I pad_flash_io0_oe VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput220 _4096_/ZN mgmt_gpio_out[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput231 _7350_/Z mgmt_gpio_out[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5357_ _5357_/A1 _5495_/A1 _5359_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_142_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput286 _6717_/Q pll_trim[23] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput264 _6924_/Q pll_div[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput275 _6723_/Q pll_trim[13] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5288_ _5369_/A2 _4947_/C _5290_/B _5288_/A4 _5381_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_102_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4308_ _5528_/A2 _5535_/B _5573_/A3 _5856_/A2 _4310_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_839 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput297 _6936_/Q pwr_ctrl_out VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_114_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7027_ _7027_/D _7302_/RN _7027_/CLK _7027_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_75_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4239_ hold424/Z hold5/Z _4243_/S _4239_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_71_802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_898 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_879 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4590_ _4759_/C _4686_/B _5307_/B _4694_/B _5503_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_147_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3610_ _6998_/Q _3953_/A2 _3939_/B1 input32/Z _3612_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_174_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3541_ _5534_/A1 _3827_/A2 _3496_/B _5534_/A2 _3938_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_6_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3472_ _6863_/Q hold7/Z _3472_/B _3507_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_131_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6260_ _6892_/Q _6260_/A2 _6260_/B1 _6834_/Q _6263_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5211_ _5347_/A1 _5211_/A2 _5211_/B _5212_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xnet533_190 net433_54/I _7079_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_170_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6191_ _6788_/Q _6191_/A2 _6192_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_43_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5142_ _5330_/A2 _5252_/A4 _5152_/B _5330_/B1 _5397_/A1 _5335_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_69_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5073_ _5073_/A1 _5073_/A2 _5073_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_84_426 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4024_ hold284/Z _4026_/C _5564_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_65_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_898 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5975_ _7280_/Q _6311_/A1 _5975_/B _5979_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_80_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4926_ _4951_/A1 _4951_/A2 _4926_/B _4926_/C _5091_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_33_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4857_ _5439_/C _4857_/A2 _4857_/B _4857_/C _5438_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_20_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3808_ _6832_/Q _5784_/A3 _5546_/A2 _5573_/A3 _3855_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_118_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4788_ _4667_/Z _5244_/A2 _4693_/Z _5255_/B _5426_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6527_ _7095_/Q _6578_/A2 _6310_/Z _6983_/Q _6578_/C1 _7177_/Q _6529_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_3739_ _6940_/Q _5544_/S _3681_/Z _6925_/Q _3740_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6458_ _7101_/Q _6563_/A3 _6561_/A3 _6563_/A4 _6471_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_69_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5409_ _4947_/C _5409_/A2 _5409_/B _5409_/C _5415_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_133_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6389_ _7204_/Q _6573_/A2 _6288_/Z _7196_/Q _6297_/Z _7042_/Q _6390_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_0_614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_25__1374_ clkbuf_4_12_0__1374_/Z net433_77/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_105__1374_ clkbuf_4_1_0__1374_/Z net833_480/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_87_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_88__1374_ clkbuf_4_4_0__1374_/Z net483_129/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_47_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_868 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet783_411 net783_411/I _6807_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet783_433 net783_433/I _6781_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet783_444 net783_445/I _6765_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_70_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet783_422 net783_425/I _6796_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_184_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_184_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5760_ hold25/Z hold497/Z _5765_/S _7132_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_15_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5691_ _4227_/B _5718_/A3 _5902_/A3 _5866_/A3 _5699_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_4711_ _4822_/A4 _5250_/C _5241_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4642_ _4642_/A1 _5230_/C _5081_/C _4650_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_175_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4573_ _5466_/B _3380_/I _3379_/I _5034_/A2 _5079_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_7361_ _7361_/I _7361_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold703 _6736_/Q hold703/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_162_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3524_ _3644_/A2 _5534_/A2 _3460_/B _3534_/C _4243_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xhold725 _6946_/Q hold725/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6312_ _7281_/Q _6563_/A3 _6563_/A4 _6312_/A4 _6312_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_7_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold736 _4221_/Z _6770_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7292_ _7292_/D _7302_/RN _7302_/CLK _7292_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold714 _4198_/Z _6755_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_170_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3455_ _6863_/Q hold20/Z _3455_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xhold747 _5507_/Z _6910_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_115_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold758 _4162_/Z _6727_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6243_ _6107_/B _6107_/C _6829_/Q _7275_/Q _6244_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
Xhold769 _6766_/Q hold769/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_170_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3386_ _5307_/B _5312_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_16
XFILLER_130_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6174_ _6990_/Q _6260_/B1 _6258_/C1 hold82/I _6176_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_97_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5125_ _5128_/A1 _5476_/A1 _5148_/B1 _5484_/A4 _5125_/C _5130_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_97_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5056_ _5347_/A1 _5330_/B2 _5435_/A1 _4568_/Z _5056_/B2 _5420_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_4007_ _3475_/Z _4006_/B _4007_/B _4009_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_38_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_879 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5958_ _7277_/Q _7276_/Q _6321_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_4909_ _5290_/C _3380_/I _3379_/I _5034_/A2 _5087_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_179_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_214 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5889_ hold164/Z hold371/Z _5892_/S _7246_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_138_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet733_363 net433_67/I _6891_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet733_374 net733_381/I _6869_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet733_352 _4109__3/I _6902_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet733_396 net783_426/I _6822_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet733_385 net783_445/I _6833_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_1_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold30 hold30/I hold30/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_152_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold41 hold41/I hold41/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_121_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold74 hold74/I hold74/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold52 hold52/I hold52/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold63 hold63/I hold63/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold85 hold85/I hold85/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_17_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold96 hold96/I hold96/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_16_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_7__f_wb_clk_i clkbuf_0_wb_clk_i/Z _4103_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_90_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6930_ _6930_/D _7262_/RN _6930_/CLK _6930_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6861_ _6861_/D _6862_/CLK _6861_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5812_ hold391/Z hold849/Z _5819_/S _5812_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6792_ _6792_/D _7281_/RN _6792_/CLK _6792_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_90_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5743_ hold62/Z hold58/Z _5744_/S hold63/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5674_ hold391/Z hold859/Z _5681_/S _7056_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4625_ _5082_/C _5435_/A1 _4454_/B _5187_/B _5077_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_135_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4556_ _4443_/Z _5459_/A3 _5439_/A1 _5389_/A2 _5213_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_163_537 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold511 _5825_/Z _7190_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold500 _6986_/Q hold500/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7344_ _7344_/D _6696_/Z _4111_/I1 _7344_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3507_ _6863_/Q _5326_/B2 hold12/Z _3511_/B2 _3507_/C hold13/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
Xhold522 _6899_/Q hold522/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold533 _7156_/Q hold533/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold544 _4298_/Z _6820_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4487_ _3379_/I _3380_/I _4487_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_4
Xhold555 _7235_/Q hold555/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold588 _4292_/Z _6814_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_171_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold577 _6882_/Q hold577/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7275_ _7275_/D _7302_/RN _7304_/CLK _7275_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_1_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold566 _7340_/Q hold566/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3438_ hold138/Z hold24/Z _3440_/S _7330_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6226_ _6864_/Q _6257_/A2 _6258_/C1 _6889_/Q _6893_/Q _6256_/B1 _6229_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_89_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold599 _4263_/Z _6798_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6157_ _7021_/Q _6259_/A2 _6261_/A2 _7005_/Q _6161_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3369_ _7019_/Q _3369_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_66_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_871 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5108_ _5373_/A1 _5108_/A2 _5110_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6088_ _6088_/I0 _7287_/Q _6559_/S _7287_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5039_ _5039_/A1 _5235_/A1 _5253_/A1 _5091_/B _5041_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_66_790 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2749 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput120 wb_adr_i[3] _4718_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
Xinput131 wb_dat_i[12] _6627_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput153 wb_dat_i[3] _6624_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput142 wb_dat_i[22] _6636_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_88_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput164 wb_sel_i[3] _6648_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_49_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_865 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_82_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_842 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4410_ _4840_/A1 _4777_/A2 _4960_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_5390_ _5390_/A1 _5404_/A2 _5390_/B _5390_/C _5391_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_99_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4341_ _4343_/S _6851_/Q _4342_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7060_ _7060_/D _7265_/RN _7060_/CLK _7060_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4272_ _4271_/Z hold556/Z _4282_/S _4272_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_125_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6011_ _6036_/A3 _6103_/A1 _6211_/B _7274_/Q _6262_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_39_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_749 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_790 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6913_ _6913_/D _6671_/Z _7346_/CLK _6913_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_54_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6844_ _6844_/D _7262_/RN _6844_/CLK _6844_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_22_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3987_ _3991_/A2 _6707_/Q _3990_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6775_ _6775_/D _6666_/Z _7346_/CLK _6775_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_50_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5726_ hold2/Z _7103_/Q hold22/Z hold23/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_10_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_868 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5657_ hold388/Z hold842/Z _5663_/S _7041_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4608_ _5459_/A3 _5225_/A2 _5225_/A1 _5225_/A3 _4608_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_5588_ hold5/Z hold396/Z _5590_/S _5588_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4539_ _5262_/A4 _5315_/A4 _5301_/A2 _4661_/C _5372_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_144_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold352 _7029_/Q hold352/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold330 _5644_/Z _7030_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7327_ _7327_/D _6681_/Z _7346_/CLK _7327_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold341 _7137_/Q hold341/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7258_ _7258_/D _7341_/RN _7258_/CLK _7258_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
Xhold363 _7051_/Q hold363/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_132_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold374 _7133_/Q hold374/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold396 _6981_/Q hold396/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold385 _7207_/Q hold385/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6209_ hold32/I _6262_/A2 _6262_/B1 _7153_/Q _6210_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_89_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7189_ _7189_/D _7341_/RN _7189_/CLK _7189_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_131_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_640 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_896 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2535 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2568 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1823 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1801 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1867 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1856 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1845 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1878 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_835 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_823 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3910_ _6833_/Q _5745_/A4 _4378_/A1 _4405_/A2 _3937_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4890_ _4423_/Z _5177_/A3 _5153_/B _5321_/A3 _4891_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_51_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3841_ input21/Z _3977_/A2 _3939_/A2 _6985_/Q _3841_/C _3886_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_20_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6560_ _6911_/Q _6563_/A2 _6562_/A3 _6563_/A4 _6572_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3772_ _6712_/Q _3942_/A2 _3975_/A2 _7220_/Q _3773_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_158_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5511_ hold388/Z hold678/Z _5511_/S _5511_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_185_470 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6491_ _6491_/A1 _6491_/A2 _6491_/A3 _6491_/A4 _6491_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_5442_ _5442_/I _5487_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_172_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_827 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5373_ _5373_/A1 _5373_/A2 _5373_/A3 _5373_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_99_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4324_ _6599_/A1 _4328_/S _4324_/B _6839_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7112_ _7112_/D _7302_/RN _7112_/CLK _7112_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_86_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7043_ _7043_/D _7302_/RN _7043_/CLK _7043_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_113_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4255_ hold621/Z _4254_/Z _4263_/S _4255_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_86_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_863 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4186_ hold164/Z hold183/Z _4189_/S _4186_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_94_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6827_ _6827_/D _7304_/RN _6827_/CLK _6827_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_11_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6758_ _6758_/D _7262_/RN _6758_/CLK _6758_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_164_610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5709_ _4227_/B _5718_/A3 hold13/Z _5866_/A3 _5717_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_6689_ input75/Z _6994_/Q _4026_/C _6689_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_164_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_827 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold171 hold171/I hold171/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold160 _6962_/Q hold160/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold193 _7038_/Q hold193/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_105_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold182 _5732_/Z _7108_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_120_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1642 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1675 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_796 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_654 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4040_ _4019_/Z _5930_/A1 _5930_/A2 _6789_/Q _4041_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_94_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_652 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5991_ _5917_/B _6587_/A2 _7285_/Q _6033_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4942_ _4963_/B _4995_/A4 _5025_/A3 _4922_/B _4942_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_80_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_793 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6612_ _6878_/Q _6612_/A2 _6612_/B1 _6640_/B2 _6613_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4873_ _4423_/Z _5177_/A3 _5153_/B _5180_/B _4874_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_20_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3824_ _3496_/B _4246_/A1 _4227_/A2 _3477_/Z _3942_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xnet583_250 net583_250/I _7019_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6543_ _6540_/Z _6543_/A2 _6543_/A3 _6543_/A4 _6555_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3755_ _6929_/Q _5745_/A4 _5518_/A1 _5552_/A2 _3784_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6474_ _6468_/Z _6474_/A2 _6474_/A3 _6474_/A4 _6481_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3686_ _6988_/Q _3939_/A2 _3939_/B1 input30/Z _3687_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_160_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5425_ _5457_/A2 _5425_/A2 _5458_/A2 _5450_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_146_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput210 _4088_/Z mgmt_gpio_out[10] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_106_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput232 _7371_/Z mgmt_gpio_out[30] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput221 _7361_/Z mgmt_gpio_out[20] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput243 _4091_/Z mgmt_gpio_out[6] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5356_ _5356_/A1 _5356_/A2 _5356_/A3 _5495_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_114_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput254 _7374_/Z pad_flash_io1_do VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput276 _6724_/Q pll_trim[14] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput265 _6925_/Q pll_div[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5287_ _5318_/A2 _5290_/B _5287_/B1 _5426_/B1 _5287_/C _5386_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_101_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4307_ hold2/Z hold197/Z _4307_/S _4307_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xoutput298 _3892_/Z reset VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput287 _6933_/Q pll_trim[24] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_102_757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4238_ hold674/Z _4237_/Z _4244_/S _4238_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7026_ _7026_/D _7281_/RN _7026_/CLK _7026_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_75_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4169_ _4405_/A3 _5535_/B _6653_/A2 _6653_/A3 _4171_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_70_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_48__1374_ clkbuf_4_15_0__1374_/Z net633_277/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_139_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_183_248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_711 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3540_ _3833_/A2 _3477_/Z _3496_/B _5534_/A2 _3945_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_143_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5210_ _5404_/B2 _5372_/A1 _5210_/B _5210_/C _5211_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3471_ _3472_/B _3470_/Z _3511_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_4
Xnet533_191 _4109__28/I _7078_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_130_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6190_ _6107_/B _6107_/C _6974_/Q _7275_/Q _6191_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
Xnet533_180 net583_233/I _7089_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5141_ _5141_/A1 _5141_/A2 _5490_/A1 _5141_/A4 _5144_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_36_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5072_ _4443_/Z _5459_/A3 _5225_/A2 _5285_/A1 _5073_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4023_ _4107_/A1 hold725/Z input67/Z _4246_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_38_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5974_ _6789_/Q _5973_/Z _5974_/B1 _6312_/A4 _7280_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4925_ _4951_/B1 _4995_/A4 _4951_/B2 _5288_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_100_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4856_ _4690_/C _5466_/B _5392_/A1 _5170_/B1 _4857_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_33_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3807_ _6869_/Q _4378_/A1 _5838_/A2 _5546_/A2 _3870_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_4787_ _5250_/B _4787_/A2 _4787_/A3 _4922_/B _5260_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_6526_ _7257_/Q _6580_/B1 _6309_/Z _7241_/Q _6749_/Q _6579_/A2 _6529_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_174_782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3738_ _7125_/Q _3956_/A2 _3956_/B1 _7157_/Q _6971_/Q _3559_/Z _3740_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_134_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6457_ _7231_/Q _6563_/A2 _6457_/A3 _6563_/A4 _6469_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_3669_ _3669_/A1 _3669_/A2 _3669_/A3 _3669_/A4 _3669_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_69_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5408_ _5408_/A1 _5408_/A2 _5408_/A3 _5408_/A4 _6906_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6388_ _7106_/Q _6285_/Z _6294_/Z _7034_/Q _6564_/C1 _7082_/Q _6390_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_88_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5339_ _5473_/A1 _5492_/A4 _5336_/Z _5338_/Z _5339_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_130_863 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7009_ _7009_/D _7302_/RN _7009_/CLK _7009_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_28_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_3_6__f_wb_clk_i clkbuf_0_wb_clk_i/Z _7281_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_44_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet783_434 net783_435/I _6780_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet783_412 net783_415/I _6806_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_140_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet783_423 net783_424/I _6795_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_156_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet783_445 net783_445/I _6764_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_156_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_4_15_0__1374_ clkbuf_3_7_0__1374_/Z clkbuf_4_15_0__1374_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_38_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5690_ hold2/Z _7071_/Q hold42/Z hold43/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4710_ _4787_/A3 _4787_/A2 _4710_/B _4710_/C _5250_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_91_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4641_ _4443_/Z _4454_/B _5050_/A2 _4960_/C _5081_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_147_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7360_ _7360_/I _7360_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_31__1374_ clkbuf_4_11_0__1374_/Z net433_58/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_116_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4572_ _4469_/B _4686_/B _5312_/B _4922_/B _5170_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_7_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_111__1374_ net733_398/I net783_408/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_155_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold726 _5547_/Z _6946_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold737 _6911_/Q hold737/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6311_ _6311_/A1 _6562_/A4 _6311_/B _6311_/C _6318_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
Xhold715 _6734_/Q hold715/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xclkbuf_leaf_94__1374_ clkbuf_4_3_0__1374_/Z _4109__3/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xhold704 _6741_/Q hold704/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3523_ _3519_/Z _3534_/C _3460_/B _4246_/A1 _3942_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_7291_ _7291_/D _7302_/RN _7302_/CLK _7291_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold748 _7179_/Q hold748/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3454_ _3450_/Z _3534_/B _3454_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_4
X_6242_ _7275_/Q _6229_/Z _6242_/B _6242_/C _6246_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
Xhold759 _6752_/Q hold759/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3385_ _4684_/B _4686_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_20
X_6173_ hold89/I _6260_/A2 _6257_/A2 _7014_/Q _6176_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_111_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5124_ _5349_/A1 _5369_/A1 _5267_/C _5327_/B _5125_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_69_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5055_ _5215_/B _5053_/Z _5055_/A3 _5058_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_69_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4006_ _6703_/Q _4073_/B1 _4006_/B _4007_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_26_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_3_0_0__1374_ clkbuf_0__1374_/Z clkbuf_4_1_0__1374_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_52_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5957_ _6310_/A4 _6306_/A3 _6562_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_80_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4908_ _5290_/A1 _5369_/A2 _5200_/B _5290_/C _4910_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5888_ hold139/Z hold376/Z _5892_/S _7245_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4839_ _5466_/B _4694_/B _4759_/C _4869_/A3 _4841_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_107_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet733_364 net733_373/I _6890_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet733_353 _4109__3/I _6901_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6509_ _6788_/Q _4019_/Z _6509_/B _7302_/Q _6533_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_136_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_145 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xnet733_375 net833_474/I _6868_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet733_397 net733_397/I _6821_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet733_386 net833_470/I _6832_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_96_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold31 hold31/I hold31/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold20 hold20/I hold20/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_188_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold64 hold64/I hold64/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold42 hold42/I hold42/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold53 hold53/I hold53/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_88_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold86 hold86/I hold86/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold75 hold75/I hold75/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_29_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold97 hold97/I hold97/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_56_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_184_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_185_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_284 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_577 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6860_ _6860_/D _6862_/CLK _6860_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5811_ _5866_/A3 _5820_/A2 _3527_/Z _4227_/B _5819_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_62_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_474 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6791_ _6791_/D _7304_/RN _6791_/CLK _6791_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_188_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5742_ hold439/Z hold5/Z _5744_/S _7117_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5673_ _4227_/B _5718_/A3 _5820_/A2 _5866_/A3 _5681_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_175_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4624_ _4661_/C _4624_/A2 _5436_/A4 _5399_/B _5229_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4555_ _4555_/A1 _4555_/A2 _5051_/A1 _5230_/A2 _4555_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_128_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold501 _5594_/Z _6986_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7343_ _7343_/D _6695_/Z _4111_/I1 _7343_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold523 _6806_/Q hold523/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_144_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold545 _7162_/Q hold545/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3506_ _3507_/C _3833_/A2 _3811_/A1 _3473_/B _3962_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_104_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold512 _7090_/Q hold512/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold534 _7034_/Q hold534/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold556 _6801_/Q hold556/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4486_ _3379_/I _3380_/I _5484_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_131_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold578 _4377_/Z _6882_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7274_ _7274_/D _7302_/RN _7304_/CLK _7274_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
Xhold567 _6654_/Z _7340_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3437_ hold163/Z hold138/Z _3440_/S _7331_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_103_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6225_ _6225_/A1 _6225_/A2 _6225_/A3 _6225_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
Xhold589 _6890_/Q hold589/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3368_ _3368_/I _5641_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6156_ _7037_/Q _6258_/A2 _6258_/B1 _6997_/Q _6260_/A2 _7077_/Q _6162_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XTAP_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_861 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5107_ _5107_/A1 _5279_/A3 _5107_/B _5108_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_100_833 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_872 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_894 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6087_ _6788_/Q _6087_/A2 _6087_/A3 _6087_/B _6088_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XTAP_2728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5038_ _5087_/A2 _5039_/A1 _5038_/B _5291_/B _5041_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_38_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6989_ _6989_/D _7281_/RN _6989_/CLK _6989_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_13_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput110 wb_adr_i[23] _4916_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_163_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput154 wb_dat_i[4] _6628_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput143 wb_dat_i[23] _6640_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput132 wb_dat_i[13] _6631_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput121 wb_adr_i[4] _4684_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
XFILLER_76_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput165 wb_stb_i _4062_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_57_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_182 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4340_ _6600_/I0 _6850_/Q _4343_/S _6850_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4271_ hold160/Z hold25/Z _4281_/S _4271_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_4_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6010_ _6036_/A3 _6211_/C _6211_/B _7271_/Q _6256_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_67_533 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_750 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6912_ _6912_/D _6670_/Z _7346_/CLK _6912_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_63_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6843_ _6843_/D _7262_/RN _6843_/CLK _6843_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_51_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3986_ _6594_/A1 _3986_/A2 _3986_/B _6912_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6774_ _6774_/D _6665_/Z _4111_/I1 _6774_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_5725_ hold58/Z hold64/Z hold22/Z hold65/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_719 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5656_ hold391/Z hold858/Z _5663_/S _7040_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4607_ _4481_/C _5062_/A3 _4502_/B _4922_/B _5225_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_163_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold320 _7224_/Q hold320/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_5587_ hold164/Z hold238/Z _5590_/S _5587_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4538_ _5347_/A2 _5230_/A1 _5050_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xhold331 _7229_/Q hold331/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold353 _5643_/Z _7029_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_2_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7326_ _7326_/D _6680_/Z _7346_/CLK _7326_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold342 _5765_/Z _7137_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4469_ _4690_/B _5098_/A2 _4469_/B _4951_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_131_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold364 _7011_/Q hold364/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold375 _5761_/Z _7133_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_435 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7257_ _7257_/D _7281_/RN _7257_/CLK _7257_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold386 _5844_/Z _7207_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_132_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6208_ _7137_/Q _6257_/A2 _6258_/B1 _6749_/Q _6210_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold397 _5588_/Z _6981_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7188_ _7188_/D _7265_/RN _7188_/CLK _7188_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_133_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6139_ _6232_/C _6139_/A2 _6139_/B _6142_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2569 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1857 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1835 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1879 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1868 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_3_0__1374_ clkbuf_4_3_0__1374_/I clkbuf_4_3_0__1374_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_1_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3840_ _3840_/A1 _3840_/A2 _3841_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3771_ _7050_/Q _3973_/A2 _3980_/A2 _7066_/Q _3773_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_158_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5510_ hold391/Z hold632/Z _5511_/S _5510_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_185_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6490_ hold89/I _6292_/Z _6571_/C1 hold78/I _6490_/C _6491_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_145_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5441_ _5441_/A1 _5441_/A2 _5442_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_66_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5372_ _5372_/A1 _5376_/A1 _5372_/B _5373_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4323_ _4328_/S _6839_/Q _4324_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7111_ _7111_/D _7304_/RN _7111_/CLK _7111_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_7042_ _7042_/D _7302_/RN _7042_/CLK _7042_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_99_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4254_ hold255/Z hold139/Z _4262_/S _4254_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4185_ hold139/Z hold280/Z _4189_/S _4185_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6826_ _6826_/D _7304_/RN _6826_/CLK _6826_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_51_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6757_ _6757_/D _7262_/RN _6757_/CLK _6757_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_50_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5708_ hold2/Z hold228/Z _5708_/S _5708_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3969_ _7112_/Q _3969_/A2 _3969_/B1 _6742_/Q _3970_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6688_ _7265_/RN _6994_/Q _4026_/C _6688_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_164_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5639_ hold410/Z hold25/Z _5645_/S _5639_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_128_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_827 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold161 _6815_/Q hold161/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold150 _5604_/Z _6995_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_132_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7309_ _7309_/D _7313_/CLK _7309_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold172 _3484_/B hold172/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_144_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold194 _5653_/Z _7038_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_78_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold183 _6746_/Q hold183/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_120_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_867 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2322 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2355 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2399 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1654 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1687 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_606 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5990_ _6788_/Q _4019_/Z _6509_/B _6559_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_4941_ _4963_/B _4995_/A4 _5025_/A3 _4922_/B _5370_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_80_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4872_ _5502_/A2 _5468_/A1 _4667_/Z _5244_/A2 _4874_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6611_ _6880_/Q _6611_/A2 _6611_/B1 _6879_/Q _6613_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_178_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3823_ _3827_/A1 _4227_/A2 _3477_/Z _3496_/B _3854_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
Xnet583_251 net433_58/I _7018_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_158_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6542_ _6891_/Q _6292_/Z _6571_/B1 _6833_/Q _6571_/C1 _6770_/Q _6543_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
Xnet583_240 net783_420/I _7029_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3754_ _3753_/Z hold882/Z _3888_/S _6915_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3685_ _7166_/Q _3878_/A2 _3980_/B1 _6980_/Q _3687_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6473_ _7207_/Q _6573_/A2 _6288_/Z _7199_/Q _6297_/Z _7045_/Q _6474_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_9_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput200 _4082_/ZN mgmt_gpio_oeb[36] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5424_ _5424_/A1 _5424_/A2 _5424_/A3 _5424_/A4 _5458_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_173_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput233 _7372_/Z mgmt_gpio_out[31] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput211 _7355_/Z mgmt_gpio_out[11] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput222 _7362_/Z mgmt_gpio_out[21] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput244 _7354_/Z mgmt_gpio_out[7] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5355_ _5404_/B2 _5355_/A2 _5355_/B _5356_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput255 _4113_/I pad_flash_io1_ie VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput277 _6725_/Q pll_trim[15] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput266 _6926_/Q pll_div[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_160_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5286_ _5286_/A1 _5452_/A2 _5368_/A2 _5289_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_102_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput288 _6934_/Q pll_trim[25] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4306_ hold58/Z hold206/Z _4307_/S _4306_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xoutput299 _4121_/Z ser_rx VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_7025_ _7025_/D _7302_/RN _7025_/CLK _7025_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4237_ hold479/Z hold164/Z _4243_/S _4237_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_74_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_3_5__f_wb_clk_i clkbuf_0_wb_clk_i/Z _7323_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_67_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4168_ hold2/Z hold273/Z _4168_/S _4168_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4099_ _6971_/Q _4246_/A3 _4099_/B _4099_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6809_ _6809_/D input75/Z _6809_/CLK _7373_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_11_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1462 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3470_ _6863_/Q hold7/Z _3470_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_115_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet533_170 net433_58/I _7099_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet533_181 net433_76/I _7088_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet533_192 net633_277/I _7077_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_142_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5140_ _5376_/A1 _5489_/A2 _5502_/B1 _5502_/A2 _5141_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_69_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5071_ _5071_/A1 _5223_/B _5071_/A3 _5071_/A4 _5071_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_111_533 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4022_ input67/Z _6946_/Q _4026_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_56_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_845 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_54__1374_ clkbuf_4_12_0__1374_/Z net783_419/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_80_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5973_ _6312_/A4 _6311_/A1 _5973_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_64_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_837 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4924_ _4951_/B1 _4951_/B2 _4926_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_21_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4855_ _5294_/B _5294_/C _5466_/B _5258_/A3 _4857_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_159_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4786_ _4706_/Z _4825_/A4 _5476_/A1 _5255_/B _4791_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3806_ input12/Z _5748_/A3 _5532_/A3 _5528_/A2 _3849_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_181_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6525_ _7161_/Q _6286_/Z _6311_/C hold87/I _6581_/B1 hold47/I _6530_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_3737_ _3737_/A1 _3737_/A2 _3737_/A3 _3737_/A4 _3737_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_162_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3668_ _7207_/Q _3938_/A2 _3980_/A2 _7069_/Q _7053_/Q _3973_/A2 _3669_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6456_ _6788_/Q _4019_/Z _6509_/B _7300_/Q _6483_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5407_ _5407_/A1 _5406_/Z hold7/I _4365_/C _5408_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6387_ _7188_/Q _6274_/Z _6567_/B1 _7140_/Q _6311_/B _7228_/Q _6390_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_3599_ _6918_/Q _3597_/Z _3887_/S _3599_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_161_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5338_ _5338_/A1 _5338_/A2 _5338_/A3 _5338_/A4 _5338_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5269_ _5344_/B _5344_/C _5343_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7008_ _7008_/D _7302_/RN _7008_/CLK _7008_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_87_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet783_402 net783_433/I _6816_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet783_435 net783_435/I _6779_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet783_413 net783_417/I _6805_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet783_424 net783_424/I _6794_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_184_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet783_446 _4109__2/I _6763_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_109_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_164_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_829 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_853 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4640_ _5046_/C _5360_/C _5285_/A1 _5078_/A2 _5082_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_175_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_249 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6310_ _7276_/Q _6563_/A4 _6562_/A4 _6310_/A4 _6310_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_4571_ _4759_/C _4684_/B _5307_/B _4694_/B _5437_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_143_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3522_ _3454_/Z _3498_/B _4227_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xhold727 _6868_/Q hold727/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold716 _4170_/Z _6734_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold705 _4180_/Z _6741_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7290_ _7290_/D _7302_/RN _7302_/CLK _7290_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_171_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold749 _5813_/Z _7179_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3453_ _6863_/Q hold16/Z _3534_/B _3460_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xhold738 _5508_/Z _6911_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6241_ _6241_/A1 _7275_/Q _6241_/B1 _6241_/B2 _6242_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_170_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6172_ _7022_/Q _6259_/A2 _6261_/A2 _7006_/Q _6176_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3384_ _4922_/B _4759_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_16
X_5123_ _5123_/A1 _5293_/A2 _5123_/B _5206_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_124_691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5054_ _5351_/A1 _5351_/A2 _5463_/A1 _5350_/B _5055_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_57_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4005_ _4004_/Z hold901/Z _4015_/S _6704_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5956_ _6789_/Q _7276_/Q _5956_/B _7276_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_80_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4907_ _4661_/C _5445_/A3 _5194_/C _5253_/A1 _5479_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_52_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5887_ hold25/Z hold536/Z _5892_/S _7244_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4838_ _5177_/A3 _5437_/A4 _5468_/A1 _5428_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_147_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4769_ _4661_/C _5253_/A1 _5255_/B _5468_/B _5256_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_174_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet733_354 net433_74/I _6900_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet733_365 net783_445/I _6889_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_20_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6508_ _6508_/A1 _6508_/A2 _6508_/B _7301_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_161_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6439_ _7076_/Q _6292_/Z _6571_/B1 _6988_/Q _6571_/C1 _7182_/Q _6440_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
Xnet733_376 net783_445/I _6867_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet733_387 net833_480/I _6831_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet733_398 net733_398/I _6820_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_134_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold32 hold32/I hold32/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold21 hold21/I hold21/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold10 hold10/I hold10/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_102_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold54 hold54/I hold54/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold65 hold65/I hold65/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold43 hold43/I hold43/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold87 hold87/I hold87/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_75_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold76 hold76/I hold76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold98 hold98/I hold98/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_83_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_829 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_101_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_364 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_399 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6790_ _6790_/D _7302_/RN _7281_/CLK _6790_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_5810_ hold2/Z hold133/Z _5810_/S _5810_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_23_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5741_ hold487/Z hold164/Z _5744_/S _7116_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_867 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5672_ hold2/Z _7055_/Q hold30/Z hold31/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4623_ _5484_/A2 _5445_/A2 _5439_/C _5399_/B _4627_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_129_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4554_ _5389_/A2 _5226_/A1 _5323_/A1 _5484_/A4 _4555_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_129_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold502 _7002_/Q hold502/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7342_ _7342_/D _6694_/Z _7346_/CLK _7342_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold524 _4282_/Z _6806_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold513 _7165_/Q hold513/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3505_ _3511_/C _3604_/A2 _5534_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_7273_ _7273_/D _7302_/RN _7304_/CLK _7273_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
Xhold535 _5649_/Z _7034_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold546 _6804_/Q hold546/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold557 _4272_/Z _6801_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4485_ _5201_/C _6879_/Q _4683_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6224_ _6881_/Q _6258_/A2 _6259_/A2 _6866_/Q _6261_/B1 _6883_/Q _6225_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
Xhold579 _6853_/Q hold579/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold568 _6757_/Q hold568/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3436_ hold4/Z hold163/Z _3440_/S _7332_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_106_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3367_ _7035_/Q _3367_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6155_ _7053_/Q _6256_/A2 _6262_/B1 _7029_/Q _6162_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5106_ _5412_/A1 _5106_/A2 _5106_/A3 _5106_/A4 _5107_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_100_823 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6086_ _6788_/Q _7286_/Q _6087_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_873 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5037_ _5037_/A1 _5290_/C _4718_/C _5290_/B _5291_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_85_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6988_ _6988_/D _7281_/RN _6988_/CLK _6988_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_40_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5939_ _6107_/B _6789_/Q _6235_/A1 _5940_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_182_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput111 wb_adr_i[24] _4060_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput100 wb_adr_i[14] _4413_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_163_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput144 wb_dat_i[24] _6611_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput122 wb_adr_i[5] _5307_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
Xinput133 wb_dat_i[14] _6635_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_76_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xinput166 wb_we_i _6648_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput155 wb_dat_i[5] _6632_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_797 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4270_ _4269_/Z hold866/Z _4282_/S _4270_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6911_ _6911_/D _7341_/RN _6911_/CLK _6911_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_48_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6842_ _6842_/D _7313_/CLK _6842_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3985_ _7338_/Q _6776_/Q _3887_/S _3986_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6773_ _6773_/D _7262_/RN _6773_/CLK _6773_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5724_ hold5/Z hold120/Z hold22/Z _5724_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5655_ _4227_/B hold29/Z _5727_/A3 _5655_/A4 _5663_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_175_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4606_ _4606_/A1 _4606_/A2 _5223_/C _5071_/A4 _4610_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_164_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold310 _5632_/Z _7020_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5586_ hold139/Z hold418/Z _5590_/S _5586_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7325_ _7325_/D _6679_/Z _7346_/CLK _7325_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnsnq_1
Xhold332 _7098_/Q hold332/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4537_ _4454_/B _5225_/A3 _5225_/A1 _4960_/C _5230_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
Xhold321 _5864_/Z _7224_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold343 _7225_/Q hold343/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold354 _7050_/Q hold354/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold387 _7328_/Q hold387/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4468_ _5046_/A1 _5046_/A2 _5078_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
Xhold365 _5622_/Z _7011_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_117_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold376 _7245_/Q hold376/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7256_ _7256_/D _7281_/RN _7256_/CLK _7256_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_7187_ _7187_/D _7341_/RN _7187_/CLK _7187_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
Xhold398 _7368_/I hold398/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_89_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6207_ _7209_/Q _6256_/B1 _6257_/B1 hold50/I _6259_/B1 _7111_/Q _6210_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_3419_ _6709_/Q _6707_/Q _6774_/Q _3442_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6138_ _6138_/A1 _6232_/C _6138_/B _6138_/C _6139_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4399_ _4405_/A3 _5535_/B _6653_/A2 _5838_/A2 _4401_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_58_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6069_ _7090_/Q _6262_/A2 _6260_/B1 _6986_/Q _6070_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_73_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2537 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1825 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1847 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1836 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_179_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_789 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_177_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3770_ _7212_/Q _3940_/A2 _3950_/B1 _7042_/Q _3953_/B1 _7188_/Q _3773_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_157_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5440_ _5440_/A1 _5440_/A2 _5440_/A3 _5440_/A4 _5441_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_8_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5371_ _5371_/A1 _5371_/A2 _5371_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_114_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4322_ _6597_/I0 _6838_/Q _4328_/S _6838_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7110_ hold61/Z _7304_/RN _7110_/CLK hold60/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_141_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4253_ hold619/Z _4252_/Z _4263_/S _4253_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7041_ _7041_/D _7302_/RN _7041_/CLK _7041_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_141_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4184_ hold25/Z hold326/Z _4189_/S _6744_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_3_4__f_wb_clk_i clkbuf_0_wb_clk_i/Z _7322_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_82_356 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6825_ _6825_/D _7304_/RN _6825_/CLK _6825_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3968_ _7104_/Q _3968_/A2 _3968_/B1 _6766_/Q _3968_/C _3970_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_6756_ _6756_/D _7262_/RN _6756_/CLK _6756_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_137_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5707_ hold58/Z hold215/Z _5708_/S _5707_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6687_ _7265_/RN _6994_/Q _4026_/C _6687_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_149_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3899_ _5534_/A1 _3519_/Z _3473_/B hold462/Z _5535_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_163_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5638_ hold669/Z hold388/Z _5645_/S _5638_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5569_ hold164/Z hold185/Z hold38/Z _6964_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_152_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold162 _4293_/Z _6815_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold151 _7199_/Q hold151/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7308_ _7308_/D _7313_/CLK _7308_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold140 _5806_/Z _7173_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold173 hold173/I hold173/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold195 _6943_/Q hold195/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold184 _4186_/Z _6746_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7239_ _7239_/D _7265_/RN _7239_/CLK _7239_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_144_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_832 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2356 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1644 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1677 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4940_ _4684_/B _4425_/Z _5026_/B _5025_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_64_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4871_ _4871_/A1 _4871_/A2 _4871_/A3 _4874_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_60_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6610_ _6610_/A1 _6610_/A2 _4362_/Z _6642_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_3822_ _7049_/Q hold21/I _5745_/A4 _4405_/A3 _3873_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_60_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6541_ _6754_/Q _6570_/A2 _6570_/B1 _6887_/Q _6570_/C1 _6843_/Q _6543_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_146_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet583_230 net633_289/I _7039_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet583_241 net633_281/I _7028_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3753_ _6914_/Q _6597_/I0 _3887_/S _3753_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3684_ _7052_/Q _3973_/A2 _3950_/B1 _7044_/Q _3950_/A2 _7100_/Q _3687_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6472_ _7191_/Q _6274_/Z _6294_/Z _7037_/Q _6472_/C _6474_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
Xoutput201 _4080_/ZN mgmt_gpio_oeb[37] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_173_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5423_ _5422_/Z _5457_/A3 _5458_/A1 _5425_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_145_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_14__1374_ clkbuf_4_8_0__1374_/Z net683_314/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5354_ _5464_/A3 _5352_/Z _5357_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput234 _4085_/Z mgmt_gpio_out[32] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_145_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput212 _7356_/Z mgmt_gpio_out[12] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput223 _7363_/Z mgmt_gpio_out[22] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xclkbuf_leaf_77__1374_ clkbuf_4_5_0__1374_/Z net833_464/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_114_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput245 _4090_/Z mgmt_gpio_out[8] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput267 _6920_/Q pll_ena VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput256 _4113_/ZN pad_flash_io1_oe VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4305_ hold5/Z hold224/Z _4307_/S _4305_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5285_ _5285_/A1 _5451_/A1 _5091_/C _5285_/B2 _5285_/C _5368_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_99_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput289 _6728_/Q pll_trim[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput278 _6710_/Q pll_trim[16] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4236_ hold553/Z _4235_/Z _4244_/S _4236_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7024_ _7024_/D _7281_/RN _7024_/CLK _7024_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_68_640 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4167_ hold58/Z hold383/Z _4168_/S _4167_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_28_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4098_ _6994_/Q _7325_/Q _4026_/C _4099_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_43_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6808_ _6808_/D input75/Z _6808_/CLK _6808_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_168_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6739_ _6739_/D _7262_/RN _6739_/CLK _6739_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_149_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1474 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet533_171 net433_86/I _7098_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet533_182 net633_273/I _7087_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet533_160 net533_163/I _7109_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet533_193 net433_89/I _7076_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_123_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5070_ _5071_/A4 _5071_/A3 _5419_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4021_ _7342_/Q hold44/I _4025_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_111_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5972_ _6310_/A4 _6306_/A3 _6324_/A1 _6323_/A1 _6311_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_92_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_1__1374_ clkbuf_4_2_0__1374_/Z net783_430/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4923_ _4922_/B _4951_/A1 _5502_/B2 _4425_/Z _4961_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_178_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4854_ _5466_/A1 _5466_/A2 _5294_/B _5294_/C _4857_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_60_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4785_ _5253_/A1 _5257_/B1 _4785_/B _4791_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_21_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3805_ _6761_/Q _5784_/A2 _5838_/A2 _5518_/A1 _3855_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6524_ _6517_/Z _6524_/A2 _6523_/Z _6531_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3736_ _7173_/Q _3966_/A2 _3958_/B1 _6721_/Q _3737_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_180_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3667_ input49/Z _4243_/S _3975_/B1 _7376_/I _3669_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6455_ _6455_/A1 _6455_/A2 _6455_/B _7299_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5406_ _5444_/B _5444_/A2 _5479_/A2 _4362_/Z _5406_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_115_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6386_ _6383_/Z _6386_/A2 _6386_/A3 _6386_/A4 _6397_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3598_ _7338_/Q _6776_/Q _3888_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_125_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5337_ _5489_/A1 _5337_/A2 _5489_/B1 _5399_/B _5338_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5268_ _5199_/B _5376_/A1 _5471_/C _5343_/C _5270_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_102_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7007_ hold88/Z _7281_/RN _7007_/CLK hold87/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4219_ hold388/Z hold691/Z _4219_/S _6769_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5199_ _5093_/B _5199_/A2 _5199_/B _5344_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_29_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet783_403 net783_433/I _6815_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_169_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet783_414 net783_414/I _6804_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_11_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet783_425 net783_425/I _6793_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_34_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet783_447 net833_470/I _6762_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet783_436 net833_469/I _6773_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_156_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_60__1374_ _4109__12/I net433_62/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_121_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1293 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4570_ _5420_/A1 _5315_/A4 _5262_/A4 _4423_/Z _4576_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_155_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3521_ _3460_/B _3534_/C _5548_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_183_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold728 _4373_/Z _6868_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold706 _6844_/Q hold706/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_7_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold717 _6761_/Q hold717/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_170_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3452_ _4016_/A2 _6777_/Q _3452_/B _3498_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_6240_ _6240_/A1 _6240_/A2 _6240_/A3 _6240_/A4 _6241_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xhold739 _6936_/Q hold739/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3383_ _4694_/B _4469_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_12
X_6171_ _7038_/Q _6258_/A2 _6262_/B1 _7030_/Q _6261_/B1 _7046_/Q _6177_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_41_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5122_ _5410_/A2 _5026_/C _3379_/I _5153_/A2 _5293_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_69_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5053_ _5421_/A1 _5053_/A2 _5053_/A3 _5211_/B _5053_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_4004_ hold171/I _4004_/A2 _4004_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_1_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5955_ _6787_/Q _6789_/Q _7276_/Q _5956_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_179_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5886_ hold388/Z hold741/Z _5892_/S _7243_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4906_ _5290_/C _4916_/A3 _4916_/A2 _4959_/A2 _5404_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_40_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4837_ _5466_/B _3379_/I _5315_/A4 _5037_/A1 _5489_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_181_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4768_ _3379_/I _5489_/A2 _5315_/A4 _5445_/A2 _4770_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_5_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet733_355 net433_75/I _6899_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4699_ _4767_/A3 _4723_/A2 _5152_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_3719_ _3716_/Z _3719_/A2 _3719_/B _6916_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6507_ _7300_/Q _6587_/A2 _6532_/B _6532_/C _6508_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_6438_ _7214_/Q _6570_/A2 _6570_/B1 _7060_/Q _6570_/C1 _6996_/Q _6440_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_105_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet733_366 net433_74/I _6888_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet733_377 _4109__16/I _6866_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet733_388 net783_427/I _6830_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet733_399 net783_411/I _6819_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_161_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6369_ _7089_/Q _6578_/A2 _6310_/Z _6977_/Q _6578_/C1 _7171_/Q _6371_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_29_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold11 hold11/I hold11/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold22 hold22/I hold22/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_130_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_640 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold33 hold33/I hold33/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold55 hold55/I hold55/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold44 hold44/I hold44/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_75_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold66 hold66/I hold66/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold77 hold77/I hold77/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold88 hold88/I hold88/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold99 hold99/I hold99/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_72_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_101_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_0_mgmt_gpio_in[4] mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_31_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5740_ hold263/Z hold139/Z _5744_/S _5740_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_188_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1090 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5671_ hold58/Z hold67/Z hold30/Z _7054_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4622_ _4469_/B _4759_/C _4684_/B _5307_/B _5187_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_4553_ _5466_/C _4661_/C _4718_/B _4487_/Z _5351_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_128_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7341_ _7341_/D _7341_/RN _7341_/CLK _7341_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4484_ _5078_/A2 _5360_/C _4437_/Z _5046_/C _5081_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3504_ hold462/Z _3473_/B _5902_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold514 _7189_/Q hold514/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold503 _5612_/Z _7002_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold525 _7257_/Q hold525/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7272_ _7272_/D _7302_/RN _7281_/CLK _7272_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_7_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold536 _7244_/Q hold536/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3435_ hold57/Z hold4/Z _3440_/S _7333_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold547 _4278_/Z _6804_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold558 _7261_/Q hold558/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6223_ _6885_/Q _6256_/A2 _6259_/B1 _6831_/Q _6225_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold569 _4201_/Z _6757_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_143_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3366_ _7043_/Q _3366_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6154_ _6989_/Q _6260_/B1 _6261_/B1 _7045_/Q _6162_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_830 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_852 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5105_ _5105_/A1 _5272_/B _4437_/Z _5454_/B1 _5105_/C _5106_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_112_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6085_ _6107_/B _6107_/C _6970_/Q _7275_/Q _6087_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XTAP_874 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_863 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5036_ _5226_/A1 _5036_/A2 _5039_/A1 _5312_/B _5293_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_85_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_896 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2719 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6987_ _6987_/D _7302_/RN _6987_/CLK _6987_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_53_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5938_ _6036_/A3 _6103_/A1 _6107_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_41_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5869_ hold467/Z hold25/Z _5874_/S _7228_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_166_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput101 wb_adr_i[15] _4413_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput145 wb_dat_i[25] _6615_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput134 wb_dat_i[15] _6639_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput123 wb_adr_i[6] _4694_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_16
Xinput112 wb_adr_i[25] _3338_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_103_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput156 wb_dat_i[6] _6636_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_102_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_173_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_3_3__f_wb_clk_i clkbuf_0_wb_clk_i/Z _7304_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_94_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6910_ _6910_/D _7341_/RN _6910_/CLK _6910_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_54_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6841_ _6841_/D _7313_/CLK _6841_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3984_ _3984_/A1 _3984_/A2 _3984_/A3 _3983_/Z _6594_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_23_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6772_ _6772_/D _7262_/RN _6772_/CLK _6772_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_188_481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5723_ hold164/Z hold316/Z hold22/Z _5723_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5654_ hold2/Z hold85/Z _5654_/S hold86/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4605_ _4443_/Z _5459_/A3 _5323_/A1 _5180_/B _5071_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_148_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5585_ hold25/Z hold400/Z _5590_/S _5585_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold311 _6712_/Q hold311/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold300 _5730_/Z _7106_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7324_ _7324_/D _6678_/Z _7346_/CLK hold44/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
Xhold322 _7099_/Q hold322/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold333 _5721_/Z _7098_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4536_ _4469_/B _4759_/C _4686_/B _5312_/B _5290_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_104_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold344 _5865_/Z _7225_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4467_ _3380_/I _5011_/A2 _4578_/B _5062_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xhold366 _6963_/Q hold366/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_132_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold377 _6989_/Q hold377/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_117_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7255_ _7255_/D _7281_/RN _7255_/CLK _7255_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold355 _6982_/Q hold355/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold388 _4137_/Z hold388/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7186_ _7186_/D _7341_/RN _7186_/CLK _7186_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
Xhold399 _5559_/Z _6955_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6206_ _6206_/A1 _6206_/A2 _6206_/A3 _6206_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_4398_ hold388/Z hold602/Z _4398_/S _4398_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3418_ input58/Z _7338_/Q _3418_/S _7338_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3349_ _7173_/Q _3349_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_98_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6137_ _7158_/Q _6258_/A2 _6137_/B _6137_/C _6138_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6068_ _7058_/Q _6257_/B1 _6259_/B1 _6978_/Q _6070_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_73_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5019_ _5353_/A3 _4947_/C _4963_/B _5288_/A4 _5020_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XTAP_2527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_165_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1848 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1837 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_182_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_827 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_877 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5370_ _5370_/A1 _5498_/B1 _5370_/B _5371_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_126_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4321_ _3790_/Z _6837_/Q _4328_/S _6837_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4252_ hold269/Z hold25/Z _4262_/S _4252_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7040_ _7040_/D _7302_/RN _7040_/CLK _7040_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_68_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4183_ hold388/Z hold699/Z _4189_/S _6743_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_94_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_37__1374_ clkbuf_4_14_0__1374_/Z net433_53/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_36_796 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6824_ _6824_/D _7304_/RN _6824_/CLK _6824_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_63_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3967_ _3967_/A1 _3967_/A2 _3967_/A3 _3971_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6755_ _6755_/D _7262_/RN _6755_/CLK _6755_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5706_ hold5/Z hold204/Z _5708_/S _5706_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6686_ _7265_/RN _6994_/Q _4026_/C _6686_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_164_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3898_ _6864_/Q _4378_/A1 _5893_/A3 _5546_/A2 _3937_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5637_ hold634/Z hold391/Z _5645_/S _5637_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_151_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5568_ hold139/Z hold366/Z hold38/Z _6963_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4519_ _4469_/B _4922_/B _4684_/B _5307_/B _5208_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
Xhold152 _7059_/Q hold152/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold130 _7022_/Q hold130/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7307_ _7307_/D _7313_/CLK _7307_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold141 _6749_/Q hold141/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold163 _7331_/Q hold163/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold185 _6964_/Q hold185/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7238_ _7238_/D _7341_/RN _7238_/CLK _7238_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5499_ _5373_/Z _5411_/Z _5455_/Z _5499_/A4 _5500_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_144_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold174 hold174/I _5551_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold196 _5542_/Z _6943_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7169_ hold10/Z _7265_/RN _7169_/CLK _7169_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_58_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2324 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1612 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_749 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1678 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_652 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4870_ _5034_/A2 _5466_/B _5392_/A1 _5503_/A1 _4871_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_177_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3821_ _7171_/Q _5856_/A1 _5802_/A2 _3527_/Z _3853_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6540_ _6540_/A1 _6540_/A2 _6540_/A3 _6540_/A4 _6540_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_186_782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet583_220 net433_59/I _7049_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_146_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3752_ _3752_/A1 _3752_/A2 _3752_/A3 _6597_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
Xnet583_231 net633_290/I _7038_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet583_242 net783_420/I _7027_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_71_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6471_ _6471_/A1 _6471_/A2 _6472_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3683_ input16/Z _5748_/A3 _5532_/A3 _5528_/A2 _3691_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5422_ _5462_/A1 _5462_/A2 _5421_/Z _5422_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_146_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput235 _4086_/Z mgmt_gpio_out[33] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_161_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5353_ _5051_/B _4454_/B _5353_/A3 _4959_/C _5360_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
Xoutput213 _4104_/Z mgmt_gpio_out[13] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput224 _7364_/Z mgmt_gpio_out[23] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput202 _3372_/ZN mgmt_gpio_oeb[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_126_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput246 _4089_/Z mgmt_gpio_out[9] VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_1
Xoutput257 _6930_/Q pll90_sel[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput268 _6927_/Q pll_sel[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4304_ hold164/Z hold313/Z _4307_/S _4304_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_142_896 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5284_ _5378_/A1 _5498_/A2 _5452_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput279 _6711_/Q pll_trim[17] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4235_ hold147/Z hold139/Z _4243_/S _4235_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7023_ hold53/Z _7265_/RN _7023_/CLK hold52/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_101_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4166_ hold5/Z hold412/Z _4168_/S _4166_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4097_ _6791_/Q input3/Z input1/Z _4097_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_55_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_711 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6807_ _6807_/D input75/Z _6807_/CLK _6807_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4999_ _4661_/C _4956_/B _5279_/B _5002_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6738_ _6738_/D _7262_/RN _6738_/CLK _6738_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_137_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6669_ input75/Z _6994_/Q _4026_/C _6669_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_152_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_847 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_20__1374_ _4109__51/I net433_82/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_2165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1431 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_100__1374_ clkbuf_4_4_0__1374_/Z net833_498/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_159_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1464 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_83__1374_ clkbuf_4_4_0__1374_/Z net433_97/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_15_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1497 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_170_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet533_172 net433_56/I _7097_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_108_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet533_161 net833_498/I _7108_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet533_194 net583_214/I _7075_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_124_896 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet533_183 net583_245/I _7086_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_151_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4020_ _4020_/A1 _4020_/A2 _3421_/B _3387_/Z _6774_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_77_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5971_ _5971_/A1 _5971_/A2 _7279_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4922_ _5136_/A2 _5098_/A2 _4922_/B _4951_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_4853_ _5389_/B _4853_/A2 _4853_/B _4858_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4784_ _4784_/A1 _4784_/A2 _5334_/B _4785_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_20_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3804_ _3496_/B _5534_/A2 _4246_/A2 _3477_/Z _3955_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_158_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6523_ _6523_/A1 _6523_/A2 _6523_/A3 _6523_/A4 _6523_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_3735_ _7115_/Q _3969_/A2 _3959_/A2 _6729_/Q _3969_/B1 _6745_/Q _3737_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_134_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_145 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6454_ _7298_/Q _6587_/A2 _6532_/B _6532_/C _6455_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5405_ _5480_/A2 _5405_/A2 _5482_/A1 _5479_/A3 _5407_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_118_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3666_ _7135_/Q _3945_/A2 _3953_/A2 _6997_/Q _3786_/B1 _5546_/A2 _3669_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_161_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6385_ _7074_/Q _6292_/Z _6571_/B1 _6986_/Q _6571_/C1 _7180_/Q _6386_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_3597_ _3597_/A1 _3597_/A2 _3597_/A3 _3597_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_142_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5336_ _5336_/A1 _5490_/A3 _5470_/A1 _5336_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_5267_ _5290_/A1 _5353_/A3 _5267_/B _5267_/C _5471_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_88_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7006_ _7006_/D _7281_/RN _7006_/CLK _7006_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_85_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4218_ hold391/Z hold784/Z _4219_/S _6768_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5198_ _5084_/C _5295_/A1 _5290_/C _5198_/B _5424_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_4149_ hold1/Z _7321_/Q _6863_/Q hold2/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_95_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet783_404 net783_433/I _6814_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet783_415 net783_415/I _6803_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_157_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet783_426 net783_426/I _6792_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_70_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet783_437 net783_437/I _6772_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet783_448 net833_454/I _6761_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_7_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_711 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_116_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3520_ _3604_/A2 _3519_/Z _3511_/C _3833_/A2 _3977_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xhold707 _4331_/Z _6844_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_6_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold718 _4207_/Z _6761_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_170_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3451_ hold11/Z _6777_/Q _3491_/B _3452_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold729 _7203_/Q hold729/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3382_ _4661_/C _5235_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_16
X_6170_ hold67/I _6256_/A2 _6256_/B1 _7086_/Q _6177_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5121_ _5355_/A2 _5381_/A2 _5121_/B _5291_/B _5123_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_69_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5052_ _5351_/A1 _5052_/A2 _5463_/A1 _5463_/B _5052_/C _5053_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_4003_ _6777_/Q _3993_/Z _6703_/Q _4004_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_93_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5954_ _5954_/A1 _5954_/A2 _7275_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_178_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4905_ _4905_/A1 _4905_/A2 _4905_/A3 _4910_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5885_ hold391/Z hold863/Z _5892_/S _7242_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4836_ _5177_/A3 _5153_/A2 _5153_/B _5502_/A2 _5256_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4767_ _5327_/B _4922_/B _4767_/A3 _4822_/A4 _5489_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_6506_ _6506_/A1 _6506_/A2 _6974_/Q _6584_/A1 _6584_/B _6508_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_4698_ _4767_/A3 _4723_/A2 _5468_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_107_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet733_356 _4109__3/I _6898_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3718_ _3888_/S _6916_/Q _3719_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_162_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3649_ _7013_/Q _3962_/A2 _3981_/A2 _7247_/Q _7263_/Q _3964_/C1 _3654_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
Xnet733_367 net433_67/I _6887_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6437_ _6437_/A1 _6437_/A2 _6437_/A3 _6437_/A4 _6446_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xnet733_378 net833_474/I _6865_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet733_389 net783_427/I _6829_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6368_ _7251_/Q _6580_/B1 _6309_/Z _7235_/Q _6743_/Q _6579_/A2 _6371_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_161_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5319_ _5319_/A1 _5481_/A1 _5481_/A2 _5322_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_102_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold12 hold12/I hold12/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold23 hold23/I hold23/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6299_ _7279_/Q _7278_/Q _6563_/A3 _6562_/A4 _6299_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_88_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold56 hold56/I hold56/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold45 hold45/I hold45/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold34 hold34/I hold34/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_103_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold67 hold67/I hold67/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold89 hold89/I hold89/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold78 hold78/I hold78/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_152_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_43_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_322 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_500 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_355 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_541 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_180_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_3_2__f_wb_clk_i clkbuf_0_wb_clk_i/Z _7302_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_121_674 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_187_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5670_ hold5/Z hold114/Z hold30/Z _7053_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1091 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4621_ _4686_/B _5312_/B _4694_/B _4922_/B _5399_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_176_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4552_ _5262_/A4 _5315_/A4 _5301_/A2 _5235_/A1 _5435_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_7340_ _7340_/D _7341_/RN _7340_/CLK _7340_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_183_390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4483_ _4437_/Z _4682_/A2 _5051_/B _5459_/A3 _5201_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
Xhold515 _5824_/Z _7189_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3503_ _3515_/A2 _3827_/A2 _3811_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xhold504 _7366_/I hold504/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7271_ _7271_/D _7302_/RN _7281_/CLK _7271_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_7_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold526 _6924_/Q hold526/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold548 _7234_/Q hold548/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3434_ hold1/Z hold57/Z _3440_/S _7334_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_171_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold559 _5906_/Z _7261_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6222_ _6833_/Q _6260_/B1 _6257_/B1 _6887_/Q _6225_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold537 _6931_/Q hold537/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_143_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3365_ _7051_/Q _3365_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6153_ _6232_/C _7101_/Q _6211_/B _6211_/C _6163_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_820 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_831 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_842 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_853 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5104_ _4926_/C _5288_/A4 _5271_/A4 _5104_/B1 _4965_/C _5272_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_111_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6084_ _6084_/A1 _6084_/A2 _6084_/B _6087_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_875 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_864 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5035_ _5235_/A1 _5294_/A1 _5290_/C _5290_/B _5038_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_73_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6986_ _6986_/D _7281_/RN _6986_/CLK _6986_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_179_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5937_ _7272_/Q _7271_/Q _6266_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_25_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5868_ hold519/Z hold388/Z _5874_/S _7227_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5799_ hold5/Z hold106/Z hold9/Z _7167_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4819_ _4690_/C _4487_/Z _5267_/B _4819_/A4 _5432_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_31_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput102 wb_adr_i[16] _4418_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_103_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput135 wb_dat_i[16] _6612_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput124 wb_adr_i[7] _4922_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
Xinput113 wb_adr_i[26] _4057_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_130_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput146 wb_dat_i[26] _6619_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput157 wb_dat_i[7] _6640_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_102_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_750 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_606 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet633_300 net833_464/I _6969_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_36_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6840_ _6840_/D _7313_/CLK _6840_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6771_ _6771_/D _7262_/RN _6771_/CLK _6771_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_188_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5722_ hold139/Z hold322/Z hold22/Z _5722_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3983_ _3983_/A1 _3983_/A2 _3983_/A3 _3983_/A4 _3983_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_176_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5653_ hold58/Z hold193/Z _5654_/S _5653_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4604_ _4443_/Z _5459_/A3 _5226_/A1 _5180_/B _5223_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5584_ hold388/Z hold676/Z _5590_/S _5584_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7323_ _7323_/D _7323_/RN _7323_/CLK _7323_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4535_ _4694_/B _4922_/B _4684_/B _5307_/B _5445_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xhold301 _7232_/Q hold301/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_7_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold323 _5722_/Z _7099_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold312 _4140_/Z _6712_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold334 _7158_/Q hold334/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4466_ _4686_/B _5223_/A1 _5046_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xhold367 _7082_/Q hold367/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold345 _7231_/Q hold345/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_132_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold378 _5597_/Z _6989_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7254_ _7254_/D _7341_/RN _7254_/CLK _7254_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_89_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold356 _5589_/Z _6982_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7185_ hold51/Z _7265_/RN _7185_/CLK hold50/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold389 _4404_/Z _6900_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6205_ _7161_/Q _6258_/A2 _6259_/A2 _7145_/Q _6260_/A2 _7201_/Q _6206_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_3417_ _6707_/Q _6774_/Q _3417_/A3 _3418_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4397_ hold391/Z hold600/Z _4398_/S _4397_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3348_ _7181_/Q _3348_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_97_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6136_ _6136_/A1 _6136_/A2 _6136_/A3 _6137_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_867 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6067_ _7050_/Q _6256_/A2 _6261_/B1 _7042_/Q _6070_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_27_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5018_ _5018_/A1 _5016_/Z _5018_/A3 _5020_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_2517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1816 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1827 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6969_ _6969_/D _7304_/RN _6969_/CLK _6969_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_41_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_827 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold890 _7336_/Q _3428_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_89_661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4320_ _6595_/I0 _6836_/Q _4328_/S _6836_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_114_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4251_ hold861/Z _4250_/Z _4263_/S _4251_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_4_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_867 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4182_ hold391/Z hold805/Z _4189_/S _6742_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_675 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6823_ _6823_/D _7304_/RN _6823_/CLK _6823_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_149_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6754_ _6754_/D _7262_/RN _6754_/CLK _6754_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_11_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3966_ _7170_/Q _3966_/A2 _3966_/B _3966_/C _3967_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_50_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6685_ _7265_/RN _6994_/Q _4026_/C _6685_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_5705_ hold164/Z hold379/Z _5708_/S _5705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_10_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5636_ _5646_/A2 _4227_/B hold13/Z _5727_/A3 _5645_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3897_ _6866_/Q _4378_/A1 _5838_/A2 _4405_/A2 _3937_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_128_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5567_ hold25/Z hold160/Z hold38/Z _6962_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_145_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4518_ _4759_/C _4686_/B _5312_/B _4694_/B _5389_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_5498_ _5372_/B _5498_/A2 _5498_/B1 _5279_/B _5498_/C _5499_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
Xhold120 _7101_/Q hold120/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold153 _7091_/Q hold153/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold131 _5634_/Z _7022_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7306_ _7306_/D _7313_/CLK _7306_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold142 _4189_/Z _6749_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_2_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7237_ _7237_/D _7341_/RN _7237_/CLK _7237_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold175 _5549_/Z _6947_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold186 _7019_/Q hold186/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4449_ _4451_/B _4774_/B _4778_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_1
Xhold164 _4143_/Z hold164/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_5_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold197 _6828_/Q hold197/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_58_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7168_ _7168_/D _7265_/RN _7168_/CLK _7168_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_113_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_642 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7099_ _7099_/D _7265_/RN _7099_/CLK _7099_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_85_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6119_ _6988_/Q _6260_/B1 _6261_/B1 _7044_/Q _6125_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_74_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2358 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1679 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_43__1374_ clkbuf_4_15_0__1374_/Z net783_433/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_68_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_797 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3820_ _3827_/A1 _4246_/A2 _3477_/Z _3496_/B _3846_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_3751_ _3751_/A1 _3751_/A2 _3751_/A3 _3751_/A4 _3752_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_185_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet583_221 net433_59/I _7048_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_174_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet583_210 net783_414/I _7059_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet583_232 _4109__14/I _7037_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet583_243 net633_289/I _7026_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_173_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6470_ hold93/I _6285_/Z _6564_/C1 _7085_/Q _6471_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3682_ _7206_/Q hold21/I _5838_/A2 _3527_/Z _3687_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5421_ _5421_/A1 _5421_/A2 _5421_/A3 _5421_/A4 _5421_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_173_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5352_ _5421_/A1 _5421_/A2 _5421_/A3 _5352_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_173_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_160_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput225 _7365_/Z mgmt_gpio_out[24] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput214 _4103_/Z mgmt_gpio_out[14] VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_1
XFILLER_99_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput203 _3371_/ZN mgmt_gpio_oeb[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput236 _7373_/Z mgmt_gpio_out[34] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_160_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput258 _6931_/Q pll90_sel[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4303_ hold139/Z hold255/Z _4307_/S _4303_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xoutput247 _4111_/Z pad_flash_clk VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_1
X_5283_ _5282_/B _5498_/A2 _5283_/B _5286_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_142_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7022_ _7022_/D _7265_/RN _7022_/CLK _7022_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_114_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput269 _6928_/Q pll_sel[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4234_ hold560/Z _4233_/Z _4244_/S _4234_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_114_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_249 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4165_ hold164/Z hold446/Z _4168_/S _4165_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4096_ _7343_/Q _4118_/A1 _4096_/B _4096_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_83_689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6806_ _6806_/D _7281_/RN _6806_/CLK _6806_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_24_789 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_3_0__1374_ clkbuf_0__1374_/Z clkbuf_4_7_0__1374_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_51_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4998_ _4998_/A1 _5109_/A1 _4998_/A3 _5002_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_11_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3949_ _3949_/A1 _3949_/A2 _3949_/A3 _3949_/A4 _3984_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_6737_ _6737_/D _7262_/RN _6737_/CLK _6737_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_176_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6668_ input75/Z _6994_/Q _4026_/C _6668_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_136_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5619_ hold391/Z hold816/Z _5626_/S _5619_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6599_ _6599_/A1 _6603_/S _6599_/B _7310_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_837 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_175_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1498 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet533_173 net433_91/I _7096_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_135_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xnet533_162 net633_301/I _7107_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet533_195 _4109__29/I _7074_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_124_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet533_184 net633_289/I _7085_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_69_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_612 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_837 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5970_ _5966_/Z _7279_/Q _5971_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_18_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_829 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4921_ _4951_/A1 _4951_/A2 _4995_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_92_497 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4852_ _5375_/A1 _3380_/I _4852_/B1 _5466_/A2 _4853_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_61_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3803_ _7089_/Q _3951_/B1 _3803_/B1 _6902_/Q _3861_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_165_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4783_ _4706_/Z _4825_/A4 _5489_/A1 _5255_/B _5334_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_20_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6522_ _7153_/Q _6575_/A2 _6566_/C1 hold52/I _6523_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_9_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3734_ input14/Z _3971_/A2 _3850_/B1 input6/Z _3737_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3665_ input17/Z _3971_/A2 _3665_/B _3665_/C _3678_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_6453_ _6972_/Q _6584_/A1 _6453_/B _6584_/B _6455_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_161_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5404_ _5194_/C _5404_/A2 _5404_/B1 _5404_/B2 _5482_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_118_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6384_ _7212_/Q _6570_/A2 _6570_/B1 _7058_/Q _6570_/C1 _6994_/Q _6386_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_3596_ _3596_/A1 _3586_/Z _3595_/Z _3597_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_125_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5335_ _5335_/A1 _5335_/A2 _5335_/A3 _5470_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_5266_ _5468_/A1 _5266_/A2 _5266_/B _5270_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_130_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_867 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7005_ _7005_/D _7281_/RN _7005_/CLK _7005_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4217_ _5535_/B _5528_/A2 _5784_/A3 _5784_/A2 _4219_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_5197_ _4056_/B _4777_/B _5445_/A2 _5445_/A3 _5444_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_56_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4148_ hold58/Z hold220/Z _4150_/S _4148_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4079_ _4078_/S input92/Z _4080_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet783_405 net783_435/I _6813_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet783_416 net783_419/I _6802_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_138_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet783_427 net783_427/I _6791_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet783_449 net833_469/I _6760_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet783_438 _4109__2/I _6771_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_165_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_842 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_1__f_wb_clk_i clkbuf_0_wb_clk_i/Z _7313_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_78_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_431 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1284 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_797 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold719 _7096_/Q hold719/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold708 _6737_/Q hold708/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_7_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3450_ _6863_/Q hold16/Z _3450_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3381_ _4718_/B _5301_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_16
XFILLER_130_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5120_ _5120_/A1 _5287_/C _5120_/A3 _5382_/A2 _5121_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_112_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5051_ _5051_/A1 _5165_/A1 _5051_/B _5051_/C _5052_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_123_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4002_ _4002_/I0 _6705_/Q _4015_/S _6705_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_112_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_464 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5953_ _6107_/B _6107_/C _5974_/B1 _7275_/Q _5954_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_4904_ _5436_/A4 _5194_/B _5194_/C _5235_/A1 _4905_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5884_ hold37/Z _5884_/A2 _5893_/A3 _5535_/B _5892_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_34_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4835_ _5466_/B _5392_/A1 _4718_/B _4661_/C _5502_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_61_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4766_ _5327_/B _4822_/A4 _5152_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_181_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6505_ _6584_/A1 _6505_/A2 _6505_/A3 _6504_/Z _6506_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3717_ hold882/Z _3887_/S _6776_/Q _7338_/Q _3719_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4697_ _4710_/C _4710_/B _4723_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_106_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6436_ _7166_/Q _6279_/Z _6299_/Z _7068_/Q _6437_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xnet733_368 net733_373/I _6886_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet733_379 net833_474/I _6864_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet733_357 net833_473/I _6897_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3648_ input31/Z _5748_/A3 _5532_/A3 _5546_/A2 _3669_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_20_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3579_ _7047_/Q _3950_/B1 _3943_/C1 hold56/I _3580_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6367_ _7155_/Q _6286_/Z _6311_/C _7001_/Q _6312_/Z _7219_/Q _6372_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_5318_ _5200_/B _5318_/A2 _5318_/B _5481_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_96_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold13 hold13/I hold13/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6298_ _6308_/A3 _7278_/Q _7279_/Q _6321_/A4 _6570_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_29_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold46 hold46/I hold46/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold24 hold24/I hold24/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold35 hold35/I hold35/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_5249_ _5249_/A1 _5428_/A1 _5251_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_612 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold57 hold57/I hold57/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold79 hold79/I hold79/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_152_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold68 hold68/I hold68/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_71_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_101_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_356 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_101_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_832 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_6_0__1374_ clkbuf_4_7_0__1374_/I net583_226/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_120_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_642 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1092 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1070 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1081 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4620_ _4620_/A1 _4620_/A2 _4620_/A3 _4627_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_148_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4551_ _3379_/I _3380_/I _4718_/B _4661_/C _5323_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_144_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4482_ _5078_/A2 _5360_/C _4437_/Z _5046_/C _5082_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xhold516 _7197_/Q hold516/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3502_ _3608_/A4 _3477_/Z hold28/Z _5646_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
Xhold505 _5557_/Z _6953_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold527 _7042_/Q hold527/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7270_ _7270_/D _7302_/RN _7304_/CLK _7270_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold538 _6948_/Q hold538/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_144_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3433_ _4119_/B _6774_/Q _6777_/Q _3440_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_6221_ _6901_/Q _6232_/C _6266_/B _6266_/C _6242_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
Xhold549 _7251_/Q hold549/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6152_ _6152_/A1 _6152_/A2 _6152_/A3 _6151_/Z _6164_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5103_ _4690_/C _5290_/C _4963_/B _3379_/I _5105_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_3364_ _7059_/Q _3364_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_97_342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_821 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_832 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_843 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_898 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6083_ _6083_/A1 _6232_/C _6107_/B _6083_/B2 _6083_/C _6084_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
XTAP_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_876 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_865 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5034_ _4487_/Z _5034_/A2 _5290_/C _5290_/B _5385_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XTAP_887 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_898 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6985_ _6985_/D _7302_/RN _6985_/CLK _6985_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_5936_ _7272_/Q _7271_/Q _6235_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5867_ hold518/Z hold391/Z _5874_/S _7226_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5798_ hold164/Z hold283/Z hold9/Z _7166_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4818_ _4661_/C _5153_/B _5266_/A2 _5301_/A2 _5342_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_182_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4749_ _5098_/A2 _5250_/C _5247_/B _3380_/I _4755_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_162_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6419_ _6413_/Z _6417_/Z _6419_/A3 _6426_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_107_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_832 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput103 wb_adr_i[17] _4418_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput114 wb_adr_i[27] _4058_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput136 wb_dat_i[17] _6616_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput125 wb_adr_i[8] _4064_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput147 wb_dat_i[27] _6623_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput158 wb_dat_i[8] _6611_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_57_762 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_153_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_356 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet633_301 net633_301/I _6968_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_94_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3982_ _3982_/A1 _3982_/A2 _3982_/A3 _3982_/A4 _3983_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_90_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_6770_ _6770_/D _7262_/RN _6770_/CLK _6770_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5721_ hold25/Z hold332/Z hold22/Z _5721_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_149_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5652_ hold5/Z hold213/Z _5654_/S _5652_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4603_ _5484_/A2 _5445_/A2 _5439_/C _5180_/B _4606_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_117_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5583_ hold391/Z hold801/Z _5590_/S _5583_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7322_ _7322_/D _7323_/RN _7322_/CLK _7322_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_144_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4534_ _4694_/B _4922_/B _4684_/B _5036_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_129_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold302 _7136_/Q hold302/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_117_723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold324 _7076_/Q hold324/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_117_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold313 _6825_/Q hold313/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold335 _7209_/Q hold335/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4465_ _3380_/I _4425_/Z _4684_/B _4578_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_144_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold368 _5703_/Z _7082_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7253_ _7253_/D _7262_/RN _7253_/CLK _7253_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
Xhold346 _6714_/Q hold346/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold357 _7094_/Q hold357/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7184_ hold79/Z _7265_/RN _7184_/CLK hold78/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold379 _7084_/Q hold379/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_132_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6204_ _7119_/Q _6260_/B1 _6258_/C1 _7193_/Q _6206_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xclkbuf_leaf_7__1374_ clkbuf_4_3_0__1374_/Z net733_381/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4396_ _5535_/B _6653_/A2 _5893_/A3 hold37/Z _4398_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_3416_ input58/Z hold888/Z _3416_/S _7339_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3347_ _7189_/Q _3347_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_98_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6135_ _7116_/Q _6260_/B1 _6256_/B1 _7206_/Q _6136_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_640 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6066_ _7066_/Q _6258_/C1 _6262_/B1 _7026_/Q _6070_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5017_ _3379_/I _3380_/I _4423_/Z _5378_/A1 _5018_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_2518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1839 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1828 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1817 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6968_ _6968_/D _7304_/RN _6968_/CLK _6968_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_53_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6899_ _6899_/D _7341_/RN _6899_/CLK _6899_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5919_ _5918_/B _5931_/A1 _5919_/B _7267_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_22_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_174_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_726 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold880 _6914_/Q hold880/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_3_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold891 hold891/I _7337_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_122_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_66__1374_ _4109__12/I net783_420/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_8_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_512 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4250_ hold630/Z hold388/Z _4262_/S _4250_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4181_ _5784_/A2 _5727_/A3 _5748_/A3 _5535_/B _4189_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_55_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6822_ _6822_/D _7281_/RN _6822_/CLK _6822_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_90_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6753_ _6753_/D _7302_/RN _6753_/CLK _6753_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3965_ _3965_/A1 _3965_/A2 _3965_/A3 _3965_/A4 _3966_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6684_ _7265_/RN _6994_/Q _4026_/C _6684_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_149_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5704_ hold139/Z hold360/Z _5708_/S _5704_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3896_ _6740_/Q _5856_/A2 _5546_/A2 _3527_/Z _3937_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5635_ hold2/Z hold52/Z _5635_/S hold53/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold110 _5817_/Z _7183_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_5566_ hold388/Z hold673/Z hold38/Z _6961_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5497_ _5421_/Z _5496_/Z _5497_/B _5500_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xhold132 _7239_/Q hold132/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7305_ _7305_/D _7323_/RN _7323_/CLK _7305_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold121 _5724_/Z _7101_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_145_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold143 _6998_/Q hold143/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4517_ _4469_/B _4922_/B _5307_/B _4852_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_117_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7236_ _7236_/D _7265_/RN _7236_/CLK _7236_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_171_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold176 _7075_/Q hold176/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold154 _7077_/Q hold154/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4448_ _5166_/A4 _4451_/B _4450_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold165 _5753_/Z _7126_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold187 _5631_/Z _7019_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_144_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold198 _4307_/Z _6828_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7167_ _7167_/D _7265_/RN _7167_/CLK _7167_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_100_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4379_ hold391/Z hold612/Z _4380_/S _4379_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7098_ _7098_/D _7265_/RN _7098_/CLK _7098_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_100_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_431 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6118_ _7052_/Q _6256_/A2 _6259_/B1 _6980_/Q _6125_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_86_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_470 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6049_ _6045_/Z _6049_/A2 _6049_/A3 _6049_/A4 _6049_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_58_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_497 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3750_ _3750_/A1 _3750_/A2 _3750_/A3 _3750_/A4 _3751_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_60_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet583_211 net433_87/I _7058_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet583_222 net433_62/I _7047_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet583_233 net583_233/I _7036_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_185_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet583_244 net783_420/I _7025_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3681_ _3534_/C _5802_/A2 _5573_/A3 _3454_/Z _3681_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_5420_ _5420_/A1 _5459_/A1 _5420_/B _5420_/C _5421_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_161_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5351_ _5351_/A1 _5351_/A2 _5351_/B1 _5463_/B _5351_/C _5421_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
Xoutput226 _7366_/Z mgmt_gpio_out[25] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput215 _4102_/Z mgmt_gpio_out[15] VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_1
XFILLER_57_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput204 _3370_/ZN mgmt_gpio_oeb[5] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput237 _4087_/Z mgmt_gpio_out[35] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_154_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5282_ _5285_/A1 _5476_/A1 _5282_/B _5379_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput259 _6932_/Q pll90_sel[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput248 _4128_/Z pad_flash_clk_oe VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4302_ hold25/Z hold269/Z _4307_/S _4302_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7021_ _7021_/D _7265_/RN _7021_/CLK _7021_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4233_ hold161/Z hold25/Z _4243_/S _4233_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4164_ hold139/Z hold429/Z _4168_/S _4164_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_687 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4095_ _7345_/Q input38/Z _4095_/B _7343_/Q _4096_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_70_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6805_ _6805_/D _7281_/RN _6805_/CLK _6805_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4997_ _5369_/A1 _4947_/C _4963_/B _5007_/A4 _4998_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_6736_ _6736_/D _7341_/RN _6736_/CLK _6736_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_23_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3948_ _6920_/Q _3948_/A2 _3948_/B _3949_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_164_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3879_ input62/Z _3975_/B1 _3879_/B _3879_/C _3883_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_6667_ input75/Z _6994_/Q _4026_/C _6667_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_118_840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5618_ _5646_/A2 _4227_/B _5902_/A3 _5866_/A3 _5626_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_6598_ _6603_/S _7310_/Q _6599_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5549_ hold25/Z _6947_/Q _5551_/S _5549_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_155_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_3_0__f_wb_clk_i clkbuf_0_wb_clk_i/Z _6862_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_105_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7219_ _7219_/D _7262_/RN _7219_/CLK _7219_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_171_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2145 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1466 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet533_163 net533_163/I _7106_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet533_152 net433_65/I _7117_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet533_196 net433_56/I _7073_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet533_185 net683_320/I _7084_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet533_174 net633_280/I _7095_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_123_342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_827 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4920_ _4690_/B _5098_/A2 _4920_/B _5410_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_80_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4851_ _5435_/A1 _5084_/B _5330_/A2 _5290_/C _5389_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3802_ _3454_/Z _3802_/A2 _3534_/C _4246_/A1 _3803_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_4782_ _5327_/B _5307_/B _4794_/A2 _5252_/A4 _5257_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_158_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6521_ _7137_/Q _6287_/Z _6300_/Z _7015_/Q _6319_/Z _7129_/Q _6523_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_3733_ _7141_/Q _3958_/A2 _3968_/A2 _7107_/Q _3737_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_118_147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6452_ _6452_/A1 _6452_/A2 _6452_/A3 _6451_/Z _6453_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3664_ _3664_/A1 _3664_/A2 _3664_/A3 _3665_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_173_253 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5403_ _5481_/A2 _5403_/A2 _5405_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_173_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_832 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6383_ _6383_/A1 _6383_/A2 _6383_/A3 _6383_/A4 _6383_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_3595_ _3595_/A1 _3595_/A2 _3595_/A3 _3594_/Z _3595_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_115_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5334_ _5466_/B _5397_/A1 _5466_/A2 _5334_/B _5335_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_142_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5265_ _5261_/Z _5340_/A2 _5263_/Z _5492_/A4 _5266_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5196_ _5301_/A2 _5290_/C _5200_/B _4661_/C _5204_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_7004_ _7004_/D _7281_/RN _7004_/CLK _7004_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4216_ hold388/Z hold651/Z _4216_/S _4216_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4147_ hold57/Z _7320_/Q _6863_/Q hold58/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_84_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4078_ _6811_/Q input89/Z _4078_/S _4078_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet783_417 net783_417/I _6801_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet783_406 net783_411/I _6812_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_52_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet783_428 net783_431/I _6786_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_11_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet783_439 _4109__2/I _6770_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_177_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6719_ _6719_/D _7304_/RN _6719_/CLK _6719_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_149_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_713 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_898 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_830 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1285 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold709 _6764_/Q hold709/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_7_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3380_ _3380_/I _5315_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_20
XFILLER_171_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5050_ _5351_/A1 _5050_/A2 _5050_/B _5211_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4001_ _4000_/Z _6777_/Q _4001_/B _4002_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_38_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5952_ _6787_/Q _6789_/Q _5952_/B _5954_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4903_ _5194_/C _5417_/A1 _4903_/B _4903_/C _4905_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_18_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5883_ _7241_/Q hold2/Z _5883_/S hold46/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4834_ _5445_/A2 _5177_/A3 _5153_/B _5321_/A3 _5469_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_178_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4765_ _4765_/A1 _4765_/A2 _4765_/B _5327_/B _5468_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_119_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6504_ _6504_/A1 _6504_/A2 _6504_/A3 _6504_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_3716_ _3887_/S _4354_/A1 _3716_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4696_ _5136_/A2 _4759_/B1 _4759_/C _4710_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
Xnet733_369 net433_74/I _6885_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6435_ _7052_/Q _6575_/B1 _6566_/C1 _7020_/Q _6437_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xnet733_358 net833_473/I _6896_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3647_ _7045_/Q _5655_/A4 _5727_/A3 hold29/I _3672_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_161_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3578_ _7071_/Q _3980_/A2 _3950_/A2 _7103_/Q _3580_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6366_ _6366_/A1 _6366_/A2 _6366_/A3 _6372_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_5317_ _5230_/C _5469_/A4 _5317_/A3 _5317_/A4 _5481_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
Xhold14 hold14/I hold14/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6297_ _7279_/Q _6457_/A3 _6562_/A4 _6323_/A1 _6297_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_76_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold47 hold47/I hold47/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold25 hold25/I hold25/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold36 hold36/I hold36/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_130_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5248_ _5329_/A2 _5376_/A1 _5502_/B1 _5394_/C _5248_/C _5428_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_2
Xhold58 hold58/I hold58/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_102_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5179_ _5179_/A1 _5176_/Z _5179_/A3 _5397_/C _5181_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xhold69 hold69/I hold69/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_28_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_324 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_137_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1060 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1071 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1082 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1093 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4550_ _5262_/A4 _3380_/I _4718_/B _4661_/C _5416_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_171_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4481_ _5046_/A1 _5046_/A2 _4628_/B _4481_/C _4682_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_143_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3501_ hold28/I _3608_/A4 _3515_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xhold517 _7254_/Q hold517/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold506 _7365_/I hold506/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold539 _6805_/Q hold539/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6220_ _6559_/S _6220_/A2 _6220_/B _7292_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3432_ _3432_/A1 _3432_/A2 _4072_/A3 _3431_/B _7335_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
Xhold528 _7220_/Q hold528/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3363_ _7067_/Q _3363_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6151_ _6151_/A1 _6151_/A2 _6151_/A3 _6151_/A4 _6151_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XTAP_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5102_ _5454_/A2 _5374_/A2 _5102_/A3 _5279_/A3 _5489_/A1 _5106_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_106_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_833 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_844 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6082_ _7098_/Q _6232_/C _6266_/B _6266_/C _6083_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_855 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_877 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5033_ _5033_/A1 _5033_/A2 _5041_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_111_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_888 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6984_ _6984_/D _7281_/RN _6984_/CLK _6984_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_179_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5935_ _6103_/A1 _7272_/Q _6233_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_15_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5866_ hold37/Z _4227_/B _5866_/A3 hold8/Z _5874_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_22_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_844 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4817_ _5471_/B2 _5468_/C _4825_/A4 _5001_/A1 _5472_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5797_ hold139/Z hold513/Z hold9/Z _7165_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4748_ _4748_/A1 _4748_/A2 _4748_/A3 _4748_/A4 _4755_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_174_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4679_ _4828_/C _4679_/A2 _4681_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6418_ _7205_/Q _6573_/A2 _6288_/Z _7197_/Q _6297_/Z _7043_/Q _6419_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_7282__382 _7282_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_150_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6349_ _6349_/A1 _6349_/A2 _7295_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput115 wb_adr_i[28] _4058_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput104 wb_adr_i[18] _4418_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput126 wb_adr_i[9] _4064_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_163_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput137 wb_dat_i[18] _6620_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput159 wb_dat_i[9] _6615_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput148 wb_dat_i[28] _6627_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_17_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_608 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_26__1374_ clkbuf_4_14_0__1374_/Z _4109__6/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_95_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_106__1374_ clkbuf_4_1_0__1374_/Z net833_470/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_95_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_89__1374_ net583_226/I net433_65/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_35_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3981_ _7242_/Q _3981_/A2 _3981_/B1 _7250_/Q _3981_/C _3982_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_90_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5720_ hold388/Z hold724/Z hold22/Z _7097_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5651_ hold164/Z hold422/Z _5654_/S _5651_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_163_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4602_ _4759_/C _5312_/B _4684_/B _4694_/B _5397_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_5582_ _4227_/B _5646_/A2 _5727_/A3 _5655_/A4 _5590_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_7321_ _7321_/D _7323_/RN _4103_/I1 _7321_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_163_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4533_ _4684_/B _5307_/B _5210_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold325 _5696_/Z _7076_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_156_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold303 _5764_/Z _7136_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7252_ _7252_/D _7302_/RN _7252_/CLK _7252_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold314 _4304_/Z _6825_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4464_ _5223_/A1 _5294_/B _5048_/B _4481_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_131_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6203_ _7177_/Q _6256_/A2 _6261_/B1 _7169_/Q _6206_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold358 _7205_/Q hold358/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold347 _4144_/Z _6714_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold369 _6819_/Q hold369/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold336 _5846_/Z _7209_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7183_ _7183_/D _7265_/RN _7183_/CLK _7183_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_89_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4395_ hold388/Z hold657/Z _4395_/S _4395_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3415_ _6774_/Q _3887_/S _3416_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3346_ _7197_/Q _3346_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_112_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6134_ _7198_/Q _6260_/A2 _6256_/A2 _7174_/Q _6136_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_652 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6065_ _7018_/Q _6233_/A2 _6233_/B1 _7010_/Q _6266_/B _7002_/Q _6071_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XTAP_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_674 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5016_ _5271_/A1 _4963_/B _5288_/A4 _4951_/C _5016_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_86_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1829 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6967_ hold39/Z _7281_/RN _6967_/CLK _6967_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5918_ _4019_/Z _6788_/Q _5918_/B _5918_/C _5919_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_6898_ _6898_/D _7341_/RN _6898_/CLK _6898_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5849_ hold388/Z hold711/Z _5855_/S _5849_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_167_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold870 _7194_/Q hold870/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_89_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold881 _6917_/Q hold881/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_107_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold892 _7346_/Q hold892/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_76_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_186_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_616 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4180_ hold388/Z hold704/Z _4180_/S _4180_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_571 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6821_ _6821_/D _7304_/RN _6821_/CLK _6821_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_51_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3964_ _7226_/Q _3964_/A2 _4264_/A1 input52/Z _3964_/C1 _7258_/Q _3965_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_6752_ _6752_/D _7262_/RN _6752_/CLK _6752_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6683_ _7265_/RN _6994_/Q _4026_/C _6683_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_148_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5703_ hold25/Z hold367/Z _5708_/S _5703_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3895_ _6895_/Q hold37/I _5748_/A3 _5546_/A2 _3981_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_164_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5634_ hold58/Z hold130/Z _5635_/S _5634_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_12_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold100 _7200_/Q hold100/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_5565_ hold391/Z hold754/Z hold38/Z _6960_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_129_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7304_ _7304_/D _7304_/RN _7304_/CLK _7304_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5496_ _5464_/Z _5496_/A2 _5496_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xhold122 _6997_/Q hold122/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold144 _5607_/Z _6998_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold111 _7223_/Q hold111/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_117_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4516_ _4759_/C _5312_/B _4694_/B _5393_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_2
Xhold133 _7177_/Q hold133/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7235_ _7235_/D _7341_/RN _7235_/CLK _7235_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
Xhold155 _5697_/Z _7077_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold177 _5695_/Z _7075_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4447_ _4669_/B _4774_/B _4777_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xhold166 _7142_/Q hold166/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold188 _7347_/Q _3313_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold199 _7233_/Q hold199/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7166_ _7166_/D _7265_/RN _7166_/CLK _7166_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_120_719 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4378_ _4378_/A1 _5856_/A2 _6653_/A2 hold45/Z _4380_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_6117_ _6211_/B _6266_/B _7036_/Q _7274_/Q _6125_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_58_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_7097_ _7097_/D _7265_/RN _7097_/CLK _7097_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XTAP_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3329_ _6788_/Q _6584_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_160_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6048_ _6993_/Q _6258_/B1 _6259_/B1 _6977_/Q _6049_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_58_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_72__1374_ clkbuf_4_5_0__1374_/Z net783_425/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_37_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1604 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_169_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_844 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_185_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet583_212 net433_56/I _7057_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_158_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet583_234 net633_290/I _7035_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet583_223 net433_62/I _7046_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_185_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet583_245 net583_245/I _7024_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3680_ _3679_/Z hold881/Z _3888_/S _6917_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5350_ _5502_/A1 _5463_/A1 _5493_/B2 _5350_/B _5421_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
Xoutput216 _7357_/Z mgmt_gpio_out[16] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput205 _3369_/ZN mgmt_gpio_oeb[6] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput238 _4078_/Z mgmt_gpio_out[36] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5281_ _5281_/A1 _5371_/A1 _5414_/A4 _5283_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xoutput227 _7367_/Z mgmt_gpio_out[26] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4301_ hold388/Z hold630/Z _4307_/S _4301_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput249 _4110_/Z pad_flash_csb VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4232_ hold853/Z _4231_/Z _4244_/S _4232_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7020_ _7020_/D _7265_/RN _7020_/CLK _7020_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_141_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4163_ hold25/Z hold432/Z _4168_/S _4163_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4094_ _4094_/A1 _4094_/A2 _7345_/Q _4095_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_95_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6804_ _6804_/D _7281_/RN _6804_/CLK _6804_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_168_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4996_ _5262_/A4 _4995_/Z input95/Z _5034_/A2 _5109_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_24_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3947_ _3947_/A1 _3947_/A2 _3947_/A3 _3948_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6735_ _6735_/D _7341_/RN _6735_/CLK _6735_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_51_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3878_ _7163_/Q _3878_/A2 _3945_/A2 _7131_/Q _3878_/C _3883_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_6666_ input75/Z _6994_/Q _4026_/C _6666_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_137_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5617_ hold2/Z hold87/Z _5617_/S hold88/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6597_ _6597_/I0 _7309_/Q _6603_/S _7309_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_151_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5548_ _4227_/B hold173/Z _5548_/A3 _5902_/A3 hold174/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_155_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7218_ _7218_/D _7341_/RN _7218_/CLK _7218_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_5479_ _4362_/Z _5479_/A2 _5479_/A3 _5479_/A4 _5479_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_78_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7149_ _7149_/D _7341_/RN _7149_/CLK _7149_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_120_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_875 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet533_164 net833_498/I _7105_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet533_153 _4109__9/I _7116_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet533_197 net433_90/I _7072_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_151_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet533_186 net683_320/I _7083_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_123_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet533_175 net633_292/I _7094_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_145_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4850_ _4425_/Z _5210_/C _5210_/B _5315_/A4 _5165_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XTAP_2691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3801_ _3827_/A2 _3496_/B _3831_/A2 _4246_/A2 _3968_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XTAP_1990 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6520_ _7193_/Q _6274_/Z _6284_/Z _7103_/Q _6523_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4781_ _3379_/I _5489_/A2 _5315_/A4 _4423_/Z _4784_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3732_ _7229_/Q _3964_/A2 _3732_/B _3732_/C _3752_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_119_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6451_ _6584_/A1 _6451_/A2 _6451_/A3 _6451_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_3663_ _7143_/Q _3958_/A2 _3959_/A2 _6731_/Q _3643_/Z _6932_/Q _3664_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_174_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5402_ _5402_/A1 _5402_/A2 _5316_/Z _5400_/Z _5403_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6382_ _7164_/Q _6279_/Z _6299_/Z _7066_/Q _6383_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3594_ _3594_/A1 _3594_/A2 _3594_/A3 _3594_/A4 _3594_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_114_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5333_ _5333_/A1 _5333_/A2 _5333_/A3 _5333_/A4 _5490_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_5264_ _5471_/B2 _4487_/Z _5445_/A2 _5264_/A4 _5340_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_130_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5195_ _5190_/Z _5435_/B _5318_/B _5480_/A2 _5204_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_7003_ _7003_/D _7302_/RN _7003_/CLK _7003_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_68_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4215_ hold391/Z hold769/Z _4216_/S _4215_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4146_ hold5/Z hold265/Z _4150_/S _4146_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4077_ _6812_/Q input91/Z _4078_/S _4077_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_37_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_853 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet783_407 net783_408/I _6811_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4979_ _4979_/A1 _4979_/A2 _4979_/A3 _4982_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xnet783_418 net783_419/I _6800_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet783_429 net783_430/I _6785_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_11_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6718_ _6718_/D _7304_/RN _6718_/CLK _6718_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_6649_ _6649_/A1 _6649_/A2 _6649_/A3 _6652_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_20_794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_842 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1253 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4000_ _6705_/Q _4000_/A2 _4000_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_111_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5951_ _6107_/B _6107_/C _7275_/Q _6789_/Q _5952_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_65_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4902_ _5330_/A2 _4694_/B _5294_/B _4922_/B _5417_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_80_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_853 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5882_ hold74/Z hold58/Z _5883_/S _7240_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_61_650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4833_ _3380_/I _5445_/A2 _5177_/A3 _5262_/A4 _5330_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_21_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4764_ _3379_/I _5253_/A2 _5315_/A4 _4423_/Z _4770_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_159_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6503_ hold80/I _6581_/B1 _6312_/Z _7224_/Q _6504_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3715_ _3715_/A1 _3715_/A2 _3715_/A3 _3715_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_4695_ _5136_/A2 _4690_/C _5484_/A2 _4759_/A2 _4694_/B _4767_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_4
X_6434_ _7134_/Q _6287_/Z _6300_/Z _7012_/Q _6319_/Z _7126_/Q _6437_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_162_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet733_359 net833_473/I _6895_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3646_ input8/Z _5700_/A1 _5748_/A3 _5532_/A3 _3664_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_20_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3577_ _5534_/A1 _3827_/A2 _3496_/B _3831_/A2 _3953_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_6365_ _6365_/A1 _6365_/A2 _6365_/A3 _6365_/A4 _6366_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_142_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5316_ _5230_/C _5469_/A4 _5317_/A3 _5317_/A4 _5316_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_114_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6296_ _7280_/Q _6296_/A2 _7281_/Q _6324_/A1 _6578_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_88_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5247_ _5416_/A1 _5271_/A4 _5247_/B _5250_/C _5248_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_2
Xhold15 hold15/I hold15/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold37 hold37/I hold37/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold26 hold26/I hold26/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_57_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold59 hold59/I hold59/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold48 hold48/I hold48/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_5178_ _5502_/A1 _5180_/B _5502_/B1 _5502_/A2 _5397_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_69_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4129_ _4131_/A1 _6878_/Q _6875_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_28_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_358 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_101_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_185_839 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_71 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_466 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1061 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1050 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1083 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_49__1374_ clkbuf_4_15_0__1374_/Z net633_271/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1094 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_872 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3500_ _6863_/Q _3500_/A2 hold35/Z _3500_/C _3608_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_30_399 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4480_ _5315_/A4 _4951_/B1 _4480_/B _4502_/B _4628_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_144_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold518 _7226_/Q hold518/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold507 _5556_/Z _6952_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3431_ _4072_/A3 _6774_/Q _3431_/B _3432_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold529 _5859_/Z _7220_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3362_ _7075_/Q _3362_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_124_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6150_ _7175_/Q _6256_/A2 _6261_/A2 hold91/I _6151_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_801 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5101_ _4963_/B _4955_/B _4951_/C _5111_/A2 _5102_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_151_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_823 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_878 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6081_ _6211_/C _7273_/Q _7124_/Q _7275_/Q _6083_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_845 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_867 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_856 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5032_ _5262_/A4 _5287_/B1 _3380_/I _5235_/A1 _5033_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_111_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_399 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_878 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6983_ _6983_/D _7281_/RN _6983_/CLK _6983_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_19_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5934_ _6036_/A3 _7271_/Q _6233_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_40_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5865_ hold343/Z hold2/Z _5865_/S _5865_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4816_ _5369_/A1 _5426_/B1 _5001_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5796_ hold25/Z hold458/Z hold9/Z _7164_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4747_ _4706_/Z _4709_/Z _4825_/A4 _5093_/B _4748_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4678_ _5459_/A3 _4682_/A2 _5355_/A2 _5051_/B _4679_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3629_ hold83/I _3940_/A2 _3950_/A2 hold64/I _3875_/A2 hold78/I _3630_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6417_ _6417_/A1 _6417_/A2 _6417_/A3 _6417_/A4 _6417_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_162_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6348_ _6968_/Q _6584_/A1 _6348_/B _6509_/B _6349_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_163_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput105 wb_adr_i[19] _4418_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput116 wb_adr_i[29] _4057_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput127 wb_cyc_i _4062_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_130_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6279_ _7276_/Q _6561_/A3 _6406_/A4 _6310_/A4 _6279_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_88_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput149 wb_dat_i[29] _6631_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput138 wb_dat_i[19] _6624_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_102_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_188_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3980_ _7064_/Q _3980_/A2 _3980_/B1 _6976_/Q _3980_/C _3982_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XPHY_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5650_ hold139/Z hold247/Z _5654_/S _5650_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4601_ _4469_/B _4686_/B _5307_/B _4922_/B _5180_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_157_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5581_ hold2/Z hold98/Z _5581_/S hold99/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7320_ _7320_/D _7323_/RN _4103_/I1 _7320_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4532_ _4694_/B _4922_/B _5210_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_7_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4463_ _4437_/Z _5436_/A1 _4463_/B _5046_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xhold304 _7192_/Q hold304/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold315 _7124_/Q hold315/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold326 _6744_/Q hold326/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7251_ _7251_/D _7341_/RN _7251_/CLK _7251_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_172_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold348 _7371_/I hold348/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6202_ _6198_/Z _6202_/A2 _6202_/A3 _6202_/A4 _6202_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
Xhold359 _5842_/Z _7205_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3414_ _6709_/Q _6708_/Q _6707_/Q _3887_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
Xhold337 _7161_/Q hold337/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7182_ _7182_/D _7265_/RN _7182_/CLK _7182_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4394_ hold391/Z hold581/Z _4395_/S _4394_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3345_ _7205_/Q _3345_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_86_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6133_ _7134_/Q _6257_/A2 _6258_/B1 _6746_/Q _6257_/B1 _7182_/Q _6136_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XTAP_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_642 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6064_ _6064_/A1 _6064_/A2 _6232_/C _6064_/A4 _6071_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_58_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_675 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5015_ _5015_/A1 _5015_/A2 _5015_/A3 _5018_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_86_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6966_ hold59/Z _7281_/RN _6966_/CLK _6966_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_1819 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5917_ _6790_/Q _6788_/Q _6789_/Q _5917_/B _5927_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_6897_ _6897_/D _7341_/RN _6897_/CLK _6897_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_42_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5848_ hold391/Z hold811/Z _5855_/S _5848_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_32__1374_ clkbuf_4_10_0__1374_/Z net433_56/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5779_ hold139/Z hold449/Z hold14/Z _7149_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_158_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_95__1374_ clkbuf_4_3_0__1374_/Z _4109__2/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_108_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold860 _7131_/Q hold860/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold871 _6799_/Q hold871/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_123_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold882 _6915_/Q hold882/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_115_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold893 _6778_/Q hold893/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_853 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6820_ _6820_/D input75/Z _6820_/CLK _6820_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_91_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6751_ _6751_/D _7262_/RN _6751_/CLK _6751_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3963_ _3963_/A1 _3963_/A2 _3963_/A3 _3966_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_50_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6682_ _7265_/RN _6994_/Q _4026_/C _6682_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_149_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5702_ hold388/Z hold661/Z _5708_/S _5702_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3894_ _6768_/Q _5784_/A2 _5784_/A3 _5528_/A2 _3965_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5633_ hold5/Z hold115/Z _5635_/S _5633_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5564_ hold37/Z _5640_/A2 _5564_/A3 _4227_/B hold38/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
Xhold101 _7191_/Q hold101/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_144_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4515_ _4690_/C _4487_/Z _5466_/B _5466_/C _4564_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_7303_ _7303_/D _7304_/RN _7304_/CLK _7303_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5495_ _5495_/A1 _5495_/A2 _5496_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xhold123 _5606_/Z _6997_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_144_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold112 _5863_/Z _7223_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold134 _5810_/Z _7177_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7234_ _7234_/D _7341_/RN _7234_/CLK _7234_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
Xhold156 _7215_/Q hold156/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_160_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4446_ _4669_/B _4774_/B _4959_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_104_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold145 _7015_/Q hold145/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold167 _5771_/Z _7142_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold178 _7067_/Q hold178/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_160_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7165_ _7165_/D _7341_/RN _7165_/CLK _7165_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold189 _3498_/C _3534_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_144_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4377_ hold388/Z hold577/Z _4377_/S _4377_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3328_ _7269_/Q _5925_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6116_ _6116_/I0 _7288_/Q _6559_/S _7288_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7096_ _7096_/D _7341_/RN _7096_/CLK _7096_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_112_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6047_ _7089_/Q _6262_/A2 _6261_/A2 _7001_/Q _6049_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_27_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1616 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6949_ _6949_/D _7281_/RN _6949_/CLK _6949_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_81_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_831 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold690 _6934_/Q hold690/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_78_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_877 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet583_213 net433_88/I _7056_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet583_202 net583_214/I _7067_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_13_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet583_224 net433_62/I _7045_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_185_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet583_246 net583_250/I _7023_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet583_235 _4109__44/I _7034_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput217 _7358_/Z mgmt_gpio_out[17] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_160_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput206 _5641_/A2 mgmt_gpio_oeb[7] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput239 _4077_/Z mgmt_gpio_out[37] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5280_ _5370_/A1 _5498_/A2 _5414_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_153_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput228 _7368_/Z mgmt_gpio_out[27] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4300_ hold391/Z hold700/Z _4307_/S _4300_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4231_ hold587/Z hold388/Z _4243_/S _4231_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4162_ hold388/Z hold757/Z _4168_/S _4162_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4093_ _6919_/Q _6994_/Q _4026_/C _4094_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_83_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4995_ _4963_/B _4922_/B _4947_/C _4995_/A4 _4995_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
X_6803_ _6803_/D _7281_/RN _6803_/CLK _7356_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_90_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3946_ _7016_/Q _3946_/A2 _3946_/B1 _6881_/Q _3947_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6734_ _6734_/D _7341_/RN _6734_/CLK _6734_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_176_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3877_ _3877_/A1 _3877_/A2 _3877_/A3 _3877_/A4 _3884_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6665_ _7262_/RN _6994_/Q _4026_/C _6665_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_149_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5616_ hold58/Z hold200/Z _5617_/S _5616_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6596_ _3790_/Z _7308_/Q _6603_/S _7308_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_129_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5547_ hold391/Z hold725/Z _5547_/S _5547_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5478_ hold27/I _4365_/C _5488_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7217_ hold33/Z _7265_/RN _7217_/CLK hold32/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4429_ _4759_/C _5136_/A2 _5098_/A2 _4957_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_120_506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7148_ _7148_/D _7265_/RN _7148_/CLK _7148_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_101_731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7079_ hold55/Z _7265_/RN _7079_/CLK hold54/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_100_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1435 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_898 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet533_154 net633_301/I _7115_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet533_187 net633_271/I _7082_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_124_867 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet533_165 net683_331/I _7104_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet533_176 net533_176/I _7093_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet533_198 net583_214/I _7071_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_124_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_464 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3800_ _3802_/A2 _3534_/C _3460_/B _4246_/A1 _3973_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_4780_ _5093_/B _5489_/A2 _4780_/B _4784_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_33_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1991 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1980 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3731_ _3731_/I _3732_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_158_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6450_ _7254_/Q _6580_/B1 _6309_/Z _7238_/Q _7158_/Q _6286_/Z _6451_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_3662_ _6973_/Q _3559_/Z _3969_/B1 _6747_/Q _3664_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_173_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3593_ input70/Z _4262_/S _3981_/A2 hold49/I _3594_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5401_ _5401_/A1 _5401_/A2 _5401_/A3 _5401_/A4 _5487_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6381_ _7050_/Q _6575_/B1 _6566_/C1 _7018_/Q _6383_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_62_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5332_ _5332_/A1 _5332_/A2 _5333_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5263_ _5263_/A1 _5263_/A2 _5263_/A3 _5263_/A4 _5263_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_5194_ _5439_/A1 _5226_/A1 _5194_/B _5194_/C _5480_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_7002_ _7002_/D _7302_/RN _7002_/CLK _7002_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4214_ _5535_/B _5518_/A1 _3527_/Z _5748_/A3 _4216_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_4145_ hold4/Z _7319_/Q _6863_/Q hold5/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_96_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4076_ _4076_/A1 _4076_/A2 _6876_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet783_408 net783_408/I _6810_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4978_ _4963_/B _4661_/C _4718_/B _5235_/A2 _5209_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xnet783_419 net783_419/I _6799_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_165_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6717_ _6717_/D _7304_/RN _6717_/CLK _6717_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_3929_ _6762_/Q _5748_/A3 _5546_/A2 _3527_/Z _3957_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6648_ _6880_/Q _6648_/A2 _6648_/A3 _6649_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_164_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6579_ _7121_/Q _6579_/A2 _6309_/Z _6737_/Q _6582_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_145_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1287 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5950_ _6211_/C _6211_/B _6107_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_1_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4901_ _5349_/A1 _5084_/B _5200_/B _5435_/A2 _5435_/A1 _4903_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_18_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5881_ hold132/Z hold5/Z _5883_/S _7239_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4832_ _5301_/A2 _5466_/B _5392_/A1 _4661_/C _5148_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xclkbuf_4_11_0__1374_ clkbuf_3_5_0__1374_/Z clkbuf_4_11_0__1374_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_147_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4763_ _5253_/A1 _5253_/A2 _4763_/B _4770_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_174_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4694_ _4689_/Z _4487_/Z _4694_/B _4787_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_6502_ hold96/I _6286_/Z _6311_/C _7006_/Q _6504_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3714_ _3714_/A1 _3711_/Z _3714_/A3 _3714_/A4 _3715_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_119_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6433_ _6433_/I _6441_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_174_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3645_ input57/Z hold21/I hold37/I _5902_/A3 _3654_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_106_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3576_ hold87/I _3961_/A2 _3961_/B1 _7031_/Q hold32/I _3940_/A2 _3582_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6364_ _7203_/Q _6573_/A2 _6288_/Z _7195_/Q _6297_/Z _7041_/Q _6365_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_130_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6295_ _6325_/A2 _7278_/Q _7279_/Q _6321_/A4 _6579_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_5315_ _5394_/A2 _5445_/A3 _5390_/A1 _5315_/A4 _5317_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
Xclkbuf_0__1374_ _4108_/ZN clkbuf_0__1374_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5246_ _5429_/A1 _5328_/A2 _5467_/A2 _5249_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
Xhold38 hold38/I hold38/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold16 hold16/I hold16/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold27 hold27/I hold27/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_102_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold49 hold49/I hold49/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_5177_ _5177_/A1 _5312_/C _5177_/A3 _5307_/B _5179_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_68_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4128_ _7343_/Q input75/Z _4128_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_4059_ input97/Z input96/Z input99/Z input98/Z _4065_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_28_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_832 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_101_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_868 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_180_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1040 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1062 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1051 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1073 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1095 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1084 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold508 _7027_/Q _3368_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_7_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold519 _7227_/Q hold519/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_109_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3430_ _3421_/B input58/Z _3432_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_171_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3361_ _7083_/Q _3361_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5100_ _5489_/A1 _5107_/A1 _5374_/A2 _4437_/Z _5412_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6080_ _7272_/Q _6080_/A2 _7271_/Q _6232_/C _6129_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XTAP_802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_835 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5031_ _4425_/Z _5026_/B _5026_/C _5315_/A4 _5433_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_111_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_868 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_857 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_879 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6982_ _6982_/D _7302_/RN _6982_/CLK _6982_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_80_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5933_ _6789_/Q _5974_/B1 _7271_/Q _7271_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_15_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_640 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5864_ hold320/Z hold58/Z _5865_/S _5864_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4815_ _5471_/A1 _4823_/A2 _5266_/A2 _5439_/A2 _5472_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_178_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5795_ hold388/Z hold611/Z hold9/Z _7163_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_175_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4746_ _5315_/A4 _5301_/A2 _5235_/A1 _3379_/I _5271_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_175_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_512 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4677_ _5210_/C _5210_/B _5468_/A1 _5194_/C _4828_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_119_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3628_ _7224_/Q _3975_/A2 _3938_/A2 _7208_/Q _7168_/Q _3878_/A2 _3630_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6416_ _7157_/Q _6286_/Z _6528_/A2 _7027_/Q _6417_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_134_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6347_ _6347_/A1 _6584_/A1 _6334_/Z _6347_/A4 _6348_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_89_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3559_ _3534_/C _5784_/A3 _5573_/A3 _3454_/Z _3559_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
Xinput117 wb_adr_i[2] _4661_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
Xinput106 wb_adr_i[1] _5004_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
X_6278_ _6324_/A1 _7278_/Q _6406_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xinput128 wb_dat_i[0] _6612_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput139 wb_dat_i[1] _6616_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_5229_ _5229_/A1 _5229_/A2 _5229_/A3 _5461_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_88_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_55__1374_ clkbuf_4_13_0__1374_/Z net783_426/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_84_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_145 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_512 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4600_ _4600_/A1 _5067_/C _4600_/A3 _4606_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_148_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5580_ hold58/Z hold217/Z _5581_/S _6974_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4531_ _5360_/C _5312_/B _4686_/B _4437_/Z _5347_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_157_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold316 _7100_/Q hold316/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_144_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold305 _5827_/Z _7192_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4462_ _5312_/B _4684_/B _5294_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_7250_ _7250_/D _7341_/RN _7250_/CLK _7250_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
Xhold338 _7074_/Q hold338/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold349 _5562_/Z _6958_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6201_ hold54/I _6260_/A2 _6260_/B1 _6991_/Q _6202_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold327 _7172_/Q hold327/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3413_ _6709_/Q _6708_/Q _3417_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7181_ _7181_/D _7341_/RN _7181_/CLK _7181_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4393_ hold45/Z _4405_/A2 _4405_/A3 _5838_/A2 _4395_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_3344_ _7213_/Q _3344_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_98_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6132_ _6132_/A1 _6132_/A2 _6137_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6063_ _6994_/Q _7272_/Q _7271_/Q _6266_/C _6064_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_654 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5014_ _5353_/A3 _4963_/B _5288_/A4 _4951_/C _5015_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_85_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_687 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6965_ _6965_/D _7281_/RN _6965_/CLK _6965_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5916_ _4019_/Z _6788_/Q _5918_/C _5920_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6896_ _6896_/D _7341_/RN _6896_/CLK _6896_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_167_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5847_ _4227_/B _3527_/Z hold13/Z _5866_/A3 _5855_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
Xclkbuf_3_6_0__1374_ clkbuf_0__1374_/Z clkbuf_3_6_0__1374_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_22_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5778_ hold25/Z hold452/Z hold14/Z _7148_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_158_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4729_ _5267_/C _5327_/B _4729_/A3 _4729_/B _4737_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_181_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold850 _5812_/Z _7178_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold872 _4268_/Z _6799_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_122_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold861 _6792_/Q hold861/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_1_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold894 _7327_/Q hold894/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold883 _6775_/Q _3322_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_130_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6750_ _6750_/D _7262_/RN _6750_/CLK _6750_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_188_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5701_ hold391/Z hold794/Z _5708_/S _5701_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3962_ _7008_/Q _3962_/A2 _3962_/B1 _7080_/Q _3967_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_92_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6681_ input75/Z _6994_/Q _4026_/C _6681_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_3893_ _3892_/Z _6653_/A2 _5532_/A3 _5838_/A2 _3938_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_5632_ hold164/Z hold309/Z _5635_/S _5632_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5563_ hold2/Z hold243/Z _5563_/S _5563_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_129_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4514_ _4469_/B _4686_/B _5307_/B _4922_/B _5466_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_145_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7302_ _7302_/D _7302_/RN _7302_/CLK _7302_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5494_ _5494_/A1 _5219_/Z _5494_/A3 _5495_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_172_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold135 _7061_/Q hold135/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold113 _7151_/Q hold113/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold102 _5826_/Z _7191_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_117_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold124 _6991_/Q hold124/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_105_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold157 _5853_/Z _7215_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4445_ _5166_/A4 _4451_/B _4777_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_132_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7233_ _7233_/D _7341_/RN _7233_/CLK _7233_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_105_729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold146 _5626_/Z _7015_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold168 _7174_/Q hold168/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7164_ _7164_/D _7265_/RN _7164_/CLK _7164_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_104_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4376_ hold391/Z hold590/Z _4377_/S _4376_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold179 _6725_/Q hold179/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_112_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3327_ _7268_/Q _5985_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
X_6115_ _6788_/Q _6115_/A2 _6115_/A3 _6115_/B _6116_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_7095_ _7095_/D _7281_/RN _7095_/CLK _7095_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_59_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_462 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6046_ _7065_/Q _6258_/C1 _6257_/B1 _7057_/Q _6985_/Q _6260_/B1 _6049_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XTAP_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1606 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1639 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6948_ _6948_/D _7281_/RN _6948_/CLK _6948_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6879_ _6879_/D _7323_/RN _7323_/CLK _6879_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_155_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold680 _7121_/Q hold680/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_762 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold691 _6769_/Q hold691/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_103_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet583_203 net433_89/I _7066_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet583_214 net583_214/I _7055_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_41_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet583_225 _4109__49/I _7044_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet583_247 net583_250/I _7022_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet583_236 net433_66/I _7033_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_185_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_640 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput207 _3367_/ZN mgmt_gpio_oeb[8] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput218 _7359_/Z mgmt_gpio_out[18] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput229 _7369_/Z mgmt_gpio_out[28] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_99_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4230_ hold864/Z _4229_/Z _4244_/S _4230_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_142_868 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4161_ hold391/Z hold838/Z _4168_/S _4161_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_122_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4092_ _5564_/A3 _6792_/Q _4094_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6802_ _6802_/D _7281_/RN _6802_/CLK _7355_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_36_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4994_ _4963_/B _4922_/B _4947_/C _4995_/A4 _5279_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_17_790 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3945_ _7130_/Q _3945_/A2 _3945_/B1 _6756_/Q _3945_/C _3949_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_6733_ _6733_/D _7262_/RN _6733_/CLK _6733_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_23_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6664_ input75/Z _6994_/Q _4026_/C _6664_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_32_782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5615_ hold5/Z hold202/Z _5617_/S _5615_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3876_ _7187_/Q _3953_/B1 _3942_/B1 _7341_/Q _3877_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6595_ _6595_/I0 _7307_/Q _6603_/S _7307_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5546_ hold45/Z _5546_/A2 _5856_/A2 hold37/Z _5547_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_160_610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5477_ _5477_/A1 _5500_/A2 _5477_/B _5477_/C _5488_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_2_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7216_ hold84/Z _7265_/RN _7216_/CLK hold83/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4428_ _4421_/Z _4425_/Z _4951_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_132_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_2_3__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/Z _4089_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4359_ _6878_/Q _6879_/Q _6880_/Q _6640_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_7147_ _7147_/D _7341_/RN _7147_/CLK _7147_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_113_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7078_ hold90/Z _7265_/RN _7078_/CLK hold89/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_74_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6029_ _6211_/B _6028_/Z _6233_/B1 _7274_/Q _6031_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_46_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1403 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_833 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet533_155 _4109__9/I _7114_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet533_166 net433_68/I _7103_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet533_188 net783_417/I _7081_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_135_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet533_177 net433_76/I _7092_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet533_199 _4109__29/I _7070_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_151_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_9_0__1374_ clkbuf_4_9_0__1374_/I _4109__51/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_65_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_830 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1970 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1981 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3730_ _7011_/Q _3962_/A2 _3961_/A2 _7003_/Q _4262_/S input67/Z _3731_/I VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_159_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3661_ _3661_/A1 _3661_/A2 _3661_/A3 _3665_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3592_ _7233_/Q _3964_/A2 _4264_/A1 input60/Z _3594_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5400_ _5401_/A1 _5401_/A2 _5401_/A3 _5401_/A4 _5400_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_6380_ _7132_/Q _6287_/Z _6300_/Z _7010_/Q _6319_/Z _7124_/Q _6383_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_173_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5331_ _5429_/A1 _5328_/Z _5429_/A2 _5336_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_55_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5262_ _3380_/I _4423_/Z _5337_/A2 _5262_/A4 _5263_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_7001_ _7001_/D _7302_/RN _7001_/CLK _7001_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_141_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5193_ _5439_/A2 _5476_/A1 _5194_/C _5194_/B _5318_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_114_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4213_ hold639/Z hold388/Z _4213_/S _4213_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4144_ hold164/Z hold346/Z _4150_/S _4144_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4075_ _6870_/Q _4075_/A2 _4065_/Z _4076_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_37_830 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4977_ _5004_/A1 input95/Z _5153_/A2 _5374_/A2 _4979_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xnet783_409 net783_411/I _6809_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6716_ _6716_/D _7304_/RN _6716_/CLK _6716_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_3928_ _6829_/Q _5856_/A2 _5528_/A2 _5573_/A3 _3965_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6647_ _6879_/Q _6648_/A3 _6647_/A3 _6649_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_165_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3859_ _7227_/Q _3964_/A2 _3962_/B1 _7081_/Q _3981_/A2 _7243_/Q _3861_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_165_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6578_ _6898_/Q _6578_/A2 _6310_/Z _6832_/Q _6578_/C1 _6773_/Q _6583_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_118_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5529_ hold391/Z hold786/Z _5529_/S _5529_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_145_481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_844 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5880_ hold431/Z hold164/Z _5883_/S _7238_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4900_ _5436_/A4 _5321_/A3 _5194_/C _5235_/A1 _5480_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_2490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4831_ _5436_/A1 _5439_/A1 _5210_/C _5194_/C _4905_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_61_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4762_ _4762_/A1 _4762_/A2 _4762_/A3 _5332_/A1 _4763_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4693_ _4794_/A2 _4765_/B _4693_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_3713_ _7150_/Q _3866_/A2 _3946_/A2 _7020_/Q _3940_/A2 _7214_/Q _3714_/A4 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_6501_ _7256_/Q _6580_/B1 _6309_/Z hold74/I hold72/I _6579_/A2 _6504_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_186_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3644_ _3454_/Z _3644_/A2 _5534_/A2 _3534_/C _3975_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_6432_ _7108_/Q _6285_/Z _6564_/C1 _7084_/Q _6433_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_161_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3575_ _7015_/Q _3962_/A2 _4281_/S input42/Z _3981_/B1 _7257_/Q _3582_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6363_ _7147_/Q _6575_/A2 _6566_/C1 _7017_/Q _6365_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5314_ _5310_/Z _5314_/A2 _5483_/B _5319_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6294_ _7279_/Q _6563_/A3 _6562_/A4 _6323_/A1 _6294_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_170_782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5245_ _5245_/A1 _5369_/A2 _5245_/B1 _5327_/B _5245_/C _5467_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_88_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold28 hold28/I hold28/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold17 hold17/I hold17/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold39 hold39/I hold39/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_5176_ _5176_/A1 _5388_/A1 _5308_/A4 _5176_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_29_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4127_ _7344_/Q input75/Z _4127_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_4058_ _4058_/A1 _4058_/A2 _4058_/A3 _4062_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_45_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_78__1374_ clkbuf_4_5_0__1374_/Z net633_301/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_152_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_188_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1030 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1041 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1052 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1096 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1085 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_830 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold509 hold509/I _7027_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_143_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3360_ _7091_/Q _3360_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_112_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_825 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5030_ _5024_/Z _5030_/A2 _5120_/A3 _5033_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_97_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_836 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_847 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6981_ _6981_/D _7302_/RN _6981_/CLK _6981_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5932_ _6787_/Q _6789_/Q _5974_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_93_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet833_490 net833_491/I _6719_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_19_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5863_ hold111/Z hold5/Z _5865_/S _5863_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_178_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5794_ hold391/Z hold545/Z hold9/Z _7162_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4814_ _3380_/I _4423_/Z _5266_/A2 _5262_/A4 _5431_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_178_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4745_ _5262_/A4 _3380_/I _4718_/B _4661_/C _5093_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_21_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4676_ _4443_/Z _5051_/C _5290_/C _5466_/A2 _5343_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_3627_ _3627_/A1 _3627_/A2 _3627_/A3 _3627_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_6415_ _7165_/Q _6279_/Z _6310_/Z _6979_/Q _6417_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3558_ hold172/Z _3608_/A4 _3482_/Z _3827_/A2 hold173/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_6346_ _7048_/Q _6575_/B1 _6312_/Z _7218_/Q _6346_/C _6347_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_89_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput107 wb_adr_i[20] _4774_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xinput118 wb_adr_i[30] _4063_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3489_ _4073_/B1 _6706_/Q _3489_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_130_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6277_ _6312_/A4 _5975_/B _6308_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_102_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput129 wb_dat_i[10] _6619_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_5228_ _4437_/Z _5360_/C _5360_/B _4956_/C _5229_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5159_ _5285_/A1 _5199_/B _5202_/B _5344_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_84_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_2__1374_ clkbuf_4_2_0__1374_/Z net783_431/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_72_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_122_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4530_ _4628_/B _5307_/B _5078_/A2 _5086_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_117_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_844 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold317 _5723_/Z _7100_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold306 _7150_/Q hold306/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_156_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4461_ _4686_/B _5307_/B _5436_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_7_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold339 _5694_/Z _7074_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7180_ _7180_/D _7265_/RN _7180_/CLK _7180_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_171_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6200_ _7087_/Q _6256_/B1 _6257_/B1 hold56/I _6202_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold328 _5805_/Z _7172_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3412_ _4073_/B2 _3412_/A2 _3412_/A3 hold898/Z _3412_/B2 hold899/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_4392_ hold388/Z hold491/Z _4392_/S _4392_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_98_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6131_ _7190_/Q _6258_/C1 _6259_/B1 _7108_/Q _6132_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3343_ _7221_/Q _5861_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6062_ _7074_/Q _6260_/A2 _6256_/B1 _7082_/Q _6064_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_58_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_644 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_677 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5013_ _5369_/A1 _4963_/B _5288_/A4 _4951_/C _5015_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_100_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_894 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6964_ _6964_/D _7281_/RN _6964_/CLK _6964_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_81_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6895_ _6895_/D _7341_/RN _6895_/CLK _6895_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_34_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5915_ _6790_/Q _6788_/Q _6789_/Q _5918_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_34_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5846_ hold2/Z hold335/Z _5846_/S _5846_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5777_ hold388/Z hold796/Z hold14/Z _7147_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4728_ _4690_/C _5392_/A1 _4819_/A4 _4808_/A2 _5127_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_162_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4659_ _5315_/A4 _5235_/A1 _4718_/B _3379_/I _5468_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_162_332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold873 _7218_/Q hold873/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold862 _4251_/Z _6792_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold840 _6922_/Q hold840/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold851 _6772_/Q hold851/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_115_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6329_ _7258_/Q _6581_/B1 _6580_/B1 _7250_/Q _7096_/Q _6284_/Z _6334_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
Xhold884 hold884/I _6775_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold895 _7335_/Q _3316_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_103_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_71 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_533 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3961_ _7000_/Q _3961_/A2 _3961_/B1 _7024_/Q _3967_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_90_374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5700_ _5700_/A1 _5902_/A3 _5718_/A3 _4227_/B _5708_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_16_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6680_ input75/Z _6994_/Q _4026_/C _6680_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_3892_ _7344_/Q _7327_/Q _6937_/Q _3892_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_31_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5631_ hold139/Z hold186/Z _5635_/S _5631_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_85_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5562_ hold58/Z hold348/Z _5563_/S _5562_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4513_ _4759_/C _5312_/B _4684_/B _4694_/B _5484_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_157_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7301_ _7301_/D _7302_/RN _7304_/CLK _7301_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5493_ _5502_/A1 _5502_/A2 _5493_/B1 _5493_/B2 _5494_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold114 _7053_/Q hold114/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold103 _7263_/Q hold103/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7232_ _7232_/D _7265_/RN _7232_/CLK _7232_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold125 _5599_/Z _6991_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold147 _6816_/Q hold147/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold136 _6965_/Q hold136/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4444_ _5225_/A1 _5225_/A3 _5051_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_145_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold158 _6717_/Q hold158/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7163_ _7163_/D _7341_/RN _7163_/CLK _7163_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4375_ hold45/Z _4405_/A2 _5856_/A2 _4378_/A1 _4377_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
Xhold169 _5807_/Z _7174_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_113_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6114_ _6788_/Q _7287_/Q _6115_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3326_ _7267_/Q _5918_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_7094_ _7094_/D _7302_/RN _7094_/CLK _7094_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_86_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6045_ _6045_/A1 _6045_/A2 _6045_/A3 _6045_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_58_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_474 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2319 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6947_ _6947_/D _7281_/RN _6947_/CLK _6947_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_81_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6878_ _6878_/D _7323_/RN _7323_/CLK _6878_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_139_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5829_ _4227_/B _3527_/Z _5902_/A3 _5884_/A2 hold18/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_22_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold670 _5638_/Z _7025_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_1_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold681 _5747_/Z _7121_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_89_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold692 _6753_/Q hold692/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_77_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_842 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_186_711 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet583_215 _4109__29/I _7054_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet583_204 net433_71/I _7065_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_9_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet583_248 net433_68/I _7021_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_158_468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet583_237 _4109__49/I _7032_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_13_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet583_226 net583_226/I _7043_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_173_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput208 _3366_/ZN mgmt_gpio_oeb[9] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput219 _7360_/Z mgmt_gpio_out[19] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_175_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4160_ _5838_/A4 _5518_/A1 _5532_/A3 _6653_/A3 _4168_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_150_891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4091_ _6797_/Q input77/Z _4091_/S _4091_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6801_ _6801_/D _7281_/RN _6801_/CLK _6801_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_91_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4993_ _5223_/A1 _4963_/B _5007_/A4 _4951_/C _5109_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_91_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3944_ _3937_/Z _3941_/Z _3944_/A3 _3944_/A4 _3984_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_6732_ _6732_/D _7262_/RN _6732_/CLK _6732_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_20_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_177_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3875_ _7179_/Q _3875_/A2 _3757_/Z _6948_/Q _3877_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6663_ input75/Z _6994_/Q _4026_/C _6663_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_32_794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5614_ hold164/Z hold259/Z _5617_/S _5614_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6594_ _6594_/A1 _6603_/S _6594_/B _7306_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_145_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_844 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5545_ _4227_/B hold763/Z _6945_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_172_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5476_ _5476_/A1 _5476_/A2 _5476_/B _5476_/C _5500_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_117_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7215_ _7215_/D _7265_/RN _7215_/CLK _7215_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4427_ _5262_/A4 _5301_/A2 _5235_/A1 _4686_/B _5011_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_7146_ _7146_/D _7341_/RN _7146_/CLK _7146_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_87_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4358_ _3597_/Z _6862_/Q _4358_/S _6862_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7077_ _7077_/D _7265_/RN _7077_/CLK _7077_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_171_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4289_ hold427/Z hold5/Z _4289_/S _4289_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_104_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6028_ _7040_/Q _7162_/Q _7275_/Q _6028_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_73_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1426 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_183_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet533_167 net433_86/I _7102_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_150_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet533_178 net783_417/I _7091_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_123_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet533_156 net683_331/I _7113_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_145_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet533_189 _4109__14/I _7080_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_78_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_466 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1982 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1971 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_186_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3660_ _5544_/S _3642_/Z _3660_/B _3661_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_173_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3591_ _7095_/Q _3951_/B1 _3964_/C1 hold47/I _3594_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5330_ _5330_/A1 _5330_/A2 _5330_/B1 _5330_/B2 _5330_/C _5429_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_5261_ _5338_/A1 _5261_/A2 _5338_/A3 _5261_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_7000_ _7000_/D _7281_/RN _7000_/CLK _7000_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4212_ hold709/Z hold391/Z _4213_/S _4212_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_69_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5192_ _5192_/A1 _5402_/A2 _5192_/A3 _5435_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_87_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4143_ hold163/Z _7318_/Q _6863_/Q _4143_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_96_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4074_ _6876_/Q _4074_/A2 _4076_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_18_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_842 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_801 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4976_ _4661_/C _4956_/B _5374_/A2 _4979_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6715_ _6715_/D _7304_/RN _6715_/CLK _6715_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_52_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3927_ _6897_/Q _5838_/A2 _4405_/A3 _5546_/A2 _3947_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_20_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6646_ _6878_/Q _6648_/A3 _6646_/A3 _6649_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_164_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3858_ _3858_/A1 _3855_/Z _3858_/A3 _3858_/A4 _3885_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_50_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6577_ _6577_/A1 _6577_/A2 _6577_/A3 _6577_/A4 _6585_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_3789_ _3789_/A1 _3789_/A2 _3789_/A3 _3789_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_173_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5528_ _5535_/B _5528_/A2 _5532_/A3 _5838_/A2 _5529_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_5459_ _5459_/A1 _5459_/A2 _5459_/A3 _4443_/Z _5460_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_160_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_880 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7129_ _7129_/D _7304_/RN _7129_/CLK _7129_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_115_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_38__1374_ clkbuf_4_14_0__1374_/Z net433_86/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_28_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1289 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4830_ _4830_/A1 _4830_/A2 _5416_/A1 _4830_/B2 _6880_/Q _5043_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_73_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1790 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4761_ _3379_/I _5253_/A2 _5315_/A4 _5445_/A2 _5332_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_14_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4692_ _4690_/B _4690_/C _5484_/A2 _4720_/A2 _5307_/B _4765_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_4
X_3712_ _7238_/Q _3943_/A2 _4243_/S input48/Z _3975_/B1 _7375_/I _3714_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6500_ _7094_/Q _6578_/A2 _6310_/Z _6982_/Q _6578_/C1 hold68/I _6505_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6431_ _7246_/Q _6563_/A2 _6562_/A3 _6563_/A4 _6440_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3643_ _3460_/B _5573_/A3 _3498_/B _5745_/A4 _3643_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_162_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6362_ _7131_/Q _6287_/Z _6300_/Z _7009_/Q _6319_/Z _7123_/Q _6365_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_155_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5313_ _5313_/A1 _5399_/B _5313_/B _5483_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3574_ _3574_/A1 _3574_/A2 _3574_/A3 _3597_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_142_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6293_ _6308_/A3 _7276_/Q _7277_/Q _6324_/A1 _6313_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_170_794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5244_ _4667_/Z _5244_/A2 _5244_/A3 _5257_/B2 _5245_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_69_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold18 hold18/I hold18/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold29 hold29/I hold29/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_5175_ _4421_/Z _5177_/A1 _5177_/A3 _4759_/C _5308_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_69_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4126_ _4131_/A1 _6880_/Q _6871_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_28_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4057_ _4057_/A1 _4057_/A2 _4058_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xnet433_100 _4109__6/I _7169_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_71_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_642 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4959_ _4958_/B _4959_/A2 _4959_/B _4959_/C _5091_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_61_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_178_894 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6629_ _6629_/A1 _6629_/A2 _6630_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1020 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1042 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1053 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1097 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1086 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_837 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_848 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6980_ _6980_/D _7281_/RN _6980_/CLK _6980_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_81_726 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet833_480 net833_480/I _6729_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_53_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5931_ _5931_/A1 _5929_/Z _5931_/A3 _5931_/B _7270_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
Xclkbuf_leaf_21__1374_ _4109__51/I _4109__8/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_84__1374_ clkbuf_4_4_0__1374_/Z net833_497/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_101__1374_ clkbuf_4_4_0__1374_/Z net833_499/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xnet833_491 net833_491/I _6718_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_179_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5862_ hold208/Z hold164/Z _5865_/S _5862_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5793_ _4227_/B _3527_/Z _5866_/A3 hold8/Z hold9/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_4813_ _5267_/B _5152_/C _4822_/A4 _5266_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_178_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4744_ _5327_/B _5307_/B _4794_/A2 _5369_/A2 _5257_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_31_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4675_ _4056_/B _4669_/B _4774_/B _5200_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_135_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3626_ _7038_/Q _3977_/B1 _3946_/A2 _7022_/Q _3980_/B1 _6982_/Q _3627_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6414_ _7133_/Q _6287_/Z _6300_/Z _7011_/Q _6319_/Z _7125_/Q _6417_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_131_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6345_ _6345_/A1 _6345_/A2 _6345_/A3 _6346_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_1_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3557_ _3604_/A2 _3519_/Z _4246_/A2 _3511_/C _3971_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_143_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6276_ _7280_/Q _7281_/Q _6562_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xinput108 wb_adr_i[21] _4451_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
X_5227_ _5073_/Z _5227_/A2 _5361_/A3 _5232_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3488_ _6863_/Q _3500_/A2 hold35/Z hold36/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_115_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput119 wb_adr_i[31] _4063_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_102_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5158_ _5199_/B _5376_/A1 _5158_/B _5343_/C _5202_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_29_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5089_ _5201_/C _4828_/C _6879_/Q _5424_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_57_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_188_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_642 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_5 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_43_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_801 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4460_ _5046_/A1 _5307_/B _5048_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
Xhold307 _7068_/Q hold307/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_8_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold318 _7014_/Q hold318/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4391_ hold391/Z hold493/Z _4392_/S _4391_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold329 _7030_/Q hold329/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3411_ _7342_/Q _7338_/Q _3421_/B _3412_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3342_ _7229_/Q _3342_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_125_794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6130_ _7142_/Q _6259_/A2 _6261_/B1 _7166_/Q _6132_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_97_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_612 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6061_ _6211_/B _6266_/B _7034_/Q _7274_/Q _6064_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5012_ _5012_/A1 _5012_/A2 _5012_/A3 _5015_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_678 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6963_ _6963_/D _7281_/RN _6963_/CLK _6963_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_81_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6894_ _6894_/D _7341_/RN _6894_/CLK _6894_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5914_ _6790_/Q _6788_/Q _5917_/B _5931_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5845_ hold58/Z hold414/Z _5846_/S _5845_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_179_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5776_ hold391/Z hold813/Z hold14/Z _7146_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4727_ _4667_/Z _4727_/A2 _4727_/A3 _4960_/C _4808_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_148_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4658_ _4658_/A1 _4658_/A2 _5366_/A4 _4658_/A4 _4681_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xhold830 _5693_/Z _7073_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_123_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput90 spimemio_flash_io2_oeb input90/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3609_ _3534_/C _5655_/A4 _5532_/A3 _3454_/Z _3861_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_4589_ _4469_/B _5312_/B _4684_/B _4922_/B _5502_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xhold863 _7242_/Q hold863/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_122_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold841 _7122_/Q hold841/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold852 _4224_/Z _6772_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold874 _5857_/Z _7218_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_107_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6328_ _7186_/Q _6274_/Z _6528_/A2 _7024_/Q _6573_/A2 _7202_/Q _6334_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
Xhold896 _7327_/Q hold896/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold885 _7345_/Q _3314_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6259_ _6867_/Q _6259_/A2 _6259_/B1 _6832_/Q _6263_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_103_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_569 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3960_ _3960_/A1 _3960_/A2 _3960_/A3 _3960_/A4 _3960_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_51_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3891_ _6750_/Q _5784_/A3 _3527_/Z _5528_/A2 _3960_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5630_ hold25/Z hold454/Z _5635_/S _5630_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5561_ hold5/Z _7370_/I _5563_/S hold6/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_78_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4512_ _4686_/B _5307_/B _4869_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5492_ _5492_/A1 _5473_/Z _5432_/B _5492_/A4 _5500_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_7300_ _7300_/D _7304_/RN _7304_/CLK _7300_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold115 _7021_/Q hold115/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold104 _5908_/Z _7263_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7231_ _7231_/D _7265_/RN _7231_/CLK _7231_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_105_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold126 _7129_/Q hold126/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold148 _4294_/Z _6816_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_171_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold137 _7247_/Q hold137/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_160_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4443_ _5225_/A1 _5225_/A3 _4443_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_104_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold159 _4150_/Z _6717_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7162_ _7162_/D _7265_/RN _7162_/CLK _7162_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4374_ hold643/Z hold388/Z _4374_/S _4374_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3325_ _6787_/Q _5966_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_431 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_7093_ _7093_/D _7302_/RN _7093_/CLK _7093_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6113_ _6107_/B _6107_/C _6971_/Q _7275_/Q _6115_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_6044_ _7033_/Q _6258_/A2 _6257_/A2 _7009_/Q _6261_/B1 _7041_/Q _6045_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XTAP_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_464 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_497 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6946_ _6946_/D _7341_/RN _6946_/CLK _6946_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XTAP_1608 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6877_ _6877_/D _7323_/RN _7323_/CLK _6877_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_149_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5828_ hold2/Z hold222/Z _5828_/S _5828_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5759_ hold388/Z hold860/Z _5765_/S _7131_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_154_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_823 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold671 _6813_/Q hold671/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold660 _5602_/Z _6993_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_151_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold693 _7250_/Q hold693/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_1_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold682 _6751_/Q hold682/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_77_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet583_205 net433_56/I _7064_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet583_216 net433_68/I _7053_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_40_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_159_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet583_249 net433_71/I _7020_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet583_238 _4109__14/I _7031_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet583_227 _4109__9/I _7042_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_173_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_642 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput209 _4097_/Z mgmt_gpio_out[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_153_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4090_ _6799_/Q input67/Z _7346_/Q _4090_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_49_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6800_ _6800_/D _7281_/RN _6800_/CLK _6800_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_84_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4992_ _4992_/A1 _4992_/A2 _4992_/A3 _4998_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_91_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3943_ _7234_/Q _3943_/A2 _3943_/B1 _7194_/Q _3943_/C1 _7056_/Q _3944_/A4 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_6731_ _6731_/D _7304_/RN _6731_/CLK _6731_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_23_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3874_ _7195_/Q _3943_/B1 _3978_/B1 _6765_/Q _3945_/B1 _6757_/Q _3877_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6662_ input75/Z _6994_/Q _4026_/C _6662_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_5613_ hold139/Z hold249/Z _5617_/S _5613_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6593_ _6603_/S _7306_/Q _6594_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_182 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5544_ hold762/Z hold391/Z _5544_/S _5544_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5475_ _5491_/A2 _5470_/Z _5475_/B _5477_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7214_ _7214_/D _7265_/RN _7214_/CLK _7214_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4426_ _3379_/I _4718_/B _4661_/C _5098_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_133_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7145_ hold3/Z _7304_/RN _7145_/CLK _7145_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_101_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4357_ _6602_/A1 _4358_/S _4357_/B _6861_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_48_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7076_ _7076_/D _7265_/RN _7076_/CLK _7076_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_140_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4288_ hold495/Z hold164/Z _4289_/S _4288_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_100_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6027_ _6103_/A1 _6211_/C _7273_/Q _7272_/Q _6261_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XTAP_2117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6929_ _6929_/D _7262_/RN _6929_/CLK _6929_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_80_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet533_168 net433_68/I _7101_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_135_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet533_179 net633_288/I _7090_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_8_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet533_157 net683_331/I _7112_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_145_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold490 _4287_/Z _6810_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_89_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2640 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_898 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1961 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1950 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1983 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1994 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1972 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3590_ hold54/I _3951_/A2 _3962_/B1 _7087_/Q _3594_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_126_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5260_ _5439_/A2 _5093_/B _5260_/B _5338_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_142_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4211_ hold45/Z _6653_/A2 _5838_/A2 hold299/Z _4213_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_5191_ _4661_/C _5436_/A4 _5321_/A3 _5194_/C _5192_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_141_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4142_ hold139/Z hold292/Z _4150_/S _4142_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4073_ _4073_/A1 _4119_/B _4073_/B1 _4073_/B2 _6776_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_95_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4975_ _4975_/A1 _5374_/C _4975_/B _4979_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_91_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6714_ _6714_/D _7304_/RN _6714_/CLK _6714_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_3926_ _6936_/Q _5856_/A1 hold37/I _5784_/A3 _3965_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_51_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6645_ _5323_/C _6877_/Q _6874_/Q _6652_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_165_726 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3857_ _6727_/Q _3959_/A2 _3958_/B1 _6719_/Q _6773_/Q _3955_/C2 _3858_/A4 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_164_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3788_ _3788_/A1 _3788_/A2 _3788_/A3 _3788_/A4 _3789_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6576_ _6576_/A1 _6576_/A2 _6576_/A3 _6577_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_117_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5527_ hold388/Z hold690/Z _5527_/S _6934_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5458_ _5458_/A1 _5458_/A2 _5457_/Z _5497_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_132_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4409_ _4451_/B _4774_/B _4916_/A2 _4916_/A3 _4777_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_5389_ _5439_/A1 _5389_/A2 _5389_/B _5391_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_99_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7128_ hold76/Z _7304_/RN _7128_/CLK hold75/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_7059_ _7059_/D _7281_/RN _7059_/CLK _7059_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_101_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_654 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2470 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4760_ _5327_/B _4922_/B _4767_/A3 _5252_/A3 _5253_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_61_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4691_ _4686_/B _4759_/B1 _5312_/B _4719_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_3711_ _3711_/A1 _3711_/A2 _3711_/A3 _3711_/A4 _3711_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_174_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6430_ _7150_/Q _6562_/A2 _6562_/A3 _6561_/A3 _6437_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3642_ _7294_/Q _6942_/Q _6944_/Q _3642_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_146_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6361_ _7163_/Q _6279_/Z _6299_/Z _7065_/Q _6575_/B1 _7049_/Q _6365_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_60_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5312_ _5312_/A1 _5313_/A1 _5312_/B _5312_/C _5314_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3573_ _6983_/Q _3980_/B1 _3875_/A2 hold50/I _3574_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xclkbuf_leaf_44__1374_ clkbuf_4_15_0__1374_/Z net783_435/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6292_ _7279_/Q _7278_/Q _6457_/A3 _6562_/A4 _6292_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
X_5243_ _5267_/C _5327_/B _5243_/A3 _5243_/B _5328_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_102_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold19 hold19/I hold19/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_114_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5174_ _5502_/B2 _5502_/A1 _5302_/B _5199_/A2 _5388_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_111_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4125_ _6951_/Q input39/Z _4125_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_83_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4056_ _4669_/B _5166_/A4 _4056_/B _4840_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_84_768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet433_101 _4109__4/I _7168_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4958_ _4451_/B _5166_/A4 _4958_/B _4959_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_61_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3909_ _7146_/Q hold299/I _5727_/A3 _5856_/A2 _3942_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_4889_ _5177_/A3 _5153_/A2 _5153_/B _5399_/B _5263_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6628_ _6878_/Q _6628_/A2 _6628_/B1 _6640_/B2 _6629_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_153_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6559_ _6559_/I0 _7303_/Q _6559_/S _7303_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_105_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_640 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1010 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1021 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1032 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1065 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1054 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1098 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1087 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_816 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_827 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet833_481 net833_483/I _6728_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet833_470 net833_470/I _6739_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5930_ _5930_/A1 _5930_/A2 _6790_/Q _5930_/B1 _7270_/Q _5931_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
Xnet833_492 net433_97/I _6717_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5861_ _5865_/S _5861_/A2 _5861_/B hold465/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_827 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4812_ _4819_/A4 _4667_/Z _4959_/C _4451_/B _4823_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_21_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5792_ hold2/Z hold337/Z _5792_/S _7161_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4743_ _4706_/Z _4709_/Z _4825_/A4 _5376_/A1 _4748_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_175_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4674_ _5166_/A4 _4916_/A2 _4916_/A3 _4451_/B _5194_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_135_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6413_ _6410_/Z _6413_/A2 _6413_/A3 _6413_/A4 _6413_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_3625_ _7192_/Q _5700_/A1 _5820_/A2 _3527_/Z _3627_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_134_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3556_ _3811_/A1 _3511_/C _3473_/B _3833_/A2 _3980_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_6344_ _7040_/Q _6297_/Z _6300_/Z _7008_/Q _6345_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_143_762 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6275_ _7279_/Q _7278_/Q _6563_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_103_604 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput109 wb_adr_i[22] _4916_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_5226_ _5226_/A1 _5226_/A2 _5225_/Z _5459_/A3 _5361_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3487_ _6863_/Q hold34/Z hold35/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_5157_ _5157_/A1 _5472_/A3 _5472_/A4 _5158_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_56_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4108_ _6863_/Q _4108_/A2 _4108_/B1 _4108_/B2 _4108_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5088_ _5088_/A1 _5366_/A1 _5236_/B _5201_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_96_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4039_ _6788_/Q _6789_/Q _6532_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_112_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_762 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_90__1374_ net583_226/I _4109__44/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_94_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_568 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_71 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_871 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold308 _7198_/Q hold308/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_117_729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold319 _5625_/Z _7014_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4390_ _4405_/A3 hold45/Z _6653_/A2 hold41/Z _4392_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_3410_ _4073_/B1 _3421_/B _7342_/Q _3412_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3341_ _7237_/Q _3341_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_124_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6060_ _6060_/I0 _7286_/Q _6559_/S _7286_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5011_ _4963_/B _5011_/A2 _4773_/B _5288_/A4 _5378_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_112_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_679 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6962_ _6962_/D _7281_/RN _6962_/CLK _6962_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_81_535 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6893_ _6893_/D _7341_/RN _6893_/CLK _6893_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5913_ _4019_/Z _6788_/Q _5917_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_50_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5844_ hold5/Z hold385/Z _5846_/S _5844_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5775_ hold299/I _5866_/A3 hold13/Z _4227_/B hold14/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_4726_ _5235_/A1 _4718_/B _3380_/I _4729_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_163_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4657_ _5459_/A3 _5445_/A3 _5471_/A1 _5051_/B _4658_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_162_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3608_ _3827_/A1 _3477_/Z _3483_/Z _3608_/A4 _3786_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xinput91 spimemio_flash_io3_do input91/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_7376_ _7376_/I _7376_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput80 spi_sck input80/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold820 _6758_/Q hold820/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold831 _7057_/Q hold831/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold853 _7358_/I hold853/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold864 _7357_/I hold864/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_162_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4588_ _4469_/B _4922_/B _4684_/B _5312_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_6327_ _7130_/Q _6287_/Z _6564_/C1 _7080_/Q _6339_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_89_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold842 _7041_/Q hold842/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold897 _6703_/Q hold897/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_143_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3539_ _3827_/A2 _3496_/B _3833_/A2 _4246_/A1 _3940_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_115_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold886 hold886/I _7345_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold875 _6912_/Q hold875/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6258_ _6882_/Q _6258_/A2 _6258_/B1 _6844_/Q _6258_/C1 _6890_/Q _6264_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_5209_ _5209_/A1 _5351_/A1 _5209_/B1 _5346_/A4 _5464_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6189_ _7275_/Q _6177_/Z _6189_/B _6189_/C _6192_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_85_830 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_844 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_754 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3890_ _6899_/Q hold37/I hold41/I hold190/I _3974_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_148_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5560_ hold164/Z hold394/Z _5563_/S _5560_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_157_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4511_ _5350_/B _5394_/A2 _5439_/C _5315_/A4 _4565_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5491_ _5491_/A1 _5491_/A2 _5490_/Z _5492_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4442_ _4957_/A4 _4417_/Z _4452_/A2 _5166_/A4 _5225_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
Xhold116 _5633_/Z _7021_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_145_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold105 _7168_/Q hold105/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7230_ _7230_/D _7265_/RN _7230_/CLK _7230_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_117_537 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold138 _7330_/Q hold138/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_172_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold149 _6995_/Q hold149/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold127 _5756_/Z _7129_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_144_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4373_ hold727/Z hold391/Z _4374_/S _4373_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7161_ _7161_/D _7302_/RN _7161_/CLK _7161_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3324_ _6994_/Q _4107_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_7092_ _7092_/D _7281_/RN _7092_/CLK _7092_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_86_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6112_ _6112_/A1 _6112_/A2 _6112_/B _6112_/C _6115_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6043_ _7073_/Q _6260_/A2 _6256_/B1 _7081_/Q _6045_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_58_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_498 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6945_ _6945_/D _7281_/RN _6945_/CLK _6945_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_1609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_719 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6876_ _6876_/D _7323_/RN _7323_/CLK _6876_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_179_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5827_ hold58/Z hold304/Z _5828_/S _5827_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_10_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5758_ hold391/Z hold740/Z _5765_/S _7130_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4709_ _4710_/C _4767_/A3 _4710_/B _4709_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_175_481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5689_ hold58/Z hold82/Z hold42/Z _7070_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7359_ _7359_/I _7359_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold672 _4291_/Z _6813_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold661 _7081_/Q hold661/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_78_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xmax_cap380 input75/Z _7262_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
Xhold650 _6951_/Q hold650/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold694 _7105_/Q hold694/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_2_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold683 _4192_/Z _6751_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_134_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet583_206 net633_277/I _7063_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_9_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet583_217 net433_87/I _7052_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_159_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet583_239 net783_420/I _7030_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet583_228 _4109__49/I _7041_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_127_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_181_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_391 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_719 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4991_ _5004_/A1 input95/Z _5153_/A2 _5372_/B _4992_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_90_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6730_ _6730_/D _7304_/RN _6730_/CLK _6730_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_189_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3942_ _6710_/Q _3942_/A2 _3942_/B1 _7340_/Q _3942_/C _3944_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_16_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6661_ _7341_/RN _6994_/Q _4026_/C _6661_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_90_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3873_ _3873_/A1 _3873_/A2 _3873_/A3 _3873_/A4 _3884_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6592_ _6877_/D _7323_/RN _6603_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_149_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5612_ hold25/Z hold502/Z _5617_/S _5612_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_14_0__1374_ clkbuf_3_7_0__1374_/Z clkbuf_4_14_0__1374_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_118_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5543_ hold388/Z hold615/Z _5543_/S _5543_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_129_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5474_ _5492_/A4 _5432_/B _5473_/Z _5475_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_7213_ _7213_/D _7265_/RN _7213_/CLK _7213_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4425_ _3379_/I _4718_/B _4661_/C _4425_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
X_7144_ hold71/Z _7304_/RN _7144_/CLK hold70/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4356_ _4358_/S _6861_/Q _4357_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7075_ _7075_/D _7265_/RN _7075_/CLK _7075_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_140_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4287_ hold489/Z hold139/Z _4289_/S _4287_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6026_ _6026_/A1 _6026_/A2 _6026_/B1 _6026_/B2 _6031_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_2107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6928_ _6928_/D _7262_/RN _6928_/CLK _6928_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_167_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6859_ _6859_/D _7313_/CLK _6859_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_654 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet533_169 net433_90/I _7100_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_108_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_8__1374_ clkbuf_4_3_0__1374_/Z net783_445/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_2_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet533_158 net433_94/I _7111_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold480 _4295_/Z _6817_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold491 _6892_/Q hold491/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_1_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2652 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2674 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1951 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1940 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_847 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1984 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1995 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1973 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1962 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4210_ hold388/Z hold655/Z _4210_/S _4210_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4109__50 net433_66/I _7219_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_141_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5190_ _5190_/A1 _5483_/C _5230_/C _5469_/A4 _5190_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_4141_ hold138/Z _7317_/Q _6863_/Q _4141_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_122_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4072_ _4073_/B2 _7337_/Q _4072_/A3 _7336_/Q _4073_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_48_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4974_ _5374_/A2 _5454_/A1 _4975_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3925_ _6901_/Q _5856_/A2 _4405_/A3 _4405_/A2 _3947_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xclkbuf_leaf_67__1374_ _4109__12/I net633_288/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6713_ _6713_/D _7304_/RN _6713_/CLK _6713_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_51_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6644_ _6872_/Q _6644_/A2 _4363_/Z _7322_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_60_880 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3856_ input53/Z _4264_/A1 _3643_/Z _6928_/Q _3856_/C _3858_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_3787_ _7148_/Q _3866_/A2 _3943_/C1 _7058_/Q _7010_/Q _3962_/A2 _3788_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6575_ _6765_/Q _6575_/A2 _6575_/B1 _6886_/Q _6576_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_20_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5526_ hold391/Z hold785/Z _5527_/S _6933_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_172_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5457_ _5457_/A1 _5457_/A2 _5457_/A3 _4647_/C _5457_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_4408_ _5323_/C _6876_/Q hold20/I _5043_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_105_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5388_ _5388_/A1 _5388_/A2 _5388_/A3 _5388_/A4 _5504_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_87_722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4339_ _4354_/A1 _4343_/S _4339_/B _6849_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7127_ hold92/Z _7302_/RN _7127_/CLK hold91/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_7058_ _7058_/D _7265_/RN _7058_/CLK _7058_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_101_543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6009_ _6992_/Q _6258_/B1 _6261_/A2 _7000_/Q _6016_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_87_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1214 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1781 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3710_ _7182_/Q _3875_/A2 _3953_/B1 _7190_/Q _3711_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_81_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_571 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4690_ _5262_/A4 _5315_/A4 _4690_/B _4690_/C _4759_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_3641_ _3888_/S _3641_/A2 _3641_/B hold877/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3572_ _7055_/Q _3973_/A2 _3946_/A2 hold52/I _6991_/Q _3939_/A2 _3574_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6360_ _6360_/A1 _6360_/A2 _6360_/A3 _6366_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_115_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5311_ _5323_/A1 _5468_/A1 _5439_/B _5439_/C _5401_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_53_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6291_ _6306_/A3 _6324_/A1 _6308_/A3 _7277_/Q _6317_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_114_145 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5242_ _5242_/A1 _5242_/A2 _5429_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5173_ _5437_/A4 _5312_/A1 _5173_/B _5176_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4124_ _6950_/Q input70/Z _4124_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_110_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput1 debug_mode input1/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4055_ _4916_/A2 _4916_/A3 _4056_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_37_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_319 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_828 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4957_ _4959_/A2 _4957_/A2 _4417_/Z _4957_/A4 _4960_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_51_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4888_ _5399_/B _5489_/B1 _4888_/B _4891_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3908_ _6927_/Q _5745_/A4 _5518_/A1 _5552_/A2 _3960_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6627_ _6880_/Q _6627_/A2 _6627_/B1 _6879_/Q _6629_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_137_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3839_ _6934_/Q _5802_/A2 _5727_/A3 _5552_/A2 _3867_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_134_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6558_ _6558_/A1 _6558_/A2 _6558_/B _6559_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_152_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6489_ _6990_/Q _6511_/A2 _6563_/A4 _6562_/A4 _6490_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_5509_ _5838_/A4 _5532_/A3 _5838_/A2 _5884_/A2 _5511_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_3_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1011 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1022 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_15_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1033 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1055 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_830 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_50__1374_ clkbuf_4_15_0__1374_/Z net583_250/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1099 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1088 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1066 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1077 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_167_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_817 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_828 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_839 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet833_460 net833_464/I _6749_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_18_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet833_471 net833_471/I _6738_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5860_ _3527_/Z hold463/Z _4227_/B hold139/Z hold464/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xnet833_482 net833_483/I _6727_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet833_493 net433_97/I _6716_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_179_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4811_ _4811_/A1 _4811_/A2 _4811_/A3 _4811_/A4 _4811_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XTAP_2290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_474 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5791_ hold58/Z hold96/Z _5792_/S hold97/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4742_ _5315_/A4 _5301_/A2 _4661_/C _3379_/I _5369_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_174_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4673_ _4451_/B _4916_/A2 _4916_/A3 _4667_/Z _5267_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_2
XFILLER_119_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_4_2_0__1374_ clkbuf_4_3_0__1374_/I clkbuf_4_2_0__1374_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_174_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3624_ _7136_/Q _3945_/A2 _4281_/S input41/Z _3964_/C1 hold80/I _3627_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6412_ _7075_/Q _6292_/Z _6571_/B1 _6987_/Q _6571_/C1 _7181_/Q _6413_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_175_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3555_ _3498_/B _4246_/A1 _3802_/A2 _3460_/B _3950_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_6343_ _6976_/Q _6457_/A3 _6563_/A4 _6562_/A4 _6345_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3486_ hold170/Z _6777_/Q _6705_/Q _3500_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_6274_ _7279_/Q _7278_/Q _6563_/A3 _6561_/A3 _6274_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_0_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5225_ _5225_/A1 _5225_/A2 _5225_/A3 _4437_/Z _5225_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_103_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5156_ _5156_/A1 _5239_/B _5156_/A3 _5157_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_56_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5087_ _5087_/A1 _5087_/A2 _5087_/B _5236_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4107_ _4107_/A1 _6946_/Q input67/Z _6863_/Q _4108_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_110_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4038_ _5925_/B _7270_/Q _5930_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5989_ _6584_/B _6789_/Q _6587_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_52_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_847 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput190 _3348_/ZN mgmt_gpio_oeb[27] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_121_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_754 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_153_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_188_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_474 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold309 _7020_/Q hold309/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_171_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5010_ _3379_/I input95/Z _4423_/Z _5282_/B _5012_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6961_ _6961_/D _7281_/RN _6961_/CLK _6961_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_47_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6892_ _6892_/D _7341_/RN _6892_/CLK _6892_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5912_ _6790_/Q _4051_/B _5912_/B _7266_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5843_ hold164/Z hold485/Z _5846_/S _5843_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_844 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5774_ hold2/Z _7145_/Q _5774_/S hold3/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_175_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4725_ _4667_/Z _5244_/A2 _4693_/Z _5468_/C _4725_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_174_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4656_ _5262_/A4 _5235_/A1 _4718_/B _3380_/I _5466_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_107_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4587_ _5082_/C _4454_/B _4587_/A3 _5435_/A1 _5063_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_163_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_847 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold810 _5821_/Z _7186_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7375_ _7375_/I _7375_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3607_ _7046_/Q _5655_/A4 _5727_/A3 hold29/I _3612_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xinput70 mgmt_gpio_in[7] input70/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput81 spi_sdo input81/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold821 _4203_/Z _6758_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold854 _4232_/Z _6780_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold832 _7072_/Q hold832/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3538_ _5534_/A1 _3827_/A2 _3496_/B _4246_/A1 _3975_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_6326_ _7088_/Q _6578_/A2 _6309_/Z _7234_/Q _6341_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_107_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput92 spimemio_flash_io3_oeb input92/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold843 _6927_/Q hold843/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold865 _4230_/Z _6779_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold887 _6706_/Q hold887/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_143_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold876 _6918_/Q hold876/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold898 _6776_/Q hold898/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3469_ hold460/Z _3469_/A2 _6863_/Q _3473_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_89_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6257_ _6865_/Q _6257_/A2 _6257_/B1 _6888_/Q _6264_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_77_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5208_ _5223_/A1 _5048_/C _5208_/A3 _5295_/A1 _5208_/B2 _5209_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_131_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6188_ _6188_/A1 _6188_/A2 _7275_/Q _6189_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5139_ _5476_/A1 _5253_/A2 _5148_/B1 _5502_/A2 _5490_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_177_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_1_1__f__1033_ clkbuf_0__1033_/Z _6599_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_153_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_188_265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_184_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4510_ _5177_/A3 _5315_/A4 _5262_/A4 _4423_/Z _5186_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_5490_ _5490_/A1 _5490_/A2 _5490_/A3 _5490_/A4 _5490_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_8_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4441_ _4774_/A1 _4451_/A2 _4774_/B _5225_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
Xhold106 _7167_/Q hold106/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold117 _7031_/Q hold117/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_171_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold139 _4141_/Z hold139/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold128 _7111_/Q hold128/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7160_ hold97/Z _7302_/RN _7160_/CLK hold96/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6111_ _7275_/Q _6111_/A2 _6111_/B _6112_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4372_ _5535_/B _6653_/A2 _5838_/A2 _4378_/A1 _4374_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XTAP_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_7091_ _7091_/D _7281_/RN _7091_/CLK _7091_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3323_ _6874_/Q _4068_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_112_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6042_ _7017_/Q _6259_/A2 _6256_/A2 _7049_/Q _6045_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_466 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_867 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6944_ _6944_/D _7304_/RN _6944_/CLK _6944_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_23_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6875_ _6875_/D _7323_/RN _7323_/CLK _6875_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_34_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5826_ hold5/Z hold101/Z _5828_/S _5826_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5757_ hold299/Z _5884_/A2 _5838_/A2 _5535_/B _5765_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_147_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4708_ _4720_/A3 _4720_/A2 _4690_/B _4759_/B1 _4719_/B _4822_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_4
X_5688_ hold5/Z hold119/Z hold42/Z _7069_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4639_ _4481_/C _4628_/B _5271_/A1 _5062_/A3 _5050_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_151_828 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xmax_cap381 _5004_/A1 _3379_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
X_7358_ _7358_/I _7358_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold662 _5702_/Z _7081_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_118_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold640 _4213_/Z _6765_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_78_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold651 _6767_/Q hold651/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold673 _6961_/Q hold673/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6309_ _6511_/A2 _6312_/A4 _7281_/Q _6563_/A4 _6309_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_104_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold695 _7171_/Q hold695/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold684 _6739_/Q hold684/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7289_ _7289_/D _7302_/RN _7304_/CLK _7289_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_104_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet583_207 _4109__29/I _7062_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_9_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet583_218 net683_320/I _7051_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_139_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet583_229 _4109__9/I _7040_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_166_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_801 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4990_ _4661_/C _4956_/B _5372_/B _4992_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_90_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3941_ _3941_/A1 _3941_/A2 _3941_/A3 _3941_/A4 _3941_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_32_731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6660_ _7341_/RN _6994_/Q _4026_/C _6660_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_3872_ _3861_/Z _3872_/A2 _3872_/A3 _3871_/Z _3884_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_31_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6591_ _6591_/I _7305_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_176_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5611_ hold388/Z hold744/Z _5617_/S _5611_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5542_ hold58/Z hold195/Z _5543_/S _5542_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_185_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5473_ _5473_/A1 _5473_/A2 _5473_/A3 _5472_/Z _5473_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_7212_ _7212_/D _7265_/RN _7212_/CLK _7212_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4424_ _4718_/B _4661_/C _4690_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_160_614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_828 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_27__1374_ clkbuf_4_14_0__1374_/Z _4109__4/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_7143_ _7143_/D _7262_/RN _7143_/CLK _7143_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xclkbuf_leaf_107__1374_ net733_398/I net783_437/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4355_ _6600_/I0 _6860_/Q _4358_/S _6860_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7074_ _7074_/D _7265_/RN _7074_/CLK _7074_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_58_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4286_ hold475/Z hold25/Z _4289_/S _4286_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_100_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6025_ _6025_/A1 _6025_/A2 _6025_/A3 _6025_/A4 _6026_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_2108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1429 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6927_ _6927_/D _7262_/RN _6927_/CLK _6927_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6858_ _6858_/D _6862_/CLK _6858_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_168_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5809_ hold58/Z hold68/Z _5810_/S hold69/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_13_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6789_ _6789_/D _7281_/RN _7281_/CLK _6789_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_13_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet533_159 net533_163/I _7110_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold470 _7180_/Q hold470/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold481 _7044_/Q hold481/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_150_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold492 _4392_/Z _6892_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_77_403 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2642 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2675 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1952 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1930 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1985 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1974 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1963 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4109__40 net433_71/I _7229_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_141_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4109__51 _4109__51/I _7218_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_79_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4140_ hold25/Z hold311/Z _4150_/S _4140_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4071_ _4071_/A1 hold896/Z _3446_/B _4073_/B1 _3387_/Z _6777_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_83_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4973_ _5106_/A4 _4973_/A2 _5374_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3924_ input71/Z hold37/I _5884_/A2 _5856_/A2 _3982_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6712_ _6712_/D _7304_/RN _6712_/CLK _6712_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_6643_ _4362_/Z _6877_/Q _6870_/Q _6643_/A4 _6644_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_137_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3855_ _3855_/A1 _3855_/A2 _3855_/A3 _3855_/A4 _3855_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_118_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3786_ _7090_/Q _3951_/B1 _3786_/B1 _3786_/B2 _3788_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6574_ _6757_/Q _6287_/Z _6300_/Z _6865_/Q _6319_/Z _6753_/Q _6576_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_161_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5525_ _5535_/B _5552_/A2 _5727_/A3 _5802_/A2 _5527_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_173_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5456_ _5456_/A1 _5455_/Z _5477_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_172_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4407_ hold388/Z hold562/Z _4407_/S _6902_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_132_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5387_ _5439_/A1 _5439_/A2 _5439_/C _5503_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4338_ _4343_/S _6849_/Q _4339_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7126_ _7126_/D _7302_/RN _7126_/CLK _7126_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_7057_ _7057_/D _7265_/RN _7057_/CLK _7057_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4269_ hold673/Z hold388/Z _4281_/S _4269_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_86_255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6008_ _6211_/B _7274_/Q _7271_/Q _7272_/Q _6261_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_28_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_188_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_319 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_861 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_10__1374_ clkbuf_4_8_0__1374_/Z net433_74/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_49_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_73__1374_ clkbuf_4_5_0__1374_/Z net783_424/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_38_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_845 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1793 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_159_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3640_ _3888_/S hold876/Z _3641_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3571_ input28/Z _3977_/A2 _3942_/A2 _6717_/Q _7137_/Q _3945_/A2 _3574_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_161_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6290_ _6324_/A1 _6308_/A3 _7278_/Q _6321_/A4 _6570_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_5310_ _5440_/A3 _5308_/Z _5440_/A1 _5310_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_5241_ _4667_/Z _5244_/A2 _5241_/A3 _5257_/B2 _5242_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_69_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5172_ _5172_/A1 _5172_/A2 _5172_/A3 _5173_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_114_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4123_ input1/Z input36/Z _4123_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_110_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput2 debug_oeb input2/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4054_ _4054_/A1 _7327_/Q _4054_/B hold884/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_848 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_678 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4956_ _4967_/A2 _4956_/A2 _4956_/B _4956_/C _4969_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_178_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3907_ _6843_/Q _5745_/A4 _4378_/A1 _5546_/A2 _3949_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4887_ _4887_/A1 _4887_/A2 _4887_/A3 _4887_/A4 _4888_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_20_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6626_ _6626_/I0 _7317_/Q _6642_/S _7317_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_165_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3838_ _6886_/Q _5745_/A4 _4405_/A3 _4405_/A2 _3873_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_153_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6557_ _6788_/Q _7302_/Q _6558_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3769_ _3766_/Z _3769_/A2 _3769_/A3 _3769_/A4 _3790_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_118_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5508_ hold737/Z hold388/Z _5508_/S _5508_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6488_ hold83/I _6570_/A2 _6570_/B1 hold66/I _6570_/C1 _6998_/Q _6491_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_106_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5439_ _5439_/A1 _5439_/A2 _5439_/B _5439_/C _5440_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_133_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7109_ hold94/Z _7304_/RN _7109_/CLK hold93/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_102_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1001 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1023 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1034 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1056 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1045 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1089 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_878 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_183_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_829 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet833_472 net833_472/I _6737_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet833_461 net433_93/I _6748_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_34_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet833_494 net433_93/I _6715_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet833_483 net833_483/I _6726_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_46_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4810_ _5439_/A2 _4693_/Z _5468_/C _4706_/Z _4811_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_18_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5790_ hold5/Z hold438/Z _5792_/S _7159_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4741_ _5262_/A4 _5235_/A1 _4718_/B _3380_/I _5376_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_187_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4672_ _4451_/B _4916_/A2 _4916_/A3 _4667_/Z _5471_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_174_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3623_ hold95/I _3981_/A2 _4264_/A1 input59/Z _3635_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6411_ _7213_/Q _6570_/A2 _6570_/B1 _7059_/Q _6570_/C1 _6995_/Q _6413_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_174_399 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3554_ _5534_/A1 _3802_/A2 _3473_/B _3507_/C _3962_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_6342_ _7146_/Q _6575_/A2 _6285_/Z _7104_/Q _6342_/C _6347_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_3485_ _6704_/Q _6777_/Q _4001_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6273_ _5917_/B _6587_/A2 _7295_/Q _6349_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5224_ _5224_/A1 _5358_/B _5419_/B _5227_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_170_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5155_ _5473_/A1 _5473_/A2 _5156_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5086_ _5087_/A1 _5086_/A2 _4956_/B _5366_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_84_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4106_ _7284_/Q _6940_/Q _6944_/Q _4106_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4037_ _5985_/A3 _7267_/Q _5930_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5988_ _6584_/B _6789_/Q _6509_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_184_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4939_ _4963_/B _4926_/C _4995_/A4 _4922_/B _5282_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_166_823 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6609_ _6876_/Q _6651_/A2 _6609_/B1 _6879_/Q _6610_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_165_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_750 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_403 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput180 _3357_/ZN mgmt_gpio_oeb[18] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput191 _3347_/ZN mgmt_gpio_oeb[28] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_101_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_877 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_604 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_789 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6960_ _6960_/D _7281_/RN _6960_/CLK _6960_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_38_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5911_ _5966_/I0 _6790_/Q _5911_/B _7266_/Q _5912_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_93_375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6891_ _6891_/D _7341_/RN _6891_/CLK _6891_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_62_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5842_ hold139/Z hold358/Z _5846_/S _5842_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_61_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5773_ hold58/Z hold70/Z _5774_/S hold71/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_166_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_823 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4724_ _4722_/Z _4750_/A4 _4750_/A3 _4960_/C _4729_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_159_182 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4655_ _5315_/A4 _5301_/A2 _4661_/C _3379_/I _5471_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xhold811 _7210_/Q hold811/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4586_ _5136_/A2 _5466_/B _5295_/A1 _4922_/B _4592_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
Xinput60 mgmt_gpio_in[31] input60/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3606_ _7200_/Q _5884_/A2 _5902_/A3 _3527_/Z _3630_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xinput71 mgmt_gpio_in[8] input71/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_7374_ _7374_/I _7374_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold800 _4136_/Z _6710_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xinput82 spi_sdoenb input82/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold855 _7064_/Q hold855/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold833 _5692_/Z _7072_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3537_ _3460_/B _3498_/B _3604_/A2 hold462/Z hold463/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_131_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6325_ _6325_/A1 _6325_/A2 _7279_/Q _7278_/Q _6568_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_89_604 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold844 _6807_/Q hold844/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xinput93 trap input93/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold822 _6760_/Q hold822/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold866 _6800_/Q hold866/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold877 hold877/I _6918_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold888 _7339_/Q hold888/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3468_ _4073_/B1 hold297/Z _3469_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6256_ _6886_/Q _6256_/A2 _6256_/B1 _6894_/Q _6264_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold899 hold899/I _7342_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_5207_ _5207_/A1 _5207_/A2 _5207_/B _6904_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_103_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6187_ _6187_/A1 _6187_/A2 _6187_/A3 _6187_/A4 _6188_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3399_ _4071_/A1 hold892/Z _3401_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5138_ _5376_/A1 _5253_/A2 _5502_/B1 _5502_/B2 _5141_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_57_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5069_ _4443_/Z _5459_/A3 _5372_/A1 _5225_/A2 _5071_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_72_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_189_789 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4440_ _3380_/I _4922_/B _4421_/Z _4425_/Z _4451_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_156_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold107 _6983_/Q hold107/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_172_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold118 _5645_/Z _7031_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold129 _5735_/Z _7111_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_113_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6110_ _7275_/Q _6110_/A2 _6108_/Z _6262_/A2 _6109_/Z _6261_/A2 _6111_/B VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_4371_ hold641/Z hold388/Z _4371_/S _4371_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_112_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7090_ _7090_/D _7302_/RN _7090_/CLK _7090_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XTAP_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3322_ _3322_/I _4054_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_79_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6041_ _7272_/Q _7271_/Q _6041_/A3 _6041_/B1 _6041_/B2 _6056_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XTAP_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_640 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6943_ _6943_/D _7304_/RN _6943_/CLK _6943_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6874_ _6877_/Q _7323_/RN _7323_/CLK _6874_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_179_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_762 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5825_ hold164/Z hold510/Z _5828_/S _5825_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_167_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_754 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5756_ hold2/Z hold126/Z _5756_/S _5756_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5687_ hold164/Z hold307/Z hold42/Z _7068_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4707_ _4707_/A1 _4665_/Z _4750_/A3 _4960_/C _5327_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_4638_ _5301_/A2 _5235_/A1 _3379_/I _3380_/I _5271_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_163_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold630 _6822_/Q hold630/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_2_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4569_ _5051_/B _4568_/Z _4454_/B _4959_/C _5420_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_7357_ _7357_/I _7357_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold663 _7355_/I hold663/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xmax_cap360 _5646_/A2 _4378_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
Xhold641 _6867_/Q hold641/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold652 _4216_/Z _6767_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6308_ _6323_/A1 _6325_/A1 _6308_/A3 _7279_/Q _6566_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xhold674 _7361_/I hold674/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold696 _5804_/Z _7171_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold685 _7139_/Q hold685/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7288_ _7288_/D _7302_/RN _7302_/CLK _7288_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_134_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6239_ _6760_/Q _6259_/A2 _6262_/A2 _6754_/Q _6240_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_58_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_990 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet583_219 _4109__28/I _7050_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet583_208 net583_214/I _7061_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_185_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_843 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_865 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3940_ _7210_/Q _3940_/A2 _3940_/B _3941_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_91_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3871_ _3868_/Z _3871_/A2 _3871_/A3 _3871_/A4 _3871_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_6590_ _6590_/A1 _7305_/Q _6877_/D _6589_/B _6591_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5610_ hold391/Z hold797/Z _5617_/S _5610_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5541_ hold5/Z hold218/Z _5543_/S _5541_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_145_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7211_ _7211_/D _7265_/RN _7211_/CLK _7211_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_129_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5472_ _5472_/A1 _5472_/A2 _5472_/A3 _5472_/A4 _5472_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_4423_ _4718_/B _4661_/C _4423_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_141_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4354_ _4354_/A1 _4358_/S _4354_/B _6859_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7142_ _7142_/D _7302_/RN _7142_/CLK _7142_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_7073_ _7073_/D _7265_/RN _7073_/CLK _7073_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_141_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6024_ _7112_/Q _6260_/B1 _6257_/B1 _7178_/Q _6025_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4285_ hold781/Z hold388/Z _4289_/S _4285_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_100_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_687 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6926_ _6926_/D _7262_/RN _6926_/CLK _6926_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_35_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6857_ _6857_/D _6862_/CLK _6857_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5808_ hold5/Z hold240/Z _5810_/S _5808_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6788_ _6788_/D _7304_/RN _7304_/CLK _6788_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
X_5739_ hold530/Z hold25/Z _5744_/S _7114_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_109_848 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold471 _5814_/Z _7180_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold460 _4011_/B hold460/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold493 _6891_/Q hold493/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold482 _6926_/Q hold482/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_145_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2654 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2687 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1942 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1931 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1986 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1975 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1964 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1953 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1997 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_33__1374_ clkbuf_4_11_0__1374_/Z net433_87/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_13_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_96__1374_ clkbuf_4_1_0__1374_/Z net833_471/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_113__1374_ clkbuf_4_2_0__1374_/Z net833_469/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_2_2__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/Z _4108_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_126_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4109__30 net433_53/I _7239_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4109__41 net433_71/I _7228_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_142_659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_512 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4070_ hold893/Z _4069_/Z _6778_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_95_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_462 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4972_ _5001_/A1 _5374_/A2 _4973_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6711_ _6711_/D _7304_/RN _6711_/CLK _6711_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_3923_ _6831_/Q _5784_/A3 _6653_/A2 _5552_/A2 _3960_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6642_ _6642_/I0 _7321_/Q _6642_/S _7321_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_149_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_573 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3854_ _7155_/Q _3956_/B1 _3968_/B1 _6767_/Q _3854_/C1 _7121_/Q _3858_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_177_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3785_ _7002_/Q _3961_/A2 _3951_/A2 _7074_/Q _7082_/Q _3962_/B1 _3788_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6573_ _6759_/Q _6573_/A2 _6288_/Z _6763_/Q _6297_/Z _6884_/Q _6576_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_9_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5524_ hold5/Z hold233/Z _5524_/S _6932_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_172_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5455_ _5455_/A1 _5455_/A2 _5455_/A3 _5455_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_117_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4406_ hold391/Z hold563/Z _4407_/S _6901_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5386_ _5386_/A1 _5380_/Z _5386_/A3 _5386_/B _5408_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_7125_ _7125_/D _7262_/RN _7125_/CLK _7125_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_141_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4337_ _6597_/I0 _6848_/Q _4343_/S _6848_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7056_ _7056_/D _7341_/RN _7056_/CLK _7056_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_140_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4268_ _4267_/Z hold871/Z _4282_/S _4268_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6007_ _6036_/A3 _6103_/A1 _7274_/Q _7273_/Q _6258_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_4199_ _5535_/B _5546_/A2 _5748_/A3 hold299/Z _4201_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_27_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6909_ _6909_/D _7323_/RN _7322_/CLK hold34/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_1249 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold290 _5852_/Z _7214_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_77_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2462 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_512 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1750 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_843 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_187_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3570_ _3604_/A2 _3802_/A2 _3511_/C _3833_/A2 _3943_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_161_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5240_ _5416_/A1 _5271_/A4 _5257_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_170_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5171_ _5199_/A2 _5298_/B _5390_/A1 _5404_/A2 _5171_/C _5172_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_39_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4122_ _4087_/S input63/Z _4122_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4053_ _4044_/Z _6325_/A1 _6307_/A1 _4053_/B _6790_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_83_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput3 debug_out input3/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_52_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4955_ _4947_/C _4951_/C _4955_/B _4963_/B _5274_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_52_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3906_ _6736_/Q _5745_/A4 hold37/I _4405_/A2 _3978_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_33_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4886_ _5445_/A2 _5177_/A3 _5153_/B _5399_/B _4887_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_32_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6625_ _6625_/A1 _6625_/A2 _6626_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3837_ _6844_/Q _5745_/A4 _4378_/A1 _5546_/A2 _3886_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_3768_ input45/Z _4243_/S _3975_/B1 input63/Z _3945_/A2 _7132_/Q _3769_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6556_ _6584_/A1 _6829_/Q _6584_/B _6558_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_173_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5507_ hold746/Z hold391/Z _5508_/S _5507_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_145_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6487_ _7208_/Q _6573_/A2 _6288_/Z _7200_/Q _6297_/Z _7046_/Q _6491_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_3699_ _7076_/Q _3951_/A2 _3961_/B1 _7028_/Q _3951_/B1 _7092_/Q _3700_/I VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_10_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5438_ _5438_/A1 _5395_/Z _5438_/A3 _5438_/A4 _5504_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_105_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput340 _6862_/Q wb_dat_o[7] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5369_ _5369_/A1 _5369_/A2 _5498_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_87_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_180 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7108_ _7108_/D _7304_/RN _7108_/CLK _7108_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_102_898 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7039_ hold86/Z _7281_/RN _7039_/CLK hold85/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_74_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_opt_2_0__1374_ clkbuf_4_8_0__1374_/Z net683_310/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_28_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1002 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1013 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1024 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1046 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1057 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1068 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_167_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_819 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet833_462 net433_94/I _6747_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_19_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet833_473 net833_473/I _6736_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet833_484 net833_499/I _6725_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet833_495 net833_499/I _6714_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4740_ _4706_/Z _4709_/Z _4825_/A4 _5489_/A1 _4748_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_1591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4671_ _4727_/A2 _4727_/A3 _4959_/C _5244_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_6410_ _6410_/A1 _6410_/A2 _6410_/A3 _6410_/A4 _6410_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_3622_ _3622_/A1 _3622_/A2 _3636_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_896 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6341_ _6341_/A1 _6341_/A2 _6341_/A3 _6341_/A4 _6342_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_155_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3553_ _3811_/A1 _3460_/B _3498_/B _5534_/A2 _3946_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_142_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3484_ _6863_/Q hold27/Z _3484_/B hold28/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_6272_ _6272_/I0 _7294_/Q _6559_/S _7294_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5223_ _5223_/A1 _5223_/A2 _5223_/B _5223_/C _5419_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5154_ _5439_/A2 _4725_/Z _5199_/A2 _5266_/A2 _5473_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_111_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4105_ _7282_/Q _6941_/Q _6944_/Q _4105_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5085_ _5085_/A1 _5418_/A1 _5085_/A3 _5088_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_96_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4036_ _5966_/I0 _6945_/Q _5911_/B _6787_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_793 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5987_ _5987_/A1 _5987_/A2 _7284_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4938_ _4951_/A1 _4951_/A2 _4951_/B1 _4951_/B2 _5007_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_12_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4869_ _4869_/A1 _5466_/B _4869_/A3 _5416_/A1 _4871_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_6608_ _6648_/A3 _6647_/A3 _6609_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6539_ _6766_/Q _6274_/Z _6568_/B1 _6738_/Q _6540_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_161_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput170 _4125_/Z irq[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput181 _3356_/ZN mgmt_gpio_oeb[19] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput192 _3346_/ZN mgmt_gpio_oeb[29] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_133_297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_896 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_789 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_153_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_43_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_183_186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_616 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5910_ hold2/Z hold47/Z _5910_/S hold48/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_81_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6890_ _6890_/D _7341_/RN _6890_/CLK _6890_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_62_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5841_ hold25/Z hold531/Z _5846_/S _5841_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5772_ hold5/Z hold230/Z _5774_/S _5772_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4723_ _4767_/A3 _4723_/A2 _4825_/A4 _5439_/A2 _5327_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_175_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4654_ _4437_/Z _5459_/A3 _5086_/A2 _5051_/B _5366_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
Xhold812 _5848_/Z _7210_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4585_ _4585_/A1 _4585_/A2 _5388_/A3 _4592_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xinput61 mgmt_gpio_in[32] input61/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput50 mgmt_gpio_in[22] input50/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold801 _6976_/Q hold801/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xinput72 mgmt_gpio_in[9] input72/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_7373_ _7373_/I _7373_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3605_ _7304_/Q _6943_/Q _6944_/Q _3605_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_171_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold834 _7016_/Q hold834/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3536_ _3454_/Z _3644_/A2 _4246_/A1 _3534_/C _4262_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_115_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6324_ _6324_/A1 _6325_/A1 _6325_/A2 _7278_/Q _6578_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xinput83 spimemio_flash_clk input83/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold845 _4284_/Z _6807_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xinput94 uart_enabled _4091_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold823 _4206_/Z _6760_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_143_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold867 _4270_/Z _6800_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold856 _7202_/Q hold856/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_89_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6255_ _6251_/Z _6255_/A2 _6255_/A3 _6255_/A4 _6268_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xhold889 _7326_/Q _3446_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold878 _6919_/Q hold878/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_170_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3467_ hold459/Z _6777_/Q _4011_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5206_ _5206_/A1 _5206_/A2 _5206_/A3 _4365_/C _5207_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_130_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6186_ hold72/I _6258_/B1 _6261_/B1 _7168_/Q _6187_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3398_ _6709_/Q _6708_/Q _6707_/Q _6774_/Q _4071_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_5137_ _5137_/A1 _5333_/A1 _5333_/A2 _5141_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_84_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5068_ _5079_/A1 _5180_/B _5285_/A1 _4597_/Z _5223_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_123_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4019_ _7283_/Q _6939_/Q _6944_/Q _4019_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_16_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold108 _5590_/Z _6983_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold119 _7069_/Q hold119/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4370_ hold807/Z hold391/Z _4371_/S _4370_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_112_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3321_ _6774_/Q _3421_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_152_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6040_ _6232_/C _7097_/Q _6211_/B _6211_/C _6041_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_435 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet433_90 net433_90/I _7179_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6942_ _6942_/D _7304_/RN _6942_/CLK _6942_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6873_ _6873_/D _7323_/RN _7322_/CLK _6873_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_81_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5824_ hold139/Z hold514/Z _5828_/S _5824_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_90_891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_711 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5755_ hold58/Z hold75/Z _5756_/S hold76/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5686_ hold139/Z hold178/Z hold42/Z _7067_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4706_ _4707_/A1 _4665_/Z _4750_/A3 _4960_/C _4706_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_175_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4637_ _5262_/A4 _5315_/A4 _4718_/B _4661_/C _5285_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_147_186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold620 _4253_/Z _6793_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4568_ _4481_/C _5048_/C _5062_/A3 _4568_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
X_7356_ _7356_/I _7356_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_150_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold631 _4301_/Z _6822_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold642 _4371_/Z _6867_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_2_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold653 _6771_/Q hold653/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4499_ _5051_/B _4454_/B _5330_/B2 _4959_/C _5045_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
Xhold664 _4274_/Z _6802_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3519_ _3608_/A4 _3482_/Z hold172/Z _3477_/Z _3519_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_6307_ _6307_/A1 _7276_/Q _7277_/Q _6580_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_103_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold675 _4238_/Z _6783_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold697 _6711_/Q hold697/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold686 _5768_/Z _7139_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7287_ _7287_/D _7304_/RN _7302_/CLK _7287_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6238_ _6738_/Q _6260_/B1 _6261_/A2 _6752_/Q _6240_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6169_ _6998_/Q _6258_/B1 _6259_/B1 _6982_/Q _6177_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_980 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_182_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_991 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_825 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet583_209 net433_87/I _7060_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_159_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_896 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_56__1374_ clkbuf_4_13_0__1374_/Z net683_324/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_48_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3870_ _7017_/Q _3946_/A2 _3938_/B1 _6884_/Q _3870_/C _3871_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_71_390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_176_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5540_ hold25/Z hold253/Z _5543_/S _5540_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5471_ _5471_/A1 _5199_/B _4722_/Z _5471_/B2 _5471_/C _5473_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_7210_ _7210_/D _7341_/RN _7210_/CLK _7210_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4422_ _4694_/B _4684_/B _5307_/B _5136_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_117_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_532 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4353_ _4358_/S _6859_/Q _4354_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7141_ _7141_/D _7262_/RN _7141_/CLK _7141_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_7072_ _7072_/D _7265_/RN _7072_/CLK _7072_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4284_ hold844/Z hold391/Z _4289_/S _4284_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6023_ _7210_/Q _6262_/A2 _6256_/B1 _7202_/Q _6025_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_99_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_0__1033_ _3715_/ZN clkbuf_0__1033_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_39_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6925_ _6925_/D input75/Z _6925_/CLK _6925_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_120_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6856_ _6856_/D _6862_/CLK _6856_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_167_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3999_ _3999_/I0 hold887/Z _4015_/S _6706_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6787_ _6787_/D _7302_/RN _7281_/CLK _6787_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_5807_ hold164/Z hold168/Z _5810_/S _5807_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_13_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5738_ hold687/Z hold388/Z _5744_/S _7113_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5669_ hold164/Z hold291/Z hold30/Z _7052_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold472 _7212_/Q hold472/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold450 _7181_/Q hold450/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold461 _3473_/C _3472_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_150_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7339_ _7339_/D _6693_/Z _7346_/CLK _7339_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold483 _7237_/Q hold483/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold494 _4391_/Z _6891_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_58_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2644 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1910 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2677 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1943 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1932 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1965 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1954 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1987 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1998 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_74 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4109__20 net433_84/I _7249_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_142_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4109__31 net433_91/I _7238_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_141_115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4109__42 _4109__48/I _7227_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_123_841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4971_ _4963_/B _5025_/A3 _4955_/B _5374_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_91_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3922_ _7178_/Q _5884_/A2 hold41/I _3527_/Z _3952_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6710_ _6710_/D _7304_/RN _6710_/CLK _6710_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_189_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6641_ _6641_/A1 _6641_/A2 _6642_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_149_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3853_ _3853_/A1 _3853_/A2 _3853_/A3 _3853_/A4 _3885_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_177_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6572_ _6572_/A1 _6572_/A2 _6572_/A3 _6577_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3784_ _3784_/A1 _3784_/A2 _3784_/A3 _3784_/A4 _3789_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_117_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5523_ hold164/Z hold537/Z _5524_/S _6931_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5454_ _5454_/A1 _5454_/A2 _5454_/B1 _5498_/A2 _5455_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_145_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5385_ _5385_/A1 _5038_/B _5291_/B _5123_/B _5476_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
X_4405_ _5535_/B _4405_/A2 _4405_/A3 _5784_/A3 _4407_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_160_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_874 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7124_ _7124_/D _7304_/RN _7124_/CLK _7124_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4336_ _3790_/Z _6847_/Q _4343_/S _6847_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7055_ hold31/Z _7265_/RN _7055_/CLK _7055_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4267_ hold754/Z hold391/Z _4281_/S _4267_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6006_ _7048_/Q _6256_/A2 _6258_/C1 _7064_/Q _6016_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4198_ hold388/Z hold713/Z _4198_/S _4198_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6908_ _6908_/D _7323_/RN _7322_/CLK hold27/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xnet633_290 net633_290/I _6979_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6839_ _6839_/D _7313_/CLK _6839_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold280 _6745_/Q hold280/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold291 _7052_/Q hold291/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_78_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2474 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1784 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1762 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_284 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5170_ _5330_/B2 _5466_/B _5295_/A1 _5170_/B1 _5186_/B2 _5171_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_110_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4121_ _4091_/S input68/Z _4121_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4052_ _4052_/A1 _7270_/Q _7269_/Q _6790_/Q _4053_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_56_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput4 mask_rev_in[0] input4/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_80_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_828 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4954_ _5372_/A1 _5454_/A2 _5454_/B1 _4437_/Z _5455_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3905_ _6893_/Q _5838_/A2 hold29/I _4405_/A2 _3951_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_178_866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4885_ _4423_/Z _5177_/A3 _5153_/B _5399_/B _4887_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6624_ _6878_/Q _6624_/A2 _6624_/B1 _6640_/B2 _6625_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3836_ _6834_/Q _5655_/A4 _4378_/A1 hold190/I _3879_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_20_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3767_ _6994_/Q _3953_/A2 _3946_/A2 _7018_/Q _3757_/Z _6947_/Q _3769_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_118_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6555_ _6555_/A1 _6555_/A2 _6555_/A3 _6558_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_5506_ hold45/Z _6653_/A2 hold37/Z _5655_/A4 _5508_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_106_616 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6486_ _7030_/Q _6562_/A2 _6562_/A3 _6562_/A4 _6505_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3698_ _3698_/A1 _3698_/A2 _3698_/A3 _3698_/A4 _3715_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5437_ _4718_/B _5484_/A2 _5439_/C _5437_/A4 _5438_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_105_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput330 _7309_/Q wb_dat_o[27] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput341 _6845_/Q wb_dat_o[8] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5368_ _5092_/B _5368_/A2 _5476_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5299_ _5466_/B _5466_/C _5466_/A2 _5299_/B _5300_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_4319_ _6594_/A1 _4328_/S _4319_/B _6835_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7107_ _7107_/D _7304_/RN _7107_/CLK _7107_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_7038_ _7038_/D _7281_/RN _7038_/CLK _7038_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_101_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1003 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1014 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1025 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1058 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1069 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet833_463 net433_98/I _6746_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet833_452 _4109__3/I _6757_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet833_474 net833_474/I _6735_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet833_485 net833_499/I _6724_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet833_496 net833_497/I _6713_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_18_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2293 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_820 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4670_ _4727_/A2 _4727_/A3 _4707_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_174_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3621_ _7030_/Q _3961_/B1 _3951_/B1 _7094_/Q _3622_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_30_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3552_ _3498_/B _3644_/A2 _5534_/A2 _3460_/B _4264_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_6340_ _7032_/Q _6294_/Z _6299_/Z _7064_/Q _6340_/C _6341_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_115_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3483_ hold172/Z _3482_/Z _3483_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_115_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6271_ _6788_/Q _6271_/A2 _6271_/A3 _6271_/B _6272_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_5222_ _5222_/A1 _5222_/A2 _5222_/A3 _5358_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_102_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5153_ _4423_/Z _5153_/A2 _5153_/B _5153_/C _5473_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_4104_ _6804_/Q input93/Z _6949_/Q _4104_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_111_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5084_ _5349_/A1 _5416_/A1 _5084_/B _5084_/C _5085_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_65_750 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4035_ _7268_/Q _6790_/Q _5985_/A2 _5918_/B _5911_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_53_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5986_ _5984_/S _7284_/Q _5987_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_4937_ _5426_/B1 _5369_/A2 _5454_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4868_ _4868_/A1 _5332_/A2 _4868_/A3 _4871_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6607_ _6648_/A3 _6607_/A2 _6651_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3819_ _6993_/Q _5727_/A3 _4378_/A1 _5748_/A3 _3840_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_20_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4799_ _3379_/I _5337_/A2 _5315_/A4 _4423_/Z _5469_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_20_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_839 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_180_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6538_ _6740_/Q _6311_/B _6567_/B1 _6760_/Q _6540_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_21_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6469_ _7143_/Q _6567_/B1 _6568_/B1 _7117_/Q _6469_/C _6474_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_133_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput171 _4101_/ZN mgmt_gpio_oeb[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput182 _4099_/ZN mgmt_gpio_oeb[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput193 _3373_/ZN mgmt_gpio_oeb[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_153_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_828 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_606 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_639 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_867 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5840_ hold388/Z hold729/Z _5846_/S _5840_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2090 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5771_ hold164/Z hold166/Z _5774_/S _5771_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_175_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4722_ _4767_/A3 _4723_/A2 _4825_/A4 _5439_/A2 _4722_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_4653_ _5459_/A3 _5086_/A2 _5355_/A2 _5051_/B _4658_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_147_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput40 mgmt_gpio_in[13] input40/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput62 mgmt_gpio_in[33] input62/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_7372_ _7372_/I _7372_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_571 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput51 mgmt_gpio_in[23] input51/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3604_ _5573_/A3 _3604_/A2 _5546_/A2 hold462/Z _5544_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
X_4584_ _5439_/A1 _4759_/C _4421_/Z _5177_/A3 _5388_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
Xhold802 _5583_/Z _6976_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xinput73 pad_flash_io0_di input73/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput95 wb_adr_i[0] input95/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
Xhold835 _5628_/Z _7016_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold813 _7146_/Q hold813/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6323_ _6323_/A1 _6325_/A1 _6325_/A2 _7279_/Q _6567_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_116_766 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3535_ _3460_/B _3498_/B _4246_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xinput84 spimemio_flash_csb input84/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold846 _6937_/Q hold846/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold824 _6740_/Q hold824/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3466_ _3491_/B hold40/Z _3466_/B _3604_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_116_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold857 _5839_/Z _7202_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6254_ _6763_/Q _6260_/A2 _6256_/B1 _6759_/Q _6255_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold868 _6791_/Q hold868/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold879 _6913_/Q hold879/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_5205_ _5323_/A1 _5404_/B1 _5205_/B _5323_/C _5206_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_131_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3397_ _4016_/A2 _4015_/S _3397_/B _7347_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6185_ _7200_/Q _6260_/A2 _6257_/A2 _7136_/Q _6187_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_97_650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5136_ _4922_/B _5136_/A2 _5330_/B1 _5136_/B1 _5330_/A2 _5333_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_85_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5067_ _5372_/A1 _4597_/Z _5067_/B _5067_/C _5071_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_45_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4018_ _4018_/A1 _4018_/A2 _6700_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_84_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5969_ _6789_/Q _6562_/A3 _6324_/A1 _7278_/Q _5971_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_25_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_2_0__1374_ clkbuf_0__1374_/Z clkbuf_4_5_0__1374_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_57_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_184_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_16__1374_ clkbuf_4_10_0__1374_/Z _4109__34/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_129_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_79__1374_ net583_226/I net533_176/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xhold109 _7183_/Q hold109/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_160_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3320_ _6776_/Q _4119_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_113_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_403 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_577 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet433_80 net433_82/I _7189_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_82_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6941_ _6941_/D _7304_/RN _6941_/CLK _6941_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_19_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6872_ _6872_/D _7323_/RN _7323_/CLK _6872_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xnet433_91 net433_91/I _7178_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5823_ hold25/Z hold456/Z _5828_/S _5823_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_167_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5754_ hold5/Z hold91/Z _5756_/S hold92/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5685_ hold25/Z hold474/Z hold42/Z _7066_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_147_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4705_ _5262_/A4 _3380_/I _4718_/B _5253_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_4636_ _5301_/A2 input95/Z _5004_/A1 _5005_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_135_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7355_ _7355_/I _7355_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold610 _4380_/Z _6884_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold621 _7351_/I hold621/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4567_ _5045_/A2 _5436_/A4 _4567_/B _4576_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_162_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6306_ _6307_/A1 _7277_/Q _6306_/A3 _6581_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
Xmax_cap362 _5884_/A2 _5727_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xhold643 _6869_/Q hold643/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold632 _6920_/Q hold632/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold654 _4222_/Z _6771_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4498_ _4469_/B _5312_/B _4684_/B _4922_/B _5330_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_131_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3518_ _3608_/A4 _3482_/Z hold172/Z _3477_/Z _5532_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_104_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold676 _6977_/Q hold676/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7286_ _7286_/D _7304_/RN _7302_/CLK _7286_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold687 _7113_/Q hold687/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold665 _7033_/Q hold665/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_134_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6237_ _6211_/B _6266_/B _6768_/Q _7274_/Q _6240_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xhold698 _4138_/Z _6711_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3449_ _3449_/A1 _4073_/B2 _4119_/B _7324_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_97_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6168_ _6168_/I0 _7290_/Q _6559_/S _7290_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_970 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5119_ _3379_/I _3380_/I _5445_/A2 _5476_/A2 _5287_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_58_867 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_981 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6099_ _6745_/Q _6266_/C _6232_/B1 _7149_/Q _6232_/C _6102_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_58_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_848 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_399 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_845 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_3__1374_ clkbuf_4_2_0__1374_/Z _4109__16/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_75_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_189_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_189_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5470_ _5470_/A1 _5338_/Z _5470_/A3 _5469_/Z _5470_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_4421_ _4694_/B _4684_/B _5307_/B _4421_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_157_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7140_ _7140_/D _7302_/RN _7140_/CLK _7140_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4352_ _6597_/I0 _6858_/Q _4358_/S _6858_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7071_ hold43/Z _7265_/RN _7071_/CLK _7071_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_152_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4283_ _5838_/A4 _5518_/A1 _5838_/A2 hold37/Z _4289_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6022_ _7194_/Q _6260_/A2 _6258_/C1 _7186_/Q _6025_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_100_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6924_ _6924_/D _7262_/RN _6924_/CLK _6924_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_35_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6855_ _6855_/D _6862_/CLK _6855_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3998_ _3489_/Z _3997_/B _3998_/B _3999_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6786_ _6786_/D input75/Z _6786_/CLK _7364_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5806_ hold139/Z _7173_/Q _5810_/S _5806_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_183_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5737_ hold779/Z hold391/Z _5744_/S _7112_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_175_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5668_ hold139/Z hold363/Z hold30/Z _7051_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_62__1374_ clkbuf_4_13_0__1374_/Z _4109__14/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4619_ _4628_/B _5046_/C _5078_/A2 _5186_/B2 _4620_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_5599_ hold124/Z hold2/Z _5599_/S _5599_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_2_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold440 _7058_/Q hold440/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold451 _5815_/Z _7181_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_163_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold462 _3507_/C hold462/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7338_ _7338_/D _6692_/Z _7346_/CLK _7338_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold473 _5850_/Z _7212_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold484 _7134_/Q hold484/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold495 _6811_/Q hold495/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7269_ _7269_/D _7302_/RN _7304_/CLK _7269_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_132_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xnet683_350 net433_74/I _6911_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_57_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2612 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2678 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1911 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1977 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1966 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1944 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1999 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4109__10 _4109__48/I _7259_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4109__32 _4109__34/I _7237_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_181_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4109__21 _4109__4/I _7248_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4109__43 _4109__48/I _7226_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_126_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4970_ _4437_/Z _5454_/A2 _5106_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_189_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3921_ _6949_/Q _5902_/A3 _5548_/A3 hold173/I _3976_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_32_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6640_ _6878_/Q _6640_/A2 _6640_/B1 _6640_/B2 _6641_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_149_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3852_ _7113_/Q _3969_/A2 _3959_/B1 _6753_/Q _3853_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6571_ _6892_/Q _6292_/Z _6571_/B1 _6834_/Q _6571_/C1 _6771_/Q _6572_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_81_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5522_ hold139/Z hold468/Z _5524_/S _6930_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3783_ _7114_/Q _3969_/A2 _3969_/B1 _6744_/Q _3784_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_157_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_4_5_0__1374_ clkbuf_4_5_0__1374_/I clkbuf_4_5_0__1374_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_5453_ _5453_/A1 _5453_/A2 _5453_/A3 _5456_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_145_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5384_ _5385_/A1 _5038_/B _5291_/B _5123_/B _5433_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_114_820 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4404_ hold388/Z _6900_/Q _4404_/S _4404_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_132_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7123_ _7123_/D _7262_/RN _7123_/CLK _7123_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4335_ _6595_/I0 _6846_/Q _4343_/S _6846_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_114_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_726 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7054_ _7054_/D _7265_/RN _7054_/CLK hold67/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4266_ _4266_/A1 _4227_/B _4282_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_86_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6005_ _6211_/C _6211_/B _7272_/Q _7271_/Q _6258_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_67_461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4197_ hold391/Z hold818/Z _4198_/S _4197_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_28_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_881 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6907_ _6907_/D _7323_/RN _7322_/CLK _6907_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xnet633_280 net633_280/I _6989_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet633_291 net633_292/I _6978_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_42_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6838_ _6838_/D _7313_/CLK _6838_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6769_ _6769_/D _7262_/RN _6769_/CLK _6769_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_148_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xhold270 _4302_/Z _6823_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_172_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold281 _4185_/Z _6745_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold292 _6713_/Q hold292/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_120_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2431 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2464 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2497 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1796 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4120_ _3888_/S _4120_/A2 _7325_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4051_ _4044_/Z _4051_/A2 _4051_/B _6789_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_96_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput5 mask_rev_in[10] input5/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_92_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4953_ _4963_/B _4953_/A2 _5454_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_91_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_823 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3904_ input34/Z _5856_/A1 _5748_/A3 _5532_/A3 _3970_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_33_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6623_ _6880_/Q _6623_/A2 _6623_/B1 _6879_/Q _6625_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4884_ _5177_/A3 _5153_/A2 _5153_/B _5439_/B _4887_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_178_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3835_ _6892_/Q hold41/I hold29/I _6653_/A2 _3879_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_20_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3766_ _3766_/A1 _3766_/A2 _3766_/A3 _3766_/A4 _3766_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_6554_ _6584_/A1 _6554_/A2 _6554_/A3 _6553_/Z _6555_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6485_ hold95/I _6563_/A2 _6562_/A3 _6563_/A4 _6491_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5505_ _5505_/A1 _5505_/A2 _5505_/B _5505_/C _6909_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_161_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5436_ _5436_/A1 _5436_/A2 _5439_/C _5436_/A4 _5438_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_10_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3697_ _6939_/Q _5544_/S _3643_/Z _6931_/Q _3697_/C _3698_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_160_222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput331 _7310_/Q wb_dat_o[28] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput320 _6837_/Q wb_dat_o[18] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput342 _6846_/Q wb_dat_o[9] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5367_ _5367_/A1 _5367_/A2 _5367_/B _5408_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_120_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5298_ _5436_/A4 _5471_/A1 _5468_/A1 _5298_/B _5299_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_4318_ _4328_/S _6835_/Q _4319_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7106_ _7106_/D _7304_/RN _7106_/CLK _7106_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_102_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_867 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7037_ _7037_/D _7281_/RN _7037_/CLK _7037_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4249_ hold868/Z _4248_/Z _4263_/S _4249_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_19_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1004 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1015 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1026 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1037 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1059 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1048 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_143_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet833_453 _4109__7/I _6756_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_74_773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet833_475 _4109__3/I _6734_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet833_464 net833_464/I _6745_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet833_486 net833_489/I _6723_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet833_497 net833_497/I _6712_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_178_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1571 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_865 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3620_ hold89/I _3951_/A2 _3981_/B1 _7256_/Q _3622_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3551_ _5534_/A1 _3477_/Z _3496_/B _4246_/A1 _3956_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_143_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_797 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3482_ _6863_/Q hold27/Z _3482_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_115_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6270_ _6788_/Q _7293_/Q _6271_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5221_ _3380_/I _4425_/Z _4956_/C _5493_/B1 _5222_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_102_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5152_ _5369_/A2 _5258_/A3 _5152_/B _5152_/C _5239_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_69_545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4103_ _6805_/Q _4103_/I1 _6947_/Q _4103_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_111_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5083_ _5087_/A1 _5394_/A2 _5194_/B _5457_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_110_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4034_ _7269_/Q _7270_/Q _5985_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5985_ _7267_/Q _5985_/A2 _5985_/A3 _6790_/Q _5987_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XPHY_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_4936_ _4628_/B _5347_/A1 _5369_/A1 _4947_/C _5020_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_33_681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4867_ _5502_/B2 _5177_/A3 _5153_/A2 _5153_/B _4868_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_21_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6606_ _6880_/Q _6606_/A2 _6606_/B1 _6878_/Q _6610_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_3818_ _6900_/Q hold37/I hold41/I hold190/I _3883_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_181_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6537_ _6734_/Q _6285_/Z _6294_/Z _6881_/Q _6564_/C1 _6893_/Q _6540_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_4798_ _3379_/I _5337_/A2 _5315_/A4 _5153_/A2 _5263_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_146_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3749_ _7075_/Q _3951_/A2 _3981_/A2 _7245_/Q _7253_/Q _3981_/B1 _3750_/A4 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_118_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6468_ _6465_/Z _6468_/A2 _6468_/A3 _6468_/A4 _6468_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_106_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5419_ _4608_/Z _5459_/A1 _5419_/B _5419_/C _5462_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_6399_ _6788_/Q _7296_/Q _6400_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput194 _3345_/ZN mgmt_gpio_oeb[30] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_133_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput172 _3365_/ZN mgmt_gpio_oeb[10] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput183 _3355_/ZN mgmt_gpio_oeb[20] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_153_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_39__1374_ clkbuf_4_14_0__1374_/Z net433_84/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_46_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2091 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5770_ hold139/Z hold466/Z _5774_/S _7141_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4721_ _5468_/C _4765_/A2 _4765_/A1 _5312_/B _4819_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XTAP_1390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4652_ _5301_/A2 _4661_/C _3379_/I _3380_/I _5353_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_175_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput30 mask_rev_in[4] input30/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3603_ hold68/I _5856_/A1 _5802_/A2 _3527_/Z _3619_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4583_ _4443_/Z _5459_/A3 _5360_/B _4598_/A4 _5355_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
Xinput63 mgmt_gpio_in[34] input63/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput41 mgmt_gpio_in[14] input41/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_7371_ _7371_/I _7371_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput52 mgmt_gpio_in[24] input52/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold803 _7032_/Q hold803/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xinput96 wb_adr_i[10] input96/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_171_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold814 _7187_/Q hold814/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3534_ _6863_/Q hold16/Z _3534_/B _3534_/C hold190/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_6322_ _6984_/Q _6511_/A2 _6563_/A4 _6562_/A4 _6345_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xinput85 spimemio_flash_io0_do input85/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput74 pad_flash_io1_di _3339_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold836 _6718_/Q hold836/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold825 _4179_/Z _6740_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3465_ hold12/Z _3511_/B2 _6863_/Q _5326_/B2 _3473_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_143_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6253_ _6757_/Q _6257_/A2 _6256_/A2 _6773_/Q _6255_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold869 _4249_/Z _6791_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold847 _5533_/Z _6937_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold858 _7040_/Q hold858/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_5204_ _5262_/A4 _5204_/A2 _5204_/B1 _5445_/A3 _5204_/C _5205_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_115_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3396_ input58/Z _6777_/Q _4015_/S _3396_/C _3397_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_130_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6184_ hold62/I _6260_/B1 _6256_/B1 _7208_/Q _6187_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_96_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5135_ _5466_/B _5170_/B1 _5258_/A3 _5136_/B1 _5369_/A2 _5333_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_85_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5066_ _5347_/A1 _5435_/A1 _5503_/A1 _5223_/A2 _5369_/A1 _5358_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_111_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4017_ _4073_/B1 _6774_/Q _4017_/B _4018_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_72_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5968_ _5968_/I _7278_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4919_ _4425_/Z _5210_/B _4919_/B _4926_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_138_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5899_ hold5/Z hold212/Z _5901_/S _7255_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_165_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_839 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_188_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_829 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_426 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6940_ _6940_/D _7304_/RN _6940_/CLK _6940_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xnet433_70 net433_84/I _7199_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet433_81 net433_81/I _7188_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_19_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6871_ _6871_/D _7323_/RN _7323_/CLK _6877_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_179_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet433_92 net433_94/I _7177_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_179_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5822_ hold388/Z hold814/Z _5828_/S _5822_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5753_ hold164/Z _7126_/Q _5756_/S _5753_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4704_ _5315_/A4 _3379_/I _4718_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_5684_ hold388/Z hold750/Z hold42/Z _7065_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_147_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4635_ _5262_/A4 _5315_/A4 _4718_/B _4956_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_136_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4566_ _4661_/C _5436_/A1 _5436_/A2 _5436_/A4 _5215_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xhold611 _7163_/Q hold611/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7354_ _7354_/I _7354_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold600 _6895_/Q hold600/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_118_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6305_ _7278_/Q _6563_/A3 _6562_/A4 _6324_/A1 _6311_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold644 _4374_/Z _6869_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold622 _4255_/Z _6794_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold633 _5510_/Z _6920_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3517_ _5534_/A1 _3477_/Z _3496_/B _5534_/A2 _3958_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xmax_cap374 input95/Z _3380_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
XFILLER_144_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4497_ _4759_/C _4686_/B _5307_/B _4694_/B _5394_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xhold677 _5584_/Z _6977_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold688 _6832_/Q hold688/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7285_ _7285_/D _7304_/RN _7302_/CLK _7285_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold655 _6763_/Q hold655/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold666 _5648_/Z _7033_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6236_ _6772_/Q _6256_/A2 _6259_/B1 _6734_/Q _6257_/B1 _6770_/Q _6240_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
Xhold699 _6743_/Q hold699/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3448_ _7339_/Q hold44/Z _3449_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3379_ _3379_/I _5262_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_20
XFILLER_134_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_470 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6167_ _6788_/Q _6167_/A2 _6167_/A3 _6167_/B _6168_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XTAP_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_971 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5118_ _5118_/A1 _5118_/A2 _5285_/C _5120_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_84_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_982 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6098_ _6098_/I _6112_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_27_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5049_ _5351_/A1 _4956_/B _5346_/A4 _5235_/A1 _5053_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xclkbuf_leaf_102__1374_ clkbuf_4_1_0__1374_/Z net833_489/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_26_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_85__1374_ clkbuf_4_4_0__1374_/Z net433_98/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_25_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_835 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_356 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_790 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4420_ _4684_/B _5307_/B _4690_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_144_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4351_ _3790_/Z _6857_/Q _4358_/S _6857_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7070_ _7070_/D _7265_/RN _7070_/CLK hold82/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4282_ _4281_/Z hold523/Z _4282_/S _4282_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6021_ _7130_/Q _6257_/A2 _6259_/B1 _7104_/Q _6025_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_104_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_816 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6923_ _6923_/D _7262_/RN _6923_/CLK _6923_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_54_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6854_ _6854_/D _7341_/RN _6854_/CLK _6854_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3997_ _3489_/Z _3490_/Z _3997_/B _3998_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_10_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5805_ hold25/Z hold327/Z _5810_/S _5805_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6785_ _6785_/D input75/Z _6785_/CLK _7363_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_176_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5736_ _5856_/A1 _5802_/A2 _5784_/A2 _5535_/B _5744_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_5667_ hold25/Z hold354/Z hold30/Z _7050_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_175_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4618_ _4686_/B _5223_/A1 _5048_/B _4628_/B _5076_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_108_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5598_ hold210/Z hold58/Z _5599_/S _5598_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold441 _7213_/Q hold441/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold452 _7148_/Q hold452/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_144_681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold463 hold463/I hold463/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_89_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4549_ _5315_/A4 _5301_/A2 _5235_/A1 _3379_/I _5439_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xhold430 _4164_/Z _6729_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7337_ _7337_/D _6691_/Z _4111_/I1 _7337_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold474 _7066_/Q hold474/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold496 _4288_/Z _6811_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold485 _7206_/Q hold485/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7268_ _7268_/D _7302_/RN _7304_/CLK _7268_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6219_ _5917_/B _6587_/A2 _7292_/Q _6220_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_7199_ _7199_/D _7265_/RN _7199_/CLK _7199_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_58_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet683_340 net833_483/I _6929_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_38_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet683_351 _4109__24/I _6910_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_100_762 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_790 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2679 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1934 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1923 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1912 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1967 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1956 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1945 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1989 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1978 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4109__11 net433_91/I _7258_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_119_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4109__33 net433_87/I _7236_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_181_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4109__22 net433_53/I _7247_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4109__44 _4109__44/I _7225_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_5_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3920_ _6853_/Q _4378_/A1 hold41/I _4405_/A2 _3952_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_91_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_874 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3851_ _7139_/Q _3958_/A2 _3851_/B1 _6771_/Q _3853_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6570_ _6755_/Q _6570_/A2 _6570_/B1 _6888_/Q _6570_/C1 _6844_/Q _6572_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_20_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3782_ _7172_/Q _3966_/A2 _3968_/A2 _7106_/Q _3784_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_185_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5521_ hold25/Z hold279/Z _5524_/S _6929_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_172_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5452_ _5452_/A1 _5452_/A2 _5452_/A3 _5453_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_173_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5383_ _5038_/B _5291_/B _5123_/B _5386_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_4403_ hold391/Z hold522/Z _4404_/S _6899_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7122_ _7122_/D _7302_/RN _7122_/CLK _7122_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4334_ _6594_/A1 _4343_/S _4334_/B _6845_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7053_ _7053_/D _7265_/RN _7053_/CLK _7053_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_113_375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4265_ _5640_/A2 _5564_/A3 _4265_/B _4266_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_6004_ _6036_/A3 _6211_/C _7273_/Q _7271_/Q _6256_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_101_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4196_ _6653_/A2 _5535_/B _3527_/Z _5838_/A2 _4198_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_67_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet633_270 net683_320/I _6999_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_70_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6906_ _6906_/D _7323_/RN _7322_/CLK hold7/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xnet633_281 net633_281/I _6988_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_82_498 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xnet633_292 net633_292/I _6977_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6837_ _6837_/D _7313_/CLK _6837_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6768_ _6768_/D _7262_/RN _6768_/CLK _6768_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_176_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6699_ _7341_/RN _6994_/Q _4026_/C _6699_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_5719_ hold391/Z hold719/Z hold22/Z _7096_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_163_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold260 _5614_/Z _7004_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold271 _7157_/Q hold271/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_132_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_898 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold293 _4142_/Z _6713_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_2_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold282 _6972_/Q hold282/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_172_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2498 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1797 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1786 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_167_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4050_ _6310_/A4 _6307_/A1 _7276_/Q _4051_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_84_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput6 mask_rev_in[11] input6/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_64_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4952_ _4952_/A1 _4926_/B _4995_/A4 _4953_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3903_ _6758_/Q _5902_/A3 _3527_/Z _4405_/A2 _3952_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4883_ _4883_/A1 _4883_/A2 _4887_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_32_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6622_ _6622_/I0 _7316_/Q _6642_/S _7316_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_60_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3834_ _6755_/Q _5838_/A2 _5546_/A2 _3527_/Z _3865_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_20_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3765_ _7236_/Q _3943_/A2 _3875_/A2 _7180_/Q _3766_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6553_ _6553_/A1 _6553_/A2 _6553_/A3 _6553_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_145_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5504_ _5504_/A1 _5504_/A2 _5486_/Z _5504_/A4 _5505_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_3696_ _3696_/I _3697_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6484_ _6788_/Q _4019_/Z _6509_/B _7301_/Q _6508_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_145_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5435_ _5435_/A1 _5435_/A2 _5435_/B _5443_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput310 _7305_/Q wb_ack_o VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_160_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput332 _7311_/Q wb_dat_o[29] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput321 _6838_/Q wb_dat_o[19] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5366_ _5366_/A1 _5457_/A2 _5366_/A3 _5366_/A4 _5367_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_114_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4317_ _6875_/Q _7323_/RN _4328_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_5297_ _4690_/C _5466_/B _5290_/C _3379_/I _5390_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_59_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7105_ _7105_/D _7304_/RN _7105_/CLK _7105_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4248_ hold700/Z hold391/Z _4262_/S _4248_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7036_ _7036_/D _7302_/RN _7036_/CLK _7036_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_142_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4179_ hold391/Z hold824/Z _4180_/S _4179_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_82_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1005 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1016 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1038 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1049 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet833_454 net833_454/I _6755_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet833_476 net833_491/I _6733_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet833_487 net833_489/I _6722_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet833_465 net433_97/I _6744_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_34_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet833_498 net833_498/I _6711_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2284 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_187_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3550_ _7111_/Q _5802_/A2 _5784_/A2 _5727_/A3 _3586_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_182_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5220_ _5220_/A1 _5356_/A2 _5219_/Z _5224_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3481_ hold171/Z _3481_/A2 _6863_/Q _3484_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_142_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_833 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5151_ _5151_/A1 _5469_/A4 _5469_/A3 _5156_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_69_535 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4102_ _6806_/Q user_clock _6948_/Q _4102_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5082_ _5082_/A1 _5082_/A2 _5082_/B1 _5082_/B2 _5082_/C _5362_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_110_142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4033_ _5918_/B _7268_/Q _4052_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5984_ _6532_/B _7283_/Q _5984_/S _7283_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4935_ _5051_/B _5051_/C _5369_/A1 _5288_/A4 _5074_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_178_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4866_ _4421_/Z _5177_/A3 _5468_/A1 _4759_/C _5332_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_60_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6605_ _6648_/A3 _6646_/A3 _6606_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4797_ _4661_/C _5253_/A1 _5337_/A2 _5263_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3817_ _6759_/Q _5838_/A2 _3527_/Z _4405_/A2 _3871_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3748_ _7237_/Q _3943_/A2 _3950_/A2 _7099_/Q _3750_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6536_ _6868_/Q _6562_/A2 _6562_/A3 _6562_/A4 _6554_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_20_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6467_ _7077_/Q _6292_/Z _6571_/B1 _6989_/Q _6571_/C1 _7183_/Q _6468_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_3679_ _6916_/Q _6600_/I0 _3887_/S _3679_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5418_ _5418_/A1 _5418_/A2 _5418_/A3 _5458_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_6398_ _6584_/A1 _6970_/Q _6584_/B _6400_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5349_ _5349_/A1 _5353_/A3 _5459_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput195 _3344_/ZN mgmt_gpio_oeb[31] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput173 _3364_/ZN mgmt_gpio_oeb[11] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput184 _3354_/ZN mgmt_gpio_oeb[21] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7019_ _7019_/D _7265_/RN _7019_/CLK _7019_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_46_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_877 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_608 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2070 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2092 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2081 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4720_ _5152_/C _4720_/A2 _4720_/A3 _5307_/B _5264_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XTAP_1391 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4651_ _5262_/A4 _5315_/A4 _5235_/A1 _4718_/B _5355_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_148_827 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput20 mask_rev_in[24] input20/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput31 mask_rev_in[5] input31/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3602_ input18/Z _5748_/A3 _5532_/A3 _5528_/A2 _3616_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xinput64 mgmt_gpio_in[35] input64/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4582_ _5062_/A3 _5502_/A1 _4598_/A4 _4481_/C _4585_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_162_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput42 mgmt_gpio_in[15] input42/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_7370_ _7370_/I _7370_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput53 mgmt_gpio_in[25] input53/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xinput97 wb_adr_i[11] input97/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xhold815 _5822_/Z _7187_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6321_ _6324_/A1 _6325_/A2 _7278_/Q _6321_/A4 _6571_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_116_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput86 spimemio_flash_io0_oeb input86/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold826 _6843_/Q hold826/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold804 _5647_/Z _7032_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xinput75 porb input75/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_16
Xhold837 _4152_/Z _6718_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3533_ _5534_/A1 _3827_/A1 _3827_/A2 _3496_/B _3966_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xhold859 _7056_/Q hold859/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3464_ _3511_/B2 hold12/Z _3466_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6252_ _6739_/Q _6260_/B1 _6262_/B1 _6765_/Q _7341_/Q _6261_/B1 _6255_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
Xhold848 _6928_/Q hold848/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_5203_ _5200_/B _4718_/B _3379_/I _5235_/A1 _5204_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_6183_ hold77/I _6262_/B1 _6257_/B1 hold78/I _6187_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3395_ _7347_/Q _6777_/Q _3396_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_97_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5134_ _5134_/A1 _5134_/A2 _5428_/A4 _5137_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_97_674 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5065_ _5061_/Z _5494_/A1 _5222_/A1 _5067_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_85_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4016_ _4016_/A1 _4016_/A2 _6774_/Q _4018_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_16_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5967_ _5966_/Z _7278_/Q _6789_/Q _5967_/B2 _5968_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_166_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4918_ _4690_/B _4661_/C _4718_/B _3379_/I _4919_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_5898_ hold164/Z hold517/Z _5901_/S _7254_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4849_ _5466_/B _4849_/A2 _4853_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6519_ _7111_/Q _6285_/Z _6294_/Z hold85/I _6564_/C1 _7087_/Q _6523_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
Xclkbuf_leaf_45__1374_ clkbuf_4_15_0__1374_/Z net783_415/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_122_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_790 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_674 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet433_71 net433_71/I _7198_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_93_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet433_60 net433_65/I _7209_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6870_ _6870_/D _7323_/RN _7323_/CLK _6870_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
Xnet433_82 net433_82/I _7187_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet433_93 net433_93/I _7176_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_179_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5821_ hold391/Z hold809/Z _5828_/S _5821_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5752_ hold139/Z hold267/Z _5756_/S _5752_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4703_ _5416_/A1 _4830_/B2 _6880_/Q _5202_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5683_ hold391/Z hold855/Z hold42/Z _7064_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_175_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4634_ _4661_/C _5439_/C _5436_/A4 _5321_/A3 _5230_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_163_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4565_ _4565_/A1 _4565_/A2 _4565_/A3 _4565_/A4 _4567_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_116_510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold612 _6883_/Q hold612/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold601 _4397_/Z _6895_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7353_ _7353_/I _7353_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3516_ _3507_/C _3833_/A2 _3802_/A2 _3473_/B _3951_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_128_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6304_ _6324_/A1 _6308_/A3 _7278_/Q _6325_/A1 _6575_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xhold634 _7024_/Q hold634/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold623 _6969_/Q hold623/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold645 _6759_/Q hold645/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_171_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xmax_cap375 _7341_/RN _7265_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
X_4496_ _4469_/B _4922_/B _5294_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_103_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold678 _6921_/Q hold678/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7284_ _7284_/D _7304_/RN _7304_/CLK _7284_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold656 _4210_/Z _6763_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold667 _7362_/I hold667/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6235_ _6235_/A1 _6235_/A2 _6235_/B1 _6235_/B2 _6235_/C _6241_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_3447_ _6707_/Q _3447_/A2 _3447_/B _7326_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold689 _4313_/Z _6832_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3378_ _7273_/Q _6211_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XFILLER_57_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_961 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_950 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6166_ _6788_/Q _7289_/Q _6167_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5117_ _5117_/A1 _5452_/A1 _5118_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6097_ _7027_/Q _6262_/B1 _7275_/Q _6098_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_972 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_983 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_994 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5048_ _4686_/B _5223_/A1 _5048_/B _5048_/C _5346_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_58_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6999_ _6999_/D _7281_/RN _6999_/CLK _6999_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_154_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_844 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_293 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4350_ _6595_/I0 _6856_/Q _4358_/S _6856_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_125_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4281_ _6967_/Q hold2/Z _4281_/S _4281_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_140_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_91__1374_ net583_226/I _4109__49/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_141_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6020_ _6020_/A1 _6020_/A2 _6020_/A3 _6026_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_67_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6922_ _6922_/D _7262_/RN _6922_/CLK _6922_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_120_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6853_ _6853_/D _7341_/RN _6853_/CLK _6853_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_23_714 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5804_ hold388/Z hold695/Z _5810_/S _5804_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3996_ _6705_/Q _6704_/Q _6703_/Q _3993_/Z _3997_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6784_ _6784_/D input75/Z _6784_/CLK _7362_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5735_ hold2/Z hold128/Z _5735_/S _5735_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5666_ hold388/Z hold585/Z hold30/Z _7049_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4617_ _5082_/C _5435_/A1 _4454_/B _5426_/A1 _4620_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_135_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5597_ hold377/Z hold5/Z _5599_/S _5597_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold420 _6721_/Q hold420/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold442 _5851_/Z _7213_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold453 _7196_/Q hold453/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold431 _7238_/Q hold431/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_89_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4548_ _5262_/A4 _3380_/I _5392_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_7336_ _7336_/D _6690_/Z _7346_/CLK _7336_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4479_ _4951_/A2 _4479_/A2 _4479_/B _4479_/C _5360_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_145_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold464 hold464/I _5861_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold475 _7373_/I hold475/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7267_ _7267_/D _7304_/RN _7302_/CLK _7267_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold486 _5843_/Z _7206_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold497 _7132_/Q hold497/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_568 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6218_ _6218_/A1 _6218_/A2 _6788_/Q _7291_/Q _6220_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7198_ _7198_/D _7265_/RN _7198_/CLK _7198_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_131_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet683_330 net783_421/I _6939_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_161_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6149_ _7135_/Q _6257_/A2 _6260_/B1 _7117_/Q _6151_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xnet683_341 net683_349/I _6928_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1924 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1913 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1902 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1946 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1935 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1979 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_711 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4109__34 _4109__34/I _7235_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_135_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4109__23 _4109__24/I _7246_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4109__12 _4109__12/I _7257_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_134_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4109__45 net433_77/I _7224_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_122_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_189_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3850_ _7025_/Q _3961_/B1 _3850_/B1 input35/Z _3969_/B1 _6743_/Q _3853_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_158_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3781_ _7156_/Q _3956_/B1 _3971_/A2 input13/Z _3559_/Z _6970_/Q _3784_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_118_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5520_ hold388/Z hold848/Z _5524_/S _6928_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_158_796 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5451_ _5451_/A1 _5498_/B1 _5452_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5382_ _5382_/A1 _5382_/A2 _5433_/A1 _5386_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4402_ hold45/Z hold190/Z hold41/Z hold37/Z _4404_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_141_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7121_ _7121_/D _7262_/RN _7121_/CLK _7121_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4333_ _4343_/S _6845_/Q _4334_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7052_ _7052_/D _7265_/RN _7052_/CLK _7052_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4264_ _4264_/A1 _5564_/A3 hold37/Z _5640_/A2 _4265_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_113_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6003_ _6003_/A1 _6003_/A2 _6003_/A3 _6026_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_83_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4195_ hold388/Z hold692/Z _4195_/S _6753_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6905_ _6905_/D _7323_/RN _7322_/CLK hold40/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xnet633_260 net633_282/I _7009_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet633_271 net633_271/I _6998_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet633_293 net683_324/I _6976_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet633_282 net633_282/I _6987_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6836_ _6836_/D _6862_/CLK _6836_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_24_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6767_ _6767_/D _7262_/RN _6767_/CLK _6767_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5718_ hold21/Z hold13/Z _5718_/A3 hold45/I hold22/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_3979_ _3979_/A1 _3979_/A2 _3979_/A3 _3979_/A4 _3983_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_164_711 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6698_ input75/Z _6994_/Q _4026_/C _6698_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_164_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5649_ hold25/Z hold534/Z _5654_/S _5649_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7319_ _7319_/D _7323_/RN _4103_/I1 _7319_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_104_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold250 _5613_/Z _7003_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_2_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold261 _7107_/Q hold261/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold294 _7060_/Q hold294/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold283 _7166_/Q hold283/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold272 _5788_/Z _7157_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_172_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2466 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1710 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_836 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1754 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_853 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput7 mask_rev_in[12] input7/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_49_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4951_ _4951_/A1 _4951_/A2 _4951_/B1 _4951_/B2 _4951_/C _4956_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_36_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_825 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4882_ _5466_/B _5037_/A1 _5392_/A1 _5426_/A1 _4883_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_3902_ _6868_/Q _4378_/A1 _5838_/A2 _5546_/A2 _3941_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_60_650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_864 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6621_ _6621_/A1 _6621_/A2 _6622_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3833_ _3507_/C _3833_/A2 _3519_/Z _3473_/B _3948_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_177_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_571 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3764_ _7164_/Q _3878_/A2 _3950_/A2 _7098_/Q _3943_/B1 _7196_/Q _3766_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6552_ _6853_/Q _6311_/C _6309_/Z _6736_/Q _6553_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_9_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5503_ _5503_/A1 _5503_/A2 _5503_/B _5504_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3695_ _7108_/Q _3968_/A2 _3681_/Z _6926_/Q _3969_/B1 _6746_/Q _3696_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6483_ _6483_/A1 _6483_/A2 _6483_/B _7300_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5434_ _4437_/Z _5436_/A1 _5210_/C _5194_/C _5479_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xoutput300 _4019_/Z serial_clock VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput322 _6856_/Q wb_dat_o[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput311 _6855_/Q wb_dat_o[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput333 _6857_/Q wb_dat_o[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_160_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5365_ _5366_/A1 _5366_/A3 _5366_/A4 _5424_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_7104_ _7104_/D _7302_/RN _7104_/CLK _7104_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_5296_ _5296_/A1 _5296_/A2 _5439_/C _5303_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_113_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4316_ hold541/Z hold388/Z _4316_/S _4316_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7035_ _7035_/D _7281_/RN _7035_/CLK _7035_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4247_ _4247_/A1 _4247_/A2 _4263_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_102_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4178_ _6653_/A2 _5535_/B _3527_/Z _6653_/A3 _4180_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_27_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1006 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1017 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_853 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6819_ _6819_/D input75/Z _6819_/CLK _6819_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_50_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet833_455 net833_472/I _6754_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet833_466 net433_98/I _6743_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet833_477 net833_491/I _6732_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet833_488 net833_489/I _6721_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet833_499 net833_499/I _6710_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_18_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2285 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_842 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1573 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_159_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3480_ _6703_/Q _6777_/Q _3481_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_9__1374_ clkbuf_4_3_0__1374_/Z net733_373/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_142_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5150_ _5376_/A1 _5337_/A2 _5502_/B1 _5399_/B _5150_/C _5151_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5081_ _5081_/A1 _5082_/C _5081_/B1 _5084_/C _5081_/C _5418_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_57_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4101_ input1/Z _6971_/Q _4101_/B _4101_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4032_ _4032_/I _6880_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_110_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5983_ _5983_/I0 _5983_/I1 _6790_/Q _5984_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4934_ _4947_/C _4963_/B _5288_/A4 _5451_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_177_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4865_ _4865_/A1 _4865_/A2 _4865_/A3 _4868_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_60_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6604_ _6648_/A2 _6648_/A3 _6606_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4796_ _4796_/A1 _4796_/A2 _4796_/A3 _4796_/A4 _4800_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_3816_ _3496_/B _4246_/A1 _4246_/A2 _3477_/Z _3846_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_3747_ _7067_/Q _3980_/A2 _3975_/B1 input64/Z _3943_/B1 _7197_/Q _3750_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6535_ _6901_/Q _6563_/A3 _6561_/A3 _6563_/A4 _6540_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_20_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6466_ _7215_/Q _6570_/A2 _6570_/B1 _7061_/Q _6570_/C1 _6997_/Q _6468_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_3678_ _3654_/Z _3678_/A2 _3677_/Z _6600_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_5417_ _5417_/A1 _5051_/B _4960_/C _4669_/B _5457_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6397_ _6397_/A1 _6397_/A2 _6397_/A3 _6400_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_5348_ _5348_/A1 _5052_/C _5212_/C _5464_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
Xoutput174 _3363_/ZN mgmt_gpio_oeb[12] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput185 _3353_/ZN mgmt_gpio_oeb[22] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_114_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput196 _5861_/A2 mgmt_gpio_oeb[32] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_153_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7018_ _7018_/D _7265_/RN _7018_/CLK _7018_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_5279_ _5285_/A1 _5476_/A1 _5279_/A3 _5279_/B _5371_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_88_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_68__1374_ _4109__12/I net633_282/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_43_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2060 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2093 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2071 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2082 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4650_ _4650_/A1 _4650_/A2 _4650_/A3 _4658_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_147_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3601_ _7232_/Q _3964_/A2 _4262_/S input69/Z _3635_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xinput10 mask_rev_in[15] input10/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput21 mask_rev_in[25] input21/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4581_ _5048_/B _4502_/B _4578_/B _4922_/B _5218_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_174_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput43 mgmt_gpio_in[16] input43/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput54 mgmt_gpio_in[26] input54/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_6320_ _7016_/Q _6566_/C1 _6319_/Z _7122_/Q _6333_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xinput32 mask_rev_in[6] input32/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput98 wb_adr_i[12] input98/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput65 mgmt_gpio_in[36] _7375_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_155_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3532_ _3454_/Z _3498_/B _3811_/A1 _4246_/A1 _3961_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xhold816 _7008_/Q hold816/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xinput87 spimemio_flash_io1_do _7374_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold827 _4330_/Z _6843_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold805 _6742_/Q hold805/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xinput76 qspi_enabled _4078_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xhold849 _7178_/Q hold849/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3463_ _4073_/B1 hold459/Z _6863_/Q _3511_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_143_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6251_ _6251_/A1 _6251_/A2 _6251_/A3 _6251_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_6_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold838 _6726_/Q hold838/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_5202_ _5202_/A1 _5344_/C _5202_/B _5206_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_88_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6182_ _6182_/A1 _6182_/A2 _6182_/A3 _6188_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_69_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3394_ _6774_/Q _4016_/A1 _4015_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_4
X_5133_ _5476_/A1 _5329_/A2 _5148_/B1 _5437_/A4 _5428_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5064_ _5079_/A1 _5502_/A2 _5209_/B1 _5493_/B1 _5222_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_111_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4015_ _4015_/I0 hold459/Z _4015_/S _6701_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_25_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5966_ _5966_/I0 _6296_/A2 _6789_/Q _5966_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_12_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4917_ _4686_/B _5312_/B _5098_/A2 _4920_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5897_ hold139/Z hold488/Z _5901_/S _7253_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_52_299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_474 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4848_ _5436_/A4 _5194_/B _5390_/A1 _5235_/A1 _4849_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_32_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4779_ _4779_/A1 _4779_/A2 _5023_/A3 _4963_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_119_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6518_ _7209_/Q _6573_/A2 _6288_/Z _7201_/Q _6297_/Z _7047_/Q _6524_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_4_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6449_ _7262_/Q _6581_/B1 _6312_/Z _7222_/Q _6746_/Q _6579_/A2 _6451_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_162_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_750 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet433_72 net433_82/I _7197_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_19_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet433_61 net433_65/I _7208_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet433_83 _4109__8/I _7186_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_62_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet433_94 net433_94/I _7175_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_47_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5820_ hold21/Z _5820_/A2 _3527_/Z _4227_/B _5828_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_179_249 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_51__1374_ clkbuf_4_12_0__1374_/Z net633_273/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_97_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5751_ hold25/Z hold315/Z _5756_/S _7124_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4702_ _5471_/B2 _4693_/Z _4767_/A3 _4723_/A2 _4830_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_187_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5682_ _5700_/A1 _5820_/A2 _5718_/A3 _4227_/B hold42/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_163_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4633_ _4633_/A1 _4633_/A2 _4633_/A3 _4642_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_148_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4564_ _4564_/A1 _4564_/A2 _4565_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold602 _6896_/Q hold602/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7352_ _7352_/I _7352_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3515_ _3477_/Z _3515_/A2 _3802_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_6303_ _6324_/A1 _6323_/A1 _6325_/A1 _6308_/A3 _6564_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xhold624 _6888_/Q hold624/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold635 _5637_/Z _7024_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold613 _4379_/Z _6883_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7283_ _7283_/D _7304_/RN _7304_/CLK _7283_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4495_ _4759_/C _4694_/B _5436_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_144_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold657 _6894_/Q hold657/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6234_ _6756_/Q _6257_/A2 _6261_/B1 _7340_/Q _6235_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold679 _5511_/Z _6921_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xmax_cap376 _7262_/RN _7341_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
Xhold668 _4240_/Z _6784_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold646 _4204_/Z _6759_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3446_ _3445_/Z _3446_/A2 _3446_/B _3447_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3377_ _7274_/Q _6211_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XFILLER_69_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6165_ _6107_/B _6107_/C _6973_/Q _7275_/Q _6167_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XTAP_940 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_962 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_951 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5116_ _5489_/A1 _5451_/A1 _5378_/A1 _4437_/Z _5452_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6096_ _7035_/Q _6258_/A2 _6096_/B _6096_/C _6111_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_973 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_984 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_995 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5047_ _5351_/A1 _5047_/A2 _5209_/B1 _5463_/B _5421_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_84_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6998_ _6998_/D _7281_/RN _6998_/CLK _6998_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_53_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5949_ _7274_/Q _7273_/Q _6266_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_13_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_403 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_842 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4280_ _4279_/Z hold539/Z _4282_/S _4280_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_98_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_497 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6921_ _6921_/D _7262_/RN _6921_/CLK _6921_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_120_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6852_ _6852_/D _6862_/CLK _6852_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5803_ hold391/Z hold788/Z _5810_/S _5803_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3995_ _6704_/Q _6703_/Q _6702_/Q _3992_/Z _4000_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_149_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6783_ _6783_/D input75/Z _6783_/CLK _7361_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_22_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5734_ hold58/Z hold60/Z _5735_/S hold61/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5665_ hold391/Z hold586/Z hold30/Z _7048_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_175_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4616_ _4616_/A1 _5073_/A1 _5184_/A3 _4620_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5596_ hold277/Z hold164/Z _5599_/S _5596_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold410 _7026_/Q hold410/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7335_ _7335_/D _6689_/Z _4111_/I1 _7335_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold454 _7018_/Q hold454/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_150_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold443 _6833_/Q hold443/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4547_ _5315_/A4 _3379_/I _5153_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold432 _6728_/Q hold432/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold421 _4155_/Z _6721_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_171_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4478_ _5136_/A2 _4690_/C _5235_/A2 _4922_/B _4479_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_143_182 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold465 hold465/I _7221_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7266_ _7266_/D _7302_/RN _7281_/CLK _7266_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold476 _4286_/Z _6809_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold487 _7116_/Q hold487/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7197_ _7197_/D _7341_/RN _7197_/CLK _7197_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_132_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_867 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold498 _7010_/Q hold498/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_58_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6217_ _6788_/Q _6217_/A2 _6218_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3429_ _3429_/A1 _3429_/A2 _7336_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xnet683_320 net683_320/I _6949_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6148_ _6747_/Q _6258_/B1 _6261_/B1 _7167_/Q _6151_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet683_331 net683_331/I _6938_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_85_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet683_342 net683_347/I _6927_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_781 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_4_10_0__1374_ clkbuf_3_5_0__1374_/Z clkbuf_4_10_0__1374_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_161_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6079_ _7212_/Q _6262_/A2 _6262_/B1 _7148_/Q _6083_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_46_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2604 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1914 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1903 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1958 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1947 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1936 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1969 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4109__35 net433_59/I _7234_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_108_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4109__24 _4109__24/I _7245_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4109__13 _4109__14/I _7256_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_5_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4109__46 _4109__6/I _7223_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_123_845 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_832 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3780_ _3780_/A1 _3780_/A2 _3780_/A3 _3780_/A4 _3789_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_173_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5450_ _5450_/A1 _5450_/A2 _5450_/A3 _5450_/A4 _6907_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4401_ hold388/Z hold628/Z _4401_/S _4401_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5381_ _5489_/A1 _5381_/A2 _5381_/B _5382_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_132_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4332_ _6872_/Q _7323_/RN _4343_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_141_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7120_ _7120_/D _7262_/RN _7120_/CLK _7120_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_7051_ _7051_/D _7281_/RN _7051_/CLK _7051_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_114_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4263_ hold598/Z _4262_/Z _4263_/S _4263_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6002_ _7032_/Q _6258_/A2 _6260_/B1 _6984_/Q _7275_/Q _6003_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_4194_ hold391/Z hold759/Z _4195_/S _6752_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_94_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6904_ _6904_/D _7323_/RN _7322_/CLK hold16/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xnet633_261 net633_261/I _7008_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_82_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet633_272 net783_414/I _6997_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet633_283 net783_419/I _6986_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_70_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet633_294 net783_421/I _6975_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_168_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6835_ _6835_/D _6862_/CLK _6835_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_865 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3978_ input43/Z _4243_/S _3978_/B1 _6764_/Q _3978_/C _3979_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_23_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6766_ _6766_/D _7262_/RN _6766_/CLK _6766_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5717_ hold2/Z hold232/Z _5717_/S _7095_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6697_ input75/Z _6994_/Q _4026_/C _6697_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
Xclkbuf_2_1__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/Z _7346_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_40_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5648_ hold388/Z hold665/Z _5654_/S _5648_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_156_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_156_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5579_ hold5/Z hold237/Z _5581_/S _6973_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7318_ _7318_/D _7323_/RN _4103_/I1 _7318_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_151_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold251 _6940_/Q hold251/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold240 _7175_/Q hold240/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold262 _5731_/Z _7107_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7249_ _7249_/D _7265_/RN _7249_/CLK hold49/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold284 _6994_/Q hold284/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold273 _6733_/Q hold273/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold295 _6722_/Q hold295/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_120_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1711 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1766 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_898 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_167_572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput8 mask_rev_in[13] input8/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_76_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4950_ _4773_/B _5011_/A2 _4951_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_91_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_821 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3901_ _6754_/Q _5838_/A2 _5546_/A2 _3527_/Z _3940_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_4881_ _4881_/A1 _5143_/B _4881_/A3 _5184_/A4 _4883_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_33_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6620_ _6878_/Q _6620_/A2 _6620_/B1 _6640_/B2 _6621_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3832_ _6890_/Q _5893_/A3 _4405_/A3 _4405_/A2 _3842_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_60_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6551_ _6768_/Q _6286_/Z _6580_/B1 _6899_/Q _6553_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5502_ _5502_/A1 _5502_/A2 _5502_/B1 _5502_/B2 _5502_/C _5503_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_3763_ input22/Z _3977_/A2 _3938_/A2 _7204_/Q _3766_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3694_ _6730_/Q _3959_/A2 _3964_/C1 _7262_/Q _3698_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6482_ _7299_/Q _6587_/A2 _6532_/B _6532_/C _6483_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5433_ _5433_/A1 _5433_/A2 _5433_/A3 _5450_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xoutput301 _3642_/Z serial_data_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_160_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5364_ _5272_/C _5051_/B _4960_/C _4669_/B _5366_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_133_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput334 _7312_/Q wb_dat_o[30] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput323 _6839_/Q wb_dat_o[20] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput312 _6847_/Q wb_dat_o[10] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_7103_ hold23/Z _7265_/RN _7103_/CLK _7103_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_160_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4315_ hold443/Z hold391/Z _4316_/S _4315_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5295_ _5295_/A1 _5290_/C _5435_/A1 _5466_/C _5295_/C _5296_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_113_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4246_ _4246_/A1 _4246_/A2 _4246_/A3 hold45/Z _4247_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_7034_ _7034_/D _7302_/RN _7034_/CLK _7034_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_95_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4177_ hold684/Z hold388/Z _4177_/S _6739_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1007 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1018 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1029 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6818_ _6818_/D input75/Z _6818_/CLK _6818_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_184_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6749_ _6749_/D _7304_/RN _6749_/CLK _6749_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_167_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_714 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_28__1374_ clkbuf_4_11_0__1374_/Z net433_81/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_2_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_108__1374_ net733_398/I net683_349/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_104_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_5_0__1374_ clkbuf_0__1374_/Z clkbuf_3_5_0__1374_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_76_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet833_467 net433_98/I _6742_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet833_478 net833_491/I _6731_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_18_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet833_456 net833_456/I _6753_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2253 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet833_489 net833_489/I _6720_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1541 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_789 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_835 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5080_ _5075_/Z _5229_/A1 _5460_/A1 _5230_/B _5085_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4100_ input1/Z input2/Z _4101_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4031_ _6880_/Q _4074_/A2 _6875_/Q _4032_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_84_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5982_ _6787_/Q _6788_/Q _6789_/Q _5983_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_178_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4933_ _3379_/I _3380_/I _5445_/A2 _4956_/C _5056_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_18_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4864_ _5136_/A2 _5466_/B _5466_/A1 _4922_/B _4865_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_119_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4795_ _5152_/C _5327_/B _5252_/A3 _5426_/B1 _4796_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_6603_ _3597_/Z _7313_/Q _6603_/S _7313_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3815_ _6854_/Q _4378_/A1 _5748_/A3 _4405_/A2 _3840_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6534_ _6910_/Q _6563_/A2 _6562_/A3 _6563_/A4 _6543_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3746_ input46/Z _4243_/S _3939_/B1 input29/Z _3980_/B1 _6979_/Q _3750_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_146_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6465_ _6465_/A1 _6465_/A2 _6465_/A3 _6465_/A4 _6465_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_146_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5416_ _5416_/A1 _5084_/B _5290_/B _5416_/B _5433_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_3677_ _3669_/Z _3677_/A2 _3677_/A3 _3676_/Z _3677_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_161_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6396_ _6584_/A1 _6396_/A2 _6396_/A3 _6395_/Z _6397_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5347_ _5347_/A1 _5347_/A2 _5347_/B _5348_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput175 _3362_/ZN mgmt_gpio_oeb[13] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput186 _3352_/ZN mgmt_gpio_oeb[23] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput197 _3342_/ZN mgmt_gpio_oeb[33] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5278_ _5372_/B _5498_/A2 _5278_/B _5281_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_141_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4229_ hold671/Z hold391/Z _4243_/S _4229_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7017_ _7017_/D _7265_/RN _7017_/CLK _7017_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_101_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_640 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_678 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2061 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2050 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2094 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2083 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1393 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1360 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_175_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4580_ _4502_/B _4922_/B _4598_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xinput22 mask_rev_in[26] input22/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput11 mask_rev_in[16] input11/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_30_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3600_ _3599_/Z hold878/Z _3888_/S _6919_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_174_147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput44 mgmt_gpio_in[17] input44/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput55 mgmt_gpio_in[27] input55/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3531_ _3454_/Z _3498_/B _3827_/A1 _3644_/A2 _3964_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xinput33 mask_rev_in[7] input33/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput66 mgmt_gpio_in[37] _7376_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_183_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold828 _7195_/Q hold828/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xinput88 spimemio_flash_io1_oeb input88/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold817 _5619_/Z _7008_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold806 _6968_/Q hold806/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xinput77 ser_tx input77/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput99 wb_adr_i[13] input99/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_171_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3462_ hold11/Z _6777_/Q hold12/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_143_545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6250_ _6769_/Q _6258_/A2 _6259_/B1 _6735_/Q _6257_/B1 _6771_/Q _6251_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
Xhold839 _4161_/Z _6726_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_143_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5201_ _5201_/A1 _5424_/A2 _6879_/Q _5201_/C _5207_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_124_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_11__1374_ clkbuf_4_8_0__1374_/Z net433_67/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6181_ hold83/I _6262_/A2 _6258_/C1 _7192_/Q hold96/I _6258_/A2 _6182_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_42_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3393_ _4020_/A2 _3389_/Z _6777_/Q _4016_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_130_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5132_ _5329_/A2 _5376_/A1 _5502_/B1 _5394_/C _5134_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xclkbuf_leaf_74__1374_ clkbuf_4_5_0__1374_/Z net733_397/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_97_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5063_ _5463_/A1 _5493_/B1 _5063_/B _5494_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_84_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4014_ _6777_/Q _3992_/Z _4014_/A3 hold12/I _4015_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_52_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5965_ _7277_/Q _7276_/Q _7278_/Q _6296_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_4916_ _4451_/B _4916_/A2 _4916_/A3 _4776_/Z _5290_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_5896_ hold25/Z hold469/Z _5901_/S _7252_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4847_ _5084_/B _4661_/C _4718_/B _4487_/Z _5404_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_119_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4778_ _4960_/C _4779_/A1 _4779_/A2 _4778_/A4 _4956_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_147_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet733_400 net783_411/I _6818_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_20_186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3729_ _3729_/A1 _3729_/A2 _3729_/A3 _3732_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6517_ _6517_/A1 _6517_/A2 _6516_/Z _6517_/A4 _6517_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_134_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6448_ _7028_/Q _6528_/A2 _6311_/C _7004_/Q _6452_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_164_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6379_ _7026_/Q _6562_/A2 _6562_/A3 _6562_/A4 _6396_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_88_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_71 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_429 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet433_62 net433_62/I _7207_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet433_84 net433_84/I _7185_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet433_73 net433_81/I _7196_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_74_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet433_95 net433_99/I _7174_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_34_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_896 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5750_ hold388/Z hold753/Z _5756_/S _7123_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5681_ hold2/Z hold56/Z _5681_/S _7063_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4701_ _5267_/C _4667_/Z _4959_/C _4451_/B _5199_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XTAP_1190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4632_ _5051_/B _5051_/C _5290_/A1 _5483_/A1 _4633_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_129_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4563_ _4555_/Z _4563_/A2 _5051_/B _5051_/C _4564_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
Xhold603 _4398_/Z _6896_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7351_ _7351_/I _7351_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4494_ _5459_/A3 _5225_/A3 _5225_/A1 _5347_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_3514_ _3827_/A2 hold28/Z _3608_/A4 hold29/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
Xhold614 _6949_/Q hold614/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xclkbuf_4_8_0__1374_ clkbuf_4_9_0__1374_/I clkbuf_4_8_0__1374_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_6302_ _6312_/A4 _6563_/A4 _7277_/Q _7276_/Q _6316_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_116_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold625 _4386_/Z _6888_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7282_ _7282_/D _7304_/RN _7304_/CLK _7282_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold636 _6830_/Q hold636/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xmax_cap344 _5573_/A3 _5552_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_144_876 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold658 _4395_/Z _6894_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold669 _7025_/Q hold669/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6233_ _6758_/Q _6233_/A2 _6233_/B1 _6762_/Q _6266_/B _6766_/Q _6235_/B1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
Xmax_cap377 _7302_/RN _7281_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
Xhold647 _6735_/Q hold647/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3445_ _7327_/Q _6707_/Q _3445_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_97_462 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6164_ _7275_/Q _6164_/A2 _6164_/B _6167_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3376_ _7271_/Q _6103_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_8
XTAP_930 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_952 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5115_ _5378_/A1 _5279_/A3 _5115_/B _5117_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6095_ _6095_/A1 _6095_/A2 _6095_/A3 _6096_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_963 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_974 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_985 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5046_ _5046_/A1 _5046_/A2 _5048_/C _5046_/C _5463_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_111_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_830 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6997_ _6997_/D _7281_/RN _6997_/CLK _6997_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_13_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5948_ _6787_/Q _6789_/Q _6211_/C _5948_/B1 _6258_/A2 _7274_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_43_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5879_ hold483/Z hold139/Z _5883_/S _7237_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_138_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_896 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_284 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_185_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_364 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6920_ _6920_/D _7262_/RN _6920_/CLK _6920_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6851_ _6851_/D _6862_/CLK _6851_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5802_ _5856_/A1 _5802_/A2 _3527_/Z _5535_/B _5810_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_3994_ _7347_/Q _6702_/Q _6701_/Q hold11/I _4006_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6782_ _6782_/D _7281_/RN _6782_/CLK _7360_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_176_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5733_ hold5/Z hold93/Z _5735_/S hold94/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5664_ _5700_/A1 hold8/Z _5718_/A3 _4227_/B hold30/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_175_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4615_ _4661_/C _5439_/C _5436_/A4 _5439_/B _5184_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_5595_ hold406/Z hold139/Z _5599_/S _5595_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_175_297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7334_ _7334_/D _6688_/Z _4089_/I1 hold1/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4546_ _3380_/I _4423_/Z _5445_/A3 _5262_/A4 _5051_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_117_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold411 _5639_/Z _7026_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold400 _6978_/Q hold400/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_145_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold444 _4315_/Z _6833_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold433 _4163_/Z _6728_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_2_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold422 _7036_/Q hold422/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4477_ _3379_/I _4421_/Z _4423_/Z _4759_/C _4951_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_7265_ hold48/Z _7265_/RN _7265_/CLK hold47/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold455 _5630_/Z _7018_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold466 _7141_/Q hold466/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold477 _7260_/Q hold477/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7196_ _7196_/D _7265_/RN _7196_/CLK _7196_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_143_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold499 _5621_/Z _7010_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_86_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold488 _7253_/Q hold488/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6216_ _6107_/B _6107_/C hold98/I _7275_/Q _6217_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_3428_ _6774_/Q _3431_/B _3428_/B _3429_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3359_ _7099_/Q _6107_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
Xnet683_321 net783_417/I _6948_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet683_310 net683_310/I _6959_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6147_ _7143_/Q _6259_/A2 _6257_/B1 _7183_/Q _6151_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet683_343 net683_347/I _6926_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet683_332 net683_347/I _6937_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_793 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6078_ _6078_/A1 _6235_/B2 _6078_/B _6078_/C _6084_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_2627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2616 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5029_ _5394_/A2 _5194_/B _5039_/A1 _5315_/A4 _5120_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_2638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1915 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1904 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1959 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1948 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1937 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1926 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_186_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4109__14 _4109__14/I _7255_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4109__25 _4109__44/I _7244_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4109__36 net433_77/I _7233_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4109__47 net433_66/I _7222_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_150_654 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_616 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_830 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4400_ hold391/Z hold722/Z _4401_/S _4400_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_8_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5380_ _5476_/B _5380_/A2 _5453_/A1 _5380_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_126_640 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4331_ hold706/Z hold388/Z _4331_/S _4331_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7050_ _7050_/D _7265_/RN _7050_/CLK _7050_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_87_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4262_ hold197/Z hold2/Z _4262_/S _4262_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6001_ _6036_/A3 _7271_/Q _7274_/Q _7273_/Q _6260_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_4193_ _5838_/A4 _5528_/A2 _5748_/A3 _5784_/A2 _4195_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_36_830 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6903_ _6903_/D _7323_/RN _7322_/CLK hold20/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_82_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet633_273 net633_273/I _6996_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet633_262 net633_289/I _7007_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet633_284 net633_292/I _6985_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet633_295 net833_464/I _6974_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_36_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6834_ _6834_/D _7341_/RN _6834_/CLK _6834_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_50_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6765_ _6765_/D _7341_/RN _6765_/CLK _6765_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3977_ input20/Z _3977_/A2 _3977_/B1 _7032_/Q _3979_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_11_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5716_ hold58/Z hold357/Z _5717_/S _7094_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_149_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6696_ input75/Z _6994_/Q _4026_/C _6696_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_163_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5647_ hold391/Z hold803/Z _5654_/S _5647_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_156_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5578_ hold164/Z hold282/Z _5581_/S _6972_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7317_ _7317_/D _7323_/RN _4103_/I1 _7317_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_144_481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4529_ _5466_/B _5037_/A1 _3379_/I _3380_/I _5218_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xhold252 _5539_/Z _6940_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold241 _5808_/Z _7175_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_2_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold230 _7143_/Q hold230/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7248_ _7248_/D _7265_/RN _7248_/CLK hold95/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold285 _5603_/Z _6994_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_132_654 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold274 _4168_/Z _6733_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold296 _4156_/Z _6722_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold263 _7115_/Q hold263/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_49_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7179_ _7179_/D _7265_/RN _7179_/CLK _7179_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_86_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2435 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_157_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1745 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1789 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput9 mask_rev_in[14] input9/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_92_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4880_ _5445_/A2 _5177_/A3 _5153_/B _5439_/B _5184_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_32_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3900_ _7349_/I _5856_/A1 _5838_/A2 _5532_/A3 _3968_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_3831_ _3496_/B _3831_/A2 _4227_/A2 _3477_/Z _3945_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_33_866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3762_ input26/Z _3939_/B1 _3977_/B1 _7034_/Q _3766_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_20_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6550_ _6895_/Q _6581_/B1 _6312_/Z _6750_/Q _7120_/Q _6579_/A2 _6553_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_5501_ hold34/I _4365_/C _5505_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3693_ _7246_/Q _3981_/A2 _3981_/B1 _7254_/Q _3698_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_9_572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6481_ _6481_/A1 _6481_/A2 _6973_/Q _6584_/A1 _6584_/B _6483_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_173_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5432_ _5432_/A1 _5432_/A2 _5432_/A3 _5432_/B _5450_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_5363_ _5363_/A1 _4647_/C _5457_/A1 _5367_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xoutput335 _7313_/Q wb_dat_o[31] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput324 _6840_/Q wb_dat_o[21] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput313 _6848_/Q wb_dat_o[11] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput302 _3605_/Z serial_data_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_7102_ hold65/Z _7265_/RN _7102_/CLK hold64/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4314_ hold45/Z hold190/Z _4378_/A1 _5655_/A4 _4316_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_5294_ _5294_/A1 _5466_/A2 _5294_/B _5294_/C _5296_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_114_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4245_ _4264_/A1 _5564_/A3 _4262_/S _4247_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_101_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7033_ _7033_/D _7302_/RN _7033_/CLK _7033_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_28_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4176_ hold771/Z hold391/Z _4177_/S _6738_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1008 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1019 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6817_ _6817_/D input75/Z _6817_/CLK _6817_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_183_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6748_ hold73/Z _7304_/RN _6748_/CLK hold72/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_176_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6679_ _7262_/RN _6994_/Q _4026_/C _6679_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_164_543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet833_468 net833_472/I _6741_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet833_457 net833_489/I _6752_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_46_446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet833_479 net833_483/I _6730_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_46_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2287 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_71 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_174_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_713 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4030_ _4030_/I _6879_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_84_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5981_ _5985_/A2 _5981_/A2 _5983_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4932_ _5369_/A1 _4963_/B _5463_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_80_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_34__1374_ clkbuf_4_11_0__1374_/Z net433_89/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4863_ _4423_/Z _5502_/B2 _5177_/A3 _5153_/B _5388_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6602_ _6602_/A1 _6603_/S _6602_/B _7312_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_114__1374_ clkbuf_4_2_0__1374_/Z net833_454/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4794_ _5312_/B _4794_/A2 _5152_/C _5327_/B _5337_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_3814_ _6896_/Q hold37/I _5748_/A3 _5546_/A2 _3862_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
Xclkbuf_leaf_97__1374_ clkbuf_4_1_0__1374_/Z net783_441/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_158_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3745_ _3745_/A1 _3745_/A2 _3745_/A3 _3751_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_21_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6533_ _6533_/A1 _6533_/A2 _6533_/B _7302_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_173_340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6464_ _7167_/Q _6279_/Z _6299_/Z _7069_/Q _6465_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_174_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5415_ _5476_/B _5415_/A2 _5415_/A3 _5453_/A2 _5416_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_133_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3676_ _3676_/A1 _3676_/A2 _3676_/A3 _3676_/A4 _3676_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_6395_ _6395_/A1 _6395_/A2 _6395_/A3 _6395_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_5346_ _4443_/Z _5459_/A3 _5355_/A2 _5346_/A4 _5347_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xoutput176 _3361_/ZN mgmt_gpio_oeb[14] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_102_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput198 _3341_/ZN mgmt_gpio_oeb[34] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5277_ _5277_/A1 _5412_/A4 _5373_/A2 _5278_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_141_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput187 _3351_/ZN mgmt_gpio_oeb[24] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_7016_ _7016_/D _7265_/RN _7016_/CLK _7016_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_141_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4228_ _4228_/A1 _4228_/A2 _4244_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_87_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4159_ hold179/Z hold2/Z _4159_/S _4159_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_46_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_714 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2051 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2040 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2095 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2073 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2084 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2062 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput12 mask_rev_in[17] input12/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput45 mgmt_gpio_in[18] input45/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3530_ _3473_/B _3802_/A2 _3511_/C _5534_/A1 _3973_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xinput23 mask_rev_in[27] input23/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_7_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput34 mask_rev_in[8] input34/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_171_833 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput56 mgmt_gpio_in[28] input56/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_115_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput89 spimemio_flash_io2_do input89/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold807 _6866_/Q hold807/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold818 _6754_/Q hold818/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_7_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput78 spi_csb input78/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput67 mgmt_gpio_in[3] input67/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xhold829 _7073_/Q hold829/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_170_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3461_ _3534_/C _3454_/Z _5534_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_5200_ _5295_/A1 _5466_/A2 _5200_/B _5290_/C _5323_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_6180_ hold70/I _6259_/A2 _6256_/A2 hold68/I _6182_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3392_ _3316_/I _3421_/A2 _4020_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5131_ _5131_/A1 _5476_/A1 _5148_/B1 _5394_/C _5131_/C _5134_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_35_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5062_ _4922_/B _5046_/C _5062_/A3 _4502_/B _5493_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_97_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4013_ _7347_/Q hold11/I _6701_/Q _4014_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_96_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5964_ _6310_/A4 _6306_/A3 _7278_/Q _5967_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_80_577 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4915_ _4451_/B _4916_/A2 _4916_/A3 _4776_/Z _5039_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_5895_ hold388/Z hold549/Z _5901_/S _7251_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4846_ _4669_/B _4774_/B _4916_/A2 _4916_/A3 _5390_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_33_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4777_ _4840_/A1 _4777_/A2 _4777_/B _4777_/C _5023_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_6516_ _6516_/A1 _6516_/A2 _6516_/A3 _6516_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
Xnet733_401 net783_411/I _6817_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_20_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3728_ _7027_/Q _3961_/B1 _3945_/A2 _7133_/Q _3729_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_173_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6447_ _7092_/Q _6578_/A2 _6310_/Z _6980_/Q _6578_/C1 _7174_/Q _6452_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_3659_ _3659_/A1 _3659_/A2 _3660_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_161_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6378_ _7148_/Q _6562_/A2 _6562_/A3 _6561_/A3 _6383_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_88_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5329_ _5489_/A1 _5329_/A2 _5489_/B1 _5394_/C _5330_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_88_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_719 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_80__1374_ clkbuf_4_4_0__1374_/Z net533_163/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_171_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_793 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_796 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet433_52 net433_53/I _7217_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet433_63 _4109__9/I _7206_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_47_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet433_85 net433_86/I _7184_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet433_74 net433_74/I _7195_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet433_96 net433_97/I _7173_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_35_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5680_ hold58/Z hold66/Z _5681_/S _7062_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4700_ _4794_/A2 _4765_/B _4767_/A3 _4723_/A2 _5267_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XTAP_1191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1180 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4631_ _4469_/B _4759_/C _4686_/B _5307_/B _5483_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_8_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4562_ _5051_/B _4454_/B _4563_/A2 _4959_/C _5351_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_8_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7350_ _7350_/I _7350_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_171_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4493_ _5051_/B _4454_/B _4959_/C _5351_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_6301_ _6325_/A1 _6308_/A3 _7279_/Q _7278_/Q _6571_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_3513_ _3811_/A1 _3460_/B _3498_/B _3831_/A2 _3961_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_7281_ _7281_/D _7281_/RN _7281_/CLK _7281_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
Xhold626 _6887_/Q hold626/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold615 _6944_/Q hold615/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold604 _7043_/Q hold604/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold659 _6993_/Q hold659/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_143_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xmax_cap367 _5655_/A4 _5745_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_89_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6232_ _7120_/Q _6266_/C _6232_/B1 _6764_/Q _6232_/C _6235_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
Xhold648 _4171_/Z _6735_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3444_ input58/Z _6709_/Q _6708_/Q _6774_/Q _3447_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xhold637 _7352_/I hold637/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xmax_cap378 _7262_/RN _7302_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
Xmax_cap356 _6653_/A3 _5784_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_103_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6163_ _7272_/Q _7271_/Q _6163_/A3 _6162_/Z _7275_/Q _6164_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_3375_ _7272_/Q _6036_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_8
XTAP_920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_931 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_942 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_953 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5114_ _5379_/A1 _5414_/A1 _5114_/A3 _5379_/A2 _5115_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_111_251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6094_ _6987_/Q _6260_/B1 _6258_/C1 _7067_/Q _6095_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_964 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_975 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_986 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5045_ _5439_/A1 _5045_/A2 _5350_/B _5209_/B1 _5215_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_97_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_997 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6996_ _6996_/D _7281_/RN _6996_/CLK _6996_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_92_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5947_ _5947_/A1 _6789_/Q _5948_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_577 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5878_ hold445/Z hold25/Z _5883_/S _7236_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_166_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4829_ _4830_/B2 _4661_/C _4718_/B _5392_/A1 _4830_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_21_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_285 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold1 hold1/I hold1/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_79_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_842 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6850_ _6850_/D _6862_/CLK _6850_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5801_ hold2/Z _7169_/Q hold9/Z hold10/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6781_ _6781_/D _7281_/RN _6781_/CLK _7359_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_90_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3993_ _7347_/Q _6702_/Q _6701_/Q hold11/I _3993_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_5732_ hold164/Z hold181/Z _5735_/S _5732_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_175_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5663_ hold2/Z hold234/Z _5663_/S _7047_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4614_ _4443_/Z _5459_/A3 _5439_/A1 _5439_/B _5073_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_135_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5594_ hold500/Z hold25/Z _5599_/S _5594_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_117_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7333_ _7333_/D _6687_/Z _4089_/I1 hold57/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4545_ _4423_/Z _5210_/C _5210_/B _5262_/A4 _5375_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_116_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold401 _5585_/Z _6978_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold445 _7236_/Q hold445/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_143_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold412 _6731_/Q hold412/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold434 _7135_/Q hold434/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold423 _5651_/Z _7036_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4476_ _4759_/C _4684_/B _5307_/B _4694_/B _4587_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_7264_ hold81/Z _7265_/RN _7264_/CLK hold80/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold456 _7188_/Q hold456/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold467 _7228_/Q hold467/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold478 _5905_/Z _7260_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7195_ _7195_/D _7341_/RN _7195_/CLK _7195_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_6215_ _7275_/Q _6202_/Z _6215_/B _6218_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold489 _6810_/Q hold489/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3427_ _3431_/B _3427_/A2 _3427_/B hold891/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3358_ _7107_/Q _3358_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet683_322 net783_417/I _6947_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet683_311 net683_314/I _6958_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_85_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6146_ _7159_/Q _6258_/A2 _6259_/B1 hold93/I _6256_/B1 _7207_/Q _6152_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XTAP_750 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xload_slew370 hold45/Z _5535_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
Xnet683_344 net683_347/I _6925_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet683_333 net433_99/I _6936_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_85_466 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6077_ _7172_/Q _6256_/A2 _6258_/B1 _6744_/Q _6261_/B1 _7164_/Q _6078_/C VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XTAP_2617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2606 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5028_ _5417_/A1 _5039_/A1 _5476_/A2 _5489_/A1 _5030_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_85_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2639 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1916 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_864 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1949 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1938 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1927 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6979_ _6979_/D _7281_/RN _6979_/CLK _6979_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_10_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4109__26 net433_58/I _7243_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_135_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4109__15 net433_75/I _7254_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_107_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4109__37 net433_77/I _7232_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4109__48 _4109__48/I _7221_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_134_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_842 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_823 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_878 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_569 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4330_ hold826/Z hold391/Z _4331_/S _4330_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_125_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4261_ hold594/Z _4260_/Z _4263_/S _4261_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6000_ _7088_/Q _6262_/A2 _6257_/A2 _7008_/Q _6003_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_86_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4192_ hold388/Z hold682/Z _4192_/S _4192_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet633_252 net433_90/I _7017_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6902_ _6902_/D _7262_/RN _6902_/CLK _6902_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xnet633_274 net783_414/I _6995_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6833_ _6833_/D _7341_/RN _6833_/CLK _6833_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xnet633_263 net633_281/I _7006_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet633_285 net633_289/I _6984_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_36_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet633_296 net633_301/I _6973_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_24_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3976_ _3976_/A1 _3976_/A2 _3976_/A3 _3976_/A4 _3983_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6764_ _6764_/D _7341_/RN _6764_/CLK _6764_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_148_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6695_ _7262_/RN _6994_/Q _4026_/C _6695_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_5715_ hold5/Z hold426/Z _5717_/S _7093_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5646_ _5700_/A1 _5646_/A2 hold13/Z _4227_/B _5654_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_176_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_156_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5577_ hold139/Z hold409/Z _5581_/S _6971_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold220 _6716_/Q hold220/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4528_ _5262_/A4 _5315_/A4 _5301_/A2 _4661_/C _5295_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_7316_ _7316_/D _7323_/RN _4103_/I1 _7316_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_144_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_836 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold242 _6970_/Q hold242/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold253 _6941_/Q hold253/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold231 _5772_/Z _7143_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7247_ _7247_/D _7265_/RN _7247_/CLK _7247_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4459_ _4684_/B _4437_/Z _5312_/B _4463_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xhold286 _7230_/Q hold286/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold275 _7028_/Q hold275/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold264 _5740_/Z _7115_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold297 _6702_/Q hold297/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7178_ _7178_/D _7341_/RN _7178_/CLK _7178_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_98_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6129_ _7126_/Q _6129_/A2 _6127_/Z _6262_/A2 _6128_/Z _6262_/B1 _6138_/C VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_85_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_403 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2403 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1713 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1746 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3830_ _6888_/Q _5655_/A4 hold29/I _5546_/A2 _3878_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_3761_ _6978_/Q _5655_/A4 _5727_/A3 _4378_/A1 _3773_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_186_861 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5500_ _5500_/A1 _5500_/A2 _5500_/B _5500_/C _5505_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_158_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6480_ _6584_/A1 _6480_/A2 _6480_/A3 _6479_/Z _6481_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3692_ _6972_/Q _3559_/Z _3692_/B _3698_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_145_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5431_ _5473_/A1 _5473_/A2 _5492_/A4 _5431_/A4 _5432_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_65_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5362_ _5362_/A1 _5362_/A2 _5418_/A2 _5461_/A2 _5363_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_114_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput325 _6841_/Q wb_dat_o[22] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput303 _4106_/Z serial_load VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput314 _6849_/Q wb_dat_o[12] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_7101_ _7101_/D _7265_/RN _7101_/CLK _7101_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4313_ hold388/Z hold688/Z _4313_/S _4313_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xoutput336 _6858_/Q wb_dat_o[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5293_ _5293_/A1 _5293_/A2 _5293_/A3 _5293_/A4 _5293_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_101_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7032_ _7032_/D _7302_/RN _7032_/CLK _7032_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_113_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_57__1374_ clkbuf_4_13_0__1374_/Z net633_290/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4244_ hold592/Z _4243_/Z _4244_/S _4244_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4175_ _5838_/A4 _5518_/A1 _5784_/A2 _5745_/A4 _4177_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_83_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1009 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6816_ _6816_/D _7281_/RN _6816_/CLK _6816_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_24_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6747_ _6747_/D _7304_/RN _6747_/CLK _6747_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_50_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3959_ _6726_/Q _3959_/A2 _3959_/B1 _6752_/Q _3960_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_167_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6678_ _7262_/RN _6994_/Q _4026_/C _6678_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_5629_ hold388/Z hold751/Z _5635_/S _5629_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet833_458 net833_470/I _6751_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet833_469 net833_469/I _6740_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_74 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1532 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_175_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_186_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_170_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_1_0__f__1033_ clkbuf_0__1033_/Z _4354_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_151_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5980_ _6787_/Q _6789_/Q _5975_/B _5980_/B _7281_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_80_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4931_ _5123_/B _5293_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4862_ _5136_/A2 _5466_/B _5416_/A1 _4922_/B _4865_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_32_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3813_ _3496_/B _5534_/A2 _4227_/A2 _3477_/Z _3978_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_6601_ _6603_/S _7312_/Q _6602_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4793_ _5250_/B _3380_/I _5098_/A2 _5252_/A4 _4796_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_21_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_500 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3744_ _7051_/Q _3973_/A2 _3946_/A2 _7019_/Q _3943_/C1 _7059_/Q _3745_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6532_ _7301_/Q _6587_/A2 _6532_/B _6532_/C _6533_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_174_875 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6463_ _7053_/Q _6575_/B1 _6566_/C1 _7021_/Q _6465_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_118_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3675_ _7077_/Q _3951_/A2 _3981_/B1 _7255_/Q _3676_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_174_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5414_ _5414_/A1 _5371_/Z _5414_/A3 _5414_/A4 _5453_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_134_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6394_ _7260_/Q _6581_/B1 _6312_/Z _7220_/Q _6395_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5345_ _5051_/B _4454_/B _5353_/A3 _4959_/C _5493_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xoutput177 _3360_/ZN mgmt_gpio_oeb[15] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_130_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_719 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput199 _4084_/ZN mgmt_gpio_oeb[35] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5276_ _4956_/C _5410_/A2 _5410_/A3 _5498_/A2 _5373_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_141_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput188 _3350_/ZN mgmt_gpio_oeb[25] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_102_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4227_ _5534_/A2 _4227_/A2 _4246_/A3 _4227_/B _4228_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_7015_ _7015_/D _7302_/RN _7015_/CLK _7015_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_68_572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4158_ hold245/Z hold58/Z _4159_/S _4158_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4089_ _6800_/Q _4089_/I1 _7345_/Q _4089_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_71_726 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_820 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_40__1374_ clkbuf_4_14_0__1374_/Z net433_68/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_47_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2052 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2041 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2030 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2085 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2096 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1395 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput13 mask_rev_in[18] input13/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput46 mgmt_gpio_in[19] input46/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput24 mask_rev_in[28] input24/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput35 mask_rev_in[9] input35/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_156_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput57 mgmt_gpio_in[29] input57/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_143_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold808 _4370_/Z _6866_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold819 _4197_/Z _6754_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xinput68 mgmt_gpio_in[5] input68/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xinput79 spi_enabled _4087_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_3460_ _6863_/Q hold20/Z _3460_/B _3460_/C hold21/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_115_249 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3391_ _7337_/Q _7336_/Q _3421_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5130_ _5130_/A1 _5242_/A1 _5243_/B _5130_/A4 _5131_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5061_ _5061_/A1 _5356_/A1 _5219_/A1 _5061_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_123_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4012_ _4012_/I0 hold903/Z _4015_/S _6702_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_111_466 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5963_ _5963_/I _7277_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_93_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4914_ _4362_/Z _4914_/A2 _5042_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5894_ hold391/Z hold693/Z _5901_/S _7250_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4845_ _4684_/B _5393_/A3 _5153_/A2 _5153_/B _5245_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_165_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4776_ _4779_/A1 _4779_/A2 _4776_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3727_ _7091_/Q _3951_/B1 _3962_/B1 _7083_/Q _3729_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6515_ hold54/I _6292_/Z _6571_/B1 _6991_/Q _6571_/C1 hold50/I _6516_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_180_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6446_ _6446_/A1 _6446_/A2 _6446_/A3 _6452_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_3658_ _7093_/Q _3951_/B1 _3958_/B1 _6723_/Q _3659_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_164_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_867 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3589_ _7169_/Q _3878_/A2 _3977_/B1 hold85/I _3595_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6377_ _7244_/Q _6563_/A2 _6562_/A3 _6563_/A4 _6386_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_130_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5328_ _5328_/A1 _5328_/A2 _5328_/A3 _5328_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_102_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5259_ _5259_/A1 _5335_/A2 _5427_/A2 _5261_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_57_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_745 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_789 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_156_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_678 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet433_53 net433_53/I _7216_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_75_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet483_150 net533_176/I _7119_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_35_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet433_86 net433_86/I _7183_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet433_75 net433_75/I _7194_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_75_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet433_64 net433_64/I _7205_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_62_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet433_97 net433_97/I _7172_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_34_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4630_ _5312_/B _4684_/B _4922_/B _4694_/B _5321_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_148_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4561_ _5307_/B _5436_/A2 _5226_/A1 _4686_/B _4563_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6300_ _6562_/A2 _6310_/A4 _7276_/Q _6562_/A4 _6300_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_183_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4492_ _4960_/C _5225_/A1 _5225_/A3 _5082_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_155_182 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold605 _7258_/Q hold605/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3512_ _3507_/C _3473_/B _3831_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_7280_ _7280_/D _7281_/RN _7281_/CLK _7280_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
Xhold627 _4385_/Z _6887_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold616 _5543_/Z _6944_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xmax_cap368 hold8/Z _5655_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_144_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6231_ _6231_/I _6241_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3443_ _6708_/Q _3443_/A2 _3443_/B _7327_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold638 _4257_/Z _6795_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold649 _6950_/Q hold649/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_103_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6162_ _6162_/A1 _6162_/A2 _6162_/A3 _6161_/Z _6162_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
Xmax_cap379 _7262_/RN _7304_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
XTAP_910 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5113_ _5355_/A2 _5093_/B _5282_/B _5379_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3374_ _7275_/Q _6232_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_4
XTAP_921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_932 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_943 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6093_ _7075_/Q _6260_/A2 _6256_/B1 _7083_/Q _6095_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_58_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_965 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_954 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_987 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5044_ _5323_/C _6876_/Q hold16/I _5207_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_111_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_998 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6995_ _6995_/D _7265_/RN _6995_/CLK _6995_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_81_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5946_ _6107_/B _7273_/Q _6211_/C _5947_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_13_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5877_ hold555/Z hold388/Z _5883_/S _7235_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_159_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4828_ _5271_/A1 _4830_/B2 _4828_/B _4828_/C _4830_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_166_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4759_ _4694_/B _4759_/A2 _4759_/B1 _5136_/A2 _4759_/C _5252_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_175_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6429_ _6788_/Q _4019_/Z _6509_/B _7299_/Q _6455_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_161_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_253 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_144_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold2 hold2/I hold2/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_66_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3992_ _7347_/Q _6701_/Q hold11/I _3992_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_5800_ hold58/Z hold105/Z hold9/Z _7168_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6780_ _6780_/D _7281_/RN _6780_/CLK _7358_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_23_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5731_ hold139/Z hold261/Z _5735_/S _5731_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5662_ hold58/Z hold362/Z _5663_/S _7046_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_175_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4613_ _5051_/B _4454_/B _5426_/A1 _4959_/C _5226_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_5593_ hold760/Z hold388/Z _5599_/S _5593_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7332_ _7332_/D _6686_/Z _4089_/I1 hold4/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_163_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4544_ _5439_/A1 _4686_/B _5307_/B _5436_/A2 _4555_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xhold402 _6996_/Q hold402/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7263_ _7263_/D _7265_/RN _7263_/CLK _7263_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_144_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold424 _6818_/Q hold424/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold413 _4166_/Z _6731_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold435 _5763_/Z _7135_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4475_ _4469_/B _4690_/B _4922_/B _5502_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
Xhold457 _5823_/Z _7188_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_144_697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6214_ _7275_/Q _6214_/A2 _6213_/Z _6261_/A2 _6214_/C _6215_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
Xhold446 _6730_/Q hold446/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold468 _6930_/Q hold468/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_132_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7194_ _7194_/D _7341_/RN _7194_/CLK _7194_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_98_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold479 _6817_/Q hold479/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3426_ _3421_/B _3426_/A2 _3428_/B _3427_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3357_ _7115_/Q _3357_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet683_312 net683_317/I _6957_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6145_ _7215_/Q _6262_/A2 _6258_/C1 _7191_/Q _6152_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xload_slew371 hold45/Z _4227_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
Xnet683_323 _4109__24/I _6946_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_97_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6076_ _7204_/Q _6233_/A2 _6233_/B1 _7196_/Q _6266_/B _7188_/Q _6078_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
Xnet683_334 net833_497/I _6935_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet683_345 net683_347/I _6924_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_762 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_784 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5027_ _4425_/Z _5194_/B _5039_/A1 _5315_/A4 _5409_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_39_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1906 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1939 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1928 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1917 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6978_ _6978_/D _7302_/RN _6978_/CLK _6978_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_179_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5929_ _7267_/Q _7268_/Q _7269_/Q _7270_/Q _5929_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_139_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_715 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_182 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4109__16 _4109__16/I _7253_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4109__38 net433_77/I _7231_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_135_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4109__27 _4109__8/I _7242_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_108_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4109__49 _4109__49/I _7220_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_123_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_865 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_358 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_71 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4260_ hold206/Z hold58/Z _4262_/S _4260_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4191_ hold391/Z hold767/Z _4192_/S _4191_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_94_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6901_ _6901_/D _7341_/RN _6901_/CLK _6901_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xnet633_275 net783_414/I _6994_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet633_253 net433_90/I _7016_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet633_286 net683_324/I _6983_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet633_264 net633_289/I _7005_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6832_ _6832_/D _7262_/RN _6832_/CLK _6832_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_51_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_537 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet633_297 net633_301/I _6972_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_50_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3975_ _7218_/Q _3975_/A2 _3975_/B1 input61/Z _3975_/C _3976_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_23_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6763_ _6763_/D _7262_/RN _6763_/CLK _6763_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xclkbuf_leaf_17__1374_ clkbuf_4_10_0__1374_/Z net433_59/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_176_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5714_ hold164/Z hold408/Z _5717_/S _7092_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6694_ _7262_/RN _6994_/Q _4026_/C _6694_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_176_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5645_ hold117/Z hold2/Z _5645_/S _5645_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_108_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold210 _6990_/Q hold210/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_5576_ hold25/Z hold242/Z _5581_/S _6970_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4527_ _5235_/A1 _4718_/B _3380_/I _3379_/I _5226_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_7315_ _7315_/D _7323_/RN _4103_/I1 _7315_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold243 _7372_/I hold243/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold232 _7095_/Q hold232/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold221 _4148_/Z _6716_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4458_ _3379_/I _3380_/I _4684_/B _4423_/Z _5046_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
Xhold287 _7182_/Q hold287/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7246_ _7246_/D _7341_/RN _7246_/CLK _7246_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_105_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold276 _5642_/Z _7028_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold265 _6715_/Q hold265/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold254 _5540_/Z _6941_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold298 _3475_/Z hold298/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3409_ _3409_/I _7343_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7177_ _7177_/D _7304_/RN _7177_/CLK _7177_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_98_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6128_ _7028_/Q _7150_/Q _7275_/Q _6128_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4389_ hold388/Z hold589/Z _4389_/S _6890_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6059_ _6788_/Q _6059_/A2 _6059_/A3 _6059_/B _6060_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_45_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2426 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1714 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_857 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_868 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_835 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3760_ _5534_/A1 _4246_/A2 _3786_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5430_ _5470_/A1 _5470_/A3 _5491_/A1 _5432_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3691_ _3691_/A1 _3691_/A2 _3691_/A3 _3691_/A4 _3692_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_173_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5361_ _5073_/Z _5361_/A2 _5361_/A3 _5361_/A4 _5461_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xoutput326 _6842_/Q wb_dat_o[23] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_58_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput304 _4105_/Z serial_resetn VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput315 _6850_/Q wb_dat_o[13] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_7100_ _7100_/D _7265_/RN _7100_/CLK _7100_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5292_ _5292_/A1 _5292_/A2 _5293_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4312_ hold391/Z hold764/Z _4313_/S _4312_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xoutput337 _6859_/Q wb_dat_o[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_113_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7031_ _7031_/D _7281_/RN _7031_/CLK _7031_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4243_ hold543/Z hold2/Z _4243_/S _4243_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_19_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4174_ hold708/Z hold388/Z _4174_/S _6737_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_4__1374_ clkbuf_4_2_0__1374_/Z net833_472/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_67_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6815_ _6815_/D _7281_/RN _6815_/CLK _6815_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_23_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6746_ _6746_/D _7304_/RN _6746_/CLK _6746_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_51_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3958_ _7138_/Q _3958_/A2 _3958_/B1 _6718_/Q _5544_/S _7266_/Q _3972_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_109_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3889_ _3888_/S hold875/Z _3986_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6677_ _7262_/RN _6994_/Q _4026_/C _6677_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_164_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5628_ hold391/Z hold834/Z _5635_/S _5628_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_137_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5559_ hold139/Z hold398/Z _5563_/S _5559_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_3_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_431 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7229_ _7229_/D _7265_/RN _7229_/CLK _7229_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_120_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet833_459 net833_480/I _6750_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1533 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1500 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2289 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_187_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1577 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_183_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_63__1374_ clkbuf_4_13_0__1374_/Z net633_289/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_123_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4930_ _5330_/A2 _5290_/B _4965_/A2 _6878_/Q _5123_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_18_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4861_ _4858_/Z _4861_/A2 _4861_/A3 _5428_/A2 _4865_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_177_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3812_ _6865_/Q _4378_/A1 _5893_/A3 _5546_/A2 _3877_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6600_ _6600_/I0 _7311_/Q _6603_/S _7311_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4792_ _5426_/B2 _4661_/C _4718_/B _4718_/C _4796_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_159_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3743_ _3743_/A1 _3743_/A2 _3743_/A3 _3743_/A4 _3751_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6531_ _6531_/A1 _6531_/A2 hold98/I _6584_/A1 _6584_/B _6533_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_146_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3674_ input68/Z _4262_/S _4281_/S input40/Z _3676_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6462_ _7135_/Q _6287_/Z _6300_/Z _7013_/Q _6319_/Z hold91/I _6465_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_5413_ _5282_/B _5498_/B1 _5414_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6393_ _7156_/Q _6286_/Z _6311_/C _7002_/Q _6395_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_161_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5344_ _5344_/A1 _5344_/A2 _5344_/B _5344_/C _5408_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_142_762 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput167 _4123_/Z debug_in VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput178 _6107_/A1 mgmt_gpio_oeb[16] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5275_ _5374_/A2 _5498_/A2 _5412_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_153_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput189 _3349_/ZN mgmt_gpio_oeb[26] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_102_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4226_ _4264_/A1 _5564_/A3 _4243_/S _4228_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_7014_ _7014_/D _7281_/RN _7014_/CLK _7014_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4157_ hold416/Z hold5/Z _4159_/S _4157_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_28_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4088_ _6801_/Q input58/Z _7346_/Q _4088_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_71_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6729_ _6729_/D _7262_/RN _6729_/CLK _6729_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_165_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2042 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2020 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2086 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2053 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2097 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_842 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput25 mask_rev_in[29] input25/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput14 mask_rev_in[19] input14/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput36 mgmt_gpio_in[0] input36/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_171_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold809 _7186_/Q hold809/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_115_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput69 mgmt_gpio_in[6] input69/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_10_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput47 mgmt_gpio_in[1] input47/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput58 mgmt_gpio_in[2] input58/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_182_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_835 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3390_ _6709_/Q _6708_/Q _6707_/Q _6776_/Q _4020_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_170_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5060_ _5502_/B2 _5079_/A1 _5218_/B1 _5209_/B1 _5219_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_123_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4011_ _6777_/Q _3993_/Z _4011_/A3 _4011_/B _4012_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_84_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_871 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5962_ _6787_/Q _6789_/Q _7277_/Q _5962_/B _5963_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_18_470 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4913_ _4913_/A1 _4913_/A2 _6640_/B2 _4914_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_178_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5893_ hold21/Z hold37/Z _5893_/A3 hold45/Z _5901_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_21_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4844_ _5393_/A3 _5148_/B1 _4844_/B _4844_/C _4858_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_60_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4775_ _4775_/A1 _4775_/A2 _5166_/A4 _4779_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_148_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6514_ hold32/I _6570_/A2 _6570_/B1 hold56/I _6570_/C1 _6999_/Q _6516_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_3726_ _7261_/Q _3964_/C1 _4281_/S input38/Z input55/Z _4264_/A1 _3729_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_174_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6445_ _6445_/A1 _6445_/A2 _6445_/A3 _6445_/A4 _6446_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3657_ hold91/I _3956_/A2 _3956_/B1 _7159_/Q _3659_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3588_ _7153_/Q _3866_/A2 _3953_/A2 _6999_/Q _3943_/B1 _7201_/Q _3595_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6376_ _7098_/Q _6284_/Z _6568_/B1 _7114_/Q _6390_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_121_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5327_ _5327_/A1 _5327_/A2 _5327_/B _5328_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_88_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5258_ _5397_/A1 _5327_/B _5258_/A3 _5258_/B _5427_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_113_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5189_ _5502_/A1 _5321_/A3 _5502_/B1 _5399_/B _5483_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_68_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4209_ hold391/Z hold774/Z _4210_/S _4209_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_4_13_0__1374_ clkbuf_3_6_0__1374_/Z clkbuf_4_13_0__1374_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_84_896 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_876 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_537 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet433_54 net433_54/I _7215_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet483_140 net433_94/I _7129_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet483_151 net533_163/I _7118_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet433_87 net433_87/I _7182_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet433_76 net433_76/I _7193_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_74_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet433_65 net433_65/I _7204_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet433_98 net433_98/I _7171_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_63_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1182 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4560_ _4560_/A1 _4560_/A2 _4565_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_129_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3511_ _6863_/Q _5326_/B2 hold12/Z _3511_/B2 _3511_/C hold41/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_143_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold606 _5903_/Z _7258_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4491_ _5262_/A4 _5315_/A4 _5235_/A1 _4718_/B _5290_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
Xhold617 _7363_/I hold617/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xmax_cap358 hold13/Z _5856_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
Xhold639 _6765_/Q hold639/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6230_ _6868_/Q _6262_/B1 _7275_/Q _6231_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xhold628 _6898_/Q hold628/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3442_ _3442_/A1 hold894/Z _3443_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_171_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6161_ _6161_/A1 _6161_/A2 _6161_/A3 _6161_/A4 _6161_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_3373_ _6987_/Q _3373_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_40_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5112_ _5279_/A3 _5370_/A1 _5112_/B _5370_/B _5114_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_58_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_911 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_944 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_253 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6092_ _7059_/Q _6257_/B1 _6261_/B1 _7043_/Q _6995_/Q _6258_/B1 _6095_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_69_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_966 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_977 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5043_ _5043_/A1 _5043_/A2 _5043_/B _6903_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_112_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_999 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_0_wbbd_sck _7322_/Q clkbuf_0_wbbd_sck/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_25_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6994_ _6994_/D _7265_/RN _6994_/CLK _6994_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_80_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5945_ _6211_/C _7273_/Q _7272_/Q _7271_/Q _6258_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_5876_ hold548/Z hold391/Z _5883_/S _7234_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_178_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4827_ _5355_/A2 _5199_/B _4722_/Z _5471_/B2 _4827_/C _4828_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_175_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4758_ _4922_/B _4787_/A3 _4787_/A2 _5255_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_135_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4689_ _4718_/B _4661_/C _4684_/B _5307_/B _4689_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_108_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3709_ _6996_/Q _3953_/A2 _3943_/B1 _7198_/Q _3711_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_107_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6428_ _6428_/A1 _6428_/A2 _6428_/B _7298_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_162_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6359_ _7073_/Q _6292_/Z _6571_/B1 _6985_/Q _6571_/C1 _7179_/Q _6360_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_68_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_124_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_844 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_719 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_287 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_184_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold3 hold3/I hold3/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_39_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_652 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3991_ _6707_/Q _3991_/A2 _6707_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5730_ hold25/Z _7106_/Q _5735_/S _5730_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_175_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5661_ hold5/Z hold393/Z _5663_/S _7045_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4612_ _4759_/C _4686_/B _5312_/B _4694_/B _5426_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_5592_ hold733/Z hold391/Z _5599_/S _5592_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4543_ _5466_/C _3379_/I _5034_/A2 _3380_/I _5047_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_128_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7331_ _7331_/D _6685_/Z _4089_/I1 _7331_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold403 _5605_/Z _6996_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold436 _6720_/Q hold436/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_7_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold425 _4296_/Z _6818_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7262_ _7262_/D _7262_/RN _7262_/CLK _7262_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold414 _7208_/Q hold414/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_144_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold458 _7164_/Q hold458/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4474_ _4759_/C _4694_/B _4869_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6213_ hold87/I _7129_/Q _7275_/Q _6213_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold469 _7252_/Q hold469/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold447 _4165_/Z _6730_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_171_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7193_ _7193_/D _7265_/RN _7193_/CLK _7193_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3425_ _4072_/A3 _7337_/Q _3426_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3356_ _6745_/Q _3356_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet683_302 net783_415/I _6967_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet683_313 net683_314/I _6956_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6144_ _7199_/Q _6260_/A2 _6262_/B1 _7151_/Q _6152_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_58_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xload_slew361 hold17/Z _5866_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xload_slew350 _5548_/A3 _5546_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
Xload_slew372 _5439_/C _5177_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xnet683_324 net683_324/I _6945_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_85_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6075_ _6075_/A1 _6075_/A2 _6075_/A3 _6078_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
Xnet683_346 net683_347/I _6923_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet683_335 net833_497/I _6934_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5026_ _4684_/B _4425_/Z _5026_/B _5026_/C _5287_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_57_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_796 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2608 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1907 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1929 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1918 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6977_ _6977_/D _7302_/RN _6977_/CLK _6977_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_53_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5928_ _5918_/B _5985_/A3 _5925_/B _5930_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_167_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5859_ hold528/Z hold25/Z _5865_/S _5859_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_181_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_868 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4109__17 _4109__49/I _7252_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4109__28 _4109__28/I _7241_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_150_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4109__39 _4109__48/I _7230_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_131_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_71 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_145 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4190_ _5838_/A4 _5518_/A1 _3527_/Z _6653_/A3 _4192_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_95_722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6900_ _6900_/D _7341_/RN _6900_/CLK _6900_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_63_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet633_276 net783_414/I _6993_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet633_265 net683_324/I _7004_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet633_254 net633_261/I _7015_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6831_ _6831_/D _7262_/RN _6831_/CLK _6831_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_35_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet633_287 net633_292/I _6982_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet633_298 net783_421/I _6971_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3974_ _3974_/A1 _3974_/A2 _3974_/A3 _3975_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6762_ _6762_/D _7262_/RN _6762_/CLK _6762_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_50_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5713_ hold139/Z hold153/Z _5717_/S _7091_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6693_ _7262_/RN _6994_/Q _4026_/C _6693_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_148_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5644_ hold329/Z hold58/Z _5645_/S _5644_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_163_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7314_ _7314_/D _7323_/RN _4103_/I1 _7314_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_163_248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_163_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_790 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold211 _5598_/Z _6990_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold200 _7006_/Q hold200/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_5575_ hold388/Z hold623/Z _5581_/S _6969_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold244 _5563_/Z _6959_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold222 _7193_/Q hold222/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_132_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4526_ _5301_/A2 _4661_/C _5037_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xhold233 _6932_/Q hold233/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_171_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4457_ _4669_/B _5051_/B _4056_/B _5084_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_132_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7245_ _7245_/D _7341_/RN _7245_/CLK _7245_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold277 _6988_/Q hold277/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold266 _4146_/Z _6715_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold255 _6824_/Q hold255/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold288 _5816_/Z _7182_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_172_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold299 hold299/I hold299/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3408_ hold893/Z _3412_/A3 _7343_/Q _3409_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7176_ hold69/Z _7304_/RN _7176_/CLK hold68/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6127_ _7092_/Q _7214_/Q _7275_/Q _6127_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4388_ hold391/Z hold574/Z _4389_/S _6889_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_85_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3339_ _3339_/I _4118_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_571 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6058_ _6788_/Q _7285_/Q _6059_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5009_ _3379_/I input95/Z _5153_/A2 _5282_/B _5012_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_2427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_4_1_0__1374_ clkbuf_4_1_0__1374_/I clkbuf_4_1_0__1374_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_26_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1715 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1748 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1726 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_23__1374_ _4109__51/I net433_75/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_77_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_103__1374_ clkbuf_4_1_0__1374_/Z net833_491/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_18_844 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_86__1374_ clkbuf_4_4_0__1374_/Z net433_99/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_91_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_177_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_896 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3690_ _7174_/Q _3966_/A2 _3958_/B1 _6722_/Q _3691_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_173_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5360_ _5502_/A1 _5360_/A2 _5360_/B _5360_/C _5361_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_154_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput305 _4122_/Z spi_sdi VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput316 _6851_/Q wb_dat_o[14] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5291_ _5355_/A2 _5381_/A2 _5291_/B _5291_/C _5292_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
Xoutput327 _7306_/Q wb_dat_o[24] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4311_ _5838_/A4 _5552_/A2 _6653_/A2 _6653_/A3 _4313_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
Xoutput338 _6860_/Q wb_dat_o[5] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_102_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7030_ _7030_/D _7302_/RN _7030_/CLK _7030_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4242_ hold617/Z _4241_/Z _4244_/S _4242_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4173_ hold703/Z hold391/Z _4174_/S _6736_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_714 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4109__2 _4109__2/I _7341_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_36_652 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6814_ _6814_/D _7281_/RN _6814_/CLK _6814_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_23_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6745_ _6745_/D _7304_/RN _6745_/CLK _6745_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3957_ _3957_/A1 _3957_/A2 _3957_/A3 _3957_/A4 _3957_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_50_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3888_ _3887_/Z hold879/Z _3888_/S _6913_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6676_ _7262_/RN _6994_/Q _4026_/C _6676_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_136_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5627_ _5700_/A1 _5646_/A2 _5902_/A3 _4227_/B _5635_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_5558_ hold25/Z _7367_/I _5563_/S hold26/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4509_ _5466_/B _3380_/I _3379_/I _4690_/C _5502_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_144_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7228_ _7228_/D _7265_/RN _7228_/CLK _7228_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_120_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5489_ _5489_/A1 _5489_/A2 _5489_/B1 _5502_/A2 _5490_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_120_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7159_ _7159_/D _7302_/RN _7159_/CLK _7159_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_100_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1512 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_836 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_74 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_186_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_284 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4860_ _5436_/A2 _5439_/C _5210_/B _5199_/A2 _4861_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3811_ _3811_/A1 _4246_/A1 _3460_/B _3534_/C _3938_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_60_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6530_ _6530_/A1 _6529_/Z _6531_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4791_ _4791_/A1 _4791_/A2 _4791_/A3 _4791_/A4 _4796_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_32_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3742_ _7149_/Q _3866_/A2 _3953_/A2 _6995_/Q _3743_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_70_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_833 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6461_ _7151_/Q _6562_/A2 _6562_/A3 _6561_/A3 _6465_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3673_ _7151_/Q _3866_/A2 _3961_/A2 _7005_/Q _3875_/A2 _7183_/Q _3676_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_173_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5412_ _5412_/A1 _5412_/A2 _5412_/A3 _5412_/A4 _5415_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6392_ _7252_/Q _6580_/B1 _6309_/Z _7236_/Q _6744_/Q _6579_/A2 _6395_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_5343_ _5199_/B _5376_/A1 _5343_/B _5343_/C _5432_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_2
Xoutput168 _7349_/Z irq[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput179 _3358_/ZN mgmt_gpio_oeb[17] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5274_ _5274_/A1 _5498_/A2 _5376_/C _5277_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_102_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7013_ _7013_/D _7281_/RN _7013_/CLK _7013_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4225_ hold388/Z hold720/Z _4225_/S _4225_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4156_ hold295/Z hold164/Z _4159_/S _4156_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4087_ _6810_/Q input81/Z _4087_/S _4087_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_55_257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_178_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4989_ _4989_/A1 _4989_/A2 _4989_/A3 _4992_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_51_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6728_ _6728_/D _7262_/RN _6728_/CLK _6728_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_177_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6659_ _7341_/RN _6994_/Q _4026_/C _6659_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_164_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2010 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2032 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2021 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2065 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2054 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2098 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2087 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1364 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_844 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput37 mgmt_gpio_in[10] input37/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput15 mask_rev_in[1] input15/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput26 mask_rev_in[2] input26/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_155_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput59 mgmt_gpio_in[30] input59/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput48 mgmt_gpio_in[20] input48/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_7_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4010_ _6702_/Q _3992_/Z _4011_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_96_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5961_ _6562_/A3 _6563_/A3 _6789_/Q _5962_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_18_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4912_ _4056_/B _4777_/B _5445_/A3 _5323_/A1 _4913_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_33_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5892_ hold2/Z hold49/Z _5892_/S _7249_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_61_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4843_ _5466_/B _5466_/C _5258_/A3 _4844_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_61_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4774_ _4774_/A1 _4774_/A2 _4774_/B _4779_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_20_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3725_ _7165_/Q _3878_/A2 _3875_/A2 _7181_/Q _7189_/Q _3953_/B1 _3752_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_6513_ _7169_/Q _6279_/Z _6299_/Z _7071_/Q _6575_/B1 _7055_/Q _6517_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_20_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6444_ _7206_/Q _6573_/A2 _6288_/Z _7198_/Q _6297_/Z _7044_/Q _6445_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_3656_ _7117_/Q _3969_/A2 _3968_/A2 hold93/I _3966_/A2 _7175_/Q _3661_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_161_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3587_ _7225_/Q _3975_/A2 _3938_/A2 _7209_/Q _3939_/B1 input33/Z _3595_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6375_ _6375_/A1 _6375_/A2 _6375_/B _7296_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5326_ _5326_/A1 _5326_/A2 _4365_/C _5326_/B2 _6905_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_115_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_435 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5257_ _5257_/A1 _5255_/B _5257_/B1 _5257_/B2 _5258_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_57_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_766 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4208_ _6653_/A2 _5838_/A4 _3527_/Z _5748_/A3 _4210_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_5188_ _5188_/A1 _5188_/A2 _5313_/B _5190_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_4139_ hold24/Z _7316_/Q _6863_/Q hold25/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_110_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet483_130 net683_331/I _7139_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_93_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet483_141 net433_93/I _7128_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet433_55 net433_87/I _7214_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet433_77 net433_77/I _7192_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_90_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet433_66 net433_66/I _7203_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet433_88 net433_88/I _7181_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet433_99 net433_99/I _7170_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_188_711 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3510_ _3833_/A2 _3477_/Z _3496_/B _4246_/A1 _3866_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_155_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4490_ _5301_/A2 _4661_/C _3379_/I _3380_/I _5439_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xhold607 _7353_/I hold607/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold618 _4242_/Z _6785_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_143_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold629 _4401_/Z _6898_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_6_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3441_ input58/Z _6709_/Q _6707_/Q _6774_/Q _3443_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_170_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3372_ _6995_/Q _3372_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6160_ _7093_/Q _6262_/A2 _6257_/A2 _7013_/Q _6161_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5111_ _4995_/Z _5111_/A2 _5111_/B _5112_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_912 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_923 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_934 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6091_ _6091_/A1 _6091_/A2 _6096_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_956 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_945 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_967 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_978 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5042_ _5042_/A1 _5293_/A4 _5042_/B _5042_/C _5043_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_97_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_989 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6993_ _6993_/D _7265_/RN _6993_/CLK _6993_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_19_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5944_ _5944_/I _7273_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_22_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5875_ hold21/Z hold8/Z hold37/Z hold45/Z _5883_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_178_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4826_ _4811_/Z _4826_/A2 _4826_/A3 _4826_/A4 _4827_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_21_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4757_ _4693_/Z _4706_/Z _4709_/Z _5476_/A1 _4762_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_21_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4688_ _4765_/A1 _4765_/A2 _4794_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_3708_ _6714_/Q _3942_/A2 _3975_/A2 _7222_/Q _3711_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_108_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6427_ _7297_/Q _6587_/A2 _6532_/B _6532_/C _6428_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3639_ _6917_/Q _3887_/S _3639_/B _3641_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_150_828 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6358_ _7211_/Q _6570_/A2 _6570_/B1 _7057_/Q _6570_/C1 _6993_/Q _6360_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_89_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5309_ _4759_/C _5313_/A1 _5436_/A1 _4694_/B _5440_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6289_ _6296_/A2 _7281_/Q _7280_/Q _7279_/Q _6528_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_103_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_149_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold4 hold4/I hold4/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_79_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_853 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_801 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_856 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3990_ _6708_/Q _3990_/A2 _6708_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_23_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5660_ hold164/Z hold481/Z _5663_/S _7044_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_188_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_175_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4611_ _4469_/B _4922_/B _4684_/B _5307_/B _5439_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_30_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5591_ _5700_/A1 _5655_/A4 _5646_/A2 _4227_/B _5599_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_30_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4542_ _5372_/A1 _4759_/C _4469_/B _5210_/B _5230_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_144_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7330_ _7330_/D _6684_/Z _4089_/I1 _7330_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4473_ _5136_/A2 _5223_/A1 _4922_/B _4480_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_143_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold404 _7012_/Q hold404/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7261_ _7261_/D _7341_/RN _7261_/CLK _7261_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_117_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold426 _7093_/Q hold426/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold415 _5845_/Z _7208_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold459 _6701_/Q hold459/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6212_ _6212_/A1 _7271_/Q _7272_/Q _6214_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
Xhold437 _4154_/Z _6720_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold448 _6925_/Q hold448/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3424_ _6774_/Q _3431_/B _7337_/Q _3427_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_171_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7192_ _7192_/D _7265_/RN _7192_/CLK _7192_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xnet683_303 net783_414/I _6966_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_112_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3355_ _7125_/Q _3355_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6143_ _6143_/I0 _7289_/Q _6559_/S _7289_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xload_slew373 _4624_/A2 _5439_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xnet683_314 net683_314/I _6955_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xload_slew351 hold29/Z _4405_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_6074_ _7156_/Q _6258_/A2 _6259_/B1 _7106_/Q _6232_/C _6075_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_57_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet683_325 net733_397/I _6944_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet683_336 net833_497/I _6933_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet683_347 net683_347/I _6922_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_786 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5025_ _5290_/B _5288_/A4 _5025_/A3 _5476_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_100_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_797 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_801 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1919 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1908 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6976_ _6976_/D _7281_/RN _6976_/CLK _6976_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_54_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5927_ _5927_/A1 _7270_/Q _5931_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5858_ hold731/Z hold388/Z _5865_/S _5858_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_154_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4809_ _5153_/C _5235_/A1 _5301_/A2 _5153_/B _4811_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5789_ hold164/Z hold334/Z _5792_/S _7158_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_181_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_175_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4109__29 _4109__29/I _7240_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_162_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4109__18 _4109__3/I _7251_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_134_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_185_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_856 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_46__1374_ clkbuf_4_15_0__1374_/Z net783_417/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_181_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_861 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet633_277 net633_277/I _6992_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet633_255 net783_419/I _7014_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet633_266 net633_281/I _7003_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_36_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6830_ _6830_/D _7304_/RN _6830_/CLK _6830_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xnet633_288 net633_288/I _6981_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_62_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet633_299 net783_421/I _6970_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6761_ _6761_/D _7262_/RN _6761_/CLK _6761_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_51_837 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3973_ _7048_/Q _3973_/A2 _3973_/B1 _6734_/Q _3976_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5712_ hold25/Z hold512/Z _5717_/S _7090_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_189_894 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6692_ input75/Z _6994_/Q _4026_/C _6692_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_31_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5643_ hold352/Z hold5/Z _5645_/S _5643_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5574_ hold391/Z hold806/Z _5581_/S _6968_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_129_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4525_ _5262_/A4 _5315_/A4 _5301_/A2 _5294_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
Xhold201 _5616_/Z _7006_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7313_ _7313_/D _7313_/CLK _7313_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_160_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold223 _5828_/Z _7193_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_105_828 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold212 _7255_/Q hold212/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold234 _7047_/Q hold234/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_171_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4456_ _4451_/B _4916_/A2 _4916_/A3 _4443_/Z _5087_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_116_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold278 _5596_/Z _6988_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold256 _4303_/Z _6824_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold245 _6724_/Q hold245/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold267 _7125_/Q hold267/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7244_ _7244_/D _7302_/RN _7244_/CLK _7244_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
Xhold289 _7214_/Q hold289/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4387_ hold45/Z _4405_/A2 _4405_/A3 _5893_/A3 _4389_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_3407_ _7344_/Q hold894/Z _3407_/S _7344_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7175_ _7175_/D _7304_/RN _7175_/CLK _7175_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3338_ _3338_/I _4060_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6126_ _7100_/Q _6232_/C _6266_/B _6266_/C _6138_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6057_ _6107_/B _6107_/C _6969_/Q _7275_/Q _6059_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_46_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5008_ _5008_/A1 _5008_/A2 _5008_/A3 _5012_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_2417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1749 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6959_ _6959_/D input75/Z _6959_/CLK _7372_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_81_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_577 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold790 _7009_/Q hold790/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_122_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_74 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_2_0__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/Z _4111_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_186_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_161_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput306 _4117_/Z spimemio_flash_io0_di VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput317 _6852_/Q wb_dat_o[15] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5290_ _5290_/A1 _5466_/A1 _5290_/B _5290_/C _5291_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
Xoutput328 _7307_/Q wb_dat_o[25] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4310_ hold388/Z hold636/Z _4310_/S _6830_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xoutput339 _6861_/Q wb_dat_o[6] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_99_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4241_ hold369/Z hold58/Z _4243_/S _4241_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_820 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4172_ hold45/Z _4405_/A2 hold37/Z _5745_/A4 _4174_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_110_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_726 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4109__3 _4109__3/I _7340_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_63_461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6813_ _6813_/D _7281_/RN _6813_/CLK _6813_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6744_ _6744_/D _7304_/RN _6744_/CLK _6744_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_3956_ _7122_/Q _3956_/A2 _3956_/B1 _7154_/Q _3957_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_167_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6675_ _7262_/RN _6994_/Q _4026_/C _6675_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_149_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5626_ hold2/Z hold145/Z _5626_/S _5626_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3887_ _6912_/Q _6595_/I0 _3887_/S _3887_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5557_ hold388/Z hold504/Z _5563_/S _5557_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_3_719 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5488_ _5505_/A1 _5488_/A2 _5488_/B _5488_/C _6908_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4508_ _4056_/B _5166_/A4 _4669_/B _5466_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_4439_ _4690_/C _4439_/A2 _5235_/A2 _4452_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_7227_ _7227_/D _7341_/RN _7227_/CLK _7227_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_104_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_92__1374_ clkbuf_4_3_0__1374_/Z net433_66/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_120_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7158_ _7158_/D _7302_/RN _7158_/CLK _7158_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6109_ _7003_/Q _7125_/Q _7275_/Q _6109_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7089_ _7089_/D _7302_/RN _7089_/CLK _7089_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XTAP_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_391 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2214 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1535 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1568 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_829 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_168_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_249 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_829 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_391 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_512 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3810_ _3454_/Z _3811_/A1 _4246_/A1 _3534_/C _3946_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_4790_ _4693_/Z _4706_/Z _5376_/A1 _5255_/B _4791_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_21_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3741_ _7205_/Q _3938_/A2 _3977_/B1 _7035_/Q _6987_/Q _3939_/A2 _3743_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_32_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6460_ _7247_/Q _6563_/A2 _6562_/A3 _6563_/A4 _6468_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_9_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3672_ input25/Z _3977_/A2 _3942_/A2 _6715_/Q _3672_/C _3676_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_174_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5411_ _5412_/A1 _5412_/A2 _5412_/A3 _5412_/A4 _5411_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_115_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6391_ _7090_/Q _6578_/A2 _6310_/Z _6978_/Q _6578_/C1 _7172_/Q _6396_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_63_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5342_ _5342_/A1 _5472_/A3 _5342_/A3 _5344_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_114_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5273_ _4963_/B _4962_/Z _5273_/B _5376_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7012_ _7012_/D _7281_/RN _7012_/CLK _7012_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_102_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput169 _4124_/Z irq[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_68_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4224_ hold391/Z hold851/Z _4225_/S _4224_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4155_ hold420/Z hold139/Z _4159_/S _4155_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4086_ _6808_/Q input78/Z _4087_/S _4086_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_102_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_829 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4988_ _5369_/A1 _4963_/B _5007_/A4 _4951_/C _4989_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_23_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3939_ _6984_/Q _3939_/A2 _3939_/B1 input4/Z _3941_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6727_ _6727_/D _7262_/RN _6727_/CLK _6727_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_6658_ _7341_/RN _6994_/Q _4026_/C _6658_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_180_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5609_ _5700_/A1 _5646_/A2 _5893_/A3 _4227_/B _5617_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_11_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6589_ _6874_/Q _6870_/Q _6877_/Q _6589_/B _6590_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_124_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2033 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2022 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2011 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2077 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2066 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2055 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2099 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2088 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_678 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_823 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput27 mask_rev_in[30] input27/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xinput16 mask_rev_in[20] input16/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_156_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput38 mgmt_gpio_in[11] input38/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput49 mgmt_gpio_in[21] input49/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_10_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5960_ _6306_/A3 _7277_/Q _6457_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5891_ hold58/Z hold95/Z _5892_/S _7248_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4911_ _5295_/A1 _5290_/C _5200_/B _4911_/B _4913_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_61_773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4842_ _5294_/B _5294_/C _5466_/B _5416_/A1 _4844_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_60_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4773_ _5307_/B _5011_/A2 _4773_/B _4947_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_147_845 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3724_ _7221_/Q _3975_/A2 _3940_/A2 _7213_/Q _3743_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6512_ _7233_/Q _6311_/B _6567_/B1 _7145_/Q _6517_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_173_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6443_ _7190_/Q _6274_/Z _6568_/B1 _7116_/Q _6445_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3655_ _7029_/Q _3961_/B1 _3962_/B1 _7085_/Q _3661_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_146_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3586_ _3586_/A1 _3586_/A2 _3586_/A3 _3586_/A4 _3586_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_6374_ _7295_/Q _6587_/A2 _6532_/B _6532_/C _6375_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5325_ _4365_/C _5325_/A2 _5293_/Z _5324_/Z _5326_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_5256_ _5256_/A1 _5256_/A2 _5256_/A3 _5335_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_69_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4207_ hold717/Z hold388/Z _4207_/S _4207_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5187_ _5295_/A1 _5466_/A1 _5187_/B _5466_/B _5313_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_84_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4138_ hold388/Z hold697/Z _4150_/S _4138_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4069_ _6709_/Q _6708_/Q _6774_/Q _3445_/Z _4069_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_189_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_180_623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet483_120 net433_88/I _7149_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_59_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet483_131 net833_498/I _7138_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet483_142 net533_163/I _7127_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_47_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet433_56 net433_56/I _7213_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet433_78 _4109__6/I _7191_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet433_67 net433_67/I _7202_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_47_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet433_89 net433_89/I _7180_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_103_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold608 _4259_/Z _6796_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3440_ hold387/Z input58/Z _3440_/S _7328_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_144_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xmax_cap349 _5546_/A2 _6653_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_16
Xhold619 _7350_/I hold619/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3371_ _7003_/Q _3371_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_170_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5110_ _5372_/B _5279_/A3 _5110_/B _5498_/C _5111_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_6090_ _7011_/Q _6257_/A2 _6256_/A2 _7051_/Q _6091_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_69_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_902 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_913 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_924 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_935 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5041_ _5041_/A1 _5041_/A2 _5041_/A3 _5042_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_112_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_946 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_979 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_0_wb_clk_i wb_clk_i clkbuf_0_wb_clk_i/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_65_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6992_ _6992_/D _7281_/RN _6992_/CLK _6992_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_25_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_537 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_179_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5943_ _5942_/Z _6789_/Q _7273_/Q _5974_/B1 _5944_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5874_ hold199/Z hold2/Z _5874_/S _7233_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_61_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4825_ _5468_/A1 _5471_/B2 _5468_/C _4825_/A4 _4826_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_21_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4756_ _4693_/Z _4706_/Z _4709_/Z _5093_/B _4762_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_146_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4687_ _4487_/Z _4684_/B _4661_/C _4718_/B _4765_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_3707_ _7134_/Q _3945_/A2 _3977_/B1 _7036_/Q input24/Z _3977_/A2 _3711_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_162_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6426_ _6426_/A1 _6426_/A2 _6971_/Q _6584_/A1 _6584_/B _6428_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_3638_ _3887_/S _6602_/A1 _3639_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_161_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6357_ _6357_/A1 _6357_/A2 _6357_/A3 _6357_/A4 _6366_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3569_ _3511_/C _3519_/Z _5534_/A1 _3604_/A2 _3850_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_103_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5308_ _5303_/Z _5397_/B _5308_/A3 _5308_/A4 _5308_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_130_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6288_ _7279_/Q _7278_/Q _6457_/A3 _6561_/A3 _6288_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_0_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5239_ _5471_/A1 _5153_/C _5239_/B _5239_/C _5492_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_187_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_289 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_130_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_678 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold5 hold5/I hold5/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_94_437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_894 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_69__1374_ _4109__12/I net633_292/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_90_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4610_ _4610_/A1 _4609_/Z _4616_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_175_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5590_ hold2/Z hold107/Z _5590_/S _5590_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4541_ _5235_/A2 _5034_/A2 _5290_/C _5272_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_117_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4472_ _4421_/Z _4437_/Z _4759_/C _4479_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_156_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold405 _5623_/Z _7012_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold427 _6812_/Q hold427/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold416 _6723_/Q hold416/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7260_ _7260_/D _7302_/RN _7260_/CLK _7260_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_171_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold449 _7149_/Q hold449/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7191_ _7191_/D _7265_/RN _7191_/CLK _7191_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_143_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6211_ _6232_/C _7103_/Q _6211_/B _6211_/C _6212_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
Xhold438 _7159_/Q hold438/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3423_ _3431_/B _4072_/A3 _3429_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_710 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6142_ _6788_/Q _6142_/A2 _6142_/A3 _6142_/B _6143_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
Xnet683_304 net783_415/I _6965_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3354_ _7133_/Q _3354_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xload_slew352 hold29/Z _5718_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xload_slew363 hold17/Z _5884_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xnet683_315 net683_317/I _6954_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_97_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6073_ _7132_/Q _6257_/A2 _6260_/B1 _7114_/Q _6075_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xnet683_337 net833_483/I _6932_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet683_326 net783_421/I _6943_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_754 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5024_ _5024_/A1 _5024_/A2 _5024_/A3 _5409_/C _5024_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_85_437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xnet683_348 net683_349/I _6921_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1909 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6975_ hold99/Z _7304_/RN _6975_/CLK hold98/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_54_868 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5926_ _5926_/A1 _5926_/A2 _7269_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_179_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5857_ hold873/Z hold391/Z _5865_/S _5857_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_166_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4808_ _5267_/C _4808_/A2 _5153_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_21_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5788_ hold139/Z hold271/Z _5792_/S _5788_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4739_ _5327_/B _5307_/B _4794_/A2 _5250_/C _5329_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_119_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6409_ _7229_/Q _6311_/B _6567_/B1 _7141_/Q _6410_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4109__19 _4109__24/I _7250_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_134_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_687 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_827 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_829 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_opt_1_0__1374_ clkbuf_4_8_0__1374_/Z clkbuf_opt_1_0__1374_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_4_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet633_256 net633_280/I _7013_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_90_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet633_267 net783_420/I _7002_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet633_278 net633_290/I _6991_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet633_289 net633_289/I _6980_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_90_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6760_ _6760_/D _7262_/RN _6760_/CLK _6760_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_93_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3972_ _3957_/Z _3972_/A2 _3960_/Z _3972_/A4 _3983_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5711_ hold388/Z hold777/Z _5717_/S _7089_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6691_ input75/Z _6994_/Q _4026_/C _6691_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_176_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5642_ hold275/Z hold164/Z _5645_/S _5642_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_163_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5573_ _5700_/A1 _5856_/A2 _5573_/A3 _5535_/B _5581_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_4524_ _3379_/I _3380_/I _4718_/B _5436_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_117_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold202 _7005_/Q hold202/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7312_ _7312_/D _7313_/CLK _7312_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold213 _7037_/Q hold213/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold235 _6747_/Q hold235/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold224 _6826_/Q hold224/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_171_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7243_ _7243_/D _7265_/RN _7243_/CLK _7243_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4455_ _4960_/C _5082_/A1 _5082_/A2 _5051_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
Xhold257 _6939_/Q hold257/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold246 _4158_/Z _6724_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold268 _5752_/Z _7125_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_113_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4386_ hold388/Z hold624/Z _4386_/S _4386_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3406_ _3446_/A2 _6707_/Q _3407_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xhold279 _6929_/Q hold279/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7174_ _7174_/D _7304_/RN _7174_/CLK _7174_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3337_ _4774_/B _5166_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_8
XFILLER_131_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6125_ _6125_/A1 _6125_/A2 _6124_/Z _6125_/A4 _6139_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_573 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6056_ _7275_/Q _6056_/A2 _6056_/B _6056_/C _6059_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5007_ _5353_/A3 _4963_/B _4926_/C _5007_/A4 _5008_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XTAP_2418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2429 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_52__1374_ clkbuf_4_12_0__1374_/Z net633_280/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6958_ _6958_/D input75/Z _6958_/CLK _7371_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5909_ hold58/Z hold80/Z _5910_/S hold81/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6889_ _6889_/D _7341_/RN _6889_/CLK _6889_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_22_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_871 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_182_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold791 _5620_/Z _7009_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold780 _7104_/Q hold780/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_89_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_189_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput307 _4118_/ZN spimemio_flash_io1_di VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_181_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput329 _7308_/Q wb_dat_o[26] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput318 _6835_/Q wb_dat_o[16] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_5_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4240_ hold667/Z _4239_/Z _4244_/S _4240_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4171_ hold388/Z hold647/Z _4171_/S _4171_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4109__4 _4109__4/I _7265_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_36_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6812_ _6812_/D input75/Z _6812_/CLK _6812_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_63_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6743_ _6743_/D _7304_/RN _6743_/CLK _6743_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_3955_ _6922_/Q _3681_/Z _3955_/B1 _6760_/Q _6772_/Q _3955_/C2 _3957_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_177_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_843 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6674_ _7262_/RN _6994_/Q _4026_/C _6674_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_50_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5625_ hold58/Z hold318/Z _5626_/S _5625_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3886_ _3886_/A1 _3845_/Z _3886_/A3 _3886_/A4 _6595_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_136_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5556_ hold391/Z hold506/Z _5563_/S _5556_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4507_ _4451_/B _4774_/B _4916_/A2 _4916_/A3 _4624_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_144_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5487_ _5487_/A1 _5487_/A2 _5487_/A3 _5486_/Z _5488_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_105_604 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4438_ _5004_/A1 input95/Z _4718_/B _4661_/C _5223_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_144_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7226_ _7226_/D _7265_/RN _7226_/CLK _7226_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_98_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4369_ hold45/Z _4405_/A2 _5838_/A2 _4378_/A1 _4371_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_7157_ _7157_/D _7302_/RN _7157_/CLK _7157_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_7088_ _7088_/D _7265_/RN _7088_/CLK _7088_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_6108_ _7091_/Q _7213_/Q _7275_/Q _6108_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6039_ _7163_/Q _6261_/B1 _6039_/B _6041_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_2226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_27_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1569 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_168_876 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet533_200 net433_68/I _7069_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_182_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_568 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3740_ _3737_/Z _3740_/A2 _3740_/A3 _3740_/A4 _3751_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_186_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3671_ _7239_/Q _3943_/A2 _3977_/B1 _7037_/Q _3980_/B1 _6981_/Q _3677_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_174_879 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5410_ _4956_/C _5410_/A2 _5410_/A3 _5498_/B1 _5412_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6390_ _6390_/A1 _6390_/A2 _6390_/A3 _6390_/A4 _6397_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_173_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5341_ _5471_/A1 _5199_/B _4722_/Z _5471_/B2 _5342_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_56_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5272_ _5445_/A3 _5489_/A1 _5272_/B _5272_/C _5273_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_114_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7011_ _7011_/D _7281_/RN _7011_/CLK _7011_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_102_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4223_ _5838_/A4 _5518_/A1 _3527_/Z _5745_/A4 _4225_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_96_863 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4154_ hold436/Z hold25/Z _4159_/S _4154_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4085_ _6807_/Q input80/Z _4087_/S _4085_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_28_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4987_ _4963_/B _4995_/A4 _4951_/C _4922_/B _5372_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_6726_ _6726_/D _7262_/RN _6726_/CLK _6726_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_3938_ _7202_/Q _3938_/A2 _3938_/B1 _6883_/Q _3938_/C _3941_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_176_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6657_ _7341_/RN _6994_/Q _4026_/C _6657_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_3869_ _7203_/Q _3938_/A2 _3980_/B1 _6977_/Q _3946_/B1 _6882_/Q _3871_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_5608_ hold2/Z hold381/Z _5608_/S _5608_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6588_ _6559_/S _6588_/A2 _6588_/B _7304_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_164_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5539_ hold139/Z hold251/Z _5543_/S _5539_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_127_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7209_ _7209_/D _7302_/RN _7209_/CLK _7209_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_47_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2001 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2034 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2023 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_160_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2056 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2045 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1322 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2089 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1355 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1399 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput28 mask_rev_in[31] input28/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput17 mask_rev_in[21] input17/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput39 mgmt_gpio_in[12] input39/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_182_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5890_ hold5/Z hold137/Z _5892_/S _7247_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4910_ _5489_/A1 _5404_/B1 _4910_/B _4910_/C _4911_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_93_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4841_ _5439_/A2 _4841_/A2 _5298_/B _5199_/A2 _5485_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_60_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4772_ _4684_/B _4425_/Z _5307_/B _4773_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_6511_ _7119_/Q _6511_/A2 _6561_/A3 _6563_/A4 _6517_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3723_ input23/Z _5727_/A3 _5748_/A3 _5532_/A3 _3743_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_174_654 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3654_ _3654_/A1 _3654_/A2 _3654_/A3 _3654_/A4 _3654_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_6442_ _7230_/Q _6311_/B _6567_/B1 _7142_/Q _6445_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_9_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3585_ _7145_/Q _3958_/A2 _3958_/B1 _6725_/Q _3969_/B1 _6749_/Q _3586_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6373_ _6969_/Q _6584_/A1 _6373_/B _6584_/B _6375_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_142_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5324_ _5479_/A2 _5324_/A2 _5444_/B _5324_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_115_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5255_ _5439_/A2 _5093_/B _5255_/B _5468_/B _5256_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_102_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4206_ hold822/Z hold391/Z _4207_/S _4206_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5186_ _5466_/B _5426_/A1 _5258_/A3 _5187_/B _5186_/B2 _5188_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_28_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4137_ hold387/Z hold900/Z _6863_/Q _4137_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_110_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4068_ _4068_/A1 _6589_/B _6870_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6709_ _6709_/D _6664_/Z _7346_/CLK _6709_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_22_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_164_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet483_121 net433_81/I _7148_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet483_110 net533_176/I _7159_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_74_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet483_143 net433_99/I _7126_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet483_132 _4109__44/I _7137_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet433_57 net433_89/I _7212_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet433_68 net433_68/I _7201_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_90_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet433_79 _4109__8/I _7190_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_179_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold609 _6884_/Q hold609/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_10_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_29__1374_ clkbuf_4_11_0__1374_/Z net433_71/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_109_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_109__1374_ net733_398/I net683_347/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3370_ _7011_/Q _3370_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_111_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_903 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_914 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5040_ _3379_/I _5026_/C _5315_/A4 _5153_/A2 _5409_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_936 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_958 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_947 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_969 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6991_ _6991_/D _7281_/RN _6991_/CLK _6991_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_93_674 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_847 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5942_ _7273_/Q _6266_/B _5942_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_34_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5873_ hold301/Z hold58/Z _5874_/S _7232_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_178_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4824_ _5372_/A1 _5471_/B2 _5468_/C _4825_/A4 _4826_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4755_ _4755_/A1 _4755_/A2 _4755_/A3 _4755_/A4 _4762_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_159_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3706_ _7004_/Q _3961_/A2 _3706_/B _3706_/C _3714_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4686_ _5262_/A4 _5315_/A4 _4686_/B _4690_/C _4720_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_6425_ _6425_/A1 _6424_/Z _6426_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3637_ _6716_/Q _3942_/A2 _3637_/B _3637_/C _6602_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_161_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6356_ _7187_/Q _6274_/Z _6568_/B1 _7113_/Q _6357_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3568_ _3833_/A2 _3477_/Z _3496_/B _3831_/A2 _3969_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_5307_ _5312_/A1 _5313_/A1 _5307_/B _5312_/C _5397_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3499_ _3460_/B _3534_/C _3833_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_6287_ _7278_/Q _6457_/A3 _6561_/A3 _6324_/A1 _6287_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_102_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5238_ _5238_/A1 _5424_/A3 _5367_/B _5326_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5169_ _5298_/B _5177_/A1 _5169_/B1 _5502_/B1 _5390_/B _5172_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_56_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold6 hold6/I hold6/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_90_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4540_ _5235_/A1 _4718_/B input95/Z _5004_/A1 _5369_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_144_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_184_793 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4471_ _4479_/A2 _4951_/A2 _4502_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_144_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold417 _4157_/Z _6723_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold406 _6987_/Q hold406/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7190_ _7190_/D _7341_/RN _7190_/CLK _7190_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_125_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6210_ _6206_/Z _6210_/A2 _6210_/A3 _6210_/A4 _6214_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xhold428 _4289_/Z _6812_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3422_ _3416_/S _3418_/S _3422_/A3 _3422_/A4 _3431_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
Xhold439 _7117_/Q hold439/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XTAP_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6141_ _6788_/Q _7288_/Q _6142_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3353_ _7141_/Q _3353_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_98_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_711 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet683_305 net783_415/I _6964_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_140_863 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet683_316 net683_317/I _6953_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_97_265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xload_slew353 _5893_/A3 _5748_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xload_slew364 hold21/Z _5856_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_6072_ _7140_/Q _6259_/A2 _6257_/B1 _7180_/Q _6075_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xnet683_338 net683_349/I _6931_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet683_327 net783_421/I _6942_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_766 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5023_ _5476_/A1 _4776_/Z _5023_/A3 _5091_/B _5409_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
Xnet683_349 net683_349/I _6920_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6974_ _6974_/D _7304_/RN _6974_/CLK _6974_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_53_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5925_ _5920_/B _5925_/A2 _5925_/B _5926_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_110_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5856_ _5856_/A1 _5856_/A2 _3527_/Z _4227_/B _5865_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_4807_ _5262_/A4 _5301_/A2 _5235_/A1 _3380_/I _5258_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_186_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5787_ hold25/Z hold533/Z _5792_/S _7156_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_175_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4738_ _5244_/A2 _4825_/A4 _4750_/A3 _4750_/A4 _5247_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_181_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_793 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4669_ _4669_/A1 _4710_/C _4669_/B _4727_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_107_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6408_ _7107_/Q _6285_/Z _6564_/C1 _7083_/Q _6408_/C _6410_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_122_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_12__1374_ clkbuf_4_8_0__1374_/Z _4109__24/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6339_ _6339_/A1 _6339_/A2 _6339_/A3 _6340_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_103_543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_75__1374_ clkbuf_4_5_0__1374_/Z net783_421/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_130_340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet633_257 net633_273/I _7012_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet633_268 net783_420/I _7001_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet633_279 net783_426/I _6990_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_90_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3971_ input11/Z _3971_/A2 _3971_/B _3971_/C _3972_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_35_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_874 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_863 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5710_ hold391/Z hold766/Z _5717_/S _7088_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_62_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6690_ input75/Z _6994_/Q _4026_/C _6690_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_86_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5641_ _5645_/S _5641_/A2 _5641_/B hold509/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5572_ hold2/Z _6967_/Q hold38/Z hold39/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_117_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4523_ _5502_/A1 _5484_/A4 _5052_/A2 _5351_/A1 _5464_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_163_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7311_ _7311_/D _7313_/CLK _7311_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7242_ _7242_/D _7341_/RN _7242_/CLK _7242_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
Xhold203 _5615_/Z _7005_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold214 _5652_/Z _7037_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold225 _4305_/Z _6826_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4454_ _4840_/A1 _4777_/A2 _4454_/B _5459_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_144_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold247 _7035_/Q hold247/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold236 _4187_/Z _6747_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold258 _5538_/Z _6939_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold269 _6823_/Q hold269/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4385_ hold391/Z hold626/Z _4386_/S _4385_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3405_ _6709_/Q _6708_/Q _6774_/Q _3446_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_7173_ _7173_/D _7304_/RN _7173_/CLK _7173_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3336_ _4451_/B _4669_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_4
XFILLER_140_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6124_ _6124_/A1 _6124_/A2 _6124_/A3 _6124_/A4 _6124_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XTAP_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_541 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6055_ _6055_/A1 _6055_/A2 _6055_/A3 _6055_/A4 _6056_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5006_ _5369_/A1 _4963_/B _4926_/C _5007_/A4 _5008_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XTAP_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6957_ hold6/Z input75/Z _6957_/CLK _7370_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_1729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5908_ hold5/Z hold103/Z _5910_/S _5908_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6888_ _6888_/D _7341_/RN _6888_/CLK _6888_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_14_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5839_ hold391/Z hold856/Z _5846_/S _5839_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_108_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_616 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold781 _6808_/Q hold781/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold770 _4215_/Z _6766_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold792 _7138_/Q hold792/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_162_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_896 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput308 _7375_/Z spimemio_flash_io2_di VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_114_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput319 _6836_/Q wb_dat_o[17] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_4_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4170_ hold391/Z hold715/Z _4171_/S _4170_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4109__5 _4109__6/I _7264_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_91_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6811_ _6811_/D input75/Z _6811_/CLK _6811_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_35_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3954_ _3954_/A1 _3954_/A2 _3954_/A3 _3954_/A4 _3984_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_6742_ _6742_/D _7304_/RN _6742_/CLK _6742_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_32_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6673_ input75/Z _6994_/Q _4026_/C _6673_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_3885_ _3885_/A1 _3885_/A2 _3885_/A3 _3884_/Z _3886_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_50_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5624_ hold5/Z hold372/Z _5626_/S _5624_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5555_ hold21/Z hold37/Z _5838_/A2 hold45/Z _5563_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_4506_ _5262_/A4 _5315_/A4 _4718_/B _4661_/C _5349_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_144_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5486_ _5486_/A1 _5486_/A2 _5486_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_104_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4437_ _5004_/A1 input95/Z _4718_/B _4661_/C _4437_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_160_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7225_ _7225_/D _7302_/RN _7225_/CLK _7225_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_99_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7156_ _7156_/D _7304_/RN _7156_/CLK _7156_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_6107_ _6107_/A1 _7275_/Q _6107_/B _6107_/C _6112_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4368_ hold388/Z hold572/Z _4368_/S _4368_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3319_ hold40/Z _5326_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_7087_ _7087_/D _7281_/RN _7087_/CLK _7087_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4299_ _4262_/S _5564_/A3 _4227_/B _4307_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_101_844 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_393 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6038_ _6235_/A1 _6038_/A2 _6038_/B1 _6235_/B2 _6038_/C _6039_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_27_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2249 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1537 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_187_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_10_500 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_183_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet533_201 net433_58/I _7068_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_136_752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_393 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2750 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3670_ _6989_/Q _3939_/A2 _3946_/A2 _7021_/Q _7191_/Q _3953_/B1 _3677_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_9_364 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_3_1_0__1374_ clkbuf_0__1374_/Z clkbuf_4_3_0__1374_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_5340_ _5339_/Z _5340_/A2 _5344_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5271_ _5271_/A1 _5353_/A3 _5330_/A2 _5271_/A4 _5498_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_99_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7010_ _7010_/D _7281_/RN _7010_/CLK _7010_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4222_ hold388/Z hold653/Z _4222_/S _4222_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4153_ hold755/Z hold388/Z _4159_/S _4153_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4084_ _4084_/I _4084_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_83_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4986_ _5223_/A1 _4963_/B _4926_/C _4955_/B _4989_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_3937_ _3937_/A1 _3937_/A2 _3937_/A3 _3937_/A4 _3937_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_6725_ _6725_/D _7304_/RN _6725_/CLK _6725_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_51_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6656_ _7341_/RN _6994_/Q _4026_/C _6656_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_3868_ _3868_/A1 _3868_/A2 _3868_/A3 _3868_/A4 _3868_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_20_853 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5607_ hold58/Z hold143/Z _5608_/S _5607_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6587_ _5917_/B _6587_/A2 _7304_/Q _6588_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3799_ _6763_/Q _5748_/A3 _5546_/A2 _3527_/Z _3855_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5538_ hold164/Z hold257/Z _5543_/S _5538_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_105_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5469_ _5263_/Z _5469_/A2 _5469_/A3 _5469_/A4 _5469_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_7208_ _7208_/D _7302_/RN _7208_/CLK _7208_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_101_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7139_ _7139_/D _7302_/RN _7139_/CLK _7139_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_143_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2024 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2013 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2002 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2068 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2057 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2046 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1356 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_168_652 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput18 mask_rev_in[22] input18/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_155_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput29 mask_rev_in[3] input29/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_171_828 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4840_ _4840_/A1 _5208_/B2 _4451_/B _4774_/B _5298_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XTAP_2591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4771_ _4684_/B _4425_/Z _5307_/B _5026_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_6510_ hold49/I _6563_/A2 _6562_/A3 _6563_/A4 _6516_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_1890 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3722_ _7043_/Q _5655_/A4 _5884_/A2 hold29/I _3745_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_146_335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3653_ _7223_/Q _3975_/A2 _3940_/A2 _7215_/Q _3653_/C _3654_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_6441_ _7100_/Q _6284_/Z _6294_/Z _7036_/Q _6441_/C _6445_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_6372_ _6372_/A1 _6372_/A2 _6371_/Z _6373_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_173_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5323_ _5323_/A1 _5404_/B1 _5323_/B _5323_/C _5444_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_3584_ _7129_/Q _3956_/A2 _3959_/A2 _6733_/Q _3850_/B1 input10/Z _3586_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_114_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5254_ _5254_/A1 _5490_/A2 _5259_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5185_ _5502_/A1 _5399_/B _5502_/B1 _5439_/B _5401_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4205_ _5838_/A4 _5518_/A1 _5838_/A2 hold299/Z _4207_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_110_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4136_ hold391/Z hold799/Z _4150_/S _4136_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_29_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4067_ _4067_/A1 _6870_/Q _6589_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4969_ _4969_/A1 _4969_/A2 _4969_/A3 _4975_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_11_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6708_ _6708_/D _6663_/Z _7346_/CLK _6708_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
X_6639_ _6880_/Q _6639_/A2 _6639_/B1 _6879_/Q _6641_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_138_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet483_111 net833_456/I _7158_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_170_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet483_122 net433_91/I _7147_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet483_133 net433_77/I _7136_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet483_144 net833_480/I _7125_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_170_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet433_58 net433_58/I _7211_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet433_69 _4109__4/I _7200_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_16_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_403 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_904 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_915 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_926 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_937 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_959 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_948 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6990_ _6990_/D _7281_/RN _6990_/CLK _6990_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_93_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5941_ _5941_/I _7272_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_19_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5872_ hold345/Z hold5/Z _5874_/S _7231_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_786 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4823_ _5471_/A1 _4823_/A2 _4823_/B _4826_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_21_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4754_ _5262_/A4 _5136_/B1 _3380_/I _5037_/A1 _4755_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_147_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3705_ _3705_/A1 _3705_/A2 _3705_/A3 _3705_/A4 _3706_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_174_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4685_ _4686_/B _4759_/B1 _4765_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_146_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6424_ _6584_/A1 _6424_/A2 _6424_/A3 _6424_/A4 _6424_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_3636_ _3636_/A1 _3636_/A2 _3636_/A3 _3636_/A4 _3637_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
X_3567_ _3644_/A2 _3460_/B _3498_/B _3831_/A2 _3981_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_108_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6355_ _7227_/Q _6311_/B _6567_/B1 _7139_/Q _6357_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_1_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6286_ _6561_/A3 _6406_/A4 _6310_/A4 _6306_/A3 _6286_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
X_5306_ _5308_/A4 _5308_/A3 _5502_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5237_ _4683_/B _5424_/A2 _5343_/C _5367_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_3498_ _6863_/Q hold16/Z _3498_/B _3498_/C hold17/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_124_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5168_ _5347_/A1 _5295_/A1 _5466_/A1 _5327_/B _5312_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_84_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5099_ _4437_/Z _5107_/A1 _5372_/B _5489_/A1 _5373_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_72_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4119_ _6778_/Q _6775_/Q _4119_/B _4120_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_72_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_4_4_0__1374_ clkbuf_4_5_0__1374_/I clkbuf_4_4_0__1374_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_25_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_35__1374_ clkbuf_4_14_0__1374_/Z _4109__29/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_214 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_98__1374_ clkbuf_4_4_0__1374_/Z net683_331/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_138_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_149_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_874 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_801 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold7 hold7/I hold7/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_74_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_848 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4470_ _4421_/Z _4437_/Z _5315_/A4 _4469_/B _4479_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_128_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold418 _6979_/Q hold418/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold407 _5595_/Z _6987_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_171_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold429 _6729_/Q hold429/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3421_ _4020_/A1 _3421_/A2 _6777_/Q _3421_/B _3422_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_171_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3352_ _7149_/Q _3352_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_98_723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6140_ _6107_/B _6107_/C _6972_/Q _7275_/Q _6142_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XTAP_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xload_slew365 hold21/Z _5700_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_140_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet683_306 net683_320/I _6963_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_100_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet683_317 net683_317/I _6952_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_97_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xload_slew354 hold41/Z _5893_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_6071_ _6071_/A1 _6080_/A2 _6071_/B _6071_/C _6084_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
Xnet683_328 net733_397/I _6941_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_745 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xload_slew343 hold299/Z _5784_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_5022_ _5253_/A1 _5091_/B _5091_/C _5235_/A1 _5024_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_140_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet683_339 net683_349/I _6930_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_789 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6973_ _6973_/D _7304_/RN _6973_/CLK _6973_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5924_ _7269_/Q _5931_/A1 _5918_/B _5985_/A3 _5926_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_5855_ hold2/Z hold32/Z _5855_/S hold33/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4806_ _5315_/A4 _4718_/B _4661_/C _3379_/I _5199_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_5786_ hold388/Z hold776/Z _5792_/S _7155_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_163_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4737_ _4737_/A1 _4737_/A2 _5467_/A1 _4737_/A4 _4748_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_175_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4668_ _4922_/B _4775_/A1 _4778_/A4 _4787_/A3 _4727_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_134_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6407_ _7099_/Q _6563_/A3 _6561_/A3 _6563_/A4 _6408_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_3619_ _3619_/A1 _3619_/A2 _3619_/A3 _3636_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4599_ _5223_/A2 _3380_/I _3379_/I _4690_/C _4600_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_134_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6338_ _7194_/Q _6288_/Z _6567_/B1 _7138_/Q _6339_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_103_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6269_ _6107_/B _6107_/C _6830_/Q _7275_/Q _6271_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_48_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_185_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_820 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_726 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet633_258 net783_419/I _7011_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_62_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_831 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet633_269 net683_324/I _7000_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3970_ _3970_/A1 _3970_/A2 _3970_/A3 _3970_/A4 _3971_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_35_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_842 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5640_ _5646_/A2 _5640_/A2 _4227_/B hold139/Z _5641_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xclkbuf_leaf_81__1374_ clkbuf_4_5_0__1374_/Z net433_94/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5571_ hold58/Z _6966_/Q hold38/Z hold59/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_145_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4522_ _5208_/B2 _4661_/C _3380_/I _3379_/I _5052_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_163_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7310_ _7310_/D _7313_/CLK _7310_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7241_ hold46/Z _7265_/RN _7241_/CLK _7241_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4453_ _5082_/A1 _5082_/A2 _4454_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_156_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold215 _7086_/Q hold215/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold204 _7085_/Q hold204/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold226 _7262_/Q hold226/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold248 _5650_/Z _7035_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold259 _7004_/Q hold259/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold237 _6973_/Q hold237/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3404_ _3991_/A2 _6778_/Q _4054_/B _3404_/B hold886/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_131_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4384_ _4405_/A3 hold45/Z _5546_/A2 _5655_/A4 _4386_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_7172_ _7172_/D _7304_/RN _7172_/CLK _7172_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_3335_ _7281_/Q _5975_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_4
X_6123_ _7068_/Q _6258_/C1 _6261_/A2 _7004_/Q _6124_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6054_ _7211_/Q _6262_/A2 _6257_/B1 _7179_/Q _6055_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_85_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5005_ _5005_/A1 _4942_/Z _5005_/B _5005_/C _5008_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_100_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3340__1 _3340__1/I _6643_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6956_ _6956_/D input75/Z _6956_/CLK _7369_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_1719 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5907_ hold164/Z hold226/Z _5910_/S _5907_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_179_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6887_ _6887_/D _7341_/RN _6887_/CLK _6887_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5838_ _5856_/A1 _5838_/A2 _3527_/Z _5838_/A4 _5846_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_136_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5769_ hold25/Z hold350/Z _5774_/S _5769_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_163_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold760 _6985_/Q hold760/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold782 _4285_/Z _6808_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold771 _6738_/Q hold771/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_122_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold793 _5767_/Z _7138_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput309 _7376_/Z spimemio_flash_io3_di VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_5_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_796 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_867 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4109__6 _4109__6/I _7263_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_75_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6810_ _6810_/D input75/Z _6810_/CLK _6810_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_35_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3953_ _6992_/Q _3953_/A2 _3953_/B1 _7186_/Q _3953_/C _3954_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_6741_ _6741_/D _7262_/RN _6741_/CLK _6741_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_188_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3884_ _3884_/A1 _3884_/A2 _3884_/A3 _3884_/A4 _3884_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
X_6672_ input75/Z _6994_/Q _4026_/C _6672_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_5623_ hold164/Z hold404/Z _5626_/S _5623_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5554_ hold388/Z hold650/Z _5554_/S _6951_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4505_ _5301_/A2 _5235_/A1 _3379_/I _3380_/I _5404_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_5485_ _5485_/A1 _5299_/B _5485_/A3 _5486_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4436_ _3379_/I _3380_/I _5235_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_7224_ _7224_/D _7341_/RN _7224_/CLK _7224_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_117_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4367_ hold391/Z hold575/Z _4368_/S _4367_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7155_ _7155_/D _7262_/RN _7155_/CLK _7155_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_6106_ _6106_/A1 _6106_/A2 _6106_/A3 _6110_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_99_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3318_ _6777_/Q _4073_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_4
X_7086_ _7086_/D _7281_/RN _7086_/CLK _7086_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_86_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4298_ hold2/Z hold543/Z _4298_/S _4298_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_100_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6037_ _7203_/Q _6233_/A2 _6233_/B1 _7195_/Q _6266_/B _7187_/Q _6038_/B1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XTAP_2217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6939_ _6939_/D _7304_/RN _6939_/CLK _6939_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XPHY_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_179_182 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold590 _6881_/Q hold590/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_173_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2762 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_403 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5270_ _5270_/A1 _5270_/A2 _5343_/B _5325_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4221_ hold391/Z hold735/Z _4222_/S _4221_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4152_ hold836/Z hold391/Z _4159_/S _4152_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4083_ _7245_/Q input82/Z _4087_/S _4084_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_102_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_431 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4985_ _4985_/A1 _4985_/A2 _4985_/A3 _4989_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_168_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3936_ _6946_/Q hold37/I _5856_/A2 _5546_/A2 _3974_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6724_ _6724_/D _7304_/RN _6724_/CLK _6724_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_20_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3867_ _7211_/Q _3940_/A2 _3867_/B _3868_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6655_ hold388/Z hold583/Z _6655_/S _6655_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_165_848 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5606_ hold5/Z hold122/Z _5608_/S _5606_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6586_ _6788_/Q _7303_/Q _6586_/B _6588_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3798_ _6751_/Q _5784_/A3 _3527_/Z _5518_/A1 _3855_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_180_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5537_ _5535_/B _5573_/A3 _5546_/A2 _5802_/A2 _5543_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_133_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_160_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5468_ _5468_/A1 _5489_/A1 _5468_/B _5468_/C _5469_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_7207_ _7207_/D _7302_/RN _7207_/CLK _7207_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4419_ _4412_/Z _4414_/Z _4417_/Z _4774_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_160_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5399_ _5439_/A1 _5439_/A2 _5399_/B _5439_/C _5401_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_101_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7138_ _7138_/D _7304_/RN _7138_/CLK _7138_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_143_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7069_ _7069_/D _7265_/RN _7069_/CLK _7069_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_74_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2025 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2014 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2003 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2058 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2069 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1324 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput19 mask_rev_in[23] input19/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_136_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_285 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1880 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4770_ _4770_/A1 _4770_/A2 _4770_/A3 _5256_/A1 _4780_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_174_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3721_ _6930_/Q _5745_/A4 _5518_/A1 _5552_/A2 _3740_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_147_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3652_ _3652_/I _3653_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6440_ _6440_/A1 _6440_/A2 _6440_/A3 _6446_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_173_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6371_ _6584_/A1 _6371_/A2 _6371_/A3 _6371_/A4 _6371_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_61_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3583_ _7177_/Q _3966_/A2 _3956_/B1 _7161_/Q _7119_/Q _3969_/A2 _3596_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_5322_ _5322_/A1 _5479_/A3 _5444_/A2 _5324_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_115_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5253_ _5253_/A1 _5253_/A2 _5502_/B1 _5502_/B2 _5253_/C _5490_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_102_439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5184_ _5184_/A1 _5440_/A4 _5184_/A3 _5184_/A4 _5188_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_69_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4204_ hold388/Z hold645/Z _4204_/S _4204_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4135_ input58/Z hold390/Z _6863_/Q _4135_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_96_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4066_ _4075_/A2 _4065_/Z _4067_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4968_ _5262_/A4 _5315_/A4 _4690_/C _4963_/B _5351_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_51_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4899_ _5307_/B _4056_/B _4777_/B _5036_/A2 _5435_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_3919_ _6910_/Q _5655_/A4 hold37/I _5546_/A2 _3974_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6707_ _6707_/D _6662_/Z _7346_/CLK _6707_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
X_6638_ _6638_/I0 _7320_/Q _6642_/S _7320_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_177_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6569_ _6569_/A1 _6569_/A2 _6569_/A3 _6577_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_3_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_789 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_58__1374_ clkbuf_4_13_0__1374_/Z net583_245/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_120_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet483_112 net833_480/I _7157_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet483_123 net433_88/I _7146_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet483_145 net833_497/I _7124_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet483_134 net433_65/I _7135_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet433_59 net433_59/I _7210_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_101_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_356 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_916 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_927 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_938 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_949 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5940_ _6787_/Q _6789_/Q _7272_/Q _5940_/B _5941_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_18_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5871_ hold286/Z hold164/Z _5874_/S _7230_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4822_ _5416_/A1 _5267_/B _5152_/C _4822_/A4 _4823_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_33_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4753_ _4693_/Z _4706_/Z _4709_/Z _5489_/A1 _5428_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_147_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3704_ _4108_/B2 _4262_/S _4281_/S input39/Z _3705_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6423_ _7091_/Q _6578_/A2 _6312_/Z _7221_/Q _6424_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4684_ _4487_/Z _4423_/Z _4684_/B _4720_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_3635_ _3635_/A1 _3635_/A2 _3627_/Z _3635_/A4 _3636_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_143_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3566_ _3802_/A2 _3511_/C _3473_/B _3833_/A2 _3950_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_6354_ _7105_/Q _6285_/Z _6564_/C1 _7081_/Q _6354_/C _6357_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_6285_ _6561_/A3 _6310_/A4 _7276_/Q _6563_/A4 _6285_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_115_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5305_ _4759_/C _5313_/A1 _4421_/Z _5308_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3497_ _5534_/A1 _3827_/A1 _3477_/Z _3496_/B _3969_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_5236_ _5084_/C _5267_/C _5243_/A3 _5236_/B _5424_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_130_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5167_ _5223_/A1 _5295_/A1 _5290_/C _5466_/B _5390_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_130_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5098_ _5315_/A4 _5098_/A2 _4995_/Z _4942_/Z _5426_/B1 _5370_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_84_643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4118_ _4118_/A1 _7343_/Q _4118_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4049_ _6324_/A1 _6312_/A4 _7281_/Q _7278_/Q _6307_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_84_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_842 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold8 hold8/I hold8/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_94_429 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_857 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_868 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold408 _7092_/Q hold408/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_144_648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold419 _5586_/Z _6979_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_7_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3420_ _6708_/Q _6707_/Q _6774_/Q _6709_/Q _3422_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3351_ _7157_/Q _3351_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_97_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_713 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xload_slew355 hold41/Z _5820_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xnet683_307 net783_417/I _6962_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_151_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6070_ _6070_/A1 _6070_/A2 _6070_/A3 _6070_/A4 _6071_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
Xnet683_329 net733_397/I _6940_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_746 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet683_318 net783_437/I _6951_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_leaf_41__1374_ clkbuf_4_15_0__1374_/Z net583_214/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5021_ _3379_/I _3380_/I _5153_/A2 _5451_/A1 _5024_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_24_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xload_slew366 _5745_/A4 _5802_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_66_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6972_ _6972_/D _7304_/RN _6972_/CLK _6972_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_80_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5923_ _5985_/A3 _5923_/A2 _5925_/A2 _5920_/B _7268_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5854_ hold58/Z hold83/Z _5855_/S hold84/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4805_ _5468_/C _5253_/A1 _5468_/B _5235_/A1 _4811_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_21_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5785_ hold391/Z hold778/Z _5792_/S _7154_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4736_ _5327_/B _4822_/A4 _5250_/C _5330_/A2 _4737_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_174_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4667_ _4750_/A3 _4750_/A4 _4667_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_119_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6406_ _7035_/Q _6563_/A3 _6562_/A4 _6406_/A4 _6410_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3618_ _6974_/Q _3559_/Z _3958_/B1 _6724_/Q _3969_/B1 hold72/I _3619_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_4598_ _4443_/Z _5459_/A3 _4598_/A3 _4598_/A4 _5223_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_6337_ _7056_/Q _6570_/B1 _6579_/A2 _6742_/Q _6339_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_135_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3549_ _3827_/A1 _3833_/A2 _3477_/Z _3496_/B _3968_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_131_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6268_ _7275_/Q _6268_/A2 _6268_/B _6271_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5219_ _5219_/A1 _5219_/A2 _5219_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_103_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6199_ hold52/I _6259_/A2 _6259_/B1 _6983_/Q _6258_/C1 _7071_/Q _6202_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_57_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet633_259 net783_419/I _7010_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_75_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_679 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_865 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5570_ hold5/Z hold136/Z hold38/Z _6965_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_172_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4521_ _4718_/B _4661_/C _5153_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_7240_ _7240_/D _7265_/RN _7240_/CLK hold74/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4452_ _4452_/A1 _4452_/A2 _4417_/Z _4957_/A4 _5082_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
Xhold216 _5707_/Z _7086_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold205 _5706_/Z _7085_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold238 _6980_/Q hold238/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold249 _7003_/Q hold249/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3403_ _4073_/B1 _4119_/B _3421_/B _3991_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
Xhold227 _5907_/Z _7262_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_171_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4383_ _4137_/Z _6886_/Q _4383_/S _4383_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7171_ _7171_/D _7304_/RN _7171_/CLK _7171_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_113_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3334_ _7280_/Q _6312_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_4
X_6122_ _7076_/Q _6260_/A2 _6257_/B1 _7060_/Q _6124_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_86_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_532 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6053_ _7139_/Q _6259_/A2 _6261_/A2 _7123_/Q _6055_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5004_ _5004_/A1 input95/Z _4423_/Z _5370_/A1 _5005_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6955_ _6955_/D input75/Z _6955_/CLK _7368_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_1709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5906_ hold139/Z hold558/Z _5910_/S _5906_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6886_ _6886_/D _7341_/RN _6886_/CLK _6886_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_34_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5837_ hold2/Z _7201_/Q hold18/Z hold19/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5768_ hold388/Z hold685/Z _5774_/S _5768_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_175_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4719_ _4686_/B _4759_/B1 _4719_/B _4825_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_5699_ hold2/Z hold54/Z _5699_/S hold55/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_147_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold750 _7065_/Q hold750/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7369_ _7369_/I _7369_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold761 _5593_/Z _6985_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_1_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold772 _7120_/Q hold772/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold794 _7080_/Q hold794/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold783 _6923_/Q hold783/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_162_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4109__7 _4109__7/I _7262_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_91_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6740_ _6740_/D _7262_/RN _6740_/CLK _6740_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3952_ _3952_/A1 _3952_/A2 _3952_/A3 _3953_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_16_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3883_ _3883_/A1 _3883_/A2 _3883_/A3 _3883_/A4 _3884_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_91_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6671_ _7262_/RN _6994_/Q _4026_/C _6671_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_5622_ hold139/Z hold364/Z _5626_/S _5622_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5553_ hold391/Z hold649/Z _5554_/S _6950_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_129_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4504_ _5301_/A2 _5235_/A1 _3379_/I _5394_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_145_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5484_ _4718_/B _5484_/A2 _5439_/C _5484_/A4 _5485_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4435_ _4759_/C _5136_/A2 _5098_/A2 _4775_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_7223_ _7223_/D _7265_/RN _7223_/CLK _7223_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_132_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4366_ _4378_/A1 _5893_/A3 _6653_/A2 _5535_/B _4368_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_7154_ _7154_/D _7302_/RN _7154_/CLK _7154_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_3317_ _6863_/Q _3491_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_4
XFILLER_140_470 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6105_ _7157_/Q _6258_/A2 _6260_/B1 _7115_/Q _6259_/B1 _7107_/Q _6106_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_59_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7085_ _7085_/D _7281_/RN _7085_/CLK _7085_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4297_ hold58/Z hold369/Z _4298_/S _4297_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6036_ _7131_/Q _6232_/B1 _6036_/A3 _7271_/Q _6038_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_395 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_6938_ _6938_/D _7262_/RN _6938_/CLK _7349_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XPHY_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_6869_ _6869_/D _7341_/RN _6869_/CLK _6869_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_41_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold580 _4345_/Z _6853_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold591 _4376_/Z _6881_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_2_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4220_ _6653_/A2 _5535_/B _3527_/Z _5745_/A4 _4222_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_4151_ _5856_/A1 _5784_/A3 _5532_/A3 _5838_/A4 _4159_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_110_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4082_ _4078_/S _7253_/Q _4082_/B _4082_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_95_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4984_ _5285_/A1 _4956_/C _5410_/A2 _5410_/A3 _4985_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3935_ _6889_/Q _5893_/A3 _4405_/A3 _4405_/A2 _3979_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6723_ _6723_/D _7304_/RN _6723_/CLK _6723_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_189_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6654_ hold391/Z hold566/Z _6655_/S _6654_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5605_ hold164/Z hold402/Z _5608_/S _5605_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3866_ _7147_/Q _3866_/A2 _3977_/B1 _7033_/Q _3866_/C _3868_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_118_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3797_ _3496_/B _3831_/A2 _4246_/A2 _3477_/Z _3959_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_6585_ _6585_/A1 _6583_/Z _6585_/B _6586_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_173_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5536_ hold551/Z _5536_/A2 hold552/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_160_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5467_ _5467_/A1 _5467_/A2 _5328_/Z _5467_/A4 _5491_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_4418_ _4418_/A1 _4418_/A2 _4418_/A3 _4418_/A4 _4432_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_172_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7206_ _7206_/D _7302_/RN _7206_/CLK _7206_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5398_ _5504_/A1 _5486_/A1 _5398_/A3 _5441_/A1 _5402_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_87_844 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4349_ _6594_/A1 _4358_/S _4349_/B _6855_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7137_ _7137_/D _7302_/RN _7137_/CLK _7137_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_7068_ _7068_/D _7265_/RN _7068_/CLK _7068_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6019_ _7154_/Q _6258_/A2 _6261_/A2 _7122_/Q _6232_/C _6020_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_86_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2015 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2004 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2059 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2048 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2037 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2026 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_796 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1358 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_18__1374_ clkbuf_4_10_0__1374_/Z net433_88/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_10_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_827 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_877 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2571 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_654 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1881 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1892 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3720_ _6713_/Q _5784_/A3 _5532_/A3 _5546_/A2 _3745_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_9_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3651_ _7101_/Q _3950_/A2 _3943_/C1 _7061_/Q _3943_/B1 _7199_/Q _3652_/I VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_155_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3582_ _3582_/A1 _3582_/A2 _3582_/A3 _3597_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6370_ _7025_/Q _6528_/A2 _6581_/B1 _7259_/Q _6371_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_161_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5321_ _5484_/A2 _5445_/A2 _5321_/A3 _5194_/C _5479_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_127_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5252_ _5416_/A1 _5327_/B _5252_/A3 _5252_/A4 _5253_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_5183_ _5226_/A1 _5471_/A1 _5439_/B _5439_/C _5401_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_87_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4203_ hold391/Z hold820/Z _4204_/S _4203_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4134_ _5535_/B _5546_/A2 _5532_/A3 _5784_/A3 _4150_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_113_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4065_ _4056_/B _4065_/A2 _4065_/A3 _4065_/A4 _4065_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_84_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4967_ _5463_/A1 _4967_/A2 _5454_/B1 _4437_/Z _4969_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_51_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6706_ _6706_/D _6661_/Z _4108_/B2 _6706_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4898_ _4423_/Z _5436_/A1 _5484_/A2 _5210_/C _5318_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_3918_ input36/Z hold37/I _5784_/A3 _5528_/A2 _3982_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6637_ _6637_/A1 _6637_/A2 _6638_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3849_ _3849_/A1 _3849_/A2 _3849_/A3 _3849_/A4 _3885_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_180_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6568_ _6767_/Q _6274_/Z _6568_/B1 _6739_/Q _6569_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_152_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5519_ hold391/Z hold843/Z _5524_/S _6927_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6499_ _6491_/Z _6499_/A2 _6499_/A3 _6498_/Z _6506_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_160_340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet483_102 _4109__6/I _7167_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_87_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_5__1374_ clkbuf_4_3_0__1374_/Z net833_473/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_59_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet483_135 _4109__49/I _7134_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet483_124 net533_163/I _7145_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet483_113 net533_176/I _7156_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_170_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet483_146 net833_489/I _7123_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_47_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_906 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_917 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_928 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_939 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5870_ hold331/Z hold139/Z _5874_/S _7229_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_18_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4821_ _5471_/B2 _5301_/A2 _5153_/B _5264_/A4 _5472_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XTAP_2390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4752_ _5262_/A4 _5136_/B1 _3380_/I _5034_/A2 _4755_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_159_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4683_ _4683_/A1 _5198_/B _4683_/B _5042_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3703_ _7230_/Q _3964_/A2 _4264_/A1 input56/Z _3705_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_119_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_64__1374_ clkbuf_4_13_0__1374_/Z net633_281/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_162_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3634_ hold82/I _3980_/A2 _3634_/B _3634_/C _3635_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_6422_ _7067_/Q _6299_/Z _6566_/C1 _7019_/Q _6578_/C1 _7173_/Q _6424_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_161_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6353_ _7097_/Q _6563_/A3 _6561_/A3 _6563_/A4 _6354_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_3565_ _3498_/B _4246_/A1 _3519_/Z _3460_/B _3958_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_3496_ _3491_/B hold298/Z _3496_/B _3496_/C hold299/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_115_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5304_ _5347_/A1 _5435_/A1 _5466_/A2 _5327_/B _5313_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_6284_ _7280_/Q _6563_/A3 _6563_/A4 _5975_/B _6284_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_88_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5235_ _5235_/A1 _5235_/A2 _4487_/Z _4718_/B _5243_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_142_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5166_ _4056_/B _5166_/A2 _4669_/B _5166_/A4 _5172_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_96_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5097_ _5489_/A1 _5282_/B _5370_/A1 _4437_/Z _5414_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_57_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4117_ _4117_/A1 input73/Z _4117_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_17_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4048_ _6323_/A1 _7279_/Q _6562_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_72_828 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_249 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5999_ _6103_/A1 _6211_/B _7274_/Q _7272_/Q _6257_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_12_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_863 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_161_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_896 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput290 _6729_/Q pll_trim[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xhold9 hold9/I hold9/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_47_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold409 _6971_/Q hold409/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_109_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3350_ _7165_/Q _3350_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_124_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_714 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5020_ _5020_/A1 _5020_/A2 _5020_/A3 _5024_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
Xload_slew345 hold173/Z _5573_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xnet683_308 net783_419/I _6961_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_97_257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet683_319 net783_437/I _6950_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6971_ _6971_/D _7304_/RN _6971_/CLK _6971_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_0_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5922_ _5918_/B _5985_/A3 _6790_/Q _6788_/Q _5925_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_53_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5853_ hold5/Z hold156/Z _5855_/S _5853_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4804_ _5152_/C _5327_/B _4822_/A4 _5271_/A4 _5239_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_5784_ _5856_/A1 _5784_/A2 _5784_/A3 _5838_/A4 _5792_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_22_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4735_ _5245_/A1 _5330_/A2 _4735_/B _5467_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4666_ _4922_/B _4775_/A1 _4787_/A3 _5166_/A4 _4750_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_107_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4597_ _4443_/Z _5459_/A3 _4598_/A3 _4598_/A4 _4597_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_135_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6405_ _7149_/Q _6562_/A2 _6562_/A3 _6561_/A3 _6417_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3617_ hold62/I _3969_/A2 _3959_/A2 _6732_/Q _3968_/A2 hold60/I _3619_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6336_ _7226_/Q _6311_/B _6292_/Z _7072_/Q _6341_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3548_ _3454_/Z _3519_/Z _3534_/C _4246_/A1 _3959_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_143_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3479_ _4073_/B1 hold170/Z hold171/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_130_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6267_ _7275_/Q _6264_/Z _6267_/B1 _6107_/B _6267_/C _6268_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5218_ _5502_/B2 _5218_/A2 _5218_/B1 _5351_/B1 _5219_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_97_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6198_ _6198_/A1 _6198_/A2 _6198_/A3 _6198_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_5149_ _5149_/A1 _5149_/A2 _5338_/A1 _5338_/A2 _5150_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_69_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_877 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4520_ _4684_/B _5484_/A2 _5445_/A2 _5393_/A3 _4558_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_172_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4451_ _4774_/A1 _4451_/A2 _4451_/B _5082_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_117_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold217 _6974_/Q hold217/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_8_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold206 _6827_/Q hold206/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold228 _7087_/Q hold228/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold239 _5587_/Z _6980_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7170_ _7170_/D _7302_/RN _7170_/CLK _7170_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_3402_ _6777_/Q _6776_/Q _6774_/Q _3412_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_6121_ _6996_/Q _6258_/B1 _6256_/B1 _7084_/Q _6124_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4382_ hold391/Z _6885_/Q _4383_/S _4382_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_500 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3333_ _7278_/Q _6323_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_4
XFILLER_112_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_533 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6052_ _6211_/B _6266_/B _7155_/Q _7274_/Q _6055_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5003_ _5003_/A1 _5003_/A2 _5005_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_577 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6954_ hold26/Z input75/Z _6954_/CLK _7367_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_81_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_500 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5905_ hold25/Z hold477/Z _5910_/S _5905_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_179_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6885_ _6885_/D _7341_/RN _6885_/CLK _6885_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_179_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5836_ hold58/Z hold100/Z hold18/Z _7200_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_14_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5767_ hold391/Z hold792/Z _5774_/S _5767_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5698_ hold58/Z hold89/Z _5699_/S hold90/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_108_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4718_ _5330_/A1 _5245_/A1 _4718_/B _4718_/C _4737_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4649_ _4443_/Z _5051_/C _5416_/A1 _5084_/B _4650_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_107_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold751 _7017_/Q hold751/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_146_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7368_ _7368_/I _7368_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold762 _6945_/Q hold762/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_89_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold773 _5746_/Z _7120_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold740 _7130_/Q hold740/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6319_ _7280_/Q _6562_/A2 _6563_/A3 _5975_/B _6319_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
Xhold795 _5701_/Z _7080_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_89_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold784 _6768_/Q hold784/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7299_ _7299_/D _7304_/RN _7304_/CLK _7299_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_103_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_828 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_186_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_825 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4109__8 _4109__8/I _7261_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3951_ _7072_/Q _3951_/A2 _3951_/B1 _7088_/Q _3951_/C _3954_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_91_797 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3882_ _7235_/Q _3943_/A2 _4243_/S input44/Z _3882_/C _3883_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_6670_ input75/Z _6994_/Q _4026_/C _6670_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_32_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5621_ hold25/Z hold498/Z _5626_/S _5621_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5552_ _5838_/A4 _5552_/A2 _6653_/A3 _5884_/A2 _5554_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_4503_ _5048_/C _5307_/B _5078_/A2 _5350_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_5483_ _5483_/A1 _5503_/A2 _5483_/B _5483_/C _5487_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_172_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4434_ _4694_/B _4922_/B _4684_/B _5307_/B _4439_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_7222_ _7222_/D _7262_/RN _7222_/CLK _7222_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4365_ _6870_/Q _3491_/B _4365_/B _4365_/C _6863_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_160_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7153_ hold15/Z _7265_/RN _7153_/CLK _7153_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_116_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7084_ _7084_/D _7281_/RN _7084_/CLK _7084_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6104_ _7173_/Q _6256_/A2 _6257_/B1 _7181_/Q _6106_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3316_ _3316_/I _4072_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_112_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6035_ _6743_/Q _6266_/C _6232_/B1 _7147_/Q _6232_/C _6038_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_4296_ hold5/Z hold424/Z _4298_/S _4296_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_6937_ _6937_/D input75/Z _6937_/CLK _6937_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6868_ _6868_/D _7341_/RN _6868_/CLK _6868_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_167_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5819_ hold2/Z hold50/Z _5819_/S hold51/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6799_ _6799_/D _7281_/RN _6799_/CLK _6799_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_22_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold581 _6893_/Q hold581/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold570 _6854_/Q hold570/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_1_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold592 _7364_/I hold592/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_77_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4150_ hold2/Z hold158/Z _4150_/S _4150_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4081_ _4078_/S input90/Z _4082_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4983_ _5355_/A2 _4956_/C _5410_/A2 _5410_/A3 _4985_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_51_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3934_ _6891_/Q hold41/I _4405_/A3 _5546_/A2 _3979_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6722_ _6722_/D _7304_/RN _6722_/CLK _6722_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6653_ _5535_/B _6653_/A2 _6653_/A3 hold299/Z _6655_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_3865_ _7219_/Q _3975_/A2 _3865_/B _3868_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5604_ hold139/Z hold149/Z _5608_/S _5604_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_149_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3796_ _6741_/Q _5856_/A2 _5546_/A2 _3527_/Z _3845_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_20_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6584_ _6584_/A1 _6830_/Q _6584_/B _6585_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5535_ hold550/Z _5535_/A2 _5535_/B hold551/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5466_ _5466_/A1 _5466_/A2 _5466_/B _5466_/C _5467_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_105_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4417_ _4418_/A1 _4418_/A2 _4418_/A3 _4418_/A4 _4417_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_7205_ _7205_/D _7262_/RN _7205_/CLK _7205_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_120_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5397_ _5397_/A1 _5503_/A2 _5397_/B _5397_/C _5441_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_141_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7136_ _7136_/D _7341_/RN _7136_/CLK _7136_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_59_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4348_ _4358_/S _6855_/Q _4349_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7067_ _7067_/D _7265_/RN _7067_/CLK _7067_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4279_ _6966_/Q hold58/Z _4281_/S _4279_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_59_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6018_ _7170_/Q _6256_/A2 _6258_/B1 _6742_/Q _6020_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_74_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2016 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2005 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2049 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2038 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_823 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1871 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_789 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_186_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3650_ _7167_/Q _3878_/A2 _3964_/A2 _7231_/Q _3654_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_9_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3581_ _7241_/Q _3943_/A2 _3953_/B1 _7193_/Q _3581_/C _3582_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_142_500 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5320_ _5484_/A2 _5445_/A2 _5321_/A3 _5194_/C _5446_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_114_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5251_ _5333_/A1 _5251_/A2 _5333_/A3 _5254_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_170_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4202_ _5838_/A4 _5518_/A1 _3527_/Z _5838_/A2 _4204_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_142_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5182_ _5502_/A1 _5439_/B _5502_/B1 _5180_/B _5440_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_87_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4133_ hold44/Z _7323_/Q _6863_/Q hold45/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_110_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4064_ _4451_/B _4774_/B _4064_/B _4064_/C _4065_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
Xclkbuf_leaf_24__1374_ clkbuf_4_11_0__1374_/Z _4109__48/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_110_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_104__1374_ clkbuf_4_1_0__1374_/Z net833_483/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_87__1374_ net583_226/I _4109__9/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_71_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6705_ _6705_/D _6660_/Z _4108_/B2 _6705_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4966_ _5105_/A1 _4966_/A2 _4969_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_149_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4897_ _4897_/A1 _5192_/A1 _4897_/A3 _4903_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3917_ _6933_/Q _5802_/A2 _5727_/A3 _5552_/A2 _3949_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_6636_ _6878_/Q _6636_/A2 _6636_/B1 _6640_/B2 _6637_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_177_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3848_ _7123_/Q _3956_/A2 _3681_/Z _6923_/Q _3849_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_22_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6567_ _6741_/Q _6311_/B _6567_/B1 _6761_/Q _6569_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_20_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3779_ _7140_/Q _3958_/A2 _3681_/Z _6924_/Q _3964_/C1 _7260_/Q _3780_/A4 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_164_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5518_ _5518_/A1 _5838_/A4 _5552_/A2 _5745_/A4 _5524_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_6498_ _6498_/A1 _6498_/A2 _6498_/A3 _6498_/A4 _6498_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_106_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5449_ _6907_/Q _4365_/C _5449_/B _5450_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_105_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_154_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet483_103 _4109__48/I _7166_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_87_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7119_ _7119_/D _7302_/RN _7119_/CLK _7119_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xnet483_136 _4109__24/I _7133_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet483_125 net433_93/I _7144_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet483_114 net783_441/I _7155_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_101_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet483_147 net833_456/I _7122_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_103_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_786 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_1_1__f_wbbd_sck clkbuf_0_wbbd_sck/Z _3340__1/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_151_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1145 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_184_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_828 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_183_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_170_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_907 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_918 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_929 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_678 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4820_ _5404_/B2 _4823_/A2 _5266_/A2 _5468_/A1 _5472_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_2391 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4751_ _4667_/Z _5244_/A2 _4693_/Z _4709_/Z _5136_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_187_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4682_ _5459_/A3 _4682_/A2 _5285_/A1 _5051_/B _5198_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_3702_ _7068_/Q _3980_/A2 _3943_/C1 _7060_/Q _7012_/Q _3962_/A2 _3705_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_3633_ _3633_/A1 _3633_/A2 _3634_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6421_ _7253_/Q _6580_/B1 _6309_/Z _7237_/Q _6745_/Q _6579_/A2 _6424_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_146_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_894 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3564_ _3454_/Z _3498_/B _3644_/A2 _4246_/A1 _4281_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_6352_ _7033_/Q _6563_/A3 _6562_/A4 _6406_/A4 _6357_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3495_ hold28/Z hold36/Z _3500_/C _3496_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_5303_ _5303_/A1 _5388_/A2 _5303_/A3 _5303_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_6283_ _6324_/A1 _6323_/A1 _6325_/A1 _6325_/A2 _6573_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_170_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5234_ _5234_/A1 _5457_/A2 _5238_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5165_ _5165_/A1 _5295_/C _5165_/A3 _5166_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_111_750 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_675 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4116_ input85/Z input58/Z _7344_/Q _4116_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5096_ _4437_/Z _5282_/B _5378_/A1 _5489_/A1 _5379_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4047_ _5975_/B _7280_/Q _6563_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_84_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5998_ _6036_/A3 _6103_/A1 _6211_/C _6211_/B _6262_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_24_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4949_ _4773_/B _5011_/A2 _4952_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_166_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6619_ _6880_/Q _6619_/A2 _6619_/B1 _6879_/Q _6621_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_177_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput280 _6712_/Q pll_trim[18] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput291 _6730_/Q pll_trim[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_833 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_877 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_70__1374_ _4109__12/I net583_233/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_15_222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_797 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_715 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet683_309 net683_320/I _6960_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_726 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_748 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xload_slew346 _5518_/A1 _5528_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_140_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xload_slew357 _5856_/A2 _6653_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_81_604 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6970_ _6970_/D _7304_/RN _6970_/CLK _6970_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_53_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5921_ _7267_/Q _7268_/Q _5981_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5852_ hold164/Z hold289/Z _5855_/S _5852_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_726 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5783_ hold2/Z _7153_/Q hold14/Z hold15/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4803_ _4803_/A1 _4803_/A2 _4803_/A3 _4811_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_159_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4734_ _5315_/A4 _4718_/B _4661_/C _3379_/I _5330_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_162_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4665_ _4774_/A1 _4710_/C _4774_/B _4665_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_107_319 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold900 _7315_/Q hold900/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4596_ _5082_/C _5435_/A1 _4454_/B _5503_/A1 _5067_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_147_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6404_ _7245_/Q _6563_/A2 _6562_/A3 _6563_/A4 _6413_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3616_ _3616_/A1 _3616_/A2 _3616_/A3 _3616_/A4 _3636_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3547_ _3604_/A2 _3507_/C _3833_/A2 _3802_/A2 _3951_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_115_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6335_ _7210_/Q _6570_/A2 _6286_/Z _7154_/Q _6341_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_142_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3478_ _3491_/B _3475_/Z _3496_/C _3827_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_6266_ _6902_/Q _6232_/C _6266_/B _6266_/C _6267_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5217_ _4437_/Z _5420_/A1 _5302_/B _5226_/A1 _5217_/C _5356_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_6197_ hold85/I _6258_/A2 _6257_/A2 _7015_/Q _6261_/B1 _7047_/Q _6198_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_69_472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5148_ _5476_/A1 _5260_/B _5148_/B1 _5399_/B _5338_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_56_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5079_ _5079_/A1 _5321_/A3 _5209_/B1 _5459_/A2 _5230_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_151_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_403 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_878 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_399 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_604 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4450_ _4959_/A2 _4450_/A2 _4452_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold207 _4306_/Z _6827_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xclkbuf_3_4_0__1374_ clkbuf_0__1374_/Z clkbuf_4_9_0__1374_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xhold229 _5708_/Z _7087_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_109_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4381_ hold45/Z hold190/Z hold29/Z _5655_/A4 _4383_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_3401_ _3401_/A1 _4054_/A1 _7346_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold218 _6942_/Q hold218/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3332_ _7279_/Q _6324_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_12
X_6120_ _7020_/Q _6259_/A2 _6257_/A2 _7012_/Q _6124_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_98_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_512 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6051_ _7113_/Q _6260_/B1 _6259_/B1 _7105_/Q _6256_/A2 _7171_/Q _6055_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XTAP_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5002_ _5002_/A1 _5002_/A2 _5002_/A3 _5002_/A4 _5003_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6953_ _6953_/D input75/Z _6953_/CLK _7366_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_93_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5904_ hold388/Z hold520/Z _5910_/S _5904_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6884_ _6884_/D _7341_/RN _6884_/CLK _6884_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5835_ hold5/Z hold151/Z hold18/Z _7199_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5766_ _5856_/A1 _5784_/A2 _5838_/A2 _5838_/A4 _5774_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_163_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5697_ hold5/Z hold154/Z _5699_/S _5697_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4717_ _5244_/A2 _5244_/A3 _4750_/A3 _4750_/A4 _5245_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_162_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4648_ _4443_/Z _5051_/C _5084_/B _5223_/A1 _5418_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_135_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold730 _5840_/Z _7203_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4579_ _5046_/A1 _5046_/A2 _5307_/B _5208_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xhold741 _7243_/Q hold741/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold752 _5629_/Z _7017_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_122_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7367_ _7367_/I _7367_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold763 _5544_/Z hold763/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold796 _7147_/Q hold796/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_115_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6318_ _6318_/A1 _6318_/A2 _6318_/A3 _6584_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_103_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold785 _6933_/Q hold785/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7298_ _7298_/D _7304_/RN _7302_/CLK _7298_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold774 _6762_/Q hold774/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6249_ _6755_/Q _6262_/A2 _6258_/C1 _6767_/Q _6251_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_162_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_873 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_865 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet733_390 net783_420/I _6828_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_5_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold90 hold90/I hold90/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4109__9 _4109__9/I _7260_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_91_765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3950_ _7096_/Q _3950_/A2 _3950_/B1 _7040_/Q _3950_/C _3954_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_17_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3881_ _3881_/A1 _3881_/A2 _3882_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_176_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5620_ hold388/Z hold790/Z _5626_/S _5620_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5551_ hold391/Z hold614/Z _5551_/S _6949_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_77_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4502_ _4479_/B _4479_/C _4502_/B _5048_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_145_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7221_ _7221_/D _7341_/RN _7221_/CLK _7221_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5482_ _5482_/A1 _5482_/A2 _5482_/A3 _5480_/Z _5505_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4433_ _4412_/Z _4414_/Z _4417_/Z _4669_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_104_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7152_ _7152_/D _7265_/RN _7152_/CLK hold77/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4364_ _4363_/Z _6877_/Q _6872_/Q _4365_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_99_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7083_ _7083_/D _7281_/RN _7083_/CLK _7083_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_112_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6103_ _6103_/A1 _6232_/B1 _7141_/Q _7272_/Q _6106_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_59_718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3315_ _7344_/Q _4117_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4295_ hold164/Z hold479/Z _4298_/S _4295_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6034_ _7025_/Q _6262_/B1 _7275_/Q _6041_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_132_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_6936_ _6936_/D _6936_/CLK _6936_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_179_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6867_ _6867_/D _7341_/RN _6867_/CLK _6867_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_23_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5818_ hold58/Z hold78/Z _5819_/S hold79/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6798_ _6798_/D _7302_/RN _6798_/CLK _7354_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_10_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5749_ hold391/Z hold841/Z _5756_/S _7122_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_41_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold560 _7359_/I hold560/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_150_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold571 _4346_/Z _6854_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_2_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold593 _4244_/Z _6786_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold582 _4394_/Z _6893_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_1_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2710 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2754 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_185_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4080_ _4078_/S _7261_/Q _4080_/B _4080_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_96_868 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4982_ _4982_/A1 _4982_/A2 _4982_/A3 _4985_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_63_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6721_ _6721_/D _7304_/RN _6721_/CLK _6721_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_3933_ _6968_/Q _5700_/A1 _5856_/A2 _5573_/A3 _3963_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_189_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6652_ _6652_/I0 _6652_/I1 _6652_/S _7323_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3864_ _7097_/Q _3950_/A2 _3948_/A2 _6921_/Q _3868_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_32_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5603_ hold25/Z hold284/Z _5608_/S _5603_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_47__1374_ clkbuf_4_15_0__1374_/Z net783_414/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6583_ _6584_/A1 _6583_/A2 _6583_/A3 _6582_/Z _6583_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_3795_ _6951_/Q _5884_/A2 _6653_/A3 _5552_/A2 _3873_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_173_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5534_ _5534_/A1 _5534_/A2 _3519_/Z hold391/Z _5536_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_5465_ _5462_/Z _5464_/Z _5497_/B _5477_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4416_ _4432_/A1 _4432_/A2 _4957_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_160_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7204_ _7204_/D _7302_/RN _7204_/CLK _7204_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_132_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5396_ _5396_/A1 _5396_/A2 _5398_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7135_ _7135_/D _7302_/RN _7135_/CLK _7135_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4347_ _6873_/Q _7323_/RN _4358_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_100_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7066_ _7066_/D _7265_/RN _7066_/CLK _7066_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4278_ _4277_/Z hold546/Z _4282_/S _4278_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_143_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6017_ _7138_/Q _6259_/A2 _6262_/B1 _7146_/Q _6020_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_86_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2006 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2017 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_1_0__f_wbbd_sck clkbuf_0_wbbd_sck/Z _4108_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_4_7_0__1374_ clkbuf_4_7_0__1374_/I _4109__12/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_6919_ _6919_/D _6677_/Z _4111_/I1 _6919_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_167_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_163_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold390 _7314_/Q hold390/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_151_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2573 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1861 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1894 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1872 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3580_ _3580_/A1 _3580_/A2 _3580_/A3 _3581_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_142_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5250_ _5416_/A1 _5271_/A4 _5250_/B _5250_/C _5333_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_181_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4201_ hold388/Z hold568/Z _4201_/S _4201_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5181_ _5218_/A2 _5180_/B _5181_/B _5181_/C _5184_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_69_835 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4132_ _7341_/RN _6994_/Q _4026_/C _4132_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_96_643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4063_ _4063_/A1 _4063_/A2 _4063_/A3 _4075_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_110_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_573 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4965_ _5426_/B1 _4965_/A2 _3380_/I _5375_/A1 _4965_/C _4966_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_51_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6704_ _6704_/D _6659_/Z _4108_/B2 _6704_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_149_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3916_ _7162_/Q _5655_/A4 _5884_/A2 _3527_/Z _3945_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_149_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4896_ _4056_/B _4777_/C _5226_/A1 _5445_/A3 _4897_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_32_470 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6635_ _6880_/Q _6635_/A2 _6635_/B1 _6879_/Q _6637_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_177_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3847_ _6969_/Q _3559_/Z _5544_/S _6944_/Q _3847_/C _3849_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_20_654 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6566_ _7341_/Q _6279_/Z _6299_/Z _6890_/Q _6566_/C1 _6867_/Q _6569_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_3778_ _7124_/Q _3956_/A2 _3959_/A2 _6728_/Q _3958_/B1 _6720_/Q _3780_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_5517_ hold164/Z hold482/Z _5517_/S _6926_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_145_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6497_ _7192_/Q _6274_/Z _6567_/B1 hold70/I _6311_/B _7232_/Q _6498_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_161_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5448_ _5448_/A1 _5479_/A4 _5448_/B _5448_/C _5449_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_105_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5379_ _5379_/A1 _5379_/A2 _5379_/A3 _5379_/A4 _5453_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_7118_ hold63/Z _7302_/RN _7118_/CLK hold62/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_7049_ _7049_/D _7341_/RN _7049_/CLK _7049_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
Xnet483_104 net433_82/I _7165_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet483_126 net833_491/I _7143_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet483_115 net683_331/I _7154_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet483_137 net433_77/I _7132_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_101_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet483_148 net833_471/I _7121_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_27_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_30__1374_ clkbuf_4_11_0__1374_/Z net433_90/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_110__1374_ net733_398/I net783_411/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_136_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_93__1374_ clkbuf_4_3_0__1374_/Z _4109__7/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_908 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_919 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4750_ _5244_/A2 _4693_/Z _4750_/A3 _4750_/A4 _5250_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XTAP_1691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4681_ _4681_/A1 _4681_/A2 _4683_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3701_ _7084_/Q _3962_/B1 _3786_/B1 hold21/I _3705_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_174_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3632_ hold77/I _3866_/A2 _3939_/A2 _6990_/Q _3633_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6420_ _7051_/Q _6575_/B1 _6311_/C _7003_/Q _6581_/B1 _7261_/Q _6425_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6351_ _7243_/Q _6563_/A2 _6562_/A3 _6563_/A4 _6360_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3563_ _3827_/A2 _3496_/B _3833_/A2 _3831_/A2 _3875_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_5302_ _5436_/A4 _5471_/A1 _5468_/A1 _5302_/B _5388_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_143_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3494_ _5534_/A1 _3644_/A2 _3511_/C _3473_/B _3943_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_6282_ _6312_/A4 _6296_/A2 _7281_/Q _7279_/Q _6575_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_5233_ _5459_/A3 _5459_/A2 _5355_/A2 _5051_/B _5457_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_69_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5164_ _5169_/B1 _5484_/A2 _4661_/C _4718_/B _5165_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_110_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4115_ _4115_/I _4115_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5095_ _4963_/B _5111_/A2 _5288_/A4 _4947_/C _5285_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_110_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4046_ _6306_/A3 _7277_/Q _6325_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XPHY_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_64_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5997_ _7016_/Q _6259_/A2 _6260_/A2 _7072_/Q _6003_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_178_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4948_ _4947_/C _4963_/B _4955_/B _5454_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_149_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4879_ _4423_/Z _5177_/A3 _5153_/B _5439_/B _4881_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6618_ _6618_/I0 _7315_/Q _6642_/S _7315_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6549_ _6897_/Q _6578_/A2 _6310_/Z _6831_/Q _6578_/C1 _6772_/Q _6554_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_180_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput270 _6929_/Q pll_sel[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_160_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput292 _6731_/Q pll_trim[5] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput281 _6713_/Q pll_trim[19] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_75_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_183_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_868 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xload_slew347 _4405_/A2 _5518_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_749 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_816 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xload_slew369 _5535_/B _5838_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_16
XFILLER_65_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5920_ _6790_/Q _5930_/A2 _5920_/B _7267_/Q _5923_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_80_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5851_ hold139/Z hold441/Z _5855_/S _5851_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5782_ hold58/Z hold77/Z hold14/Z _7152_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4802_ _5152_/C _5327_/B _4822_/A4 _5369_/A2 _4803_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_21_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4733_ _5262_/A4 _5301_/A2 _5235_/A1 _3380_/I _5476_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_159_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4664_ _4774_/A1 _4710_/C _4774_/B _4750_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_6403_ _7189_/Q _6274_/Z _6568_/B1 _7115_/Q _6410_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4595_ _4595_/A1 _4595_/A2 _5222_/A3 _4600_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xhold901 _6704_/Q hold901/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_134_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3615_ hold70/I _3958_/A2 _3956_/B1 hold96/I _3616_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3546_ _3511_/C _3802_/A2 _5534_/A1 _3604_/A2 _3980_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_6334_ _6334_/A1 _6334_/A2 _6333_/Z _6334_/A4 _6334_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_135_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_898 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6265_ _6211_/C _7273_/Q _6753_/Q _7275_/Q _6267_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5216_ _5216_/A1 _5420_/B _5220_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_142_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3477_ hold298/Z _6907_/Q _6863_/Q _3477_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
X_6196_ _7095_/Q _6262_/A2 _6256_/A2 _7055_/Q _6198_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_111_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5147_ _5376_/A1 _5260_/B _5502_/B1 _5439_/B _5338_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_28_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5078_ _4481_/C _5078_/A2 _5360_/C _5285_/A1 _5081_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_151_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_72_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4029_ _6879_/Q _4074_/A2 _6873_/Q _4030_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_44_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet783_450 net833_473/I _6759_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_157_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold208 _7222_/Q hold208/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4380_ hold388/Z hold609/Z _4380_/S _4380_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold219 _5541_/Z _6942_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3400_ _3446_/B _6774_/Q _3387_/Z _4054_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_171_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3331_ _7276_/Q _6306_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_4
XFILLER_112_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_568 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6050_ _7275_/Q _6049_/Z _6056_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_535 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5001_ _5001_/A1 _5370_/A1 _5279_/B _4437_/Z _5002_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_112_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_568 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6952_ _6952_/D input75/Z _6952_/CLK _7365_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_81_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5903_ hold391/Z hold605/Z _5910_/S _5903_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6883_ _6883_/D _7341_/RN _6883_/CLK _6883_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5834_ hold164/Z hold308/Z hold18/Z _7198_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5765_ hold2/Z hold341/Z _5765_/S _5765_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5696_ hold164/Z hold324/Z _5699_/S _5696_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4716_ _5312_/B _4794_/A2 _5327_/B _5250_/C _5128_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_4647_ _5082_/B1 _5347_/A1 _4647_/B1 _5084_/C _4647_/C _4650_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_147_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7366_ _7366_/I _7366_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold720 _6773_/Q hold720/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4578_ _3380_/I _5011_/A2 _4578_/B _5312_/B _5360_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
Xhold742 _6992_/Q hold742/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6317_ _6317_/A1 _6571_/B1 _6317_/A3 _6570_/B1 _6318_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_116_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold753 _7123_/Q hold753/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold764 _6831_/Q hold764/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold731 _7219_/Q hold731/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_143_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3529_ _3473_/B _3811_/A1 _3511_/C _5534_/A1 _3939_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xhold797 _7000_/Q hold797/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_89_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_535 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold786 _6935_/Q hold786/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_1_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold775 _4209_/Z _6762_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7297_ _7297_/D _7302_/RN _7304_/CLK _7297_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_130_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6248_ _6761_/Q _6259_/A2 _6258_/B1 _7121_/Q _6251_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_162_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6179_ hold75/I _6261_/A2 _6259_/B1 hold60/I _6182_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_72_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet733_380 net833_473/I _6854_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet733_391 net733_397/I _6827_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_106_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold80 hold80/I hold80/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_76_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold91 hold91/I hold91/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_36_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_833 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3880_ _6911_/Q _5655_/A4 hold37/I _5546_/A2 _3881_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_188_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5550_ hold388/Z hold538/Z _5551_/S _6948_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_129_253 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4501_ _3380_/I _5011_/A2 _4578_/B _5307_/B _4598_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_145_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5481_ _5481_/A1 _5481_/A2 _5448_/C _5482_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_4432_ _4432_/A1 _4432_/A2 _4432_/A3 _4775_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_184_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7220_ _7220_/D _7302_/RN _7220_/CLK _7220_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_7151_ _7151_/D _7265_/RN _7151_/CLK _7151_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4363_ _6877_/D _6874_/Q _6873_/Q _6875_/Q _4363_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_99_844 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4294_ hold139/Z hold147/Z _4298_/S _4294_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7082_ _7082_/D _7281_/RN _7082_/CLK _7082_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_86_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6102_ _6235_/A1 _6102_/A2 _6102_/B1 _6235_/B2 _6102_/C _6112_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_59_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3314_ _3314_/I _3404_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_101_827 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6033_ _6031_/Z _6033_/A2 _6587_/A2 _6033_/B _7285_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XTAP_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_6935_ _6935_/D _7304_/RN _6935_/CLK _6935_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XPHY_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6866_ _6866_/D _7341_/RN _6866_/CLK _6866_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_22_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5817_ hold5/Z hold109/Z _5819_/S _5817_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6797_ _6797_/D _7304_/RN _6797_/CLK _6797_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5748_ _5856_/A1 _5784_/A2 _5748_/A3 _5838_/A4 _5756_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_41_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5679_ hold5/Z hold135/Z _5681_/S _7061_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_135_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold561 _4234_/Z _6781_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold572 _6865_/Q hold572/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7349_ _7349_/I _7349_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold550 _7349_/I hold550/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_173_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold594 _6797_/Q hold594/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold583 _7341_/Q hold583/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2711 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2766 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4981_ _5369_/A1 _4963_/B _4926_/C _4955_/B _4982_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_51_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3932_ _6935_/Q _5838_/A2 _5532_/A3 _5528_/A2 _3963_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6720_ _6720_/D _7304_/RN _6720_/CLK _6720_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_6651_ _6876_/Q _6651_/A2 _6651_/B _6652_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3863_ _7009_/Q _3962_/A2 _3961_/A2 _7001_/Q _3951_/A2 _7073_/Q _3872_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_20_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5602_ hold388/Z hold659/Z _5608_/S _5602_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6582_ _6582_/A1 _6582_/A2 _6582_/A3 _6582_/A4 _6582_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_164_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3794_ _6898_/Q _5838_/A2 _4405_/A3 _5546_/A2 _3873_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5533_ hold391/Z hold846/Z _5533_/S _5533_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5464_ _5464_/A1 _5464_/A2 _5464_/A3 _5464_/A4 _5464_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_117_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4415_ _4064_/B _4064_/C input97/Z input96/Z _4432_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_5395_ _5396_/A1 _5396_/A2 _5395_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7203_ _7203_/D _7302_/RN _7203_/CLK _7203_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_99_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4346_ hold388/Z hold570/Z _4346_/S _4346_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7134_ _7134_/D _7302_/RN _7134_/CLK _7134_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_101_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4277_ hold136/Z hold5/Z _4281_/S _4277_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7065_ _7065_/D _7265_/RN _7065_/CLK _7065_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_140_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6016_ _6016_/A1 _6016_/A2 _6016_/A3 _6016_/A4 _6026_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_2007 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2029 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2018 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6918_ _6918_/D _6676_/Z _4111_/I1 _6918_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_168_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6849_ _6849_/D _7313_/CLK _6849_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_863 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold380 _5705_/Z _7084_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_2_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold391 _4135_/Z hold391/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_117_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2541 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_53__1374_ clkbuf_4_12_0__1374_/Z net683_320/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_73_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1873 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4200_ hold391/Z hold596/Z _4201_/S _4200_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5180_ _5226_/A1 _5471_/A1 _5180_/B _5439_/C _5440_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4131_ _4131_/A1 _6879_/Q _6872_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4062_ _4062_/A1 _4062_/A2 _4062_/A3 _4062_/A4 _4063_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_96_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4964_ _4926_/C _5288_/A4 _5034_/A2 _4718_/C _5285_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_24_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6703_ _6703_/D _6658_/Z _4108_/B2 _6703_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_32_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3915_ _7120_/Q _5802_/A2 _5784_/A2 _5546_/A2 _3970_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4895_ _4056_/B _4777_/C _5436_/A4 _5445_/A3 _5402_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6634_ _6634_/I0 _7319_/Q _6642_/S _7319_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_165_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3846_ _7105_/Q _3968_/A2 _3846_/B1 _6769_/Q _3846_/C1 _6739_/Q _3849_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_6565_ _6565_/A1 _6565_/A2 _6577_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3777_ _7244_/Q _3981_/A2 _3981_/B1 _7252_/Q _6941_/Q _5544_/S _3780_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_118_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6496_ _7168_/Q _6279_/Z _6299_/Z hold82/I _6575_/B1 hold67/I _6498_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_5516_ hold139/Z hold448/Z _5517_/S _6925_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_161_844 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5447_ _5480_/A2 _5482_/A1 _5446_/Z _5448_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_105_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5378_ _5378_/A1 _5498_/B1 _5379_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4329_ _5535_/B _6653_/A2 _4378_/A1 _5745_/A4 _4331_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_7117_ _7117_/D _7302_/RN _7117_/CLK _7117_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_7048_ _7048_/D _7341_/RN _7048_/CLK _7048_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
Xnet483_116 _4109__6/I _7153_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet483_105 net433_81/I _7164_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_59_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet483_127 net433_99/I _7142_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_47_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet483_138 _4109__8/I _7131_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_86_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet483_149 net833_471/I _7120_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_67_390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_909 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_894 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2360 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2393 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3700_ _3700_/I _3706_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_14_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4680_ _4682_/A2 _5051_/B _5459_/A3 _5355_/A2 _5087_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_119_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3631_ hold67/I _3973_/A2 _3943_/C1 hold66/I _3633_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3562_ _3454_/Z _3498_/B _3644_/A2 _5534_/A2 _3964_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_6350_ _6788_/Q _4019_/Z _6509_/B _7296_/Q _6375_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5301_ _5389_/A2 _5301_/A2 _4661_/C _5153_/B _5327_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_52_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3493_ _3483_/Z hold36/Z _3500_/C _3827_/A2 _3644_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_6281_ _7242_/Q _6563_/A2 _6562_/A3 _6563_/A4 _6334_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5232_ _5232_/A1 _5461_/A1 _5418_/A2 _5232_/A4 _5234_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_130_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5163_ _5330_/B2 _5466_/C _5169_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4114_ _4117_/A1 input86/Z _4115_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5094_ _5353_/A3 _5271_/A4 _5279_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4045_ _6310_/A4 _7276_/Q _6511_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_92_691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5996_ _6103_/A1 _6211_/C _6211_/B _7272_/Q _6260_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_12_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4947_ _4951_/A1 _4951_/A2 _4951_/B1 _4951_/B2 _4947_/C _4967_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_80_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4878_ _5177_/A3 _5153_/A2 _5153_/B _5180_/B _5143_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6617_ _6617_/A1 _6617_/A2 _6618_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_177_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3829_ _6737_/Q _5655_/A4 hold37/I _4405_/A2 _3881_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_20_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6548_ _6548_/A1 _6548_/A2 _6548_/A3 _6548_/A4 _6555_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_161_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6479_ _6479_/A1 _6479_/A2 _6479_/A3 _6479_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_133_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput260 _6935_/Q pll_bypass VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput271 _6726_/Q pll_trim[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_160_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput293 _6732_/Q pll_trim[6] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput282 _6727_/Q pll_trim[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_711 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xload_slew348 hold190/Z _4405_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xload_slew359 _5902_/A3 _5838_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
XFILLER_78_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5850_ hold25/Z hold472/Z _5855_/S _5850_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5781_ hold5/Z hold113/Z hold14/Z _7151_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4801_ _5152_/C _5327_/B _4822_/A4 _5426_/B1 _4803_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_62_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4732_ _4667_/Z _5244_/A2 _5241_/A3 _5489_/A1 _4735_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4663_ _4421_/Z _4487_/Z _4423_/Z _4922_/B _4710_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_9_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3614_ _7014_/Q _3962_/A2 _3961_/A2 _7006_/Q _3962_/B1 _7086_/Q _3616_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6402_ _6788_/Q _4019_/Z _6509_/B _7298_/Q _6428_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4594_ _4443_/Z _5459_/A3 _5226_/A1 _5502_/A2 _5222_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xhold902 hold11/I _4017_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_143_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3545_ _3811_/A1 _3460_/B _3498_/B _4246_/A1 _3977_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_6333_ _6333_/A1 _6333_/A2 _6333_/A3 _6333_/A4 _6333_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_170_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3476_ _6863_/Q _6907_/Q _3496_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_89_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6264_ _6264_/A1 _6264_/A2 _6264_/A3 _6263_/Z _6264_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_5215_ _5347_/A1 _5215_/A2 _5215_/B _5215_/C _5420_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_131_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6195_ _6999_/Q _6258_/B1 _6262_/B1 _7031_/Q _6198_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_85_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5146_ _5330_/A2 _5247_/B _5252_/A4 _5330_/B1 _5426_/A1 _5427_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_5077_ _5459_/A2 _5463_/A1 _5077_/B _5460_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_151_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4028_ _4028_/I _6878_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_72_639 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_831 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5979_ _5979_/A1 _6570_/A2 _6789_/Q _5980_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_40_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_766 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_853 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet783_440 net783_441/I _6769_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet783_451 net833_469/I _6758_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_8_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold209 _5862_/Z _7222_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_152_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3330_ _7277_/Q _6310_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_113_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_847 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5000_ _5004_/A1 input95/Z _5153_/A2 _5279_/B _5002_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_100_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_569 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6951_ _6951_/D _7262_/RN _6951_/CLK _6951_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_53_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5902_ hold37/Z hold17/Z _5902_/A3 hold45/Z _5910_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_6882_ _6882_/D _7341_/RN _6882_/CLK _6882_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5833_ hold139/Z hold516/Z hold18/Z _7197_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_14_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5764_ hold58/Z hold302/Z _5765_/S _5764_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5695_ hold139/Z hold176/Z _5699_/S _5695_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4715_ _5250_/C _5252_/A3 _5244_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4646_ _4684_/B _4437_/Z _5210_/C _5312_/B _4647_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_148_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4577_ _5436_/A4 _5302_/B _4577_/B _4585_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_163_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7365_ _7365_/I _7365_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold710 _4212_/Z _6764_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold721 _4225_/Z _6773_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold743 _5601_/Z _6992_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold754 _6960_/Q hold754/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6316_ _6316_/A1 _6316_/A2 _6325_/A2 _6317_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xhold732 _5858_/Z _7219_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3528_ _3827_/A1 _3827_/A2 _3496_/B _3833_/A2 _3878_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_116_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold787 _5529_/Z _6935_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold765 _4312_/Z _6831_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7296_ _7296_/D _7304_/RN _7302_/CLK _7296_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold776 _7155_/Q hold776/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3459_ _3455_/Z _3460_/C _3498_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_4
XFILLER_103_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold798 _5610_/Z _7000_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_77_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6247_ _6559_/S _6247_/A2 _6247_/B _7293_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6178_ hold64/I _6232_/C _6266_/B _6266_/C _6189_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5129_ _5349_/A1 _5369_/A1 _5267_/C _5327_/B _5328_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_85_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet733_370 net733_381/I _6884_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet733_381 net733_381/I _6853_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet733_392 net783_425/I _6826_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_122_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold81 hold81/I hold81/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_91_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold70 hold70/I hold70/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_29_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold92 hold92/I hold92/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_90_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4500_ _4443_/Z _5459_/A3 _5439_/A1 _5394_/C _4565_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_129_265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5480_ _5435_/B _5480_/A2 _5479_/Z _5480_/A4 _5480_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_4431_ _4774_/A1 _4774_/A2 _4958_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_144_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4362_ _6878_/Q _6879_/Q _6880_/Q _6876_/Q _4362_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_2
X_7150_ _7150_/D _7265_/RN _7150_/CLK _7150_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_125_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4293_ hold25/Z hold161/Z _4298_/S _4293_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3313_ _3313_/I _4016_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
X_7081_ _7081_/D _7281_/RN _7081_/CLK _7081_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_113_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6101_ _7197_/Q _6260_/A2 _6257_/A2 _7133_/Q _6261_/B1 _7165_/Q _6102_/C VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_140_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6032_ _6107_/B _6107_/C _6968_/Q _7275_/Q _6033_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_79_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_399 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_6934_ _6934_/D _7304_/RN _6934_/CLK _6934_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XPHY_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6865_ _6865_/D _7341_/RN _6865_/CLK _6865_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_50_642 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5816_ hold164/Z hold287/Z _5819_/S _5816_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6796_ _6796_/D _7304_/RN _6796_/CLK _7353_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_148_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5747_ hold680/Z hold388/Z _5747_/S _5747_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_157_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5678_ hold164/Z hold294/Z _5681_/S _7060_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_157_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4629_ _4628_/B _5186_/B2 _5046_/C _5062_/A3 _4633_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_135_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold540 _4280_/Z _6805_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_150_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold551 hold551/I hold551/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold562 _6902_/Q hold562/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7279_ _7279_/D _7281_/RN _7281_/CLK _7279_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
Xhold573 _4368_/Z _6865_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold595 _4261_/Z _6797_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold584 _6655_/Z _7341_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_103_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_786 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2745 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_828 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_13__1374_ clkbuf_opt_1_0__1374_/Z net683_317/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_182_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_76__1374_ clkbuf_4_5_0__1374_/Z net783_427/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_122_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput160 wb_rstn_i _7323_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
XFILLER_49_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4980_ _5223_/A1 _4963_/B _5025_/A3 _4955_/B _4982_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_63_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3931_ _6950_/Q _5884_/A2 _6653_/A3 _5552_/A2 _3950_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_44_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6650_ _7323_/Q _6876_/Q _6651_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_149_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3862_ input47/Z _4262_/S _3981_/B1 _7251_/Q _3862_/C _3872_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_31_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5601_ hold391/Z hold742/Z _5608_/S _5601_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_82_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6581_ _6769_/Q _6286_/Z _6581_/B1 _6896_/Q _6582_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_176_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_894 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5532_ _5838_/A4 _6653_/A2 _5532_/A3 _5838_/A2 _5533_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_9_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3793_ _6830_/Q _5856_/A2 _5528_/A2 _5573_/A3 _3847_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_118_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5463_ _5463_/A1 _5493_/B2 _5463_/B _5464_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_172_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4414_ _4064_/B _4064_/C input97/Z input96/Z _4414_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_133_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5394_ _5439_/A1 _5394_/A2 _5439_/C _5394_/C _5396_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_7202_ _7202_/D _7341_/RN _7202_/CLK _7202_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_7133_ _7133_/D _7341_/RN _7133_/CLK _7133_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4345_ hold391/Z hold579/Z _4346_/S _4345_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7064_ _7064_/D _7341_/RN _7064_/CLK _7064_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4276_ _4275_/Z hold564/Z _4282_/S _4276_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_100_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6015_ _7056_/Q _6257_/B1 _6259_/B1 _6976_/Q _6016_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_100_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2019 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2008 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6917_ _6917_/D _6675_/Z _7346_/CLK _6917_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_22_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6848_ _6848_/D _6862_/CLK _6848_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_52_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6779_ _6779_/D _7281_/RN _6779_/CLK _7357_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_176_691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold381 _6999_/Q hold381/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold370 _4297_/Z _6819_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_132_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold392 _4382_/Z _6885_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1852 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1830 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_0__1374_ clkbuf_4_2_0__1374_/Z net433_64/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_60_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1874 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1863 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1896 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4130_ _4131_/A1 _6876_/Q _6873_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_123_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4061_ _4413_/A3 _4413_/A4 _4418_/A1 _4418_/A2 _4065_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_95_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4963_ _5104_/B1 _4965_/C _4963_/B _5105_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_64_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6702_ _6702_/D _6657_/Z _4108_/B2 _6702_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3914_ _6738_/Q _5745_/A4 _5784_/A2 _5528_/A2 _3957_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_189_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6633_ _6633_/A1 _6633_/A2 _6634_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4894_ _5439_/C _5436_/A4 _5445_/A3 _5235_/A1 _5192_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_20_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3845_ _3845_/A1 _3845_/A2 _3845_/A3 _3845_/A4 _3845_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_22_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3776_ _3776_/A1 _3776_/A2 _3790_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6564_ _6735_/Q _6285_/Z _6294_/Z _6882_/Q _6564_/C1 _6894_/Q _6565_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6495_ hold77/I _6575_/A2 _6566_/C1 _7022_/Q _6498_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5515_ hold25/Z hold526/Z _5517_/S _6924_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_173_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_146_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5446_ _4362_/Z _5479_/A2 _5446_/A3 _5482_/A3 _5446_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_105_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5377_ _5371_/Z _5373_/Z _5412_/A2 _5455_/A2 _5380_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_99_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4328_ _3597_/Z _6842_/Q _4328_/S _6842_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7116_ _7116_/D _7302_/RN _7116_/CLK _7116_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xnet483_117 net433_86/I _7152_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet483_106 net433_91/I _7163_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_101_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7047_ _7047_/D _7302_/RN _7047_/CLK _7047_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4259_ hold607/Z _4258_/Z _4263_/S _4259_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet483_128 net683_349/I _7141_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet483_139 net433_66/I _7130_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_83_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_533 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_823 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_569 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3630_ _3630_/A1 _3630_/A2 _3630_/A3 _3634_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3561_ _3827_/A2 _3496_/B _3833_/A2 _5534_/A2 _3943_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_143_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5300_ _5390_/A1 _5404_/A2 _5300_/B _5390_/C _5303_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_6_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3492_ _3483_/Z hold36/Z _3500_/C _3827_/A2 hold37/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6280_ _6563_/A2 _6310_/A4 _7276_/Q _6563_/A4 _6311_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_5_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5231_ _5457_/A1 _4647_/C _5232_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5162_ _5177_/A1 _5484_/A4 _5394_/C _5471_/A1 _5295_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5093_ _4661_/C _4956_/B _5093_/B _5111_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_110_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4113_ _4113_/I _4113_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_56_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4044_ _6584_/B _4019_/Z _5930_/A1 _5930_/A2 _4044_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_140_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_865 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5995_ _7274_/Q _7273_/Q _6235_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4946_ _4963_/B _4926_/C _4955_/B _5107_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_40_729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4877_ _4877_/A1 _5181_/C _4877_/A3 _4881_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_6616_ _6878_/Q _6616_/A2 _6616_/B1 _6640_/B2 _6617_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_165_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3828_ _6894_/Q _5838_/A2 _4405_/A3 _4405_/A2 _3856_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_6547_ _6758_/Q _6573_/A2 _6288_/Z _6762_/Q _6297_/Z _6883_/Q _6548_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_152_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_146_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3759_ _6986_/Q _5700_/A1 _5655_/A4 _4378_/A1 _3769_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6478_ _7263_/Q _6581_/B1 _6312_/Z _7223_/Q _6479_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_134_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5429_ _5429_/A1 _5429_/A2 _5429_/A3 _5491_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
Xoutput261 _6921_/Q pll_dco_ena VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput250 _4127_/Z pad_flash_csb_oe VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput272 _6720_/Q pll_trim[10] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput294 _6733_/Q pll_trim[7] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput283 _6714_/Q pll_trim[20] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_847 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_726 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_435 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_642 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2180 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4800_ _4800_/A1 _5263_/A1 _5263_/A2 _5469_/A3 _4803_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5780_ hold164/Z hold306/Z hold14/Z _7150_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4731_ _5315_/A4 _5235_/A1 _4718_/B _3379_/I _5426_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XTAP_1490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4662_ _4690_/B _5484_/A2 _4690_/C _4469_/B _4787_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_147_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3613_ input9/Z _3850_/B1 _3605_/Z _5544_/S hold75/I _3956_/A2 _3616_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_30_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6401_ _6401_/I0 _7297_/Q _6559_/S _7297_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4593_ _4443_/Z _5459_/A3 _5439_/A1 _5502_/A2 _4595_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xhold903 _6702_/Q hold903/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_134_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_182 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6332_ _6992_/Q _6570_/C1 _6311_/C _7000_/Q _6333_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3544_ _3519_/Z _3534_/C _3460_/B _3831_/A2 _3939_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_3475_ _6703_/Q hold297/Z _6777_/Q _3475_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_116_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_867 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6263_ _6263_/A1 _6263_/A2 _6263_/A3 _6263_/A4 _6263_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_5214_ _3380_/I _4425_/Z _5350_/B _4956_/C _5215_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_131_848 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6194_ _6559_/S _6194_/A2 _6194_/B _7291_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_96_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5145_ _5476_/A1 _5257_/B1 _5148_/B1 _5439_/B _5149_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_28_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5076_ _5079_/A1 _5399_/B _5209_/B1 _5076_/B2 _5229_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_84_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4027_ _6878_/Q _4074_/A2 _6872_/Q _4028_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_38_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5978_ _7281_/Q _6296_/A2 _6324_/A1 _6312_/A4 _6570_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_4929_ _5288_/A4 _4776_/Z _4959_/C _4451_/B _5026_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_165_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_176_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_898 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet783_441 net783_441/I _6768_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet783_430 net783_430/I _6784_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_184_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_537 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6950_ _6950_/D _7262_/RN _6950_/CLK _6950_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_93_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5901_ hold2/Z hold525/Z _5901_/S _7257_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6881_ _6881_/D _7341_/RN _6881_/CLK _6881_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_35_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5832_ hold25/Z hold453/Z hold18/Z _7196_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_62_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5763_ hold5/Z hold434/Z _5765_/S _5763_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4714_ _4765_/A2 _5307_/B _4765_/A1 _5252_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_5694_ hold25/Z hold338/Z _5699_/S _5694_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_163_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4645_ _4469_/B _4759_/C _5312_/B _4684_/B _5084_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_30_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold711 _7211_/Q hold711/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4576_ _4576_/A1 _4576_/A2 _5057_/B _4577_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_162_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7364_ _7364_/I _7364_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold700 _6821_/Q hold700/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_162_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3527_ hold28/Z hold36/Z _3500_/C _3477_/Z _3527_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_115_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6315_ _6528_/A2 _6581_/B1 _6580_/B1 _6566_/C1 _6316_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_104_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold733 _6984_/Q hold733/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold744 _7001_/Q hold744/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold722 _6897_/Q hold722/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold755 _6719_/Q hold755/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold766 _7088_/Q hold766/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_89_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold788 _7170_/Q hold788/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7295_ _7295_/D _7304_/RN _7302_/CLK _7295_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold777 _7089_/Q hold777/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3458_ _6863_/Q hold20/Z _3460_/C _3534_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_104_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold799 _6710_/Q hold799/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6246_ _6246_/A1 _6246_/A2 _6788_/Q _7292_/Q _6247_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_103_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6177_ _6177_/A1 _6177_/A2 _6177_/A3 _6176_/Z _6177_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_29_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3389_ _6709_/Q _6708_/Q _6707_/Q _6776_/Q _3389_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_5128_ _5128_/A1 _5376_/A1 _5502_/B1 _5389_/A2 _5130_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_85_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5059_ _5323_/A1 _5302_/B _5355_/B _5372_/A1 _5356_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_72_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet733_371 net733_381/I _6883_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet733_360 _4109__16/I _6894_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet733_382 net833_472/I _6844_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet733_393 net783_424/I _6825_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_20_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold82 hold82/I hold82/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold71 hold71/I hold71/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold60 hold60/I hold60/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_75_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold93 hold93/I hold93/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_29_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_36__1374_ clkbuf_4_14_0__1374_/Z _4109__28/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_16_375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_99__1374_ clkbuf_4_1_0__1374_/Z net833_456/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_726 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4430_ _4922_/B _4421_/Z _4425_/Z _4774_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_117_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4361_ _6878_/Q _6879_/Q _6880_/Q _6876_/Q _4365_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_113_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6100_ _7205_/Q _6233_/A2 _6266_/B _7189_/Q _6102_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4292_ hold388/Z hold587/Z _4298_/S _4292_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_125_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7080_ _7080_/D _7281_/RN _7080_/CLK _7080_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_140_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6031_ _6031_/A1 _6031_/A2 _6031_/A3 _6031_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_79_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_573 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_6933_ _6933_/D _7304_/RN _6933_/CLK _6933_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XPHY_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_6864_ _6864_/D _7341_/RN _6864_/CLK _6864_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_179_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5815_ hold139/Z hold450/Z _5819_/S _5815_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6795_ _6795_/D _7304_/RN _6795_/CLK _7352_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_50_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5746_ hold772/Z hold391/Z _5747_/S _5746_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5677_ hold139/Z hold152/Z _5681_/S _7059_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4628_ _5046_/A1 _5046_/A2 _4628_/B _5046_/C _5459_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_163_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold530 _7114_/Q hold530/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7347_ _7347_/D _6699_/Z _4108_/B2 _7347_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4559_ _5082_/C _5347_/A2 _4560_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold541 _6834_/Q hold541/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold563 _6901_/Q hold563/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_2_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold552 hold552/I _6938_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold585 _7049_/Q hold585/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7278_ _7278_/D _7281_/RN _7281_/CLK _7278_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
Xhold574 _6889_/Q hold574/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold596 _6756_/Q hold596/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_103_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6229_ _6225_/Z _6229_/A2 _6229_/A3 _6229_/A4 _6229_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_57_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_890 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2746 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2713 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_185_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_214 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_4_12_0__1374_ clkbuf_3_6_0__1374_/Z clkbuf_4_12_0__1374_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_134_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput161 wb_sel_i[0] _6607_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput150 wb_dat_i[2] _6620_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_64_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3930_ input93/Z _5884_/A2 _5856_/A2 _5532_/A3 _3976_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_189_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3861_ _3861_/A1 _3861_/A2 _3861_/A3 _3861_/A4 _3861_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_32_654 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5600_ _5646_/A2 _4227_/B _5820_/A2 _5866_/A3 _5608_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_6580_ _6854_/Q _6311_/C _6580_/B1 _6900_/Q _6582_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3792_ _3791_/Z hold880/Z _3888_/S _6914_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5531_ hold391/Z hold739/Z _5531_/S _6936_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_117_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5462_ _5462_/A1 _5462_/A2 _5462_/A3 _5462_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_173_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7201_ hold19/Z _7265_/RN _7201_/CLK _7201_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_105_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4413_ input99/Z input98/Z _4413_/A3 _4413_/A4 _4432_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_5393_ _5439_/C _5393_/A2 _5393_/A3 _4686_/B _5396_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_132_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7132_ _7132_/D _7341_/RN _7132_/CLK _7132_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_125_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4344_ hold45/Z _4405_/A2 _5893_/A3 _4378_/A1 _4346_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_7063_ _7063_/D _7281_/RN _7063_/CLK hold56/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_141_773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4275_ hold185/Z hold164/Z _4281_/S _4275_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_140_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6014_ _6103_/A1 _7274_/Q _7273_/Q _7272_/Q _6259_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_67_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2009 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1319 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6916_ _6916_/D _6674_/Z _4108_/B2 _6916_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_23_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6847_ _6847_/D _6862_/CLK _6847_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_149_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_82__1374_ clkbuf_4_4_0__1374_/Z net433_93/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_22_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6778_ _6778_/D _6669_/Z _7346_/CLK _6778_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_183_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5729_ hold388/Z hold694/Z _5735_/S _7105_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold360 _7083_/Q hold360/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold371 _7246_/Q hold371/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_431 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold382 _5608_/Z _6999_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_117_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold393 _7045_/Q hold393/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_18_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2532 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1842 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1831 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1820 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1875 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1864 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1853 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_827 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4060_ _4060_/A1 _4060_/A2 _4418_/A3 _4418_/A4 _4062_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_95_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4962_ _5104_/B1 _4965_/C _4962_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_51_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6701_ _6701_/D _6656_/Z _4108_/B2 _6701_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4893_ _5321_/A3 _5489_/B1 _4893_/B _4897_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_32_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3913_ _6770_/Q _5802_/A2 _5546_/A2 _3527_/Z _3963_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6632_ _6878_/Q _6632_/A2 _6632_/B1 _6640_/B2 _6633_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3844_ input15/Z _3939_/B1 _3950_/B1 _7041_/Q _3845_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_20_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3775_ _7228_/Q _3964_/A2 _4281_/S input37/Z _3776_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_118_512 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6563_ _6751_/Q _6563_/A2 _6563_/A3 _6563_/A4 _6582_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_118_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6494_ _7136_/Q _6287_/Z _6300_/Z _7014_/Q _6319_/Z hold75/I _6498_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_5514_ hold388/Z hold783/Z _5517_/S _6923_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_145_364 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5445_ _3379_/I _5445_/A2 _5445_/A3 _5194_/C _5482_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_106_718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5376_ _5376_/A1 _5454_/B1 _5376_/B1 _4956_/C _5376_/C _5455_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_7115_ _7115_/D _7304_/RN _7115_/CLK _7115_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_160_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4327_ _6602_/A1 _4328_/S _4327_/B _6841_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xnet483_118 net433_86/I _7151_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet483_107 _4109__48/I _7162_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4258_ hold224/Z hold5/Z _4262_/S _4258_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7046_ _7046_/D _7302_/RN _7046_/CLK _7046_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_170_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet483_129 net483_129/I _7140_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4189_ hold2/Z hold141/Z _4189_/S _4189_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_27_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_137_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_843 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_868 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_845 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold190 hold190/I hold190/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_104_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2395 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3560_ input19/Z _3971_/A2 _3559_/Z hold98/I _3586_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5230_ _5230_/A1 _5230_/A2 _5230_/B _5230_/C _5418_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_3491_ _3489_/Z _3490_/Z _3491_/B _3500_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_115_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_537 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_7_0__1374_ clkbuf_0__1374_/Z clkbuf_3_7_0__1374_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_69_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5161_ _5295_/A1 _5466_/A1 _5177_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5092_ _4947_/C _5409_/A2 _5092_/B _5409_/C _5118_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_96_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4112_ _7343_/Q input88/Z _4113_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_68_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4043_ _6584_/B _4019_/Z _6532_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_83_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5994_ _6036_/A3 _6211_/B _7274_/Q _7271_/Q _6259_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_64_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4945_ _4995_/A4 _4926_/B _4955_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_178_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4876_ _5466_/B _5037_/A1 _5392_/A1 _5397_/A1 _4877_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_6615_ _6880_/Q _6615_/A2 _6615_/B1 _6879_/Q _6617_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_177_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3827_ _3827_/A1 _3827_/A2 _3496_/B _4227_/A2 _3851_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_119_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6546_ _6764_/Q _6575_/A2 _6566_/C1 _6866_/Q _6548_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3758_ input5/Z _5700_/A1 _5748_/A3 _5532_/A3 _3780_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6477_ _7159_/Q _6286_/Z _6311_/C _7005_/Q _6479_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3689_ _7116_/Q _3969_/A2 _3956_/A2 _7126_/Q _3691_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5428_ _5428_/A1 _5428_/A2 _5428_/A3 _5428_/A4 _5429_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_88_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput262 _6922_/Q pll_div[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput251 _4116_/Z pad_flash_io0_do VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput240 _7351_/Z mgmt_gpio_out[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5359_ _5359_/A1 _5462_/A1 _5362_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput273 _6721_/Q pll_trim[11] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput284 _6715_/Q pll_trim[21] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_837 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput295 _6718_/Q pll_trim[8] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_102_765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7029_ _7029_/D _7302_/RN _7029_/CLK _7029_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_101_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_844 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_188_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_4_0_0__1374_ clkbuf_4_1_0__1374_/I net733_398/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_124_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_719 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4730_ _5262_/A4 _5301_/A2 _4661_/C _3380_/I _5489_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XTAP_1491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_159_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4661_ _3379_/I _3380_/I _4718_/B _4661_/C _4759_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_9_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3612_ _3612_/A1 _3612_/A2 _3612_/A3 _3861_/A2 _3637_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_6400_ _6400_/A1 _6400_/A2 _6400_/B _6401_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4592_ _4592_/A1 _4592_/A2 _5063_/B _4592_/A4 _4595_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_6331_ _7178_/Q _6571_/C1 _6568_/B1 _7112_/Q _6333_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_143_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3543_ _3604_/A2 _3811_/A1 _3511_/C _3833_/A2 _3953_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_3474_ _3604_/A2 _3507_/C _3827_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_131_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6262_ _6898_/Q _6262_/A2 _6262_/B1 _6869_/Q _6263_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5213_ _5464_/A1 _5213_/A2 _5421_/A1 _5213_/A4 _5216_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_142_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6193_ _5917_/B _6587_/A2 _7291_/Q _6194_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5144_ _5144_/A1 _5335_/A1 _5144_/A3 _5149_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_56_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5075_ _5071_/Z _5073_/Z _5361_/A2 _5075_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_84_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4026_ _7342_/Q hold44/I _6994_/Q _4026_/C _4131_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_44_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5977_ _5975_/B _7280_/Q _6325_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_52_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4928_ _4965_/A2 _4776_/Z _4959_/C _4451_/B _5381_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_100_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4859_ _5445_/A2 _5177_/A3 _5153_/B _5437_/A4 _4861_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_119_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6529_ _6584_/A1 _6529_/A2 _6529_/A3 _6529_/A4 _6529_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_134_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_188_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_674 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet783_420 net783_420/I _6798_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_70_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet783_431 net783_431/I _6783_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet783_442 _4109__2/I _6767_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_7_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_59__1374_ clkbuf_4_12_0__1374_/Z net433_76/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_98_516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5900_ hold58/Z hold192/Z _5901_/S _7256_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_19_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6880_ _6880_/D _7323_/RN _7323_/CLK _6880_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_62_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5831_ hold388/Z hold828/Z hold18/Z _7195_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5762_ hold164/Z hold484/Z _5765_/S _7134_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_188_871 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4713_ _5244_/A2 _5241_/A3 _4750_/A3 _4750_/A4 _5330_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_5693_ hold388/Z hold829/Z _5699_/S _5693_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_147_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4644_ _4686_/B _5307_/B _4694_/B _4922_/B _5194_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xhold712 _5849_/Z _7211_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4575_ _5439_/A1 _5436_/A2 _4624_/A2 _5210_/B _5057_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_146_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7363_ _7363_/I _7363_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold701 _4300_/Z _6821_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_115_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6314_ _6313_/Z _6312_/Z _6310_/Z _6575_/B1 _6318_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xhold734 _5592_/Z _6984_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold745 _5611_/Z _7001_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold723 _4400_/Z _6897_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7294_ _7294_/D _7304_/RN _7304_/CLK _7294_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3526_ _5534_/A1 _3477_/Z _3496_/B _3831_/A2 _3956_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_116_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold756 _4153_/Z _6719_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold767 _6750_/Q hold767/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6245_ _5917_/B _6587_/A2 _7293_/Q _6247_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xhold778 _7154_/Q hold778/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3457_ _4016_/A2 _4073_/B1 _3457_/B _6863_/Q _3460_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_103_359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold789 _5803_/Z _7170_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_39_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6176_ _6176_/A1 _6176_/A2 _6176_/A3 _6176_/A4 _6176_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_3388_ _6709_/Q _6708_/Q _6707_/Q _4073_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_5127_ _4725_/Z _5199_/A2 _5127_/B _5243_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5058_ _5058_/A1 _5420_/C _5217_/C _5061_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_4009_ _4015_/S _4009_/A2 _4009_/B _6703_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_44_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet733_361 net733_381/I _6893_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet733_372 net833_474/I _6882_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet733_383 net433_64/I _6843_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_4_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_793 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet733_394 net733_397/I _6824_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold50 hold50/I hold50/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_121_178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold83 hold83/I hold83/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_102_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold72 hold72/I hold72/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold61 hold61/I hold61/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_48_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_714 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold94 hold94/I hold94/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_16_332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_360 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_176_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4360_ _6878_/Q _6879_/Q _6880_/Q _5323_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_172_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4291_ hold391/Z hold671/Z _4298_/S _4291_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6030_ _7096_/Q _6232_/C _6266_/B _6266_/C _6031_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_100_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_6932_ _6932_/D _7262_/RN _6932_/CLK _6932_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_35_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6863_ _6863_/D _7323_/RN _7323_/CLK _6863_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_25_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5814_ hold25/Z hold470/Z _5819_/S _5814_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_23_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6794_ _6794_/D _7304_/RN _6794_/CLK _7351_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_148_543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5745_ _5838_/A4 _6653_/A2 _5784_/A2 _5745_/A4 _5747_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_5676_ hold25/Z hold440/Z _5681_/S _7058_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4627_ _4627_/A1 _4627_/A2 _5229_/A3 _4627_/A4 _4633_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_135_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold520 _7259_/Q hold520/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold553 _7360_/I hold553/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_173_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4558_ _4558_/A1 _4558_/A2 _5051_/B _5051_/C _4560_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
Xhold542 _4316_/Z _6834_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7346_ _7346_/D _6698_/Z _7346_/CLK _7346_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold531 _7204_/Q hold531/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_4489_ _5235_/A1 _4718_/B _5034_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xhold586 _7048_/Q hold586/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold564 _7356_/I hold564/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3509_ _3454_/Z _3498_/B _3604_/A2 hold462/Z _5640_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_7277_ _7277_/D _7281_/RN _7281_/CLK _7277_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
Xhold575 _6864_/Q hold575/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold597 _4200_/Z _6756_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xclkbuf_leaf_42__1374_ clkbuf_4_14_0__1374_/Z net433_54/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6228_ _6891_/Q _6260_/A2 _6258_/B1 _6843_/Q _6229_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_89_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6159_ _7069_/Q _6258_/C1 _6256_/B1 _7085_/Q _6161_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_58_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_880 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2714 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_844 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput151 wb_dat_i[30] _6635_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput162 wb_sel_i[1] _6647_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput140 wb_dat_i[20] _6628_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_76_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3860_ _7259_/Q _3964_/C1 _4281_/S input72/Z _3861_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_177_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3791_ _6913_/Q _3790_/Z _3887_/S _3791_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5530_ _5535_/B hold463/Z hold37/Z _7302_/RN _5531_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_5461_ _5461_/A1 _5461_/A2 _5461_/A3 _5462_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_117_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4412_ input99/Z input98/Z _4413_/A3 _4413_/A4 _4412_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_172_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7200_ _7200_/D _7265_/RN _7200_/CLK _7200_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_68_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5392_ _5392_/A1 _4423_/Z _4718_/B _4487_/Z _5393_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_172_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7131_ _7131_/D _7341_/RN _7131_/CLK _7131_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_4343_ _3597_/Z _6852_/Q _4343_/S _6852_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7062_ _7062_/D _7265_/RN _7062_/CLK hold66/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4274_ _4273_/Z hold663/Z _4282_/S _4274_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6013_ _6036_/A3 _6103_/A1 _6211_/C _7273_/Q _6257_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_67_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6915_ _6915_/D _6673_/Z _4111_/I1 _6915_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_35_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6846_ _6846_/D _6862_/CLK _6846_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_52_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6777_ _6777_/D _6668_/Z _4111_/I1 _6777_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_50_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3989_ _6709_/Q _3989_/A2 _6709_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_22_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5728_ hold391/Z hold780/Z _5735_/S _7104_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_182_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5659_ hold139/Z hold604/Z _5663_/S _7043_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_163_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7329_ _7329_/D _6683_/Z _4089_/I1 hold24/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold361 _5704_/Z _7083_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_89_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold350 _7140_/Q hold350/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold394 _7369_/I hold394/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold372 _7013_/Q hold372/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold383 _6732_/Q hold383/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2500 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2533 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2577 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1843 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1832 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1821 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1876 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1865 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1887 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1898 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_833 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4961_ _4995_/A4 _4961_/A2 _5210_/B _5476_/A1 _4965_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_92_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6700_ _6700_/D _4132_/Z _4108_/B2 hold11/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4892_ _5307_/B _5439_/C _5036_/A2 _5468_/A1 _5317_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_3912_ _6885_/Q _5655_/A4 hold29/I hold190/I _3980_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_6631_ _6880_/Q _6631_/A2 _6631_/B1 _6879_/Q _6633_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3843_ _7057_/Q _3943_/C1 _3973_/B1 _6735_/Q _3843_/C _3845_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_32_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3774_ input58/Z _4262_/S _4264_/A1 input54/Z _3776_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6562_ _6869_/Q _6562_/A2 _6562_/A3 _6562_/A4 _6583_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_173_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6493_ hold64/I _6284_/Z _6568_/B1 hold62/I _6499_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5513_ hold391/Z hold840/Z _5517_/S _6922_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_145_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5444_ _3379_/I _5444_/A2 _5444_/B _5448_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_161_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5375_ _5375_/A1 _4965_/C _5376_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7114_ _7114_/D _7302_/RN _7114_/CLK _7114_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_114_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4326_ _4328_/S _6841_/Q _4327_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4257_ hold637/Z _4256_/Z _4263_/S _4257_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xnet483_108 net533_176/I _7161_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7045_ _7045_/D _7302_/RN _7045_/CLK _7045_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xnet483_119 net433_81/I _7150_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_86_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4188_ hold58/Z hold72/Z _4189_/S hold73/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_28_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6829_ _6829_/D _7304_/RN _6829_/CLK _6829_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_51_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold180 _4159_/Z _6725_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_132_571 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold191 _4383_/Z _6886_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_77_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1640 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3490_ _6705_/Q _6777_/Q _3490_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_127_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5160_ _5502_/A1 _5502_/A2 _5502_/B1 _5502_/B2 _5179_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5091_ _5476_/A1 _5093_/B _5091_/B _5091_/C _5092_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_96_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4111_ input83/Z _4111_/I1 _7343_/Q _4111_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_111_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4042_ _6787_/Q _6945_/Q _4051_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_639 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5993_ _6211_/C _7273_/Q _6080_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_178_711 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4944_ _4951_/A1 _4951_/A2 _4951_/B1 _4951_/B2 _5410_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_64_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4875_ _5034_/A2 _5466_/B _5392_/A1 _5397_/A1 _5181_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_6614_ _6614_/I0 _7314_/Q _6642_/S _7314_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_137_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3826_ _3827_/A1 _3827_/A2 _3496_/B _4246_/A2 _3955_/C2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_137_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3757_ hold173/I _3498_/B _3454_/Z _5902_/A3 _3757_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_118_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6545_ _6756_/Q _6287_/Z _6300_/Z _6864_/Q _6319_/Z _6752_/Q _6548_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_161_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6476_ _7255_/Q _6580_/B1 _6309_/Z _7239_/Q _6747_/Q _6579_/A2 _6479_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_3688_ _7142_/Q _3958_/A2 _3850_/B1 input7/Z _3956_/B1 _7158_/Q _3691_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
Xoutput230 _7370_/Z mgmt_gpio_out[29] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_134_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5427_ _5427_/A1 _5427_/A2 _5427_/A3 _5470_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
Xoutput252 _4115_/ZN pad_flash_io0_ie VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput241 _7352_/Z mgmt_gpio_out[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5358_ _4597_/Z _5459_/A1 _5358_/B _5358_/C _5462_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_161_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput263 _6923_/Q pll_div[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput274 _6722_/Q pll_trim[12] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput285 _6716_/Q pll_trim[22] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_181_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4309_ hold391/Z hold702/Z _4310_/S _6829_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xoutput296 _6719_/Q pll_trim[9] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5289_ _5289_/A1 _5386_/A1 _5381_/B _5292_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_7028_ _7028_/D _7281_/RN _7028_/CLK _7028_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_87_466 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_639 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_19__1374_ clkbuf_4_10_0__1374_/Z net433_91/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_2193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2182 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1470 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4660_ _5262_/A4 _5301_/A2 _4661_/C _3380_/I _5466_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_3611_ hold74/I _3943_/A2 _3977_/A2 input27/Z _4243_/S input50/Z _3612_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_80_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4591_ _4690_/C _4487_/Z _5466_/B _5503_/A1 _4592_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_162_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6330_ _7162_/Q _6279_/Z _6578_/C1 _7170_/Q _6333_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3542_ _3454_/Z _3498_/B _3644_/A2 _3831_/A2 _3981_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_127_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3473_ _6863_/Q hold7/Z _3473_/B _3473_/C hold8/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_116_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6261_ _6854_/Q _6261_/A2 _6261_/B1 _6884_/Q _6263_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5212_ _5484_/A4 _5218_/A2 _5351_/B1 _5463_/B _5212_/C _5213_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_170_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6192_ _6192_/A1 _6192_/A2 _6788_/Q _7290_/Q _6194_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_124_891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5143_ _5247_/B _5369_/A2 _5252_/A4 _5143_/B _5144_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_96_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5074_ _5323_/A1 _5226_/A2 _5074_/B1 _5360_/B _5361_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_69_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4025_ _4107_/A1 _4025_/A2 input67/Z _6946_/Q _4074_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_84_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5976_ _6312_/A4 _7281_/Q _6561_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_13_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4927_ _4951_/B1 _5410_/A2 _4995_/A4 _4951_/B2 _4965_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_21_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4858_ _4858_/A1 _5438_/A1 _5485_/A1 _4858_/A4 _4858_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_60_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_166_758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3809_ _6867_/Q _4378_/A1 _5838_/A2 _4405_/A2 _3866_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_180_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4789_ _4693_/Z _4706_/Z _5489_/A1 _5255_/B _4791_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_180_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6528_ _7031_/Q _6528_/A2 _6312_/Z _7225_/Q _6529_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_4_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6459_ _7029_/Q _6562_/A2 _6562_/A3 _6562_/A4 _6480_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_133_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet783_410 net783_411/I _6808_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet783_432 net783_433/I _6782_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet783_421 net783_421/I _6797_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet783_443 net833_471/I _6766_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_144_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_6__1374_ clkbuf_4_3_0__1374_/Z net833_474/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_66_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_801 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5830_ hold391/Z hold870/Z hold18/Z _7194_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_61_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5761_ hold139/Z hold374/Z _5765_/S _5761_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_98_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4712_ _5327_/B _4822_/A4 _5250_/C _5131_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_30_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5692_ hold391/Z hold832/Z _5699_/S _5692_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_175_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4643_ _5459_/A3 _5086_/A2 _5372_/A1 _5051_/B _4647_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_162_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4574_ _5466_/B _5307_/B _4684_/B _5294_/C _5302_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_7362_ _7362_/I _7362_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold702 _6829_/Q hold702/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold724 _7097_/Q hold724/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold746 _6910_/Q hold746/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3525_ input51/Z hold37/I _5902_/A3 _6653_/A2 _3580_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6313_ _6313_/A1 _6300_/Z _6564_/C1 _6309_/Z _6313_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
Xhold713 _6755_/Q hold713/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7293_ _7293_/D _7304_/RN _7302_/CLK _7293_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold735 _6770_/Q hold735/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_171_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold757 _6727_/Q hold757/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold768 _4191_/Z _6750_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold779 _7112_/Q hold779/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_6244_ _6788_/Q _6244_/A2 _6246_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3456_ _4073_/B1 input58/Z _3457_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_143_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6175_ _7094_/Q _6262_/A2 _6257_/B1 hold66/I _6176_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_85_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3387_ _6709_/Q _6708_/Q _6707_/Q _3387_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_130_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5126_ _5131_/A1 _5376_/A1 _5502_/B1 _5484_/A4 _5242_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_57_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5057_ _5347_/A1 _4568_/Z _5271_/A1 _5057_/B _5217_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_38_650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4008_ hold897/Z _4015_/S _4009_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_856 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5959_ _7277_/Q _7276_/Q _6563_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_71_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_65__1374_ clkbuf_4_13_0__1374_/Z net633_261/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_139_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet733_362 net433_67/I _6892_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet733_373 net733_373/I _6881_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_134_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet733_384 net433_67/I _6834_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet733_395 net783_425/I _6823_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_88_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold40 hold40/I hold40/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_88_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold51 hold51/I hold51/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_76_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold73 hold73/I hold73/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_29_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold62 hold62/I hold62/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_36_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold84 hold84/I hold84/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold95 hold95/I hold95/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_63_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4290_ _4243_/S _5564_/A3 _4227_/B _4298_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_125_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_793 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6931_ _6931_/D _7262_/RN _6931_/CLK _6931_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_47_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6862_ _6862_/D _6862_/CLK _6862_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5813_ hold388/Z hold748/Z _5819_/S _5813_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_319 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6793_ _6793_/D _7304_/RN _6793_/CLK _7350_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_10_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5744_ hold340/Z hold2/Z _5744_/S _7119_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5675_ hold388/Z hold831/Z _5681_/S _7057_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_176_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4626_ _4443_/Z _5459_/A3 _5323_/A1 _5399_/B _4627_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_151_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold510 _7190_/Q hold510/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_7345_ _7345_/D _6697_/Z _7346_/CLK _7345_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold554 _4236_/Z _6782_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_150_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4557_ _4684_/B _5307_/B _5436_/A2 _5323_/A1 _4558_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_132_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold521 _5904_/Z _7259_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_116_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold543 _6820_/Q hold543/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold532 _5841_/Z _7204_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
Xhold587 _6814_/Q hold587/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_173_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold565 _4276_/Z _6803_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3508_ _3473_/B _3511_/C _4246_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_7276_ _7276_/D _7281_/RN _7281_/CLK _7276_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_4488_ _5301_/A2 _4661_/C _5445_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold576 _4367_/Z _6864_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
X_3439_ hold24/Z hold387/Z _3440_/S _7329_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_131_466 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6227_ _6897_/Q _6262_/A2 _6261_/A2 _6853_/Q _6229_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold598 _7354_/I hold598/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_131_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6158_ _7061_/Q _6257_/B1 _6259_/B1 _6981_/Q _6161_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5109_ _5109_/A1 _5109_/A2 _5498_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_100_831 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_881 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_892 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6089_ _7019_/Q _6259_/A2 _6259_/B1 _6979_/Q _6091_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_100_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2726 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2715 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2748 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput141 wb_dat_i[21] _6632_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput130 wb_dat_i[11] _6623_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput152 wb_dat_i[31] _6639_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput163 wb_sel_i[2] _6646_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_76_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_715 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3790_ _3790_/A1 _3790_/A2 _3790_/A3 _3789_/Z _3790_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_2
XFILLER_20_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_180 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5460_ _5460_/A1 _5460_/A2 _5461_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_158_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_845 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4411_ _4960_/C _4959_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_8
X_5391_ _5466_/B _5391_/A2 _5391_/B _5486_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4342_ _6602_/A1 _4343_/S _4342_/B _6851_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7130_ _7130_/D _7262_/RN _7130_/CLK _7130_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_7061_ _7061_/D _7265_/RN _7061_/CLK _7061_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_141_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4273_ hold366/Z hold139/Z _4281_/S _4273_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6012_ _7080_/Q _6256_/B1 _6262_/B1 _7024_/Q _6016_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
.ends

