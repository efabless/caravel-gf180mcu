VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 3000.000 BY 3000.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 33.040 3004.800 34.160 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 2032.800 3004.800 2033.920 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 2232.720 3004.800 2233.840 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 2432.640 3004.800 2433.760 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 2632.560 3004.800 2633.680 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 2832.480 3004.800 2833.600 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2943.920 2997.600 2945.040 3004.800 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2610.720 2997.600 2611.840 3004.800 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2276.960 2997.600 2278.080 3004.800 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1943.760 2997.600 1944.880 3004.800 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1610.560 2997.600 1611.680 3004.800 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 232.960 3004.800 234.080 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1276.800 2997.600 1277.920 3004.800 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 943.600 2997.600 944.720 3004.800 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 610.400 2997.600 611.520 3004.800 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 276.640 2997.600 277.760 3004.800 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2963.520 2.400 2964.640 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2749.040 2.400 2750.160 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2535.120 2.400 2536.240 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2320.640 2.400 2321.760 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2106.160 2.400 2107.280 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1892.240 2.400 1893.360 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 432.880 3004.800 434.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1677.760 2.400 1678.880 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1463.280 2.400 1464.400 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1249.360 2.400 1250.480 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1034.880 2.400 1036.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 820.960 2.400 822.080 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 606.480 2.400 607.600 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 392.000 2.400 393.120 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 178.080 2.400 179.200 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 632.800 3004.800 633.920 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 832.720 3004.800 833.840 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 1032.640 3004.800 1033.760 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 1232.560 3004.800 1233.680 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 1432.480 3004.800 1433.600 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 1632.960 3004.800 1634.080 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 1832.880 3004.800 1834.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 166.320 3004.800 167.440 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 2166.080 3004.800 2167.200 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 2366.000 3004.800 2367.120 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 2565.920 3004.800 2567.040 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 2765.840 3004.800 2766.960 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 2965.760 3004.800 2966.880 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2721.600 2997.600 2722.720 3004.800 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2388.400 2997.600 2389.520 3004.800 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2055.200 2997.600 2056.320 3004.800 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1721.440 2997.600 1722.560 3004.800 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1388.240 2997.600 1389.360 3004.800 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 366.240 3004.800 367.360 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1055.040 2997.600 1056.160 3004.800 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 721.280 2997.600 722.400 3004.800 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 388.080 2997.600 389.200 3004.800 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 54.880 2997.600 56.000 3004.800 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2820.720 2.400 2821.840 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2606.240 2.400 2607.360 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2392.320 2.400 2393.440 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2177.840 2.400 2178.960 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1963.360 2.400 1964.480 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1749.440 2.400 1750.560 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 566.160 3004.800 567.280 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1534.960 2.400 1536.080 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1320.480 2.400 1321.600 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1106.560 2.400 1107.680 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 892.080 2.400 893.200 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 677.600 2.400 678.720 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 463.680 2.400 464.800 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 249.200 2.400 250.320 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 35.280 2.400 36.400 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 766.080 3004.800 767.200 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 966.000 3004.800 967.120 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 1165.920 3004.800 1167.040 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 1365.840 3004.800 1366.960 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 1566.320 3004.800 1567.440 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 1766.240 3004.800 1767.360 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 1966.160 3004.800 1967.280 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 99.680 3004.800 100.800 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 2099.440 3004.800 2100.560 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 2299.360 3004.800 2300.480 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 2499.280 3004.800 2500.400 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 2699.200 3004.800 2700.320 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 2899.120 3004.800 2900.240 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2833.040 2997.600 2834.160 3004.800 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2499.280 2997.600 2500.400 3004.800 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2166.080 2997.600 2167.200 3004.800 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1832.880 2997.600 1834.000 3004.800 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1499.120 2997.600 1500.240 3004.800 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 299.600 3004.800 300.720 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1165.920 2997.600 1167.040 3004.800 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 832.720 2997.600 833.840 3004.800 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 498.960 2997.600 500.080 3004.800 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 165.760 2997.600 166.880 3004.800 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2891.840 2.400 2892.960 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2677.920 2.400 2679.040 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2463.440 2.400 2464.560 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2248.960 2.400 2250.080 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2035.040 2.400 2036.160 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1820.560 2.400 1821.680 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 499.520 3004.800 500.640 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1606.640 2.400 1607.760 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1392.160 2.400 1393.280 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1177.680 2.400 1178.800 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 963.760 2.400 964.880 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 749.280 2.400 750.400 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 534.800 2.400 535.920 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 320.880 2.400 322.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 106.400 2.400 107.520 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 699.440 3004.800 700.560 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 899.360 3004.800 900.480 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 1099.280 3004.800 1100.400 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 1299.200 3004.800 1300.320 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 1499.120 3004.800 1500.240 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 1699.600 3004.800 1700.720 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 1899.520 3004.800 1900.640 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1056.720 -4.800 1057.840 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1354.640 -4.800 1355.760 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1384.880 -4.800 1386.000 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1414.560 -4.800 1415.680 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1444.240 -4.800 1445.360 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1473.920 -4.800 1475.040 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1504.160 -4.800 1505.280 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1533.840 -4.800 1534.960 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1563.520 -4.800 1564.640 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1593.200 -4.800 1594.320 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1622.880 -4.800 1624.000 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1086.400 -4.800 1087.520 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1653.120 -4.800 1654.240 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1682.800 -4.800 1683.920 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1712.480 -4.800 1713.600 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1742.160 -4.800 1743.280 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1772.400 -4.800 1773.520 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1802.080 -4.800 1803.200 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1831.760 -4.800 1832.880 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1861.440 -4.800 1862.560 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1891.120 -4.800 1892.240 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1921.360 -4.800 1922.480 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1116.640 -4.800 1117.760 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1951.040 -4.800 1952.160 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1980.720 -4.800 1981.840 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2010.400 -4.800 2011.520 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2040.640 -4.800 2041.760 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2070.320 -4.800 2071.440 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2100.000 -4.800 2101.120 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2129.680 -4.800 2130.800 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2159.360 -4.800 2160.480 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2189.600 -4.800 2190.720 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2219.280 -4.800 2220.400 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1146.320 -4.800 1147.440 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2248.960 -4.800 2250.080 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2278.640 -4.800 2279.760 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2308.880 -4.800 2310.000 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2338.560 -4.800 2339.680 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2368.240 -4.800 2369.360 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2397.920 -4.800 2399.040 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2427.600 -4.800 2428.720 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2457.840 -4.800 2458.960 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2487.520 -4.800 2488.640 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2517.200 -4.800 2518.320 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1176.000 -4.800 1177.120 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2546.880 -4.800 2548.000 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2577.120 -4.800 2578.240 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2606.800 -4.800 2607.920 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2636.480 -4.800 2637.600 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2666.160 -4.800 2667.280 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2696.400 -4.800 2697.520 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2726.080 -4.800 2727.200 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2755.760 -4.800 2756.880 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2785.440 -4.800 2786.560 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2815.120 -4.800 2816.240 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1205.680 -4.800 1206.800 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2845.360 -4.800 2846.480 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2875.040 -4.800 2876.160 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2904.720 -4.800 2905.840 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2934.400 -4.800 2935.520 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1235.360 -4.800 1236.480 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1265.600 -4.800 1266.720 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1295.280 -4.800 1296.400 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1324.960 -4.800 1326.080 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1066.800 -4.800 1067.920 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1364.720 -4.800 1365.840 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1394.400 -4.800 1395.520 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1424.640 -4.800 1425.760 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1454.320 -4.800 1455.440 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1484.000 -4.800 1485.120 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1513.680 -4.800 1514.800 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1543.360 -4.800 1544.480 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1573.600 -4.800 1574.720 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1603.280 -4.800 1604.400 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1632.960 -4.800 1634.080 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1096.480 -4.800 1097.600 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1662.640 -4.800 1663.760 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1692.880 -4.800 1694.000 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1722.560 -4.800 1723.680 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1752.240 -4.800 1753.360 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1781.920 -4.800 1783.040 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1811.600 -4.800 1812.720 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1841.840 -4.800 1842.960 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1871.520 -4.800 1872.640 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1901.200 -4.800 1902.320 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1930.880 -4.800 1932.000 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1126.160 -4.800 1127.280 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1961.120 -4.800 1962.240 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1990.800 -4.800 1991.920 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2020.480 -4.800 2021.600 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2050.160 -4.800 2051.280 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2080.400 -4.800 2081.520 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2110.080 -4.800 2111.200 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2139.760 -4.800 2140.880 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2169.440 -4.800 2170.560 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2199.120 -4.800 2200.240 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2229.360 -4.800 2230.480 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1156.400 -4.800 1157.520 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2259.040 -4.800 2260.160 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2288.720 -4.800 2289.840 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2318.400 -4.800 2319.520 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2348.640 -4.800 2349.760 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2378.320 -4.800 2379.440 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2408.000 -4.800 2409.120 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2437.680 -4.800 2438.800 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2467.360 -4.800 2468.480 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2497.600 -4.800 2498.720 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2527.280 -4.800 2528.400 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1186.080 -4.800 1187.200 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2556.960 -4.800 2558.080 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2586.640 -4.800 2587.760 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2616.880 -4.800 2618.000 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2646.560 -4.800 2647.680 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2676.240 -4.800 2677.360 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2705.920 -4.800 2707.040 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2735.600 -4.800 2736.720 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2765.840 -4.800 2766.960 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2795.520 -4.800 2796.640 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2825.200 -4.800 2826.320 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1215.760 -4.800 1216.880 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2854.880 -4.800 2856.000 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2885.120 -4.800 2886.240 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2914.800 -4.800 2915.920 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2944.480 -4.800 2945.600 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1245.440 -4.800 1246.560 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1275.120 -4.800 1276.240 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1305.360 -4.800 1306.480 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1335.040 -4.800 1336.160 2.400 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1076.880 -4.800 1078.000 2.400 ;
    END
  END la_oenb[0]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1374.800 -4.800 1375.920 2.400 ;
    END
  END la_oenb[10]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1404.480 -4.800 1405.600 2.400 ;
    END
  END la_oenb[11]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1434.160 -4.800 1435.280 2.400 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1464.400 -4.800 1465.520 2.400 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1494.080 -4.800 1495.200 2.400 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1523.760 -4.800 1524.880 2.400 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1553.440 -4.800 1554.560 2.400 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1583.120 -4.800 1584.240 2.400 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1613.360 -4.800 1614.480 2.400 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1643.040 -4.800 1644.160 2.400 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1106.560 -4.800 1107.680 2.400 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1672.720 -4.800 1673.840 2.400 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1702.400 -4.800 1703.520 2.400 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1732.640 -4.800 1733.760 2.400 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1762.320 -4.800 1763.440 2.400 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1792.000 -4.800 1793.120 2.400 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1821.680 -4.800 1822.800 2.400 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1851.360 -4.800 1852.480 2.400 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1881.600 -4.800 1882.720 2.400 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1911.280 -4.800 1912.400 2.400 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1940.960 -4.800 1942.080 2.400 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1136.240 -4.800 1137.360 2.400 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1970.640 -4.800 1971.760 2.400 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2000.880 -4.800 2002.000 2.400 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2030.560 -4.800 2031.680 2.400 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2060.240 -4.800 2061.360 2.400 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2089.920 -4.800 2091.040 2.400 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2119.600 -4.800 2120.720 2.400 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2149.840 -4.800 2150.960 2.400 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2179.520 -4.800 2180.640 2.400 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2209.200 -4.800 2210.320 2.400 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2238.880 -4.800 2240.000 2.400 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1165.920 -4.800 1167.040 2.400 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2269.120 -4.800 2270.240 2.400 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2298.800 -4.800 2299.920 2.400 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2328.480 -4.800 2329.600 2.400 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2358.160 -4.800 2359.280 2.400 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2388.400 -4.800 2389.520 2.400 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2418.080 -4.800 2419.200 2.400 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2447.760 -4.800 2448.880 2.400 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2477.440 -4.800 2478.560 2.400 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2507.120 -4.800 2508.240 2.400 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2537.360 -4.800 2538.480 2.400 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1196.160 -4.800 1197.280 2.400 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2567.040 -4.800 2568.160 2.400 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2596.720 -4.800 2597.840 2.400 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2626.400 -4.800 2627.520 2.400 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2656.640 -4.800 2657.760 2.400 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2686.320 -4.800 2687.440 2.400 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2716.000 -4.800 2717.120 2.400 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2745.680 -4.800 2746.800 2.400 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2775.360 -4.800 2776.480 2.400 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2805.600 -4.800 2806.720 2.400 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2835.280 -4.800 2836.400 2.400 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1225.840 -4.800 1226.960 2.400 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2864.960 -4.800 2866.080 2.400 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2894.640 -4.800 2895.760 2.400 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2924.880 -4.800 2926.000 2.400 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2954.560 -4.800 2955.680 2.400 ;
    END
  END la_oenb[63]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1255.520 -4.800 1256.640 2.400 ;
    END
  END la_oenb[6]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1285.200 -4.800 1286.320 2.400 ;
    END
  END la_oenb[7]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1314.880 -4.800 1316.000 2.400 ;
    END
  END la_oenb[8]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1345.120 -4.800 1346.240 2.400 ;
    END
  END la_oenb[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2964.640 -4.800 2965.760 2.400 ;
    END
  END user_clock2
  PIN user_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2974.160 -4.800 2975.280 2.400 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2984.240 -4.800 2985.360 2.400 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2994.320 -4.800 2995.440 2.400 ;
    END
  END user_irq[2]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT -10.380 -1.420 -7.280 3000.220 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -10.380 -1.420 3010.300 1.680 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -10.380 2997.120 3010.300 3000.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 3007.200 -1.420 3010.300 3000.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 10.170 -6.220 13.270 3005.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 190.170 -6.220 193.270 3005.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 370.170 -6.220 373.270 3005.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 550.170 -6.220 553.270 3005.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 730.170 -6.220 733.270 3005.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 910.170 -6.220 913.270 3005.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1090.170 -6.220 1093.270 3005.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1270.170 -6.220 1273.270 3005.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1450.170 -6.220 1453.270 3005.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1630.170 -6.220 1633.270 3005.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1810.170 -6.220 1813.270 3005.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1990.170 -6.220 1993.270 3005.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2170.170 -6.220 2173.270 3005.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2350.170 -6.220 2353.270 3005.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2530.170 -6.220 2533.270 3005.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2710.170 -6.220 2713.270 3005.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2890.170 -6.220 2893.270 3005.020 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -15.180 19.130 3015.100 22.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -15.180 199.130 3015.100 202.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -15.180 379.130 3015.100 382.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -15.180 559.130 3015.100 562.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -15.180 739.130 3015.100 742.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -15.180 919.130 3015.100 922.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -15.180 1099.130 3015.100 1102.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -15.180 1279.130 3015.100 1282.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -15.180 1459.130 3015.100 1462.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -15.180 1639.130 3015.100 1642.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -15.180 1819.130 3015.100 1822.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -15.180 1999.130 3015.100 2002.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -15.180 2179.130 3015.100 2182.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -15.180 2359.130 3015.100 2362.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -15.180 2539.130 3015.100 2542.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -15.180 2719.130 3015.100 2722.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -15.180 2899.130 3015.100 2902.230 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT -15.180 -6.220 -12.080 3005.020 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -15.180 -6.220 3015.100 -3.120 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -15.180 3001.920 3015.100 3005.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 3012.000 -6.220 3015.100 3005.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 100.170 -6.220 103.270 3005.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 280.170 -6.220 283.270 3005.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 460.170 -6.220 463.270 3005.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 640.170 -6.220 643.270 3005.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 820.170 -6.220 823.270 3005.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1000.170 -6.220 1003.270 3005.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1180.170 -6.220 1183.270 3005.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1360.170 -6.220 1363.270 3005.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1540.170 -6.220 1543.270 3005.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1720.170 -6.220 1723.270 3005.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1900.170 -6.220 1903.270 3005.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2080.170 -6.220 2083.270 3005.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2260.170 -6.220 2263.270 3005.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2440.170 -6.220 2443.270 3005.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2620.170 -6.220 2623.270 3005.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2800.170 -6.220 2803.270 3005.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2980.170 -6.220 2983.270 3005.020 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -15.180 109.130 3015.100 112.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -15.180 289.130 3015.100 292.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -15.180 469.130 3015.100 472.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -15.180 649.130 3015.100 652.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -15.180 829.130 3015.100 832.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -15.180 1009.130 3015.100 1012.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -15.180 1189.130 3015.100 1192.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -15.180 1369.130 3015.100 1372.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -15.180 1549.130 3015.100 1552.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -15.180 1729.130 3015.100 1732.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -15.180 1909.130 3015.100 1912.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -15.180 2089.130 3015.100 2092.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -15.180 2269.130 3015.100 2272.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -15.180 2449.130 3015.100 2452.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -15.180 2629.130 3015.100 2632.230 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -15.180 2809.130 3015.100 2812.230 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3.920 -4.800 5.040 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 13.440 -4.800 14.560 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 23.520 -4.800 24.640 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 63.280 -4.800 64.400 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 400.960 -4.800 402.080 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 430.640 -4.800 431.760 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 460.880 -4.800 462.000 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 490.560 -4.800 491.680 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 520.240 -4.800 521.360 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 549.920 -4.800 551.040 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 580.160 -4.800 581.280 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 609.840 -4.800 610.960 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 639.520 -4.800 640.640 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 669.200 -4.800 670.320 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 103.040 -4.800 104.160 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 698.880 -4.800 700.000 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 729.120 -4.800 730.240 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 758.800 -4.800 759.920 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 788.480 -4.800 789.600 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 818.160 -4.800 819.280 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 848.400 -4.800 849.520 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 878.080 -4.800 879.200 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 907.760 -4.800 908.880 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 937.440 -4.800 938.560 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 967.120 -4.800 968.240 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 142.800 -4.800 143.920 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 997.360 -4.800 998.480 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1027.040 -4.800 1028.160 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 182.560 -4.800 183.680 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 222.320 -4.800 223.440 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 252.000 -4.800 253.120 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 281.680 -4.800 282.800 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 311.360 -4.800 312.480 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 341.600 -4.800 342.720 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 371.280 -4.800 372.400 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 33.600 -4.800 34.720 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 73.360 -4.800 74.480 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 411.040 -4.800 412.160 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 440.720 -4.800 441.840 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 470.400 -4.800 471.520 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 500.640 -4.800 501.760 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 530.320 -4.800 531.440 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 560.000 -4.800 561.120 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 589.680 -4.800 590.800 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 619.360 -4.800 620.480 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 649.600 -4.800 650.720 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 679.280 -4.800 680.400 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 113.120 -4.800 114.240 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 708.960 -4.800 710.080 2.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 738.640 -4.800 739.760 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 768.880 -4.800 770.000 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 798.560 -4.800 799.680 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 828.240 -4.800 829.360 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 857.920 -4.800 859.040 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 888.160 -4.800 889.280 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 917.840 -4.800 918.960 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 947.520 -4.800 948.640 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 977.200 -4.800 978.320 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 152.880 -4.800 154.000 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1006.880 -4.800 1008.000 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1037.120 -4.800 1038.240 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 192.640 -4.800 193.760 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 232.400 -4.800 233.520 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 262.080 -4.800 263.200 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 291.760 -4.800 292.880 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 321.440 -4.800 322.560 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 351.120 -4.800 352.240 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 381.360 -4.800 382.480 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 82.880 -4.800 84.000 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 421.120 -4.800 422.240 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 450.800 -4.800 451.920 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 480.480 -4.800 481.600 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 510.160 -4.800 511.280 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 540.400 -4.800 541.520 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 570.080 -4.800 571.200 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 599.760 -4.800 600.880 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 629.440 -4.800 630.560 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 659.120 -4.800 660.240 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 689.360 -4.800 690.480 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 122.640 -4.800 123.760 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 719.040 -4.800 720.160 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 748.720 -4.800 749.840 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 778.400 -4.800 779.520 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 808.640 -4.800 809.760 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 838.320 -4.800 839.440 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 868.000 -4.800 869.120 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 897.680 -4.800 898.800 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 927.360 -4.800 928.480 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 957.600 -4.800 958.720 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 987.280 -4.800 988.400 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 162.400 -4.800 163.520 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1016.960 -4.800 1018.080 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1046.640 -4.800 1047.760 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 202.160 -4.800 203.280 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 241.920 -4.800 243.040 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 272.160 -4.800 273.280 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 301.840 -4.800 302.960 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 331.520 -4.800 332.640 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 361.200 -4.800 362.320 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 390.880 -4.800 392.000 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 92.960 -4.800 94.080 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 132.720 -4.800 133.840 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 172.480 -4.800 173.600 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 212.240 -4.800 213.360 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 43.120 -4.800 44.240 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 53.200 -4.800 54.320 2.400 ;
    END
  END wbs_we_i
  OBS
      LAYER Metal1 ;
        RECT 6.720 13.870 2995.070 2983.420 ;
      LAYER Metal2 ;
        RECT 8.260 2997.300 54.580 2998.380 ;
        RECT 56.300 2997.300 165.460 2998.380 ;
        RECT 167.180 2997.300 276.340 2998.380 ;
        RECT 278.060 2997.300 387.780 2998.380 ;
        RECT 389.500 2997.300 498.660 2998.380 ;
        RECT 500.380 2997.300 610.100 2998.380 ;
        RECT 611.820 2997.300 720.980 2998.380 ;
        RECT 722.700 2997.300 832.420 2998.380 ;
        RECT 834.140 2997.300 943.300 2998.380 ;
        RECT 945.020 2997.300 1054.740 2998.380 ;
        RECT 1056.460 2997.300 1165.620 2998.380 ;
        RECT 1167.340 2997.300 1276.500 2998.380 ;
        RECT 1278.220 2997.300 1387.940 2998.380 ;
        RECT 1389.660 2997.300 1498.820 2998.380 ;
        RECT 1500.540 2997.300 1610.260 2998.380 ;
        RECT 1611.980 2997.300 1721.140 2998.380 ;
        RECT 1722.860 2997.300 1832.580 2998.380 ;
        RECT 1834.300 2997.300 1943.460 2998.380 ;
        RECT 1945.180 2997.300 2054.900 2998.380 ;
        RECT 2056.620 2997.300 2165.780 2998.380 ;
        RECT 2167.500 2997.300 2276.660 2998.380 ;
        RECT 2278.380 2997.300 2388.100 2998.380 ;
        RECT 2389.820 2997.300 2498.980 2998.380 ;
        RECT 2500.700 2997.300 2610.420 2998.380 ;
        RECT 2612.140 2997.300 2721.300 2998.380 ;
        RECT 2723.020 2997.300 2832.740 2998.380 ;
        RECT 2834.460 2997.300 2943.620 2998.380 ;
        RECT 2945.340 2997.300 2995.020 2998.380 ;
        RECT 8.260 2.700 2995.020 2997.300 ;
        RECT 8.260 2.100 13.140 2.700 ;
        RECT 14.860 2.100 23.220 2.700 ;
        RECT 24.940 2.100 33.300 2.700 ;
        RECT 35.020 2.100 42.820 2.700 ;
        RECT 44.540 2.100 52.900 2.700 ;
        RECT 54.620 2.100 62.980 2.700 ;
        RECT 64.700 2.100 73.060 2.700 ;
        RECT 74.780 2.100 82.580 2.700 ;
        RECT 84.300 2.100 92.660 2.700 ;
        RECT 94.380 2.100 102.740 2.700 ;
        RECT 104.460 2.100 112.820 2.700 ;
        RECT 114.540 2.100 122.340 2.700 ;
        RECT 124.060 2.100 132.420 2.700 ;
        RECT 134.140 2.100 142.500 2.700 ;
        RECT 144.220 2.100 152.580 2.700 ;
        RECT 154.300 2.100 162.100 2.700 ;
        RECT 163.820 2.100 172.180 2.700 ;
        RECT 173.900 2.100 182.260 2.700 ;
        RECT 183.980 2.100 192.340 2.700 ;
        RECT 194.060 2.100 201.860 2.700 ;
        RECT 203.580 2.100 211.940 2.700 ;
        RECT 213.660 2.100 222.020 2.700 ;
        RECT 223.740 2.100 232.100 2.700 ;
        RECT 233.820 2.100 241.620 2.700 ;
        RECT 243.340 2.100 251.700 2.700 ;
        RECT 253.420 2.100 261.780 2.700 ;
        RECT 263.500 2.100 271.860 2.700 ;
        RECT 273.580 2.100 281.380 2.700 ;
        RECT 283.100 2.100 291.460 2.700 ;
        RECT 293.180 2.100 301.540 2.700 ;
        RECT 303.260 2.100 311.060 2.700 ;
        RECT 312.780 2.100 321.140 2.700 ;
        RECT 322.860 2.100 331.220 2.700 ;
        RECT 332.940 2.100 341.300 2.700 ;
        RECT 343.020 2.100 350.820 2.700 ;
        RECT 352.540 2.100 360.900 2.700 ;
        RECT 362.620 2.100 370.980 2.700 ;
        RECT 372.700 2.100 381.060 2.700 ;
        RECT 382.780 2.100 390.580 2.700 ;
        RECT 392.300 2.100 400.660 2.700 ;
        RECT 402.380 2.100 410.740 2.700 ;
        RECT 412.460 2.100 420.820 2.700 ;
        RECT 422.540 2.100 430.340 2.700 ;
        RECT 432.060 2.100 440.420 2.700 ;
        RECT 442.140 2.100 450.500 2.700 ;
        RECT 452.220 2.100 460.580 2.700 ;
        RECT 462.300 2.100 470.100 2.700 ;
        RECT 471.820 2.100 480.180 2.700 ;
        RECT 481.900 2.100 490.260 2.700 ;
        RECT 491.980 2.100 500.340 2.700 ;
        RECT 502.060 2.100 509.860 2.700 ;
        RECT 511.580 2.100 519.940 2.700 ;
        RECT 521.660 2.100 530.020 2.700 ;
        RECT 531.740 2.100 540.100 2.700 ;
        RECT 541.820 2.100 549.620 2.700 ;
        RECT 551.340 2.100 559.700 2.700 ;
        RECT 561.420 2.100 569.780 2.700 ;
        RECT 571.500 2.100 579.860 2.700 ;
        RECT 581.580 2.100 589.380 2.700 ;
        RECT 591.100 2.100 599.460 2.700 ;
        RECT 601.180 2.100 609.540 2.700 ;
        RECT 611.260 2.100 619.060 2.700 ;
        RECT 620.780 2.100 629.140 2.700 ;
        RECT 630.860 2.100 639.220 2.700 ;
        RECT 640.940 2.100 649.300 2.700 ;
        RECT 651.020 2.100 658.820 2.700 ;
        RECT 660.540 2.100 668.900 2.700 ;
        RECT 670.620 2.100 678.980 2.700 ;
        RECT 680.700 2.100 689.060 2.700 ;
        RECT 690.780 2.100 698.580 2.700 ;
        RECT 700.300 2.100 708.660 2.700 ;
        RECT 710.380 2.100 718.740 2.700 ;
        RECT 720.460 2.100 728.820 2.700 ;
        RECT 730.540 2.100 738.340 2.700 ;
        RECT 740.060 2.100 748.420 2.700 ;
        RECT 750.140 2.100 758.500 2.700 ;
        RECT 760.220 2.100 768.580 2.700 ;
        RECT 770.300 2.100 778.100 2.700 ;
        RECT 779.820 2.100 788.180 2.700 ;
        RECT 789.900 2.100 798.260 2.700 ;
        RECT 799.980 2.100 808.340 2.700 ;
        RECT 810.060 2.100 817.860 2.700 ;
        RECT 819.580 2.100 827.940 2.700 ;
        RECT 829.660 2.100 838.020 2.700 ;
        RECT 839.740 2.100 848.100 2.700 ;
        RECT 849.820 2.100 857.620 2.700 ;
        RECT 859.340 2.100 867.700 2.700 ;
        RECT 869.420 2.100 877.780 2.700 ;
        RECT 879.500 2.100 887.860 2.700 ;
        RECT 889.580 2.100 897.380 2.700 ;
        RECT 899.100 2.100 907.460 2.700 ;
        RECT 909.180 2.100 917.540 2.700 ;
        RECT 919.260 2.100 927.060 2.700 ;
        RECT 928.780 2.100 937.140 2.700 ;
        RECT 938.860 2.100 947.220 2.700 ;
        RECT 948.940 2.100 957.300 2.700 ;
        RECT 959.020 2.100 966.820 2.700 ;
        RECT 968.540 2.100 976.900 2.700 ;
        RECT 978.620 2.100 986.980 2.700 ;
        RECT 988.700 2.100 997.060 2.700 ;
        RECT 998.780 2.100 1006.580 2.700 ;
        RECT 1008.300 2.100 1016.660 2.700 ;
        RECT 1018.380 2.100 1026.740 2.700 ;
        RECT 1028.460 2.100 1036.820 2.700 ;
        RECT 1038.540 2.100 1046.340 2.700 ;
        RECT 1048.060 2.100 1056.420 2.700 ;
        RECT 1058.140 2.100 1066.500 2.700 ;
        RECT 1068.220 2.100 1076.580 2.700 ;
        RECT 1078.300 2.100 1086.100 2.700 ;
        RECT 1087.820 2.100 1096.180 2.700 ;
        RECT 1097.900 2.100 1106.260 2.700 ;
        RECT 1107.980 2.100 1116.340 2.700 ;
        RECT 1118.060 2.100 1125.860 2.700 ;
        RECT 1127.580 2.100 1135.940 2.700 ;
        RECT 1137.660 2.100 1146.020 2.700 ;
        RECT 1147.740 2.100 1156.100 2.700 ;
        RECT 1157.820 2.100 1165.620 2.700 ;
        RECT 1167.340 2.100 1175.700 2.700 ;
        RECT 1177.420 2.100 1185.780 2.700 ;
        RECT 1187.500 2.100 1195.860 2.700 ;
        RECT 1197.580 2.100 1205.380 2.700 ;
        RECT 1207.100 2.100 1215.460 2.700 ;
        RECT 1217.180 2.100 1225.540 2.700 ;
        RECT 1227.260 2.100 1235.060 2.700 ;
        RECT 1236.780 2.100 1245.140 2.700 ;
        RECT 1246.860 2.100 1255.220 2.700 ;
        RECT 1256.940 2.100 1265.300 2.700 ;
        RECT 1267.020 2.100 1274.820 2.700 ;
        RECT 1276.540 2.100 1284.900 2.700 ;
        RECT 1286.620 2.100 1294.980 2.700 ;
        RECT 1296.700 2.100 1305.060 2.700 ;
        RECT 1306.780 2.100 1314.580 2.700 ;
        RECT 1316.300 2.100 1324.660 2.700 ;
        RECT 1326.380 2.100 1334.740 2.700 ;
        RECT 1336.460 2.100 1344.820 2.700 ;
        RECT 1346.540 2.100 1354.340 2.700 ;
        RECT 1356.060 2.100 1364.420 2.700 ;
        RECT 1366.140 2.100 1374.500 2.700 ;
        RECT 1376.220 2.100 1384.580 2.700 ;
        RECT 1386.300 2.100 1394.100 2.700 ;
        RECT 1395.820 2.100 1404.180 2.700 ;
        RECT 1405.900 2.100 1414.260 2.700 ;
        RECT 1415.980 2.100 1424.340 2.700 ;
        RECT 1426.060 2.100 1433.860 2.700 ;
        RECT 1435.580 2.100 1443.940 2.700 ;
        RECT 1445.660 2.100 1454.020 2.700 ;
        RECT 1455.740 2.100 1464.100 2.700 ;
        RECT 1465.820 2.100 1473.620 2.700 ;
        RECT 1475.340 2.100 1483.700 2.700 ;
        RECT 1485.420 2.100 1493.780 2.700 ;
        RECT 1495.500 2.100 1503.860 2.700 ;
        RECT 1505.580 2.100 1513.380 2.700 ;
        RECT 1515.100 2.100 1523.460 2.700 ;
        RECT 1525.180 2.100 1533.540 2.700 ;
        RECT 1535.260 2.100 1543.060 2.700 ;
        RECT 1544.780 2.100 1553.140 2.700 ;
        RECT 1554.860 2.100 1563.220 2.700 ;
        RECT 1564.940 2.100 1573.300 2.700 ;
        RECT 1575.020 2.100 1582.820 2.700 ;
        RECT 1584.540 2.100 1592.900 2.700 ;
        RECT 1594.620 2.100 1602.980 2.700 ;
        RECT 1604.700 2.100 1613.060 2.700 ;
        RECT 1614.780 2.100 1622.580 2.700 ;
        RECT 1624.300 2.100 1632.660 2.700 ;
        RECT 1634.380 2.100 1642.740 2.700 ;
        RECT 1644.460 2.100 1652.820 2.700 ;
        RECT 1654.540 2.100 1662.340 2.700 ;
        RECT 1664.060 2.100 1672.420 2.700 ;
        RECT 1674.140 2.100 1682.500 2.700 ;
        RECT 1684.220 2.100 1692.580 2.700 ;
        RECT 1694.300 2.100 1702.100 2.700 ;
        RECT 1703.820 2.100 1712.180 2.700 ;
        RECT 1713.900 2.100 1722.260 2.700 ;
        RECT 1723.980 2.100 1732.340 2.700 ;
        RECT 1734.060 2.100 1741.860 2.700 ;
        RECT 1743.580 2.100 1751.940 2.700 ;
        RECT 1753.660 2.100 1762.020 2.700 ;
        RECT 1763.740 2.100 1772.100 2.700 ;
        RECT 1773.820 2.100 1781.620 2.700 ;
        RECT 1783.340 2.100 1791.700 2.700 ;
        RECT 1793.420 2.100 1801.780 2.700 ;
        RECT 1803.500 2.100 1811.300 2.700 ;
        RECT 1813.020 2.100 1821.380 2.700 ;
        RECT 1823.100 2.100 1831.460 2.700 ;
        RECT 1833.180 2.100 1841.540 2.700 ;
        RECT 1843.260 2.100 1851.060 2.700 ;
        RECT 1852.780 2.100 1861.140 2.700 ;
        RECT 1862.860 2.100 1871.220 2.700 ;
        RECT 1872.940 2.100 1881.300 2.700 ;
        RECT 1883.020 2.100 1890.820 2.700 ;
        RECT 1892.540 2.100 1900.900 2.700 ;
        RECT 1902.620 2.100 1910.980 2.700 ;
        RECT 1912.700 2.100 1921.060 2.700 ;
        RECT 1922.780 2.100 1930.580 2.700 ;
        RECT 1932.300 2.100 1940.660 2.700 ;
        RECT 1942.380 2.100 1950.740 2.700 ;
        RECT 1952.460 2.100 1960.820 2.700 ;
        RECT 1962.540 2.100 1970.340 2.700 ;
        RECT 1972.060 2.100 1980.420 2.700 ;
        RECT 1982.140 2.100 1990.500 2.700 ;
        RECT 1992.220 2.100 2000.580 2.700 ;
        RECT 2002.300 2.100 2010.100 2.700 ;
        RECT 2011.820 2.100 2020.180 2.700 ;
        RECT 2021.900 2.100 2030.260 2.700 ;
        RECT 2031.980 2.100 2040.340 2.700 ;
        RECT 2042.060 2.100 2049.860 2.700 ;
        RECT 2051.580 2.100 2059.940 2.700 ;
        RECT 2061.660 2.100 2070.020 2.700 ;
        RECT 2071.740 2.100 2080.100 2.700 ;
        RECT 2081.820 2.100 2089.620 2.700 ;
        RECT 2091.340 2.100 2099.700 2.700 ;
        RECT 2101.420 2.100 2109.780 2.700 ;
        RECT 2111.500 2.100 2119.300 2.700 ;
        RECT 2121.020 2.100 2129.380 2.700 ;
        RECT 2131.100 2.100 2139.460 2.700 ;
        RECT 2141.180 2.100 2149.540 2.700 ;
        RECT 2151.260 2.100 2159.060 2.700 ;
        RECT 2160.780 2.100 2169.140 2.700 ;
        RECT 2170.860 2.100 2179.220 2.700 ;
        RECT 2180.940 2.100 2189.300 2.700 ;
        RECT 2191.020 2.100 2198.820 2.700 ;
        RECT 2200.540 2.100 2208.900 2.700 ;
        RECT 2210.620 2.100 2218.980 2.700 ;
        RECT 2220.700 2.100 2229.060 2.700 ;
        RECT 2230.780 2.100 2238.580 2.700 ;
        RECT 2240.300 2.100 2248.660 2.700 ;
        RECT 2250.380 2.100 2258.740 2.700 ;
        RECT 2260.460 2.100 2268.820 2.700 ;
        RECT 2270.540 2.100 2278.340 2.700 ;
        RECT 2280.060 2.100 2288.420 2.700 ;
        RECT 2290.140 2.100 2298.500 2.700 ;
        RECT 2300.220 2.100 2308.580 2.700 ;
        RECT 2310.300 2.100 2318.100 2.700 ;
        RECT 2319.820 2.100 2328.180 2.700 ;
        RECT 2329.900 2.100 2338.260 2.700 ;
        RECT 2339.980 2.100 2348.340 2.700 ;
        RECT 2350.060 2.100 2357.860 2.700 ;
        RECT 2359.580 2.100 2367.940 2.700 ;
        RECT 2369.660 2.100 2378.020 2.700 ;
        RECT 2379.740 2.100 2388.100 2.700 ;
        RECT 2389.820 2.100 2397.620 2.700 ;
        RECT 2399.340 2.100 2407.700 2.700 ;
        RECT 2409.420 2.100 2417.780 2.700 ;
        RECT 2419.500 2.100 2427.300 2.700 ;
        RECT 2429.020 2.100 2437.380 2.700 ;
        RECT 2439.100 2.100 2447.460 2.700 ;
        RECT 2449.180 2.100 2457.540 2.700 ;
        RECT 2459.260 2.100 2467.060 2.700 ;
        RECT 2468.780 2.100 2477.140 2.700 ;
        RECT 2478.860 2.100 2487.220 2.700 ;
        RECT 2488.940 2.100 2497.300 2.700 ;
        RECT 2499.020 2.100 2506.820 2.700 ;
        RECT 2508.540 2.100 2516.900 2.700 ;
        RECT 2518.620 2.100 2526.980 2.700 ;
        RECT 2528.700 2.100 2537.060 2.700 ;
        RECT 2538.780 2.100 2546.580 2.700 ;
        RECT 2548.300 2.100 2556.660 2.700 ;
        RECT 2558.380 2.100 2566.740 2.700 ;
        RECT 2568.460 2.100 2576.820 2.700 ;
        RECT 2578.540 2.100 2586.340 2.700 ;
        RECT 2588.060 2.100 2596.420 2.700 ;
        RECT 2598.140 2.100 2606.500 2.700 ;
        RECT 2608.220 2.100 2616.580 2.700 ;
        RECT 2618.300 2.100 2626.100 2.700 ;
        RECT 2627.820 2.100 2636.180 2.700 ;
        RECT 2637.900 2.100 2646.260 2.700 ;
        RECT 2647.980 2.100 2656.340 2.700 ;
        RECT 2658.060 2.100 2665.860 2.700 ;
        RECT 2667.580 2.100 2675.940 2.700 ;
        RECT 2677.660 2.100 2686.020 2.700 ;
        RECT 2687.740 2.100 2696.100 2.700 ;
        RECT 2697.820 2.100 2705.620 2.700 ;
        RECT 2707.340 2.100 2715.700 2.700 ;
        RECT 2717.420 2.100 2725.780 2.700 ;
        RECT 2727.500 2.100 2735.300 2.700 ;
        RECT 2737.020 2.100 2745.380 2.700 ;
        RECT 2747.100 2.100 2755.460 2.700 ;
        RECT 2757.180 2.100 2765.540 2.700 ;
        RECT 2767.260 2.100 2775.060 2.700 ;
        RECT 2776.780 2.100 2785.140 2.700 ;
        RECT 2786.860 2.100 2795.220 2.700 ;
        RECT 2796.940 2.100 2805.300 2.700 ;
        RECT 2807.020 2.100 2814.820 2.700 ;
        RECT 2816.540 2.100 2824.900 2.700 ;
        RECT 2826.620 2.100 2834.980 2.700 ;
        RECT 2836.700 2.100 2845.060 2.700 ;
        RECT 2846.780 2.100 2854.580 2.700 ;
        RECT 2856.300 2.100 2864.660 2.700 ;
        RECT 2866.380 2.100 2874.740 2.700 ;
        RECT 2876.460 2.100 2884.820 2.700 ;
        RECT 2886.540 2.100 2894.340 2.700 ;
        RECT 2896.060 2.100 2904.420 2.700 ;
        RECT 2906.140 2.100 2914.500 2.700 ;
        RECT 2916.220 2.100 2924.580 2.700 ;
        RECT 2926.300 2.100 2934.100 2.700 ;
        RECT 2935.820 2.100 2944.180 2.700 ;
        RECT 2945.900 2.100 2954.260 2.700 ;
        RECT 2955.980 2.100 2964.340 2.700 ;
        RECT 2966.060 2.100 2973.860 2.700 ;
        RECT 2975.580 2.100 2983.940 2.700 ;
        RECT 2985.660 2.100 2994.020 2.700 ;
      LAYER Metal3 ;
        RECT 2.400 2967.180 2998.380 2981.580 ;
        RECT 2.400 2965.460 2997.300 2967.180 ;
        RECT 2.400 2964.940 2998.380 2965.460 ;
        RECT 2.700 2963.220 2998.380 2964.940 ;
        RECT 2.400 2900.540 2998.380 2963.220 ;
        RECT 2.400 2898.820 2997.300 2900.540 ;
        RECT 2.400 2893.260 2998.380 2898.820 ;
        RECT 2.700 2891.540 2998.380 2893.260 ;
        RECT 2.400 2833.900 2998.380 2891.540 ;
        RECT 2.400 2832.180 2997.300 2833.900 ;
        RECT 2.400 2822.140 2998.380 2832.180 ;
        RECT 2.700 2820.420 2998.380 2822.140 ;
        RECT 2.400 2767.260 2998.380 2820.420 ;
        RECT 2.400 2765.540 2997.300 2767.260 ;
        RECT 2.400 2750.460 2998.380 2765.540 ;
        RECT 2.700 2748.740 2998.380 2750.460 ;
        RECT 2.400 2700.620 2998.380 2748.740 ;
        RECT 2.400 2698.900 2997.300 2700.620 ;
        RECT 2.400 2679.340 2998.380 2698.900 ;
        RECT 2.700 2677.620 2998.380 2679.340 ;
        RECT 2.400 2633.980 2998.380 2677.620 ;
        RECT 2.400 2632.260 2997.300 2633.980 ;
        RECT 2.400 2607.660 2998.380 2632.260 ;
        RECT 2.700 2605.940 2998.380 2607.660 ;
        RECT 2.400 2567.340 2998.380 2605.940 ;
        RECT 2.400 2565.620 2997.300 2567.340 ;
        RECT 2.400 2536.540 2998.380 2565.620 ;
        RECT 2.700 2534.820 2998.380 2536.540 ;
        RECT 2.400 2500.700 2998.380 2534.820 ;
        RECT 2.400 2498.980 2997.300 2500.700 ;
        RECT 2.400 2464.860 2998.380 2498.980 ;
        RECT 2.700 2463.140 2998.380 2464.860 ;
        RECT 2.400 2434.060 2998.380 2463.140 ;
        RECT 2.400 2432.340 2997.300 2434.060 ;
        RECT 2.400 2393.740 2998.380 2432.340 ;
        RECT 2.700 2392.020 2998.380 2393.740 ;
        RECT 2.400 2367.420 2998.380 2392.020 ;
        RECT 2.400 2365.700 2997.300 2367.420 ;
        RECT 2.400 2322.060 2998.380 2365.700 ;
        RECT 2.700 2320.340 2998.380 2322.060 ;
        RECT 2.400 2300.780 2998.380 2320.340 ;
        RECT 2.400 2299.060 2997.300 2300.780 ;
        RECT 2.400 2250.380 2998.380 2299.060 ;
        RECT 2.700 2248.660 2998.380 2250.380 ;
        RECT 2.400 2234.140 2998.380 2248.660 ;
        RECT 2.400 2232.420 2997.300 2234.140 ;
        RECT 2.400 2179.260 2998.380 2232.420 ;
        RECT 2.700 2177.540 2998.380 2179.260 ;
        RECT 2.400 2167.500 2998.380 2177.540 ;
        RECT 2.400 2165.780 2997.300 2167.500 ;
        RECT 2.400 2107.580 2998.380 2165.780 ;
        RECT 2.700 2105.860 2998.380 2107.580 ;
        RECT 2.400 2100.860 2998.380 2105.860 ;
        RECT 2.400 2099.140 2997.300 2100.860 ;
        RECT 2.400 2036.460 2998.380 2099.140 ;
        RECT 2.700 2034.740 2998.380 2036.460 ;
        RECT 2.400 2034.220 2998.380 2034.740 ;
        RECT 2.400 2032.500 2997.300 2034.220 ;
        RECT 2.400 1967.580 2998.380 2032.500 ;
        RECT 2.400 1965.860 2997.300 1967.580 ;
        RECT 2.400 1964.780 2998.380 1965.860 ;
        RECT 2.700 1963.060 2998.380 1964.780 ;
        RECT 2.400 1900.940 2998.380 1963.060 ;
        RECT 2.400 1899.220 2997.300 1900.940 ;
        RECT 2.400 1893.660 2998.380 1899.220 ;
        RECT 2.700 1891.940 2998.380 1893.660 ;
        RECT 2.400 1834.300 2998.380 1891.940 ;
        RECT 2.400 1832.580 2997.300 1834.300 ;
        RECT 2.400 1821.980 2998.380 1832.580 ;
        RECT 2.700 1820.260 2998.380 1821.980 ;
        RECT 2.400 1767.660 2998.380 1820.260 ;
        RECT 2.400 1765.940 2997.300 1767.660 ;
        RECT 2.400 1750.860 2998.380 1765.940 ;
        RECT 2.700 1749.140 2998.380 1750.860 ;
        RECT 2.400 1701.020 2998.380 1749.140 ;
        RECT 2.400 1699.300 2997.300 1701.020 ;
        RECT 2.400 1679.180 2998.380 1699.300 ;
        RECT 2.700 1677.460 2998.380 1679.180 ;
        RECT 2.400 1634.380 2998.380 1677.460 ;
        RECT 2.400 1632.660 2997.300 1634.380 ;
        RECT 2.400 1608.060 2998.380 1632.660 ;
        RECT 2.700 1606.340 2998.380 1608.060 ;
        RECT 2.400 1567.740 2998.380 1606.340 ;
        RECT 2.400 1566.020 2997.300 1567.740 ;
        RECT 2.400 1536.380 2998.380 1566.020 ;
        RECT 2.700 1534.660 2998.380 1536.380 ;
        RECT 2.400 1500.540 2998.380 1534.660 ;
        RECT 2.400 1498.820 2997.300 1500.540 ;
        RECT 2.400 1464.700 2998.380 1498.820 ;
        RECT 2.700 1462.980 2998.380 1464.700 ;
        RECT 2.400 1433.900 2998.380 1462.980 ;
        RECT 2.400 1432.180 2997.300 1433.900 ;
        RECT 2.400 1393.580 2998.380 1432.180 ;
        RECT 2.700 1391.860 2998.380 1393.580 ;
        RECT 2.400 1367.260 2998.380 1391.860 ;
        RECT 2.400 1365.540 2997.300 1367.260 ;
        RECT 2.400 1321.900 2998.380 1365.540 ;
        RECT 2.700 1320.180 2998.380 1321.900 ;
        RECT 2.400 1300.620 2998.380 1320.180 ;
        RECT 2.400 1298.900 2997.300 1300.620 ;
        RECT 2.400 1250.780 2998.380 1298.900 ;
        RECT 2.700 1249.060 2998.380 1250.780 ;
        RECT 2.400 1233.980 2998.380 1249.060 ;
        RECT 2.400 1232.260 2997.300 1233.980 ;
        RECT 2.400 1179.100 2998.380 1232.260 ;
        RECT 2.700 1177.380 2998.380 1179.100 ;
        RECT 2.400 1167.340 2998.380 1177.380 ;
        RECT 2.400 1165.620 2997.300 1167.340 ;
        RECT 2.400 1107.980 2998.380 1165.620 ;
        RECT 2.700 1106.260 2998.380 1107.980 ;
        RECT 2.400 1100.700 2998.380 1106.260 ;
        RECT 2.400 1098.980 2997.300 1100.700 ;
        RECT 2.400 1036.300 2998.380 1098.980 ;
        RECT 2.700 1034.580 2998.380 1036.300 ;
        RECT 2.400 1034.060 2998.380 1034.580 ;
        RECT 2.400 1032.340 2997.300 1034.060 ;
        RECT 2.400 967.420 2998.380 1032.340 ;
        RECT 2.400 965.700 2997.300 967.420 ;
        RECT 2.400 965.180 2998.380 965.700 ;
        RECT 2.700 963.460 2998.380 965.180 ;
        RECT 2.400 900.780 2998.380 963.460 ;
        RECT 2.400 899.060 2997.300 900.780 ;
        RECT 2.400 893.500 2998.380 899.060 ;
        RECT 2.700 891.780 2998.380 893.500 ;
        RECT 2.400 834.140 2998.380 891.780 ;
        RECT 2.400 832.420 2997.300 834.140 ;
        RECT 2.400 822.380 2998.380 832.420 ;
        RECT 2.700 820.660 2998.380 822.380 ;
        RECT 2.400 767.500 2998.380 820.660 ;
        RECT 2.400 765.780 2997.300 767.500 ;
        RECT 2.400 750.700 2998.380 765.780 ;
        RECT 2.700 748.980 2998.380 750.700 ;
        RECT 2.400 700.860 2998.380 748.980 ;
        RECT 2.400 699.140 2997.300 700.860 ;
        RECT 2.400 679.020 2998.380 699.140 ;
        RECT 2.700 677.300 2998.380 679.020 ;
        RECT 2.400 634.220 2998.380 677.300 ;
        RECT 2.400 632.500 2997.300 634.220 ;
        RECT 2.400 607.900 2998.380 632.500 ;
        RECT 2.700 606.180 2998.380 607.900 ;
        RECT 2.400 567.580 2998.380 606.180 ;
        RECT 2.400 565.860 2997.300 567.580 ;
        RECT 2.400 536.220 2998.380 565.860 ;
        RECT 2.700 534.500 2998.380 536.220 ;
        RECT 2.400 500.940 2998.380 534.500 ;
        RECT 2.400 499.220 2997.300 500.940 ;
        RECT 2.400 465.100 2998.380 499.220 ;
        RECT 2.700 463.380 2998.380 465.100 ;
        RECT 2.400 434.300 2998.380 463.380 ;
        RECT 2.400 432.580 2997.300 434.300 ;
        RECT 2.400 393.420 2998.380 432.580 ;
        RECT 2.700 391.700 2998.380 393.420 ;
        RECT 2.400 367.660 2998.380 391.700 ;
        RECT 2.400 365.940 2997.300 367.660 ;
        RECT 2.400 322.300 2998.380 365.940 ;
        RECT 2.700 320.580 2998.380 322.300 ;
        RECT 2.400 301.020 2998.380 320.580 ;
        RECT 2.400 299.300 2997.300 301.020 ;
        RECT 2.400 250.620 2998.380 299.300 ;
        RECT 2.700 248.900 2998.380 250.620 ;
        RECT 2.400 234.380 2998.380 248.900 ;
        RECT 2.400 232.660 2997.300 234.380 ;
        RECT 2.400 179.500 2998.380 232.660 ;
        RECT 2.700 177.780 2998.380 179.500 ;
        RECT 2.400 167.740 2998.380 177.780 ;
        RECT 2.400 166.020 2997.300 167.740 ;
        RECT 2.400 107.820 2998.380 166.020 ;
        RECT 2.700 106.100 2998.380 107.820 ;
        RECT 2.400 101.100 2998.380 106.100 ;
        RECT 2.400 99.380 2997.300 101.100 ;
        RECT 2.400 36.700 2998.380 99.380 ;
        RECT 2.700 34.980 2998.380 36.700 ;
        RECT 2.400 34.460 2998.380 34.980 ;
        RECT 2.400 34.020 2997.300 34.460 ;
  END
END user_project_wrapper
END LIBRARY

