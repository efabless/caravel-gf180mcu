magic
tech gf180mcuC
magscale 1 10
timestamp 1670265379
<< metal1 >>
rect 1120 11786 13776 11820
rect 1120 11734 4254 11786
rect 4306 11734 4358 11786
rect 4410 11734 4462 11786
rect 4514 11734 7444 11786
rect 7496 11734 7548 11786
rect 7600 11734 7652 11786
rect 7704 11734 10634 11786
rect 10686 11734 10738 11786
rect 10790 11734 10842 11786
rect 10894 11734 13776 11786
rect 1120 11700 13776 11734
rect 2158 11506 2210 11518
rect 2158 11442 2210 11454
rect 7758 11282 7810 11294
rect 7758 11218 7810 11230
rect 12462 11282 12514 11294
rect 12462 11218 12514 11230
rect 1120 11002 13776 11036
rect 1120 10950 5849 11002
rect 5901 10950 5953 11002
rect 6005 10950 6057 11002
rect 6109 10950 9039 11002
rect 9091 10950 9143 11002
rect 9195 10950 9247 11002
rect 9299 10950 12229 11002
rect 12281 10950 12333 11002
rect 12385 10950 12437 11002
rect 12489 10950 13776 11002
rect 1120 10916 13776 10950
rect 6526 10834 6578 10846
rect 1922 10782 1934 10834
rect 1986 10782 1998 10834
rect 6526 10770 6578 10782
rect 11342 10834 11394 10846
rect 11342 10770 11394 10782
rect 3054 10722 3106 10734
rect 2370 10670 2382 10722
rect 2434 10670 2446 10722
rect 12002 10670 12014 10722
rect 12066 10670 12078 10722
rect 12562 10670 12574 10722
rect 12626 10670 12638 10722
rect 3054 10658 3106 10670
rect 12798 10610 12850 10622
rect 2482 10558 2494 10610
rect 2546 10558 2558 10610
rect 7298 10558 7310 10610
rect 7362 10558 7374 10610
rect 8194 10558 8206 10610
rect 8258 10558 8270 10610
rect 12798 10546 12850 10558
rect 6962 10446 6974 10498
rect 7026 10446 7038 10498
rect 7970 10446 7982 10498
rect 8034 10446 8046 10498
rect 13134 10386 13186 10398
rect 13794 10334 13806 10386
rect 13858 10383 13870 10386
rect 14802 10383 14814 10386
rect 13858 10337 14814 10383
rect 13858 10334 13870 10337
rect 14802 10334 14814 10337
rect 14866 10334 14878 10386
rect 13134 10322 13186 10334
rect 1120 10218 13776 10252
rect 1120 10166 4254 10218
rect 4306 10166 4358 10218
rect 4410 10166 4462 10218
rect 4514 10166 7444 10218
rect 7496 10166 7548 10218
rect 7600 10166 7652 10218
rect 7704 10166 10634 10218
rect 10686 10166 10738 10218
rect 10790 10166 10842 10218
rect 10894 10166 13776 10218
rect 1120 10132 13776 10166
rect 2494 9714 2546 9726
rect 2494 9650 2546 9662
rect 7982 9714 8034 9726
rect 7982 9650 8034 9662
rect 12126 9714 12178 9726
rect 12126 9650 12178 9662
rect 1120 9434 13776 9468
rect 1120 9382 5849 9434
rect 5901 9382 5953 9434
rect 6005 9382 6057 9434
rect 6109 9382 9039 9434
rect 9091 9382 9143 9434
rect 9195 9382 9247 9434
rect 9299 9382 12229 9434
rect 12281 9382 12333 9434
rect 12385 9382 12437 9434
rect 12489 9382 13776 9434
rect 1120 9348 13776 9382
rect 1120 8650 13776 8684
rect 1120 8598 4254 8650
rect 4306 8598 4358 8650
rect 4410 8598 4462 8650
rect 4514 8598 7444 8650
rect 7496 8598 7548 8650
rect 7600 8598 7652 8650
rect 7704 8598 10634 8650
rect 10686 8598 10738 8650
rect 10790 8598 10842 8650
rect 10894 8598 13776 8650
rect 1120 8564 13776 8598
rect 2158 8482 2210 8494
rect 2158 8418 2210 8430
rect 6974 8370 7026 8382
rect 6974 8306 7026 8318
rect 7310 8258 7362 8270
rect 7310 8194 7362 8206
rect 7522 8094 7534 8146
rect 7586 8094 7598 8146
rect 8082 8094 8094 8146
rect 8146 8094 8158 8146
rect 6302 8034 6354 8046
rect 6302 7970 6354 7982
rect 8654 8034 8706 8046
rect 8654 7970 8706 7982
rect 11342 8034 11394 8046
rect 11342 7970 11394 7982
rect 1120 7866 13776 7900
rect 1120 7814 5849 7866
rect 5901 7814 5953 7866
rect 6005 7814 6057 7866
rect 6109 7814 9039 7866
rect 9091 7814 9143 7866
rect 9195 7814 9247 7866
rect 9299 7814 12229 7866
rect 12281 7814 12333 7866
rect 12385 7814 12437 7866
rect 12489 7814 13776 7866
rect 1120 7780 13776 7814
rect 7086 7698 7138 7710
rect 7086 7634 7138 7646
rect 8542 7698 8594 7710
rect 8542 7634 8594 7646
rect 5854 7586 5906 7598
rect 5854 7522 5906 7534
rect 6526 7586 6578 7598
rect 6526 7522 6578 7534
rect 7870 7586 7922 7598
rect 7870 7522 7922 7534
rect 9662 7586 9714 7598
rect 9662 7522 9714 7534
rect 10546 7422 10558 7474
rect 10610 7422 10622 7474
rect 10994 7422 11006 7474
rect 11058 7422 11070 7474
rect 10994 7198 11006 7250
rect 11058 7198 11070 7250
rect 1120 7082 13776 7116
rect 1120 7030 4254 7082
rect 4306 7030 4358 7082
rect 4410 7030 4462 7082
rect 4514 7030 7444 7082
rect 7496 7030 7548 7082
rect 7600 7030 7652 7082
rect 7704 7030 10634 7082
rect 10686 7030 10738 7082
rect 10790 7030 10842 7082
rect 10894 7030 13776 7082
rect 1120 6996 13776 7030
rect 10110 6802 10162 6814
rect 8754 6750 8766 6802
rect 8818 6750 8830 6802
rect 10110 6738 10162 6750
rect 5854 6690 5906 6702
rect 5854 6626 5906 6638
rect 6414 6690 6466 6702
rect 6414 6626 6466 6638
rect 1120 6298 13776 6332
rect 1120 6246 5849 6298
rect 5901 6246 5953 6298
rect 6005 6246 6057 6298
rect 6109 6246 9039 6298
rect 9091 6246 9143 6298
rect 9195 6246 9247 6298
rect 9299 6246 12229 6298
rect 12281 6246 12333 6298
rect 12385 6246 12437 6298
rect 12489 6246 13776 6298
rect 1120 6212 13776 6246
rect 7298 5854 7310 5906
rect 7362 5854 7374 5906
rect 6962 5742 6974 5794
rect 7026 5742 7038 5794
rect 1120 5514 13776 5548
rect 1120 5462 4254 5514
rect 4306 5462 4358 5514
rect 4410 5462 4462 5514
rect 4514 5462 7444 5514
rect 7496 5462 7548 5514
rect 7600 5462 7652 5514
rect 7704 5462 10634 5514
rect 10686 5462 10738 5514
rect 10790 5462 10842 5514
rect 10894 5462 13776 5514
rect 1120 5428 13776 5462
rect 1120 4730 13776 4764
rect 1120 4678 5849 4730
rect 5901 4678 5953 4730
rect 6005 4678 6057 4730
rect 6109 4678 9039 4730
rect 9091 4678 9143 4730
rect 9195 4678 9247 4730
rect 9299 4678 12229 4730
rect 12281 4678 12333 4730
rect 12385 4678 12437 4730
rect 12489 4678 13776 4730
rect 1120 4644 13776 4678
rect 3390 4562 3442 4574
rect 3390 4498 3442 4510
rect 10894 4562 10946 4574
rect 10894 4498 10946 4510
rect 2270 4450 2322 4462
rect 2270 4386 2322 4398
rect 6526 4226 6578 4238
rect 6526 4162 6578 4174
rect 7646 4226 7698 4238
rect 7646 4162 7698 4174
rect 12686 4226 12738 4238
rect 12686 4162 12738 4174
rect 1120 3946 13776 3980
rect 1120 3894 4254 3946
rect 4306 3894 4358 3946
rect 4410 3894 4462 3946
rect 4514 3894 7444 3946
rect 7496 3894 7548 3946
rect 7600 3894 7652 3946
rect 7704 3894 10634 3946
rect 10686 3894 10738 3946
rect 10790 3894 10842 3946
rect 10894 3894 13776 3946
rect 1120 3860 13776 3894
rect 4286 3666 4338 3678
rect 2706 3614 2718 3666
rect 2770 3614 2782 3666
rect 4286 3602 4338 3614
rect 5406 3666 5458 3678
rect 5406 3602 5458 3614
rect 12574 3666 12626 3678
rect 12574 3602 12626 3614
rect 2818 3502 2830 3554
rect 2882 3502 2894 3554
rect 7858 3502 7870 3554
rect 7922 3502 7934 3554
rect 8418 3502 8430 3554
rect 8482 3502 8494 3554
rect 10770 3502 10782 3554
rect 10834 3502 10846 3554
rect 11106 3502 11118 3554
rect 11170 3502 11182 3554
rect 12002 3502 12014 3554
rect 12066 3502 12078 3554
rect 2270 3442 2322 3454
rect 2270 3378 2322 3390
rect 3614 3330 3666 3342
rect 3614 3266 3666 3278
rect 6078 3330 6130 3342
rect 6078 3266 6130 3278
rect 6862 3330 6914 3342
rect 6862 3266 6914 3278
rect 1120 3162 13776 3196
rect 1120 3110 5849 3162
rect 5901 3110 5953 3162
rect 6005 3110 6057 3162
rect 6109 3110 9039 3162
rect 9091 3110 9143 3162
rect 9195 3110 9247 3162
rect 9299 3110 12229 3162
rect 12281 3110 12333 3162
rect 12385 3110 12437 3162
rect 12489 3110 13776 3162
rect 1120 3076 13776 3110
rect 9550 2994 9602 3006
rect 9550 2930 9602 2942
rect 10334 2994 10386 3006
rect 10334 2930 10386 2942
rect 12574 2994 12626 3006
rect 12574 2930 12626 2942
rect 13022 2994 13074 3006
rect 13022 2930 13074 2942
rect 5842 2830 5854 2882
rect 5906 2830 5918 2882
rect 8418 2830 8430 2882
rect 8482 2830 8494 2882
rect 1810 2718 1822 2770
rect 1874 2718 1886 2770
rect 2146 2718 2158 2770
rect 2210 2718 2222 2770
rect 4610 2718 4622 2770
rect 4674 2718 4686 2770
rect 5058 2718 5070 2770
rect 5122 2718 5134 2770
rect 6850 2718 6862 2770
rect 6914 2718 6926 2770
rect 7858 2718 7870 2770
rect 7922 2718 7934 2770
rect 7186 2606 7198 2658
rect 7250 2606 7262 2658
rect 8082 2606 8094 2658
rect 8146 2606 8158 2658
rect 1120 2378 13776 2412
rect 1120 2326 4254 2378
rect 4306 2326 4358 2378
rect 4410 2326 4462 2378
rect 4514 2326 7444 2378
rect 7496 2326 7548 2378
rect 7600 2326 7652 2378
rect 7704 2326 10634 2378
rect 10686 2326 10738 2378
rect 10790 2326 10842 2378
rect 10894 2326 13776 2378
rect 1120 2292 13776 2326
rect 4062 2098 4114 2110
rect 4062 2034 4114 2046
rect 6862 2098 6914 2110
rect 6862 2034 6914 2046
rect 7982 2098 8034 2110
rect 7982 2034 8034 2046
rect 5630 1874 5682 1886
rect 5630 1810 5682 1822
rect 7422 1874 7474 1886
rect 7422 1810 7474 1822
rect 2158 1762 2210 1774
rect 2158 1698 2210 1710
rect 6302 1762 6354 1774
rect 6302 1698 6354 1710
rect 8654 1762 8706 1774
rect 8654 1698 8706 1710
rect 1120 1594 13776 1628
rect 1120 1542 5849 1594
rect 5901 1542 5953 1594
rect 6005 1542 6057 1594
rect 6109 1542 9039 1594
rect 9091 1542 9143 1594
rect 9195 1542 9247 1594
rect 9299 1542 12229 1594
rect 12281 1542 12333 1594
rect 12385 1542 12437 1594
rect 12489 1542 13776 1594
rect 1120 1508 13776 1542
<< via1 >>
rect 4254 11734 4306 11786
rect 4358 11734 4410 11786
rect 4462 11734 4514 11786
rect 7444 11734 7496 11786
rect 7548 11734 7600 11786
rect 7652 11734 7704 11786
rect 10634 11734 10686 11786
rect 10738 11734 10790 11786
rect 10842 11734 10894 11786
rect 2158 11454 2210 11506
rect 7758 11230 7810 11282
rect 12462 11230 12514 11282
rect 5849 10950 5901 11002
rect 5953 10950 6005 11002
rect 6057 10950 6109 11002
rect 9039 10950 9091 11002
rect 9143 10950 9195 11002
rect 9247 10950 9299 11002
rect 12229 10950 12281 11002
rect 12333 10950 12385 11002
rect 12437 10950 12489 11002
rect 1934 10782 1986 10834
rect 6526 10782 6578 10834
rect 11342 10782 11394 10834
rect 2382 10670 2434 10722
rect 3054 10670 3106 10722
rect 12014 10670 12066 10722
rect 12574 10670 12626 10722
rect 2494 10558 2546 10610
rect 7310 10558 7362 10610
rect 8206 10558 8258 10610
rect 12798 10558 12850 10610
rect 6974 10446 7026 10498
rect 7982 10446 8034 10498
rect 13134 10334 13186 10386
rect 13806 10334 13858 10386
rect 14814 10334 14866 10386
rect 4254 10166 4306 10218
rect 4358 10166 4410 10218
rect 4462 10166 4514 10218
rect 7444 10166 7496 10218
rect 7548 10166 7600 10218
rect 7652 10166 7704 10218
rect 10634 10166 10686 10218
rect 10738 10166 10790 10218
rect 10842 10166 10894 10218
rect 2494 9662 2546 9714
rect 7982 9662 8034 9714
rect 12126 9662 12178 9714
rect 5849 9382 5901 9434
rect 5953 9382 6005 9434
rect 6057 9382 6109 9434
rect 9039 9382 9091 9434
rect 9143 9382 9195 9434
rect 9247 9382 9299 9434
rect 12229 9382 12281 9434
rect 12333 9382 12385 9434
rect 12437 9382 12489 9434
rect 4254 8598 4306 8650
rect 4358 8598 4410 8650
rect 4462 8598 4514 8650
rect 7444 8598 7496 8650
rect 7548 8598 7600 8650
rect 7652 8598 7704 8650
rect 10634 8598 10686 8650
rect 10738 8598 10790 8650
rect 10842 8598 10894 8650
rect 2158 8430 2210 8482
rect 6974 8318 7026 8370
rect 7310 8206 7362 8258
rect 7534 8094 7586 8146
rect 8094 8094 8146 8146
rect 6302 7982 6354 8034
rect 8654 7982 8706 8034
rect 11342 7982 11394 8034
rect 5849 7814 5901 7866
rect 5953 7814 6005 7866
rect 6057 7814 6109 7866
rect 9039 7814 9091 7866
rect 9143 7814 9195 7866
rect 9247 7814 9299 7866
rect 12229 7814 12281 7866
rect 12333 7814 12385 7866
rect 12437 7814 12489 7866
rect 7086 7646 7138 7698
rect 8542 7646 8594 7698
rect 5854 7534 5906 7586
rect 6526 7534 6578 7586
rect 7870 7534 7922 7586
rect 9662 7534 9714 7586
rect 10558 7422 10610 7474
rect 11006 7422 11058 7474
rect 11006 7198 11058 7250
rect 4254 7030 4306 7082
rect 4358 7030 4410 7082
rect 4462 7030 4514 7082
rect 7444 7030 7496 7082
rect 7548 7030 7600 7082
rect 7652 7030 7704 7082
rect 10634 7030 10686 7082
rect 10738 7030 10790 7082
rect 10842 7030 10894 7082
rect 8766 6750 8818 6802
rect 10110 6750 10162 6802
rect 5854 6638 5906 6690
rect 6414 6638 6466 6690
rect 5849 6246 5901 6298
rect 5953 6246 6005 6298
rect 6057 6246 6109 6298
rect 9039 6246 9091 6298
rect 9143 6246 9195 6298
rect 9247 6246 9299 6298
rect 12229 6246 12281 6298
rect 12333 6246 12385 6298
rect 12437 6246 12489 6298
rect 7310 5854 7362 5906
rect 6974 5742 7026 5794
rect 4254 5462 4306 5514
rect 4358 5462 4410 5514
rect 4462 5462 4514 5514
rect 7444 5462 7496 5514
rect 7548 5462 7600 5514
rect 7652 5462 7704 5514
rect 10634 5462 10686 5514
rect 10738 5462 10790 5514
rect 10842 5462 10894 5514
rect 5849 4678 5901 4730
rect 5953 4678 6005 4730
rect 6057 4678 6109 4730
rect 9039 4678 9091 4730
rect 9143 4678 9195 4730
rect 9247 4678 9299 4730
rect 12229 4678 12281 4730
rect 12333 4678 12385 4730
rect 12437 4678 12489 4730
rect 3390 4510 3442 4562
rect 10894 4510 10946 4562
rect 2270 4398 2322 4450
rect 6526 4174 6578 4226
rect 7646 4174 7698 4226
rect 12686 4174 12738 4226
rect 4254 3894 4306 3946
rect 4358 3894 4410 3946
rect 4462 3894 4514 3946
rect 7444 3894 7496 3946
rect 7548 3894 7600 3946
rect 7652 3894 7704 3946
rect 10634 3894 10686 3946
rect 10738 3894 10790 3946
rect 10842 3894 10894 3946
rect 2718 3614 2770 3666
rect 4286 3614 4338 3666
rect 5406 3614 5458 3666
rect 12574 3614 12626 3666
rect 2830 3502 2882 3554
rect 7870 3502 7922 3554
rect 8430 3502 8482 3554
rect 10782 3502 10834 3554
rect 11118 3502 11170 3554
rect 12014 3502 12066 3554
rect 2270 3390 2322 3442
rect 3614 3278 3666 3330
rect 6078 3278 6130 3330
rect 6862 3278 6914 3330
rect 5849 3110 5901 3162
rect 5953 3110 6005 3162
rect 6057 3110 6109 3162
rect 9039 3110 9091 3162
rect 9143 3110 9195 3162
rect 9247 3110 9299 3162
rect 12229 3110 12281 3162
rect 12333 3110 12385 3162
rect 12437 3110 12489 3162
rect 9550 2942 9602 2994
rect 10334 2942 10386 2994
rect 12574 2942 12626 2994
rect 13022 2942 13074 2994
rect 5854 2830 5906 2882
rect 8430 2830 8482 2882
rect 1822 2718 1874 2770
rect 2158 2718 2210 2770
rect 4622 2718 4674 2770
rect 5070 2718 5122 2770
rect 6862 2718 6914 2770
rect 7870 2718 7922 2770
rect 7198 2606 7250 2658
rect 8094 2606 8146 2658
rect 4254 2326 4306 2378
rect 4358 2326 4410 2378
rect 4462 2326 4514 2378
rect 7444 2326 7496 2378
rect 7548 2326 7600 2378
rect 7652 2326 7704 2378
rect 10634 2326 10686 2378
rect 10738 2326 10790 2378
rect 10842 2326 10894 2378
rect 4062 2046 4114 2098
rect 6862 2046 6914 2098
rect 7982 2046 8034 2098
rect 5630 1822 5682 1874
rect 7422 1822 7474 1874
rect 2158 1710 2210 1762
rect 6302 1710 6354 1762
rect 8654 1710 8706 1762
rect 5849 1542 5901 1594
rect 5953 1542 6005 1594
rect 6057 1542 6109 1594
rect 9039 1542 9091 1594
rect 9143 1542 9195 1594
rect 9247 1542 9299 1594
rect 12229 1542 12281 1594
rect 12333 1542 12385 1594
rect 12437 1542 12489 1594
<< metal2 >>
rect 0 13200 112 14000
rect 252 13244 1092 13300
rect 28 10836 84 13200
rect 28 10770 84 10780
rect 252 8428 308 13244
rect 1036 13076 1092 13244
rect 1344 13200 1456 14000
rect 1820 13244 2436 13300
rect 1372 13076 1428 13200
rect 1036 13020 1428 13076
rect 28 8372 308 8428
rect 28 4116 84 8372
rect 1820 7700 1876 13244
rect 2380 13076 2436 13244
rect 2688 13200 2800 14000
rect 3388 13244 3780 13300
rect 2716 13076 2772 13200
rect 2380 13020 2772 13076
rect 2156 11508 2212 11518
rect 2156 11414 2212 11452
rect 1932 10836 1988 10846
rect 1932 10742 1988 10780
rect 2380 10722 2436 10734
rect 2380 10670 2382 10722
rect 2434 10670 2436 10722
rect 2380 10052 2436 10670
rect 2492 10724 2548 10734
rect 2492 10610 2548 10668
rect 3052 10724 3108 10734
rect 3052 10630 3108 10668
rect 2492 10558 2494 10610
rect 2546 10558 2548 10610
rect 2492 10546 2548 10558
rect 2380 9716 2436 9996
rect 2492 9716 2548 9726
rect 2380 9714 2548 9716
rect 2380 9662 2494 9714
rect 2546 9662 2548 9714
rect 2380 9660 2548 9662
rect 2492 9650 2548 9660
rect 2156 8820 2212 8830
rect 2156 8482 2212 8764
rect 2156 8430 2158 8482
rect 2210 8430 2212 8482
rect 2156 8418 2212 8430
rect 1820 7634 1876 7644
rect 3388 7588 3444 13244
rect 3724 13076 3780 13244
rect 4032 13200 4144 14000
rect 5376 13200 5488 14000
rect 6720 13200 6832 14000
rect 8064 13200 8176 14000
rect 9408 13200 9520 14000
rect 10752 13200 10864 14000
rect 12096 13200 12208 14000
rect 13440 13200 13552 14000
rect 14140 13244 14532 13300
rect 4060 13076 4116 13200
rect 3724 13020 4116 13076
rect 4732 12852 4788 12862
rect 4252 11788 4516 11798
rect 4308 11732 4356 11788
rect 4412 11732 4460 11788
rect 4252 11722 4516 11732
rect 3388 7522 3444 7532
rect 3500 10724 3556 10734
rect 3500 6132 3556 10668
rect 4252 10220 4516 10230
rect 4308 10164 4356 10220
rect 4412 10164 4460 10220
rect 4252 10154 4516 10164
rect 4252 8652 4516 8662
rect 4308 8596 4356 8652
rect 4412 8596 4460 8652
rect 4252 8586 4516 8596
rect 4252 7084 4516 7094
rect 4308 7028 4356 7084
rect 4412 7028 4460 7084
rect 4252 7018 4516 7028
rect 3500 6066 3556 6076
rect 4252 5516 4516 5526
rect 4308 5460 4356 5516
rect 4412 5460 4460 5516
rect 4252 5450 4516 5460
rect 3388 5012 3444 5022
rect 3388 4562 3444 4956
rect 4060 5012 4116 5022
rect 3388 4510 3390 4562
rect 3442 4510 3444 4562
rect 3388 4498 3444 4510
rect 3500 4788 3556 4798
rect 2268 4450 2324 4462
rect 2268 4398 2270 4450
rect 2322 4398 2324 4450
rect 28 4050 84 4060
rect 1820 4116 1876 4126
rect 1372 3780 1428 3790
rect 28 1764 84 1774
rect 28 800 84 1708
rect 1372 800 1428 3724
rect 1820 2770 1876 4060
rect 2268 4116 2324 4398
rect 2268 4050 2324 4060
rect 2716 3666 2772 3678
rect 2716 3614 2718 3666
rect 2770 3614 2772 3666
rect 2268 3444 2324 3454
rect 2268 3350 2324 3388
rect 2716 3332 2772 3614
rect 2828 3556 2884 3566
rect 2828 3462 2884 3500
rect 1820 2718 1822 2770
rect 1874 2718 1876 2770
rect 1820 2706 1876 2718
rect 2156 2770 2212 2782
rect 2156 2718 2158 2770
rect 2210 2718 2212 2770
rect 2156 1764 2212 2718
rect 2156 1670 2212 1708
rect 2716 800 2772 3276
rect 3500 2884 3556 4732
rect 4060 3780 4116 4956
rect 4252 3948 4516 3958
rect 4308 3892 4356 3948
rect 4412 3892 4460 3948
rect 4252 3882 4516 3892
rect 4060 3724 4340 3780
rect 4060 3556 4116 3724
rect 4284 3666 4340 3724
rect 4284 3614 4286 3666
rect 4338 3614 4340 3666
rect 4284 3602 4340 3614
rect 4060 3490 4116 3500
rect 3612 3332 3668 3342
rect 3612 3238 3668 3276
rect 4732 2996 4788 12796
rect 5404 10052 5460 13200
rect 5847 11004 6111 11014
rect 5903 10948 5951 11004
rect 6007 10948 6055 11004
rect 5847 10938 6111 10948
rect 6524 10836 6580 10846
rect 6524 10742 6580 10780
rect 6748 10500 6804 13200
rect 7442 11788 7706 11798
rect 7498 11732 7546 11788
rect 7602 11732 7650 11788
rect 7442 11722 7706 11732
rect 7308 11284 7364 11294
rect 7308 10836 7364 11228
rect 7756 11284 7812 11294
rect 7756 11190 7812 11228
rect 8092 10836 8148 13200
rect 9037 11004 9301 11014
rect 9093 10948 9141 11004
rect 9197 10948 9245 11004
rect 9037 10938 9301 10948
rect 7308 10610 7364 10780
rect 7308 10558 7310 10610
rect 7362 10558 7364 10610
rect 7308 10546 7364 10558
rect 7868 10780 8148 10836
rect 6748 10434 6804 10444
rect 6972 10498 7028 10510
rect 6972 10446 6974 10498
rect 7026 10446 7028 10498
rect 6972 10388 7028 10446
rect 6972 10322 7028 10332
rect 7196 10388 7252 10398
rect 5404 9986 5460 9996
rect 5847 9436 6111 9446
rect 5903 9380 5951 9436
rect 6007 9380 6055 9436
rect 5847 9370 6111 9380
rect 7196 8428 7252 10332
rect 7442 10220 7706 10230
rect 7498 10164 7546 10220
rect 7602 10164 7650 10220
rect 7442 10154 7706 10164
rect 7442 8652 7706 8662
rect 7498 8596 7546 8652
rect 7602 8596 7650 8652
rect 7442 8586 7706 8596
rect 6972 8372 7252 8428
rect 6972 8370 7028 8372
rect 6972 8318 6974 8370
rect 7026 8318 7028 8370
rect 6972 8306 7028 8318
rect 6300 8260 6356 8270
rect 6300 8034 6356 8204
rect 7308 8260 7364 8270
rect 7308 8166 7364 8204
rect 6300 7982 6302 8034
rect 6354 7982 6356 8034
rect 5847 7868 6111 7878
rect 5903 7812 5951 7868
rect 6007 7812 6055 7868
rect 5847 7802 6111 7812
rect 5852 7588 5908 7598
rect 4732 2930 4788 2940
rect 4956 7364 5012 7374
rect 3500 2818 3556 2828
rect 4620 2772 4676 2782
rect 4620 2678 4676 2716
rect 4252 2380 4516 2390
rect 4308 2324 4356 2380
rect 4412 2324 4460 2380
rect 4252 2314 4516 2324
rect 4060 2098 4116 2110
rect 4060 2046 4062 2098
rect 4114 2046 4116 2098
rect 4060 800 4116 2046
rect 4956 2100 5012 7308
rect 5852 6692 5908 7532
rect 6300 7364 6356 7982
rect 7532 8146 7588 8158
rect 7532 8094 7534 8146
rect 7586 8094 7588 8146
rect 7532 8036 7588 8094
rect 7084 7700 7140 7710
rect 7084 7606 7140 7644
rect 7532 7700 7588 7980
rect 7532 7634 7588 7644
rect 6300 7298 6356 7308
rect 6524 7586 6580 7598
rect 6524 7534 6526 7586
rect 6578 7534 6580 7586
rect 6524 7364 6580 7534
rect 6524 7298 6580 7308
rect 7868 7586 7924 10780
rect 8204 10610 8260 10622
rect 8204 10558 8206 10610
rect 8258 10558 8260 10610
rect 7980 10500 8036 10510
rect 7980 10406 8036 10444
rect 8204 10500 8260 10558
rect 7980 9716 8036 9726
rect 8204 9716 8260 10444
rect 9436 10052 9492 13200
rect 10780 11956 10836 13200
rect 10780 11900 11172 11956
rect 10632 11788 10896 11798
rect 10688 11732 10736 11788
rect 10792 11732 10840 11788
rect 10632 11722 10896 11732
rect 10632 10220 10896 10230
rect 10688 10164 10736 10220
rect 10792 10164 10840 10220
rect 10632 10154 10896 10164
rect 9436 9986 9492 9996
rect 7980 9714 8260 9716
rect 7980 9662 7982 9714
rect 8034 9662 8260 9714
rect 7980 9660 8260 9662
rect 7980 9650 8036 9660
rect 9037 9436 9301 9446
rect 9093 9380 9141 9436
rect 9197 9380 9245 9436
rect 9037 9370 9301 9380
rect 9548 8820 9604 8830
rect 8092 8146 8148 8158
rect 8092 8094 8094 8146
rect 8146 8094 8148 8146
rect 8092 7700 8148 8094
rect 8652 8036 8708 8046
rect 8652 7942 8708 7980
rect 9037 7868 9301 7878
rect 9093 7812 9141 7868
rect 9197 7812 9245 7868
rect 9037 7802 9301 7812
rect 8092 7634 8148 7644
rect 8540 7700 8596 7710
rect 8540 7606 8596 7644
rect 7868 7534 7870 7586
rect 7922 7534 7924 7586
rect 7442 7084 7706 7094
rect 7498 7028 7546 7084
rect 7602 7028 7650 7084
rect 7442 7018 7706 7028
rect 5852 6598 5908 6636
rect 6412 6692 6468 6702
rect 6412 6598 6468 6636
rect 5847 6300 6111 6310
rect 5903 6244 5951 6300
rect 6007 6244 6055 6300
rect 5847 6234 6111 6244
rect 7308 5908 7364 5918
rect 7868 5908 7924 7534
rect 8764 6804 8820 6814
rect 8764 6710 8820 6748
rect 9037 6300 9301 6310
rect 9093 6244 9141 6300
rect 9197 6244 9245 6300
rect 9037 6234 9301 6244
rect 7308 5906 7924 5908
rect 7308 5854 7310 5906
rect 7362 5854 7924 5906
rect 7308 5852 7924 5854
rect 7308 5842 7364 5852
rect 6972 5794 7028 5806
rect 6972 5742 6974 5794
rect 7026 5742 7028 5794
rect 5847 4732 6111 4742
rect 5903 4676 5951 4732
rect 6007 4676 6055 4732
rect 5847 4666 6111 4676
rect 6524 4226 6580 4238
rect 6524 4174 6526 4226
rect 6578 4174 6580 4226
rect 5404 4116 5460 4126
rect 5404 3666 5460 4060
rect 5404 3614 5406 3666
rect 5458 3614 5460 3666
rect 5404 3602 5460 3614
rect 5628 4116 5684 4126
rect 5516 3444 5572 3454
rect 5068 3332 5124 3342
rect 5068 2770 5124 3276
rect 5068 2718 5070 2770
rect 5122 2718 5124 2770
rect 5068 2706 5124 2718
rect 5516 2100 5572 3388
rect 4956 2034 5012 2044
rect 5404 2044 5572 2100
rect 5628 2772 5684 4060
rect 6524 4116 6580 4174
rect 6524 4050 6580 4060
rect 6300 3556 6356 3566
rect 6076 3332 6132 3370
rect 6076 3266 6132 3276
rect 5847 3164 6111 3174
rect 5903 3108 5951 3164
rect 6007 3108 6055 3164
rect 5847 3098 6111 3108
rect 5852 2884 5908 2894
rect 5852 2790 5908 2828
rect 4732 1652 4788 1662
rect 0 0 112 800
rect 1344 0 1456 800
rect 2688 0 2800 800
rect 4032 0 4144 800
rect 4732 756 4788 1596
rect 5404 800 5460 2044
rect 5628 1874 5684 2716
rect 5628 1822 5630 1874
rect 5682 1822 5684 1874
rect 5628 1810 5684 1822
rect 6300 1764 6356 3500
rect 6972 3444 7028 5742
rect 7442 5516 7706 5526
rect 7498 5460 7546 5516
rect 7602 5460 7650 5516
rect 7442 5450 7706 5460
rect 9037 4732 9301 4742
rect 9093 4676 9141 4732
rect 9197 4676 9245 4732
rect 9037 4666 9301 4676
rect 7644 4226 7700 4238
rect 7644 4174 7646 4226
rect 7698 4174 7700 4226
rect 7644 4116 7700 4174
rect 7644 4060 7924 4116
rect 7442 3948 7706 3958
rect 7498 3892 7546 3948
rect 7602 3892 7650 3948
rect 7442 3882 7706 3892
rect 7868 3556 7924 4060
rect 7868 3462 7924 3500
rect 8428 3556 8484 3566
rect 8428 3462 8484 3500
rect 9548 3556 9604 8764
rect 10632 8652 10896 8662
rect 10688 8596 10736 8652
rect 10792 8596 10840 8652
rect 10632 8586 10896 8596
rect 11004 8036 11060 8046
rect 9660 7586 9716 7598
rect 9660 7534 9662 7586
rect 9714 7534 9716 7586
rect 9660 7476 9716 7534
rect 9660 7410 9716 7420
rect 10556 7474 10612 7486
rect 10556 7422 10558 7474
rect 10610 7422 10612 7474
rect 10108 7364 10164 7374
rect 10108 6802 10164 7308
rect 10556 7364 10612 7422
rect 11004 7474 11060 7980
rect 11004 7422 11006 7474
rect 11058 7422 11060 7474
rect 11004 7410 11060 7422
rect 10556 7298 10612 7308
rect 11004 7250 11060 7262
rect 11004 7198 11006 7250
rect 11058 7198 11060 7250
rect 10632 7084 10896 7094
rect 10688 7028 10736 7084
rect 10792 7028 10840 7084
rect 10632 7018 10896 7028
rect 10108 6750 10110 6802
rect 10162 6750 10164 6802
rect 10108 6738 10164 6750
rect 9996 6132 10052 6142
rect 9996 5012 10052 6076
rect 10632 5516 10896 5526
rect 10688 5460 10736 5516
rect 10792 5460 10840 5516
rect 10632 5450 10896 5460
rect 9996 4946 10052 4956
rect 10892 4564 10948 4574
rect 10892 4470 10948 4508
rect 10632 3948 10896 3958
rect 10688 3892 10736 3948
rect 10792 3892 10840 3948
rect 10632 3882 10896 3892
rect 6972 3378 7028 3388
rect 6860 3330 6916 3342
rect 6860 3278 6862 3330
rect 6914 3278 6916 3330
rect 6860 2772 6916 3278
rect 6300 1670 6356 1708
rect 6748 2770 6916 2772
rect 6748 2718 6862 2770
rect 6914 2718 6916 2770
rect 6748 2716 6916 2718
rect 5847 1596 6111 1606
rect 5903 1540 5951 1596
rect 6007 1540 6055 1596
rect 5847 1530 6111 1540
rect 6748 800 6804 2716
rect 6860 2706 6916 2716
rect 6972 3220 7028 3230
rect 6860 2100 6916 2110
rect 6972 2100 7028 3164
rect 9037 3164 9301 3174
rect 9093 3108 9141 3164
rect 9197 3108 9245 3164
rect 9037 3098 9301 3108
rect 7868 2996 7924 3006
rect 7868 2772 7924 2940
rect 9548 2994 9604 3500
rect 9548 2942 9550 2994
rect 9602 2942 9604 2994
rect 9548 2930 9604 2942
rect 10332 3780 10388 3790
rect 10332 3556 10388 3724
rect 10332 2994 10388 3500
rect 10780 3780 10836 3790
rect 10780 3554 10836 3724
rect 10780 3502 10782 3554
rect 10834 3502 10836 3554
rect 10780 3490 10836 3502
rect 10332 2942 10334 2994
rect 10386 2942 10388 2994
rect 10332 2930 10388 2942
rect 8428 2882 8484 2894
rect 8428 2830 8430 2882
rect 8482 2830 8484 2882
rect 7868 2770 8036 2772
rect 7868 2718 7870 2770
rect 7922 2718 8036 2770
rect 7868 2716 8036 2718
rect 7868 2706 7924 2716
rect 7196 2658 7252 2670
rect 7196 2606 7198 2658
rect 7250 2606 7252 2658
rect 7196 2548 7252 2606
rect 7196 2482 7252 2492
rect 7442 2380 7706 2390
rect 7498 2324 7546 2380
rect 7602 2324 7650 2380
rect 7442 2314 7706 2324
rect 6860 2098 7028 2100
rect 6860 2046 6862 2098
rect 6914 2046 7028 2098
rect 6860 2044 7028 2046
rect 7980 2098 8036 2716
rect 7980 2046 7982 2098
rect 8034 2046 8036 2098
rect 6860 2034 6916 2044
rect 7420 1876 7476 1886
rect 7420 1782 7476 1820
rect 7980 1876 8036 2046
rect 7980 1810 8036 1820
rect 8092 2658 8148 2670
rect 8092 2606 8094 2658
rect 8146 2606 8148 2658
rect 8092 800 8148 2606
rect 8428 1764 8484 2830
rect 10632 2380 10896 2390
rect 10688 2324 10736 2380
rect 10792 2324 10840 2380
rect 10632 2314 10896 2324
rect 11004 2212 11060 7198
rect 11116 4564 11172 11900
rect 11228 11508 11284 11518
rect 11228 10500 11284 11452
rect 11340 11172 11396 11182
rect 11340 10834 11396 11116
rect 12124 11172 12180 13200
rect 12460 12852 12516 12862
rect 12460 11284 12516 12796
rect 12460 11282 12628 11284
rect 12460 11230 12462 11282
rect 12514 11230 12628 11282
rect 12460 11228 12628 11230
rect 12460 11218 12516 11228
rect 12124 11106 12180 11116
rect 12227 11004 12491 11014
rect 12283 10948 12331 11004
rect 12387 10948 12435 11004
rect 12227 10938 12491 10948
rect 11340 10782 11342 10834
rect 11394 10782 11396 10834
rect 11340 10770 11396 10782
rect 11900 10836 11956 10846
rect 11228 10434 11284 10444
rect 11340 8036 11396 8046
rect 11340 7942 11396 7980
rect 11900 8036 11956 10780
rect 12012 10722 12068 10734
rect 12012 10670 12014 10722
rect 12066 10670 12068 10722
rect 12012 10052 12068 10670
rect 12572 10722 12628 11228
rect 12572 10670 12574 10722
rect 12626 10670 12628 10722
rect 12572 10658 12628 10670
rect 12796 11172 12852 11182
rect 12796 10610 12852 11116
rect 13468 10836 13524 13200
rect 14140 11284 14196 13244
rect 14476 13076 14532 13244
rect 14784 13200 14896 14000
rect 14812 13076 14868 13200
rect 14476 13020 14868 13076
rect 14140 11218 14196 11228
rect 13468 10770 13524 10780
rect 12796 10558 12798 10610
rect 12850 10558 12852 10610
rect 12796 10546 12852 10558
rect 13132 10388 13188 10398
rect 13804 10388 13860 10398
rect 13132 10386 13860 10388
rect 13132 10334 13134 10386
rect 13186 10334 13806 10386
rect 13858 10334 13860 10386
rect 13132 10332 13860 10334
rect 13132 10322 13188 10332
rect 13804 10322 13860 10332
rect 14812 10386 14868 10398
rect 14812 10334 14814 10386
rect 14866 10334 14868 10386
rect 12012 9716 12068 9996
rect 12124 9716 12180 9726
rect 12012 9714 12180 9716
rect 12012 9662 12126 9714
rect 12178 9662 12180 9714
rect 12012 9660 12180 9662
rect 12124 9650 12180 9660
rect 12227 9436 12491 9446
rect 12283 9380 12331 9436
rect 12387 9380 12435 9436
rect 12227 9370 12491 9380
rect 11900 7970 11956 7980
rect 12227 7868 12491 7878
rect 12283 7812 12331 7868
rect 12387 7812 12435 7868
rect 12227 7802 12491 7812
rect 12796 6804 12852 6814
rect 12227 6300 12491 6310
rect 12283 6244 12331 6300
rect 12387 6244 12435 6300
rect 12227 6234 12491 6244
rect 12684 4788 12740 4798
rect 12227 4732 12491 4742
rect 12283 4676 12331 4732
rect 12387 4676 12435 4732
rect 12227 4666 12491 4676
rect 11116 3780 11172 4508
rect 12684 4226 12740 4732
rect 12684 4174 12686 4226
rect 12738 4174 12740 4226
rect 12684 4162 12740 4174
rect 11116 3714 11172 3724
rect 11900 4116 11956 4126
rect 11116 3556 11172 3566
rect 11116 2996 11172 3500
rect 11116 2930 11172 2940
rect 10780 2156 11060 2212
rect 8652 1764 8708 1774
rect 8428 1708 8652 1764
rect 8652 1670 8708 1708
rect 9436 1764 9492 1774
rect 9037 1596 9301 1606
rect 9093 1540 9141 1596
rect 9197 1540 9245 1596
rect 9037 1530 9301 1540
rect 9436 800 9492 1708
rect 10780 800 10836 2156
rect 11900 1428 11956 4060
rect 12684 3780 12740 3790
rect 12572 3668 12628 3678
rect 12572 3574 12628 3612
rect 12012 3556 12068 3566
rect 12012 3462 12068 3500
rect 12227 3164 12491 3174
rect 12283 3108 12331 3164
rect 12387 3108 12435 3164
rect 12227 3098 12491 3108
rect 12572 2996 12628 3006
rect 12684 2996 12740 3724
rect 12572 2994 12740 2996
rect 12572 2942 12574 2994
rect 12626 2942 12740 2994
rect 12572 2940 12740 2942
rect 12572 2930 12628 2940
rect 12227 1596 12491 1606
rect 12283 1540 12331 1596
rect 12387 1540 12435 1596
rect 12227 1530 12491 1540
rect 11900 1372 12180 1428
rect 12124 800 12180 1372
rect 4732 690 4788 700
rect 5376 0 5488 800
rect 6720 0 6832 800
rect 8064 0 8176 800
rect 9408 0 9520 800
rect 10752 0 10864 800
rect 12096 0 12208 800
rect 12796 756 12852 6748
rect 13468 3556 13524 3566
rect 13020 2996 13076 3006
rect 13020 2902 13076 2940
rect 13468 800 13524 3500
rect 14812 800 14868 10334
rect 12796 690 12852 700
rect 13440 0 13552 800
rect 14784 0 14896 800
<< via2 >>
rect 28 10780 84 10836
rect 2156 11506 2212 11508
rect 2156 11454 2158 11506
rect 2158 11454 2210 11506
rect 2210 11454 2212 11506
rect 2156 11452 2212 11454
rect 1932 10834 1988 10836
rect 1932 10782 1934 10834
rect 1934 10782 1986 10834
rect 1986 10782 1988 10834
rect 1932 10780 1988 10782
rect 2492 10668 2548 10724
rect 3052 10722 3108 10724
rect 3052 10670 3054 10722
rect 3054 10670 3106 10722
rect 3106 10670 3108 10722
rect 3052 10668 3108 10670
rect 2380 9996 2436 10052
rect 2156 8764 2212 8820
rect 1820 7644 1876 7700
rect 4732 12796 4788 12852
rect 4252 11786 4308 11788
rect 4252 11734 4254 11786
rect 4254 11734 4306 11786
rect 4306 11734 4308 11786
rect 4252 11732 4308 11734
rect 4356 11786 4412 11788
rect 4356 11734 4358 11786
rect 4358 11734 4410 11786
rect 4410 11734 4412 11786
rect 4356 11732 4412 11734
rect 4460 11786 4516 11788
rect 4460 11734 4462 11786
rect 4462 11734 4514 11786
rect 4514 11734 4516 11786
rect 4460 11732 4516 11734
rect 3388 7532 3444 7588
rect 3500 10668 3556 10724
rect 4252 10218 4308 10220
rect 4252 10166 4254 10218
rect 4254 10166 4306 10218
rect 4306 10166 4308 10218
rect 4252 10164 4308 10166
rect 4356 10218 4412 10220
rect 4356 10166 4358 10218
rect 4358 10166 4410 10218
rect 4410 10166 4412 10218
rect 4356 10164 4412 10166
rect 4460 10218 4516 10220
rect 4460 10166 4462 10218
rect 4462 10166 4514 10218
rect 4514 10166 4516 10218
rect 4460 10164 4516 10166
rect 4252 8650 4308 8652
rect 4252 8598 4254 8650
rect 4254 8598 4306 8650
rect 4306 8598 4308 8650
rect 4252 8596 4308 8598
rect 4356 8650 4412 8652
rect 4356 8598 4358 8650
rect 4358 8598 4410 8650
rect 4410 8598 4412 8650
rect 4356 8596 4412 8598
rect 4460 8650 4516 8652
rect 4460 8598 4462 8650
rect 4462 8598 4514 8650
rect 4514 8598 4516 8650
rect 4460 8596 4516 8598
rect 4252 7082 4308 7084
rect 4252 7030 4254 7082
rect 4254 7030 4306 7082
rect 4306 7030 4308 7082
rect 4252 7028 4308 7030
rect 4356 7082 4412 7084
rect 4356 7030 4358 7082
rect 4358 7030 4410 7082
rect 4410 7030 4412 7082
rect 4356 7028 4412 7030
rect 4460 7082 4516 7084
rect 4460 7030 4462 7082
rect 4462 7030 4514 7082
rect 4514 7030 4516 7082
rect 4460 7028 4516 7030
rect 3500 6076 3556 6132
rect 4252 5514 4308 5516
rect 4252 5462 4254 5514
rect 4254 5462 4306 5514
rect 4306 5462 4308 5514
rect 4252 5460 4308 5462
rect 4356 5514 4412 5516
rect 4356 5462 4358 5514
rect 4358 5462 4410 5514
rect 4410 5462 4412 5514
rect 4356 5460 4412 5462
rect 4460 5514 4516 5516
rect 4460 5462 4462 5514
rect 4462 5462 4514 5514
rect 4514 5462 4516 5514
rect 4460 5460 4516 5462
rect 3388 4956 3444 5012
rect 4060 4956 4116 5012
rect 3500 4732 3556 4788
rect 28 4060 84 4116
rect 1820 4060 1876 4116
rect 1372 3724 1428 3780
rect 28 1708 84 1764
rect 2268 4060 2324 4116
rect 2268 3442 2324 3444
rect 2268 3390 2270 3442
rect 2270 3390 2322 3442
rect 2322 3390 2324 3442
rect 2268 3388 2324 3390
rect 2828 3554 2884 3556
rect 2828 3502 2830 3554
rect 2830 3502 2882 3554
rect 2882 3502 2884 3554
rect 2828 3500 2884 3502
rect 2716 3276 2772 3332
rect 2156 1762 2212 1764
rect 2156 1710 2158 1762
rect 2158 1710 2210 1762
rect 2210 1710 2212 1762
rect 2156 1708 2212 1710
rect 4252 3946 4308 3948
rect 4252 3894 4254 3946
rect 4254 3894 4306 3946
rect 4306 3894 4308 3946
rect 4252 3892 4308 3894
rect 4356 3946 4412 3948
rect 4356 3894 4358 3946
rect 4358 3894 4410 3946
rect 4410 3894 4412 3946
rect 4356 3892 4412 3894
rect 4460 3946 4516 3948
rect 4460 3894 4462 3946
rect 4462 3894 4514 3946
rect 4514 3894 4516 3946
rect 4460 3892 4516 3894
rect 4060 3500 4116 3556
rect 3612 3330 3668 3332
rect 3612 3278 3614 3330
rect 3614 3278 3666 3330
rect 3666 3278 3668 3330
rect 3612 3276 3668 3278
rect 5847 11002 5903 11004
rect 5847 10950 5849 11002
rect 5849 10950 5901 11002
rect 5901 10950 5903 11002
rect 5847 10948 5903 10950
rect 5951 11002 6007 11004
rect 5951 10950 5953 11002
rect 5953 10950 6005 11002
rect 6005 10950 6007 11002
rect 5951 10948 6007 10950
rect 6055 11002 6111 11004
rect 6055 10950 6057 11002
rect 6057 10950 6109 11002
rect 6109 10950 6111 11002
rect 6055 10948 6111 10950
rect 6524 10834 6580 10836
rect 6524 10782 6526 10834
rect 6526 10782 6578 10834
rect 6578 10782 6580 10834
rect 6524 10780 6580 10782
rect 7442 11786 7498 11788
rect 7442 11734 7444 11786
rect 7444 11734 7496 11786
rect 7496 11734 7498 11786
rect 7442 11732 7498 11734
rect 7546 11786 7602 11788
rect 7546 11734 7548 11786
rect 7548 11734 7600 11786
rect 7600 11734 7602 11786
rect 7546 11732 7602 11734
rect 7650 11786 7706 11788
rect 7650 11734 7652 11786
rect 7652 11734 7704 11786
rect 7704 11734 7706 11786
rect 7650 11732 7706 11734
rect 7308 11228 7364 11284
rect 7756 11282 7812 11284
rect 7756 11230 7758 11282
rect 7758 11230 7810 11282
rect 7810 11230 7812 11282
rect 7756 11228 7812 11230
rect 9037 11002 9093 11004
rect 9037 10950 9039 11002
rect 9039 10950 9091 11002
rect 9091 10950 9093 11002
rect 9037 10948 9093 10950
rect 9141 11002 9197 11004
rect 9141 10950 9143 11002
rect 9143 10950 9195 11002
rect 9195 10950 9197 11002
rect 9141 10948 9197 10950
rect 9245 11002 9301 11004
rect 9245 10950 9247 11002
rect 9247 10950 9299 11002
rect 9299 10950 9301 11002
rect 9245 10948 9301 10950
rect 7308 10780 7364 10836
rect 6748 10444 6804 10500
rect 6972 10332 7028 10388
rect 7196 10332 7252 10388
rect 5404 9996 5460 10052
rect 5847 9434 5903 9436
rect 5847 9382 5849 9434
rect 5849 9382 5901 9434
rect 5901 9382 5903 9434
rect 5847 9380 5903 9382
rect 5951 9434 6007 9436
rect 5951 9382 5953 9434
rect 5953 9382 6005 9434
rect 6005 9382 6007 9434
rect 5951 9380 6007 9382
rect 6055 9434 6111 9436
rect 6055 9382 6057 9434
rect 6057 9382 6109 9434
rect 6109 9382 6111 9434
rect 6055 9380 6111 9382
rect 7442 10218 7498 10220
rect 7442 10166 7444 10218
rect 7444 10166 7496 10218
rect 7496 10166 7498 10218
rect 7442 10164 7498 10166
rect 7546 10218 7602 10220
rect 7546 10166 7548 10218
rect 7548 10166 7600 10218
rect 7600 10166 7602 10218
rect 7546 10164 7602 10166
rect 7650 10218 7706 10220
rect 7650 10166 7652 10218
rect 7652 10166 7704 10218
rect 7704 10166 7706 10218
rect 7650 10164 7706 10166
rect 7442 8650 7498 8652
rect 7442 8598 7444 8650
rect 7444 8598 7496 8650
rect 7496 8598 7498 8650
rect 7442 8596 7498 8598
rect 7546 8650 7602 8652
rect 7546 8598 7548 8650
rect 7548 8598 7600 8650
rect 7600 8598 7602 8650
rect 7546 8596 7602 8598
rect 7650 8650 7706 8652
rect 7650 8598 7652 8650
rect 7652 8598 7704 8650
rect 7704 8598 7706 8650
rect 7650 8596 7706 8598
rect 6300 8204 6356 8260
rect 7308 8258 7364 8260
rect 7308 8206 7310 8258
rect 7310 8206 7362 8258
rect 7362 8206 7364 8258
rect 7308 8204 7364 8206
rect 5847 7866 5903 7868
rect 5847 7814 5849 7866
rect 5849 7814 5901 7866
rect 5901 7814 5903 7866
rect 5847 7812 5903 7814
rect 5951 7866 6007 7868
rect 5951 7814 5953 7866
rect 5953 7814 6005 7866
rect 6005 7814 6007 7866
rect 5951 7812 6007 7814
rect 6055 7866 6111 7868
rect 6055 7814 6057 7866
rect 6057 7814 6109 7866
rect 6109 7814 6111 7866
rect 6055 7812 6111 7814
rect 5852 7586 5908 7588
rect 5852 7534 5854 7586
rect 5854 7534 5906 7586
rect 5906 7534 5908 7586
rect 5852 7532 5908 7534
rect 4732 2940 4788 2996
rect 4956 7308 5012 7364
rect 3500 2828 3556 2884
rect 4620 2770 4676 2772
rect 4620 2718 4622 2770
rect 4622 2718 4674 2770
rect 4674 2718 4676 2770
rect 4620 2716 4676 2718
rect 4252 2378 4308 2380
rect 4252 2326 4254 2378
rect 4254 2326 4306 2378
rect 4306 2326 4308 2378
rect 4252 2324 4308 2326
rect 4356 2378 4412 2380
rect 4356 2326 4358 2378
rect 4358 2326 4410 2378
rect 4410 2326 4412 2378
rect 4356 2324 4412 2326
rect 4460 2378 4516 2380
rect 4460 2326 4462 2378
rect 4462 2326 4514 2378
rect 4514 2326 4516 2378
rect 4460 2324 4516 2326
rect 7532 7980 7588 8036
rect 7084 7698 7140 7700
rect 7084 7646 7086 7698
rect 7086 7646 7138 7698
rect 7138 7646 7140 7698
rect 7084 7644 7140 7646
rect 7532 7644 7588 7700
rect 6300 7308 6356 7364
rect 6524 7308 6580 7364
rect 7980 10498 8036 10500
rect 7980 10446 7982 10498
rect 7982 10446 8034 10498
rect 8034 10446 8036 10498
rect 7980 10444 8036 10446
rect 8204 10444 8260 10500
rect 10632 11786 10688 11788
rect 10632 11734 10634 11786
rect 10634 11734 10686 11786
rect 10686 11734 10688 11786
rect 10632 11732 10688 11734
rect 10736 11786 10792 11788
rect 10736 11734 10738 11786
rect 10738 11734 10790 11786
rect 10790 11734 10792 11786
rect 10736 11732 10792 11734
rect 10840 11786 10896 11788
rect 10840 11734 10842 11786
rect 10842 11734 10894 11786
rect 10894 11734 10896 11786
rect 10840 11732 10896 11734
rect 10632 10218 10688 10220
rect 10632 10166 10634 10218
rect 10634 10166 10686 10218
rect 10686 10166 10688 10218
rect 10632 10164 10688 10166
rect 10736 10218 10792 10220
rect 10736 10166 10738 10218
rect 10738 10166 10790 10218
rect 10790 10166 10792 10218
rect 10736 10164 10792 10166
rect 10840 10218 10896 10220
rect 10840 10166 10842 10218
rect 10842 10166 10894 10218
rect 10894 10166 10896 10218
rect 10840 10164 10896 10166
rect 9436 9996 9492 10052
rect 9037 9434 9093 9436
rect 9037 9382 9039 9434
rect 9039 9382 9091 9434
rect 9091 9382 9093 9434
rect 9037 9380 9093 9382
rect 9141 9434 9197 9436
rect 9141 9382 9143 9434
rect 9143 9382 9195 9434
rect 9195 9382 9197 9434
rect 9141 9380 9197 9382
rect 9245 9434 9301 9436
rect 9245 9382 9247 9434
rect 9247 9382 9299 9434
rect 9299 9382 9301 9434
rect 9245 9380 9301 9382
rect 9548 8764 9604 8820
rect 8652 8034 8708 8036
rect 8652 7982 8654 8034
rect 8654 7982 8706 8034
rect 8706 7982 8708 8034
rect 8652 7980 8708 7982
rect 9037 7866 9093 7868
rect 9037 7814 9039 7866
rect 9039 7814 9091 7866
rect 9091 7814 9093 7866
rect 9037 7812 9093 7814
rect 9141 7866 9197 7868
rect 9141 7814 9143 7866
rect 9143 7814 9195 7866
rect 9195 7814 9197 7866
rect 9141 7812 9197 7814
rect 9245 7866 9301 7868
rect 9245 7814 9247 7866
rect 9247 7814 9299 7866
rect 9299 7814 9301 7866
rect 9245 7812 9301 7814
rect 8092 7644 8148 7700
rect 8540 7698 8596 7700
rect 8540 7646 8542 7698
rect 8542 7646 8594 7698
rect 8594 7646 8596 7698
rect 8540 7644 8596 7646
rect 7442 7082 7498 7084
rect 7442 7030 7444 7082
rect 7444 7030 7496 7082
rect 7496 7030 7498 7082
rect 7442 7028 7498 7030
rect 7546 7082 7602 7084
rect 7546 7030 7548 7082
rect 7548 7030 7600 7082
rect 7600 7030 7602 7082
rect 7546 7028 7602 7030
rect 7650 7082 7706 7084
rect 7650 7030 7652 7082
rect 7652 7030 7704 7082
rect 7704 7030 7706 7082
rect 7650 7028 7706 7030
rect 5852 6690 5908 6692
rect 5852 6638 5854 6690
rect 5854 6638 5906 6690
rect 5906 6638 5908 6690
rect 5852 6636 5908 6638
rect 6412 6690 6468 6692
rect 6412 6638 6414 6690
rect 6414 6638 6466 6690
rect 6466 6638 6468 6690
rect 6412 6636 6468 6638
rect 5847 6298 5903 6300
rect 5847 6246 5849 6298
rect 5849 6246 5901 6298
rect 5901 6246 5903 6298
rect 5847 6244 5903 6246
rect 5951 6298 6007 6300
rect 5951 6246 5953 6298
rect 5953 6246 6005 6298
rect 6005 6246 6007 6298
rect 5951 6244 6007 6246
rect 6055 6298 6111 6300
rect 6055 6246 6057 6298
rect 6057 6246 6109 6298
rect 6109 6246 6111 6298
rect 6055 6244 6111 6246
rect 8764 6802 8820 6804
rect 8764 6750 8766 6802
rect 8766 6750 8818 6802
rect 8818 6750 8820 6802
rect 8764 6748 8820 6750
rect 9037 6298 9093 6300
rect 9037 6246 9039 6298
rect 9039 6246 9091 6298
rect 9091 6246 9093 6298
rect 9037 6244 9093 6246
rect 9141 6298 9197 6300
rect 9141 6246 9143 6298
rect 9143 6246 9195 6298
rect 9195 6246 9197 6298
rect 9141 6244 9197 6246
rect 9245 6298 9301 6300
rect 9245 6246 9247 6298
rect 9247 6246 9299 6298
rect 9299 6246 9301 6298
rect 9245 6244 9301 6246
rect 5847 4730 5903 4732
rect 5847 4678 5849 4730
rect 5849 4678 5901 4730
rect 5901 4678 5903 4730
rect 5847 4676 5903 4678
rect 5951 4730 6007 4732
rect 5951 4678 5953 4730
rect 5953 4678 6005 4730
rect 6005 4678 6007 4730
rect 5951 4676 6007 4678
rect 6055 4730 6111 4732
rect 6055 4678 6057 4730
rect 6057 4678 6109 4730
rect 6109 4678 6111 4730
rect 6055 4676 6111 4678
rect 5404 4060 5460 4116
rect 5628 4060 5684 4116
rect 5516 3388 5572 3444
rect 5068 3276 5124 3332
rect 4956 2044 5012 2100
rect 6524 4060 6580 4116
rect 6300 3500 6356 3556
rect 6076 3330 6132 3332
rect 6076 3278 6078 3330
rect 6078 3278 6130 3330
rect 6130 3278 6132 3330
rect 6076 3276 6132 3278
rect 5847 3162 5903 3164
rect 5847 3110 5849 3162
rect 5849 3110 5901 3162
rect 5901 3110 5903 3162
rect 5847 3108 5903 3110
rect 5951 3162 6007 3164
rect 5951 3110 5953 3162
rect 5953 3110 6005 3162
rect 6005 3110 6007 3162
rect 5951 3108 6007 3110
rect 6055 3162 6111 3164
rect 6055 3110 6057 3162
rect 6057 3110 6109 3162
rect 6109 3110 6111 3162
rect 6055 3108 6111 3110
rect 5852 2882 5908 2884
rect 5852 2830 5854 2882
rect 5854 2830 5906 2882
rect 5906 2830 5908 2882
rect 5852 2828 5908 2830
rect 5628 2716 5684 2772
rect 4732 1596 4788 1652
rect 7442 5514 7498 5516
rect 7442 5462 7444 5514
rect 7444 5462 7496 5514
rect 7496 5462 7498 5514
rect 7442 5460 7498 5462
rect 7546 5514 7602 5516
rect 7546 5462 7548 5514
rect 7548 5462 7600 5514
rect 7600 5462 7602 5514
rect 7546 5460 7602 5462
rect 7650 5514 7706 5516
rect 7650 5462 7652 5514
rect 7652 5462 7704 5514
rect 7704 5462 7706 5514
rect 7650 5460 7706 5462
rect 9037 4730 9093 4732
rect 9037 4678 9039 4730
rect 9039 4678 9091 4730
rect 9091 4678 9093 4730
rect 9037 4676 9093 4678
rect 9141 4730 9197 4732
rect 9141 4678 9143 4730
rect 9143 4678 9195 4730
rect 9195 4678 9197 4730
rect 9141 4676 9197 4678
rect 9245 4730 9301 4732
rect 9245 4678 9247 4730
rect 9247 4678 9299 4730
rect 9299 4678 9301 4730
rect 9245 4676 9301 4678
rect 7442 3946 7498 3948
rect 7442 3894 7444 3946
rect 7444 3894 7496 3946
rect 7496 3894 7498 3946
rect 7442 3892 7498 3894
rect 7546 3946 7602 3948
rect 7546 3894 7548 3946
rect 7548 3894 7600 3946
rect 7600 3894 7602 3946
rect 7546 3892 7602 3894
rect 7650 3946 7706 3948
rect 7650 3894 7652 3946
rect 7652 3894 7704 3946
rect 7704 3894 7706 3946
rect 7650 3892 7706 3894
rect 7868 3554 7924 3556
rect 7868 3502 7870 3554
rect 7870 3502 7922 3554
rect 7922 3502 7924 3554
rect 7868 3500 7924 3502
rect 8428 3554 8484 3556
rect 8428 3502 8430 3554
rect 8430 3502 8482 3554
rect 8482 3502 8484 3554
rect 8428 3500 8484 3502
rect 10632 8650 10688 8652
rect 10632 8598 10634 8650
rect 10634 8598 10686 8650
rect 10686 8598 10688 8650
rect 10632 8596 10688 8598
rect 10736 8650 10792 8652
rect 10736 8598 10738 8650
rect 10738 8598 10790 8650
rect 10790 8598 10792 8650
rect 10736 8596 10792 8598
rect 10840 8650 10896 8652
rect 10840 8598 10842 8650
rect 10842 8598 10894 8650
rect 10894 8598 10896 8650
rect 10840 8596 10896 8598
rect 11004 7980 11060 8036
rect 9660 7420 9716 7476
rect 10108 7308 10164 7364
rect 10556 7308 10612 7364
rect 10632 7082 10688 7084
rect 10632 7030 10634 7082
rect 10634 7030 10686 7082
rect 10686 7030 10688 7082
rect 10632 7028 10688 7030
rect 10736 7082 10792 7084
rect 10736 7030 10738 7082
rect 10738 7030 10790 7082
rect 10790 7030 10792 7082
rect 10736 7028 10792 7030
rect 10840 7082 10896 7084
rect 10840 7030 10842 7082
rect 10842 7030 10894 7082
rect 10894 7030 10896 7082
rect 10840 7028 10896 7030
rect 9996 6076 10052 6132
rect 10632 5514 10688 5516
rect 10632 5462 10634 5514
rect 10634 5462 10686 5514
rect 10686 5462 10688 5514
rect 10632 5460 10688 5462
rect 10736 5514 10792 5516
rect 10736 5462 10738 5514
rect 10738 5462 10790 5514
rect 10790 5462 10792 5514
rect 10736 5460 10792 5462
rect 10840 5514 10896 5516
rect 10840 5462 10842 5514
rect 10842 5462 10894 5514
rect 10894 5462 10896 5514
rect 10840 5460 10896 5462
rect 9996 4956 10052 5012
rect 10892 4562 10948 4564
rect 10892 4510 10894 4562
rect 10894 4510 10946 4562
rect 10946 4510 10948 4562
rect 10892 4508 10948 4510
rect 10632 3946 10688 3948
rect 10632 3894 10634 3946
rect 10634 3894 10686 3946
rect 10686 3894 10688 3946
rect 10632 3892 10688 3894
rect 10736 3946 10792 3948
rect 10736 3894 10738 3946
rect 10738 3894 10790 3946
rect 10790 3894 10792 3946
rect 10736 3892 10792 3894
rect 10840 3946 10896 3948
rect 10840 3894 10842 3946
rect 10842 3894 10894 3946
rect 10894 3894 10896 3946
rect 10840 3892 10896 3894
rect 9548 3500 9604 3556
rect 6972 3388 7028 3444
rect 6300 1762 6356 1764
rect 6300 1710 6302 1762
rect 6302 1710 6354 1762
rect 6354 1710 6356 1762
rect 6300 1708 6356 1710
rect 5847 1594 5903 1596
rect 5847 1542 5849 1594
rect 5849 1542 5901 1594
rect 5901 1542 5903 1594
rect 5847 1540 5903 1542
rect 5951 1594 6007 1596
rect 5951 1542 5953 1594
rect 5953 1542 6005 1594
rect 6005 1542 6007 1594
rect 5951 1540 6007 1542
rect 6055 1594 6111 1596
rect 6055 1542 6057 1594
rect 6057 1542 6109 1594
rect 6109 1542 6111 1594
rect 6055 1540 6111 1542
rect 6972 3164 7028 3220
rect 9037 3162 9093 3164
rect 9037 3110 9039 3162
rect 9039 3110 9091 3162
rect 9091 3110 9093 3162
rect 9037 3108 9093 3110
rect 9141 3162 9197 3164
rect 9141 3110 9143 3162
rect 9143 3110 9195 3162
rect 9195 3110 9197 3162
rect 9141 3108 9197 3110
rect 9245 3162 9301 3164
rect 9245 3110 9247 3162
rect 9247 3110 9299 3162
rect 9299 3110 9301 3162
rect 9245 3108 9301 3110
rect 7868 2940 7924 2996
rect 10332 3724 10388 3780
rect 10332 3500 10388 3556
rect 10780 3724 10836 3780
rect 7196 2492 7252 2548
rect 7442 2378 7498 2380
rect 7442 2326 7444 2378
rect 7444 2326 7496 2378
rect 7496 2326 7498 2378
rect 7442 2324 7498 2326
rect 7546 2378 7602 2380
rect 7546 2326 7548 2378
rect 7548 2326 7600 2378
rect 7600 2326 7602 2378
rect 7546 2324 7602 2326
rect 7650 2378 7706 2380
rect 7650 2326 7652 2378
rect 7652 2326 7704 2378
rect 7704 2326 7706 2378
rect 7650 2324 7706 2326
rect 7420 1874 7476 1876
rect 7420 1822 7422 1874
rect 7422 1822 7474 1874
rect 7474 1822 7476 1874
rect 7420 1820 7476 1822
rect 7980 1820 8036 1876
rect 10632 2378 10688 2380
rect 10632 2326 10634 2378
rect 10634 2326 10686 2378
rect 10686 2326 10688 2378
rect 10632 2324 10688 2326
rect 10736 2378 10792 2380
rect 10736 2326 10738 2378
rect 10738 2326 10790 2378
rect 10790 2326 10792 2378
rect 10736 2324 10792 2326
rect 10840 2378 10896 2380
rect 10840 2326 10842 2378
rect 10842 2326 10894 2378
rect 10894 2326 10896 2378
rect 10840 2324 10896 2326
rect 11228 11452 11284 11508
rect 11340 11116 11396 11172
rect 12460 12796 12516 12852
rect 12124 11116 12180 11172
rect 12227 11002 12283 11004
rect 12227 10950 12229 11002
rect 12229 10950 12281 11002
rect 12281 10950 12283 11002
rect 12227 10948 12283 10950
rect 12331 11002 12387 11004
rect 12331 10950 12333 11002
rect 12333 10950 12385 11002
rect 12385 10950 12387 11002
rect 12331 10948 12387 10950
rect 12435 11002 12491 11004
rect 12435 10950 12437 11002
rect 12437 10950 12489 11002
rect 12489 10950 12491 11002
rect 12435 10948 12491 10950
rect 11900 10780 11956 10836
rect 11228 10444 11284 10500
rect 11340 8034 11396 8036
rect 11340 7982 11342 8034
rect 11342 7982 11394 8034
rect 11394 7982 11396 8034
rect 11340 7980 11396 7982
rect 12796 11116 12852 11172
rect 14140 11228 14196 11284
rect 13468 10780 13524 10836
rect 12012 9996 12068 10052
rect 12227 9434 12283 9436
rect 12227 9382 12229 9434
rect 12229 9382 12281 9434
rect 12281 9382 12283 9434
rect 12227 9380 12283 9382
rect 12331 9434 12387 9436
rect 12331 9382 12333 9434
rect 12333 9382 12385 9434
rect 12385 9382 12387 9434
rect 12331 9380 12387 9382
rect 12435 9434 12491 9436
rect 12435 9382 12437 9434
rect 12437 9382 12489 9434
rect 12489 9382 12491 9434
rect 12435 9380 12491 9382
rect 11900 7980 11956 8036
rect 12227 7866 12283 7868
rect 12227 7814 12229 7866
rect 12229 7814 12281 7866
rect 12281 7814 12283 7866
rect 12227 7812 12283 7814
rect 12331 7866 12387 7868
rect 12331 7814 12333 7866
rect 12333 7814 12385 7866
rect 12385 7814 12387 7866
rect 12331 7812 12387 7814
rect 12435 7866 12491 7868
rect 12435 7814 12437 7866
rect 12437 7814 12489 7866
rect 12489 7814 12491 7866
rect 12435 7812 12491 7814
rect 12796 6748 12852 6804
rect 12227 6298 12283 6300
rect 12227 6246 12229 6298
rect 12229 6246 12281 6298
rect 12281 6246 12283 6298
rect 12227 6244 12283 6246
rect 12331 6298 12387 6300
rect 12331 6246 12333 6298
rect 12333 6246 12385 6298
rect 12385 6246 12387 6298
rect 12331 6244 12387 6246
rect 12435 6298 12491 6300
rect 12435 6246 12437 6298
rect 12437 6246 12489 6298
rect 12489 6246 12491 6298
rect 12435 6244 12491 6246
rect 12227 4730 12283 4732
rect 12227 4678 12229 4730
rect 12229 4678 12281 4730
rect 12281 4678 12283 4730
rect 12227 4676 12283 4678
rect 12331 4730 12387 4732
rect 12331 4678 12333 4730
rect 12333 4678 12385 4730
rect 12385 4678 12387 4730
rect 12331 4676 12387 4678
rect 12435 4730 12491 4732
rect 12435 4678 12437 4730
rect 12437 4678 12489 4730
rect 12489 4678 12491 4730
rect 12435 4676 12491 4678
rect 12684 4732 12740 4788
rect 11116 4508 11172 4564
rect 11116 3724 11172 3780
rect 11900 4060 11956 4116
rect 11116 3554 11172 3556
rect 11116 3502 11118 3554
rect 11118 3502 11170 3554
rect 11170 3502 11172 3554
rect 11116 3500 11172 3502
rect 11116 2940 11172 2996
rect 8652 1762 8708 1764
rect 8652 1710 8654 1762
rect 8654 1710 8706 1762
rect 8706 1710 8708 1762
rect 8652 1708 8708 1710
rect 9436 1708 9492 1764
rect 9037 1594 9093 1596
rect 9037 1542 9039 1594
rect 9039 1542 9091 1594
rect 9091 1542 9093 1594
rect 9037 1540 9093 1542
rect 9141 1594 9197 1596
rect 9141 1542 9143 1594
rect 9143 1542 9195 1594
rect 9195 1542 9197 1594
rect 9141 1540 9197 1542
rect 9245 1594 9301 1596
rect 9245 1542 9247 1594
rect 9247 1542 9299 1594
rect 9299 1542 9301 1594
rect 9245 1540 9301 1542
rect 12684 3724 12740 3780
rect 12572 3666 12628 3668
rect 12572 3614 12574 3666
rect 12574 3614 12626 3666
rect 12626 3614 12628 3666
rect 12572 3612 12628 3614
rect 12012 3554 12068 3556
rect 12012 3502 12014 3554
rect 12014 3502 12066 3554
rect 12066 3502 12068 3554
rect 12012 3500 12068 3502
rect 12227 3162 12283 3164
rect 12227 3110 12229 3162
rect 12229 3110 12281 3162
rect 12281 3110 12283 3162
rect 12227 3108 12283 3110
rect 12331 3162 12387 3164
rect 12331 3110 12333 3162
rect 12333 3110 12385 3162
rect 12385 3110 12387 3162
rect 12331 3108 12387 3110
rect 12435 3162 12491 3164
rect 12435 3110 12437 3162
rect 12437 3110 12489 3162
rect 12489 3110 12491 3162
rect 12435 3108 12491 3110
rect 12227 1594 12283 1596
rect 12227 1542 12229 1594
rect 12229 1542 12281 1594
rect 12281 1542 12283 1594
rect 12227 1540 12283 1542
rect 12331 1594 12387 1596
rect 12331 1542 12333 1594
rect 12333 1542 12385 1594
rect 12385 1542 12387 1594
rect 12331 1540 12387 1542
rect 12435 1594 12491 1596
rect 12435 1542 12437 1594
rect 12437 1542 12489 1594
rect 12489 1542 12491 1594
rect 12435 1540 12491 1542
rect 4732 700 4788 756
rect 13468 3500 13524 3556
rect 13020 2994 13076 2996
rect 13020 2942 13022 2994
rect 13022 2942 13074 2994
rect 13074 2942 13076 2994
rect 13020 2940 13076 2942
rect 12796 700 12852 756
<< metal3 >>
rect 0 12852 800 12880
rect 14200 12852 15000 12880
rect 0 12796 4732 12852
rect 4788 12796 4798 12852
rect 12450 12796 12460 12852
rect 12516 12796 15000 12852
rect 0 12768 800 12796
rect 14200 12768 15000 12796
rect 4242 11732 4252 11788
rect 4308 11732 4356 11788
rect 4412 11732 4460 11788
rect 4516 11732 4526 11788
rect 7432 11732 7442 11788
rect 7498 11732 7546 11788
rect 7602 11732 7650 11788
rect 7706 11732 7716 11788
rect 10622 11732 10632 11788
rect 10688 11732 10736 11788
rect 10792 11732 10840 11788
rect 10896 11732 10906 11788
rect 0 11508 800 11536
rect 14200 11508 15000 11536
rect 0 11452 2156 11508
rect 2212 11452 2222 11508
rect 11218 11452 11228 11508
rect 11284 11452 15000 11508
rect 0 11424 800 11452
rect 14200 11424 15000 11452
rect 7298 11228 7308 11284
rect 7364 11228 7756 11284
rect 7812 11228 14140 11284
rect 14196 11228 14206 11284
rect 11330 11116 11340 11172
rect 11396 11116 12124 11172
rect 12180 11116 12796 11172
rect 12852 11116 12862 11172
rect 5837 10948 5847 11004
rect 5903 10948 5951 11004
rect 6007 10948 6055 11004
rect 6111 10948 6121 11004
rect 9027 10948 9037 11004
rect 9093 10948 9141 11004
rect 9197 10948 9245 11004
rect 9301 10948 9311 11004
rect 12217 10948 12227 11004
rect 12283 10948 12331 11004
rect 12387 10948 12435 11004
rect 12491 10948 12501 11004
rect 18 10780 28 10836
rect 84 10780 1932 10836
rect 1988 10780 1998 10836
rect 6514 10780 6524 10836
rect 6580 10780 7308 10836
rect 7364 10780 7374 10836
rect 11890 10780 11900 10836
rect 11956 10780 13468 10836
rect 13524 10780 13534 10836
rect 2482 10668 2492 10724
rect 2548 10668 3052 10724
rect 3108 10668 3500 10724
rect 3556 10668 3566 10724
rect 6738 10444 6748 10500
rect 6804 10444 7980 10500
rect 8036 10444 8046 10500
rect 8194 10444 8204 10500
rect 8260 10444 11228 10500
rect 11284 10444 11294 10500
rect 1036 10332 6972 10388
rect 7028 10332 7038 10388
rect 7186 10332 7196 10388
rect 7252 10332 11396 10388
rect 0 10164 800 10192
rect 1036 10164 1092 10332
rect 4242 10164 4252 10220
rect 4308 10164 4356 10220
rect 4412 10164 4460 10220
rect 4516 10164 4526 10220
rect 7432 10164 7442 10220
rect 7498 10164 7546 10220
rect 7602 10164 7650 10220
rect 7706 10164 7716 10220
rect 10622 10164 10632 10220
rect 10688 10164 10736 10220
rect 10792 10164 10840 10220
rect 10896 10164 10906 10220
rect 11340 10164 11396 10332
rect 14200 10164 15000 10192
rect 0 10108 1092 10164
rect 11340 10108 15000 10164
rect 0 10080 800 10108
rect 14200 10080 15000 10108
rect 2370 9996 2380 10052
rect 2436 9996 5404 10052
rect 5460 9996 5470 10052
rect 9426 9996 9436 10052
rect 9492 9996 12012 10052
rect 12068 9996 12078 10052
rect 5837 9380 5847 9436
rect 5903 9380 5951 9436
rect 6007 9380 6055 9436
rect 6111 9380 6121 9436
rect 9027 9380 9037 9436
rect 9093 9380 9141 9436
rect 9197 9380 9245 9436
rect 9301 9380 9311 9436
rect 12217 9380 12227 9436
rect 12283 9380 12331 9436
rect 12387 9380 12435 9436
rect 12491 9380 12501 9436
rect 0 8820 800 8848
rect 14200 8820 15000 8848
rect 0 8764 2156 8820
rect 2212 8764 2222 8820
rect 9538 8764 9548 8820
rect 9604 8764 15000 8820
rect 0 8736 800 8764
rect 14200 8736 15000 8764
rect 4242 8596 4252 8652
rect 4308 8596 4356 8652
rect 4412 8596 4460 8652
rect 4516 8596 4526 8652
rect 7432 8596 7442 8652
rect 7498 8596 7546 8652
rect 7602 8596 7650 8652
rect 7706 8596 7716 8652
rect 10622 8596 10632 8652
rect 10688 8596 10736 8652
rect 10792 8596 10840 8652
rect 10896 8596 10906 8652
rect 6290 8204 6300 8260
rect 6356 8204 7308 8260
rect 7364 8204 7374 8260
rect 7522 7980 7532 8036
rect 7588 7980 8652 8036
rect 8708 7980 8718 8036
rect 10994 7980 11004 8036
rect 11060 7980 11340 8036
rect 11396 7980 11900 8036
rect 11956 7980 11966 8036
rect 5837 7812 5847 7868
rect 5903 7812 5951 7868
rect 6007 7812 6055 7868
rect 6111 7812 6121 7868
rect 9027 7812 9037 7868
rect 9093 7812 9141 7868
rect 9197 7812 9245 7868
rect 9301 7812 9311 7868
rect 12217 7812 12227 7868
rect 12283 7812 12331 7868
rect 12387 7812 12435 7868
rect 12491 7812 12501 7868
rect 1810 7644 1820 7700
rect 1876 7644 7084 7700
rect 7140 7644 7532 7700
rect 7588 7644 7598 7700
rect 8082 7644 8092 7700
rect 8148 7644 8540 7700
rect 8596 7644 10388 7700
rect 3378 7532 3388 7588
rect 3444 7532 5852 7588
rect 5908 7532 5918 7588
rect 0 7476 800 7504
rect 10332 7476 10388 7644
rect 14200 7476 15000 7504
rect 0 7420 9660 7476
rect 9716 7420 9726 7476
rect 10332 7420 15000 7476
rect 0 7392 800 7420
rect 9660 7364 9716 7420
rect 14200 7392 15000 7420
rect 4946 7308 4956 7364
rect 5012 7308 6300 7364
rect 6356 7308 6524 7364
rect 6580 7308 6590 7364
rect 9660 7308 10108 7364
rect 10164 7308 10556 7364
rect 10612 7308 10622 7364
rect 4242 7028 4252 7084
rect 4308 7028 4356 7084
rect 4412 7028 4460 7084
rect 4516 7028 4526 7084
rect 7432 7028 7442 7084
rect 7498 7028 7546 7084
rect 7602 7028 7650 7084
rect 7706 7028 7716 7084
rect 10622 7028 10632 7084
rect 10688 7028 10736 7084
rect 10792 7028 10840 7084
rect 10896 7028 10906 7084
rect 8754 6748 8764 6804
rect 8820 6748 12796 6804
rect 12852 6748 12862 6804
rect 5842 6636 5852 6692
rect 5908 6636 6412 6692
rect 6468 6636 6478 6692
rect 5837 6244 5847 6300
rect 5903 6244 5951 6300
rect 6007 6244 6055 6300
rect 6111 6244 6121 6300
rect 9027 6244 9037 6300
rect 9093 6244 9141 6300
rect 9197 6244 9245 6300
rect 9301 6244 9311 6300
rect 12217 6244 12227 6300
rect 12283 6244 12331 6300
rect 12387 6244 12435 6300
rect 12491 6244 12501 6300
rect 0 6132 800 6160
rect 14200 6132 15000 6160
rect 0 6076 3500 6132
rect 3556 6076 3566 6132
rect 9986 6076 9996 6132
rect 10052 6076 15000 6132
rect 0 6048 800 6076
rect 14200 6048 15000 6076
rect 4242 5460 4252 5516
rect 4308 5460 4356 5516
rect 4412 5460 4460 5516
rect 4516 5460 4526 5516
rect 7432 5460 7442 5516
rect 7498 5460 7546 5516
rect 7602 5460 7650 5516
rect 7706 5460 7716 5516
rect 10622 5460 10632 5516
rect 10688 5460 10736 5516
rect 10792 5460 10840 5516
rect 10896 5460 10906 5516
rect 3378 4956 3388 5012
rect 3444 4956 4060 5012
rect 4116 4956 9996 5012
rect 10052 4956 10062 5012
rect 0 4788 800 4816
rect 14200 4788 15000 4816
rect 0 4732 3500 4788
rect 3556 4732 3566 4788
rect 12674 4732 12684 4788
rect 12740 4732 15000 4788
rect 0 4704 800 4732
rect 5837 4676 5847 4732
rect 5903 4676 5951 4732
rect 6007 4676 6055 4732
rect 6111 4676 6121 4732
rect 9027 4676 9037 4732
rect 9093 4676 9141 4732
rect 9197 4676 9245 4732
rect 9301 4676 9311 4732
rect 12217 4676 12227 4732
rect 12283 4676 12331 4732
rect 12387 4676 12435 4732
rect 12491 4676 12501 4732
rect 14200 4704 15000 4732
rect 10882 4508 10892 4564
rect 10948 4508 11116 4564
rect 11172 4508 11182 4564
rect 18 4060 28 4116
rect 84 4060 1820 4116
rect 1876 4060 2268 4116
rect 2324 4060 5404 4116
rect 5460 4060 5470 4116
rect 5618 4060 5628 4116
rect 5684 4060 6524 4116
rect 6580 4060 11900 4116
rect 11956 4060 11966 4116
rect 4242 3892 4252 3948
rect 4308 3892 4356 3948
rect 4412 3892 4460 3948
rect 4516 3892 4526 3948
rect 7432 3892 7442 3948
rect 7498 3892 7546 3948
rect 7602 3892 7650 3948
rect 7706 3892 7716 3948
rect 10622 3892 10632 3948
rect 10688 3892 10736 3948
rect 10792 3892 10840 3948
rect 10896 3892 10906 3948
rect 1362 3724 1372 3780
rect 1428 3724 10332 3780
rect 10388 3724 10398 3780
rect 10770 3724 10780 3780
rect 10836 3724 11116 3780
rect 11172 3724 12684 3780
rect 12740 3724 12750 3780
rect 9548 3612 12572 3668
rect 12628 3612 12638 3668
rect 9548 3556 9604 3612
rect 2818 3500 2828 3556
rect 2884 3500 4060 3556
rect 4116 3500 4126 3556
rect 6290 3500 6300 3556
rect 6356 3500 7868 3556
rect 7924 3500 7934 3556
rect 8418 3500 8428 3556
rect 8484 3500 9548 3556
rect 9604 3500 9614 3556
rect 10322 3500 10332 3556
rect 10388 3500 11116 3556
rect 11172 3500 11182 3556
rect 12002 3500 12012 3556
rect 12068 3500 13468 3556
rect 13524 3500 13534 3556
rect 0 3444 800 3472
rect 14200 3444 15000 3472
rect 0 3388 2268 3444
rect 2324 3388 2334 3444
rect 5506 3388 5516 3444
rect 5572 3388 6972 3444
rect 7028 3388 7038 3444
rect 8372 3388 15000 3444
rect 0 3360 800 3388
rect 8372 3332 8428 3388
rect 14200 3360 15000 3388
rect 2706 3276 2716 3332
rect 2772 3276 3612 3332
rect 3668 3276 3678 3332
rect 5058 3276 5068 3332
rect 5124 3276 6076 3332
rect 6132 3276 8428 3332
rect 6972 3220 7028 3276
rect 6962 3164 6972 3220
rect 7028 3164 7038 3220
rect 5837 3108 5847 3164
rect 5903 3108 5951 3164
rect 6007 3108 6055 3164
rect 6111 3108 6121 3164
rect 9027 3108 9037 3164
rect 9093 3108 9141 3164
rect 9197 3108 9245 3164
rect 9301 3108 9311 3164
rect 12217 3108 12227 3164
rect 12283 3108 12331 3164
rect 12387 3108 12435 3164
rect 12491 3108 12501 3164
rect 4722 2940 4732 2996
rect 4788 2940 7868 2996
rect 7924 2940 7934 2996
rect 11106 2940 11116 2996
rect 11172 2940 13020 2996
rect 13076 2940 13086 2996
rect 3490 2828 3500 2884
rect 3556 2828 5852 2884
rect 5908 2828 5918 2884
rect 4610 2716 4620 2772
rect 4676 2716 5628 2772
rect 5684 2716 5694 2772
rect 7186 2492 7196 2548
rect 7252 2492 8428 2548
rect 4242 2324 4252 2380
rect 4308 2324 4356 2380
rect 4412 2324 4460 2380
rect 4516 2324 4526 2380
rect 7432 2324 7442 2380
rect 7498 2324 7546 2380
rect 7602 2324 7650 2380
rect 7706 2324 7716 2380
rect 0 2100 800 2128
rect 8372 2100 8428 2492
rect 10622 2324 10632 2380
rect 10688 2324 10736 2380
rect 10792 2324 10840 2380
rect 10896 2324 10906 2380
rect 14200 2100 15000 2128
rect 0 2044 4956 2100
rect 5012 2044 5022 2100
rect 8372 2044 15000 2100
rect 0 2016 800 2044
rect 14200 2016 15000 2044
rect 7410 1820 7420 1876
rect 7476 1820 7980 1876
rect 8036 1820 8046 1876
rect 18 1708 28 1764
rect 84 1708 2156 1764
rect 2212 1708 2222 1764
rect 5628 1708 6300 1764
rect 6356 1708 6366 1764
rect 8642 1708 8652 1764
rect 8708 1708 9436 1764
rect 9492 1708 9502 1764
rect 5628 1652 5684 1708
rect 4722 1596 4732 1652
rect 4788 1596 5684 1652
rect 5837 1540 5847 1596
rect 5903 1540 5951 1596
rect 6007 1540 6055 1596
rect 6111 1540 6121 1596
rect 9027 1540 9037 1596
rect 9093 1540 9141 1596
rect 9197 1540 9245 1596
rect 9301 1540 9311 1596
rect 12217 1540 12227 1596
rect 12283 1540 12331 1596
rect 12387 1540 12435 1596
rect 12491 1540 12501 1596
rect 0 756 800 784
rect 14200 756 15000 784
rect 0 700 4732 756
rect 4788 700 4798 756
rect 12786 700 12796 756
rect 12852 700 15000 756
rect 0 672 800 700
rect 14200 672 15000 700
<< via3 >>
rect 4252 11732 4308 11788
rect 4356 11732 4412 11788
rect 4460 11732 4516 11788
rect 7442 11732 7498 11788
rect 7546 11732 7602 11788
rect 7650 11732 7706 11788
rect 10632 11732 10688 11788
rect 10736 11732 10792 11788
rect 10840 11732 10896 11788
rect 5847 10948 5903 11004
rect 5951 10948 6007 11004
rect 6055 10948 6111 11004
rect 9037 10948 9093 11004
rect 9141 10948 9197 11004
rect 9245 10948 9301 11004
rect 12227 10948 12283 11004
rect 12331 10948 12387 11004
rect 12435 10948 12491 11004
rect 4252 10164 4308 10220
rect 4356 10164 4412 10220
rect 4460 10164 4516 10220
rect 7442 10164 7498 10220
rect 7546 10164 7602 10220
rect 7650 10164 7706 10220
rect 10632 10164 10688 10220
rect 10736 10164 10792 10220
rect 10840 10164 10896 10220
rect 5847 9380 5903 9436
rect 5951 9380 6007 9436
rect 6055 9380 6111 9436
rect 9037 9380 9093 9436
rect 9141 9380 9197 9436
rect 9245 9380 9301 9436
rect 12227 9380 12283 9436
rect 12331 9380 12387 9436
rect 12435 9380 12491 9436
rect 4252 8596 4308 8652
rect 4356 8596 4412 8652
rect 4460 8596 4516 8652
rect 7442 8596 7498 8652
rect 7546 8596 7602 8652
rect 7650 8596 7706 8652
rect 10632 8596 10688 8652
rect 10736 8596 10792 8652
rect 10840 8596 10896 8652
rect 5847 7812 5903 7868
rect 5951 7812 6007 7868
rect 6055 7812 6111 7868
rect 9037 7812 9093 7868
rect 9141 7812 9197 7868
rect 9245 7812 9301 7868
rect 12227 7812 12283 7868
rect 12331 7812 12387 7868
rect 12435 7812 12491 7868
rect 4252 7028 4308 7084
rect 4356 7028 4412 7084
rect 4460 7028 4516 7084
rect 7442 7028 7498 7084
rect 7546 7028 7602 7084
rect 7650 7028 7706 7084
rect 10632 7028 10688 7084
rect 10736 7028 10792 7084
rect 10840 7028 10896 7084
rect 5847 6244 5903 6300
rect 5951 6244 6007 6300
rect 6055 6244 6111 6300
rect 9037 6244 9093 6300
rect 9141 6244 9197 6300
rect 9245 6244 9301 6300
rect 12227 6244 12283 6300
rect 12331 6244 12387 6300
rect 12435 6244 12491 6300
rect 4252 5460 4308 5516
rect 4356 5460 4412 5516
rect 4460 5460 4516 5516
rect 7442 5460 7498 5516
rect 7546 5460 7602 5516
rect 7650 5460 7706 5516
rect 10632 5460 10688 5516
rect 10736 5460 10792 5516
rect 10840 5460 10896 5516
rect 5847 4676 5903 4732
rect 5951 4676 6007 4732
rect 6055 4676 6111 4732
rect 9037 4676 9093 4732
rect 9141 4676 9197 4732
rect 9245 4676 9301 4732
rect 12227 4676 12283 4732
rect 12331 4676 12387 4732
rect 12435 4676 12491 4732
rect 4252 3892 4308 3948
rect 4356 3892 4412 3948
rect 4460 3892 4516 3948
rect 7442 3892 7498 3948
rect 7546 3892 7602 3948
rect 7650 3892 7706 3948
rect 10632 3892 10688 3948
rect 10736 3892 10792 3948
rect 10840 3892 10896 3948
rect 5847 3108 5903 3164
rect 5951 3108 6007 3164
rect 6055 3108 6111 3164
rect 9037 3108 9093 3164
rect 9141 3108 9197 3164
rect 9245 3108 9301 3164
rect 12227 3108 12283 3164
rect 12331 3108 12387 3164
rect 12435 3108 12491 3164
rect 4252 2324 4308 2380
rect 4356 2324 4412 2380
rect 4460 2324 4516 2380
rect 7442 2324 7498 2380
rect 7546 2324 7602 2380
rect 7650 2324 7706 2380
rect 10632 2324 10688 2380
rect 10736 2324 10792 2380
rect 10840 2324 10896 2380
rect 5847 1540 5903 1596
rect 5951 1540 6007 1596
rect 6055 1540 6111 1596
rect 9037 1540 9093 1596
rect 9141 1540 9197 1596
rect 9245 1540 9301 1596
rect 12227 1540 12283 1596
rect 12331 1540 12387 1596
rect 12435 1540 12491 1596
<< metal4 >>
rect 4224 11788 4544 11820
rect 4224 11732 4252 11788
rect 4308 11732 4356 11788
rect 4412 11732 4460 11788
rect 4516 11732 4544 11788
rect 4224 10220 4544 11732
rect 4224 10164 4252 10220
rect 4308 10164 4356 10220
rect 4412 10164 4460 10220
rect 4516 10164 4544 10220
rect 4224 8652 4544 10164
rect 4224 8596 4252 8652
rect 4308 8596 4356 8652
rect 4412 8596 4460 8652
rect 4516 8596 4544 8652
rect 4224 7084 4544 8596
rect 4224 7028 4252 7084
rect 4308 7028 4356 7084
rect 4412 7028 4460 7084
rect 4516 7028 4544 7084
rect 4224 5516 4544 7028
rect 4224 5460 4252 5516
rect 4308 5460 4356 5516
rect 4412 5460 4460 5516
rect 4516 5460 4544 5516
rect 4224 5030 4544 5460
rect 4224 4974 4252 5030
rect 4308 4974 4356 5030
rect 4412 4974 4460 5030
rect 4516 4974 4544 5030
rect 4224 4926 4544 4974
rect 4224 4870 4252 4926
rect 4308 4870 4356 4926
rect 4412 4870 4460 4926
rect 4516 4870 4544 4926
rect 4224 4822 4544 4870
rect 4224 4766 4252 4822
rect 4308 4766 4356 4822
rect 4412 4766 4460 4822
rect 4516 4766 4544 4822
rect 4224 3948 4544 4766
rect 4224 3892 4252 3948
rect 4308 3892 4356 3948
rect 4412 3892 4460 3948
rect 4516 3892 4544 3948
rect 4224 2380 4544 3892
rect 4224 2324 4252 2380
rect 4308 2324 4356 2380
rect 4412 2324 4460 2380
rect 4516 2324 4544 2380
rect 4224 1508 4544 2324
rect 5819 11004 6139 11820
rect 5819 10948 5847 11004
rect 5903 10948 5951 11004
rect 6007 10948 6055 11004
rect 6111 10948 6139 11004
rect 5819 9436 6139 10948
rect 5819 9380 5847 9436
rect 5903 9380 5951 9436
rect 6007 9380 6055 9436
rect 6111 9380 6139 9436
rect 5819 7868 6139 9380
rect 5819 7812 5847 7868
rect 5903 7812 5951 7868
rect 6007 7812 6055 7868
rect 6111 7812 6139 7868
rect 5819 6388 6139 7812
rect 5819 6332 5847 6388
rect 5903 6332 5951 6388
rect 6007 6332 6055 6388
rect 6111 6332 6139 6388
rect 5819 6300 6139 6332
rect 5819 6228 5847 6300
rect 5903 6228 5951 6300
rect 6007 6228 6055 6300
rect 6111 6228 6139 6300
rect 5819 6180 6139 6228
rect 5819 6124 5847 6180
rect 5903 6124 5951 6180
rect 6007 6124 6055 6180
rect 6111 6124 6139 6180
rect 5819 4732 6139 6124
rect 5819 4676 5847 4732
rect 5903 4676 5951 4732
rect 6007 4676 6055 4732
rect 6111 4676 6139 4732
rect 5819 3164 6139 4676
rect 5819 3108 5847 3164
rect 5903 3108 5951 3164
rect 6007 3108 6055 3164
rect 6111 3108 6139 3164
rect 5819 1596 6139 3108
rect 5819 1540 5847 1596
rect 5903 1540 5951 1596
rect 6007 1540 6055 1596
rect 6111 1540 6139 1596
rect 5819 1508 6139 1540
rect 7414 11788 7734 11820
rect 7414 11732 7442 11788
rect 7498 11732 7546 11788
rect 7602 11732 7650 11788
rect 7706 11732 7734 11788
rect 7414 10220 7734 11732
rect 7414 10164 7442 10220
rect 7498 10164 7546 10220
rect 7602 10164 7650 10220
rect 7706 10164 7734 10220
rect 7414 8652 7734 10164
rect 7414 8596 7442 8652
rect 7498 8596 7546 8652
rect 7602 8596 7650 8652
rect 7706 8596 7734 8652
rect 7414 7084 7734 8596
rect 7414 7028 7442 7084
rect 7498 7028 7546 7084
rect 7602 7028 7650 7084
rect 7706 7028 7734 7084
rect 7414 5516 7734 7028
rect 7414 5460 7442 5516
rect 7498 5460 7546 5516
rect 7602 5460 7650 5516
rect 7706 5460 7734 5516
rect 7414 5030 7734 5460
rect 7414 4974 7442 5030
rect 7498 4974 7546 5030
rect 7602 4974 7650 5030
rect 7706 4974 7734 5030
rect 7414 4926 7734 4974
rect 7414 4870 7442 4926
rect 7498 4870 7546 4926
rect 7602 4870 7650 4926
rect 7706 4870 7734 4926
rect 7414 4822 7734 4870
rect 7414 4766 7442 4822
rect 7498 4766 7546 4822
rect 7602 4766 7650 4822
rect 7706 4766 7734 4822
rect 7414 3948 7734 4766
rect 7414 3892 7442 3948
rect 7498 3892 7546 3948
rect 7602 3892 7650 3948
rect 7706 3892 7734 3948
rect 7414 2380 7734 3892
rect 7414 2324 7442 2380
rect 7498 2324 7546 2380
rect 7602 2324 7650 2380
rect 7706 2324 7734 2380
rect 7414 1508 7734 2324
rect 9009 11004 9329 11820
rect 9009 10948 9037 11004
rect 9093 10948 9141 11004
rect 9197 10948 9245 11004
rect 9301 10948 9329 11004
rect 9009 9436 9329 10948
rect 9009 9380 9037 9436
rect 9093 9380 9141 9436
rect 9197 9380 9245 9436
rect 9301 9380 9329 9436
rect 9009 7868 9329 9380
rect 9009 7812 9037 7868
rect 9093 7812 9141 7868
rect 9197 7812 9245 7868
rect 9301 7812 9329 7868
rect 9009 6388 9329 7812
rect 9009 6332 9037 6388
rect 9093 6332 9141 6388
rect 9197 6332 9245 6388
rect 9301 6332 9329 6388
rect 9009 6300 9329 6332
rect 9009 6228 9037 6300
rect 9093 6228 9141 6300
rect 9197 6228 9245 6300
rect 9301 6228 9329 6300
rect 9009 6180 9329 6228
rect 9009 6124 9037 6180
rect 9093 6124 9141 6180
rect 9197 6124 9245 6180
rect 9301 6124 9329 6180
rect 9009 4732 9329 6124
rect 9009 4676 9037 4732
rect 9093 4676 9141 4732
rect 9197 4676 9245 4732
rect 9301 4676 9329 4732
rect 9009 3164 9329 4676
rect 9009 3108 9037 3164
rect 9093 3108 9141 3164
rect 9197 3108 9245 3164
rect 9301 3108 9329 3164
rect 9009 1596 9329 3108
rect 9009 1540 9037 1596
rect 9093 1540 9141 1596
rect 9197 1540 9245 1596
rect 9301 1540 9329 1596
rect 9009 1508 9329 1540
rect 10604 11788 10924 11820
rect 10604 11732 10632 11788
rect 10688 11732 10736 11788
rect 10792 11732 10840 11788
rect 10896 11732 10924 11788
rect 10604 10220 10924 11732
rect 10604 10164 10632 10220
rect 10688 10164 10736 10220
rect 10792 10164 10840 10220
rect 10896 10164 10924 10220
rect 10604 8652 10924 10164
rect 10604 8596 10632 8652
rect 10688 8596 10736 8652
rect 10792 8596 10840 8652
rect 10896 8596 10924 8652
rect 10604 7084 10924 8596
rect 10604 7028 10632 7084
rect 10688 7028 10736 7084
rect 10792 7028 10840 7084
rect 10896 7028 10924 7084
rect 10604 5516 10924 7028
rect 10604 5460 10632 5516
rect 10688 5460 10736 5516
rect 10792 5460 10840 5516
rect 10896 5460 10924 5516
rect 10604 5030 10924 5460
rect 10604 4974 10632 5030
rect 10688 4974 10736 5030
rect 10792 4974 10840 5030
rect 10896 4974 10924 5030
rect 10604 4926 10924 4974
rect 10604 4870 10632 4926
rect 10688 4870 10736 4926
rect 10792 4870 10840 4926
rect 10896 4870 10924 4926
rect 10604 4822 10924 4870
rect 10604 4766 10632 4822
rect 10688 4766 10736 4822
rect 10792 4766 10840 4822
rect 10896 4766 10924 4822
rect 10604 3948 10924 4766
rect 10604 3892 10632 3948
rect 10688 3892 10736 3948
rect 10792 3892 10840 3948
rect 10896 3892 10924 3948
rect 10604 2380 10924 3892
rect 10604 2324 10632 2380
rect 10688 2324 10736 2380
rect 10792 2324 10840 2380
rect 10896 2324 10924 2380
rect 10604 1508 10924 2324
rect 12199 11004 12519 11820
rect 12199 10948 12227 11004
rect 12283 10948 12331 11004
rect 12387 10948 12435 11004
rect 12491 10948 12519 11004
rect 12199 9436 12519 10948
rect 12199 9380 12227 9436
rect 12283 9380 12331 9436
rect 12387 9380 12435 9436
rect 12491 9380 12519 9436
rect 12199 7868 12519 9380
rect 12199 7812 12227 7868
rect 12283 7812 12331 7868
rect 12387 7812 12435 7868
rect 12491 7812 12519 7868
rect 12199 6388 12519 7812
rect 12199 6332 12227 6388
rect 12283 6332 12331 6388
rect 12387 6332 12435 6388
rect 12491 6332 12519 6388
rect 12199 6300 12519 6332
rect 12199 6228 12227 6300
rect 12283 6228 12331 6300
rect 12387 6228 12435 6300
rect 12491 6228 12519 6300
rect 12199 6180 12519 6228
rect 12199 6124 12227 6180
rect 12283 6124 12331 6180
rect 12387 6124 12435 6180
rect 12491 6124 12519 6180
rect 12199 4732 12519 6124
rect 12199 4676 12227 4732
rect 12283 4676 12331 4732
rect 12387 4676 12435 4732
rect 12491 4676 12519 4732
rect 12199 3164 12519 4676
rect 12199 3108 12227 3164
rect 12283 3108 12331 3164
rect 12387 3108 12435 3164
rect 12491 3108 12519 3164
rect 12199 1596 12519 3108
rect 12199 1540 12227 1596
rect 12283 1540 12331 1596
rect 12387 1540 12435 1596
rect 12491 1540 12519 1596
rect 12199 1508 12519 1540
<< via4 >>
rect 4252 4974 4308 5030
rect 4356 4974 4412 5030
rect 4460 4974 4516 5030
rect 4252 4870 4308 4926
rect 4356 4870 4412 4926
rect 4460 4870 4516 4926
rect 4252 4766 4308 4822
rect 4356 4766 4412 4822
rect 4460 4766 4516 4822
rect 5847 6332 5903 6388
rect 5951 6332 6007 6388
rect 6055 6332 6111 6388
rect 5847 6244 5903 6284
rect 5847 6228 5903 6244
rect 5951 6244 6007 6284
rect 5951 6228 6007 6244
rect 6055 6244 6111 6284
rect 6055 6228 6111 6244
rect 5847 6124 5903 6180
rect 5951 6124 6007 6180
rect 6055 6124 6111 6180
rect 7442 4974 7498 5030
rect 7546 4974 7602 5030
rect 7650 4974 7706 5030
rect 7442 4870 7498 4926
rect 7546 4870 7602 4926
rect 7650 4870 7706 4926
rect 7442 4766 7498 4822
rect 7546 4766 7602 4822
rect 7650 4766 7706 4822
rect 9037 6332 9093 6388
rect 9141 6332 9197 6388
rect 9245 6332 9301 6388
rect 9037 6244 9093 6284
rect 9037 6228 9093 6244
rect 9141 6244 9197 6284
rect 9141 6228 9197 6244
rect 9245 6244 9301 6284
rect 9245 6228 9301 6244
rect 9037 6124 9093 6180
rect 9141 6124 9197 6180
rect 9245 6124 9301 6180
rect 10632 4974 10688 5030
rect 10736 4974 10792 5030
rect 10840 4974 10896 5030
rect 10632 4870 10688 4926
rect 10736 4870 10792 4926
rect 10840 4870 10896 4926
rect 10632 4766 10688 4822
rect 10736 4766 10792 4822
rect 10840 4766 10896 4822
rect 12227 6332 12283 6388
rect 12331 6332 12387 6388
rect 12435 6332 12491 6388
rect 12227 6244 12283 6284
rect 12227 6228 12283 6244
rect 12331 6244 12387 6284
rect 12331 6228 12387 6244
rect 12435 6244 12491 6284
rect 12435 6228 12491 6244
rect 12227 6124 12283 6180
rect 12331 6124 12387 6180
rect 12435 6124 12491 6180
<< metal5 >>
rect 1060 6388 13836 6416
rect 1060 6332 5847 6388
rect 5903 6332 5951 6388
rect 6007 6332 6055 6388
rect 6111 6332 9037 6388
rect 9093 6332 9141 6388
rect 9197 6332 9245 6388
rect 9301 6332 12227 6388
rect 12283 6332 12331 6388
rect 12387 6332 12435 6388
rect 12491 6332 13836 6388
rect 1060 6284 13836 6332
rect 1060 6228 5847 6284
rect 5903 6228 5951 6284
rect 6007 6228 6055 6284
rect 6111 6228 9037 6284
rect 9093 6228 9141 6284
rect 9197 6228 9245 6284
rect 9301 6228 12227 6284
rect 12283 6228 12331 6284
rect 12387 6228 12435 6284
rect 12491 6228 13836 6284
rect 1060 6180 13836 6228
rect 1060 6124 5847 6180
rect 5903 6124 5951 6180
rect 6007 6124 6055 6180
rect 6111 6124 9037 6180
rect 9093 6124 9141 6180
rect 9197 6124 9245 6180
rect 9301 6124 12227 6180
rect 12283 6124 12331 6180
rect 12387 6124 12435 6180
rect 12491 6124 13836 6180
rect 1060 6096 13836 6124
rect 1060 5030 13836 5058
rect 1060 4974 4252 5030
rect 4308 4974 4356 5030
rect 4412 4974 4460 5030
rect 4516 4974 7442 5030
rect 7498 4974 7546 5030
rect 7602 4974 7650 5030
rect 7706 4974 10632 5030
rect 10688 4974 10736 5030
rect 10792 4974 10840 5030
rect 10896 4974 13836 5030
rect 1060 4926 13836 4974
rect 1060 4870 4252 4926
rect 4308 4870 4356 4926
rect 4412 4870 4460 4926
rect 4516 4870 7442 4926
rect 7498 4870 7546 4926
rect 7602 4870 7650 4926
rect 7706 4870 10632 4926
rect 10688 4870 10736 4926
rect 10792 4870 10840 4926
rect 10896 4870 13836 4926
rect 1060 4822 13836 4870
rect 1060 4766 4252 4822
rect 4308 4766 4356 4822
rect 4412 4766 4460 4822
rect 4516 4766 7442 4822
rect 7498 4766 7546 4822
rect 7602 4766 7650 4822
rect 7706 4766 10632 4822
rect 10688 4766 10736 4822
rect 10792 4766 10840 4822
rect 10896 4766 13836 4822
rect 1060 4738 13836 4766
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_spare_logic_biginv_I OpenLane/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1670211287
transform -1 0 5936 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_spare_logic_flop\[0\]_CLK
timestamp 1670211287
transform 1 0 5376 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_spare_logic_flop\[0\]_RN
timestamp 1670211287
transform -1 0 6944 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_spare_logic_flop\[0\]_SETN
timestamp 1670211287
transform -1 0 6608 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_spare_logic_flop\[1\]_CLK
timestamp 1670211287
transform -1 0 7728 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_spare_logic_flop\[1\]_D
timestamp 1670211287
transform 1 0 12544 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_spare_logic_flop\[1\]_RN
timestamp 1670211287
transform 1 0 12992 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_spare_logic_flop\[1\]_SETN
timestamp 1670211287
transform 1 0 12544 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_spare_logic_inv\[3\]_I
timestamp 1670211287
transform -1 0 6608 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_spare_logic_mux\[1\]_I1
timestamp 1670211287
transform 1 0 6272 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_spare_logic_mux\[1\]_S
timestamp 1670211287
transform 1 0 8624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_spare_logic_nand\[1\]_A2
timestamp 1670211287
transform 1 0 7952 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_spare_logic_nor\[0\]_A1
timestamp 1670211287
transform -1 0 4368 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_spare_logic_nor\[1\]_A1
timestamp 1670211287
transform -1 0 10192 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2 OpenLane/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1670211287
transform 1 0 1344 0 1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6 OpenLane/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1670211287
transform 1 0 1792 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12 OpenLane/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1670211287
transform 1 0 2464 0 1 1568
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20
timestamp 1670211287
transform 1 0 3360 0 1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24 OpenLane/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1670211287
transform 1 0 3808 0 1 1568
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29
timestamp 1670211287
transform 1 0 4368 0 1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33
timestamp 1670211287
transform 1 0 4816 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37
timestamp 1670211287
transform 1 0 5264 0 1 1568
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42
timestamp 1670211287
transform 1 0 5824 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48
timestamp 1670211287
transform 1 0 6496 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52
timestamp 1670211287
transform 1 0 6944 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54
timestamp 1670211287
transform 1 0 7168 0 1 1568
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59
timestamp 1670211287
transform 1 0 7728 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63
timestamp 1670211287
transform 1 0 8176 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69
timestamp 1670211287
transform 1 0 8848 0 1 1568
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_72 OpenLane/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1670211287
transform 1 0 9184 0 1 1568
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_104
timestamp 1670211287
transform 1 0 12768 0 1 1568
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_107
timestamp 1670211287
transform 1 0 13104 0 1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_2
timestamp 1670211287
transform 1 0 1344 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_45
timestamp 1670211287
transform 1 0 6160 0 -1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_49
timestamp 1670211287
transform 1 0 6608 0 -1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_56
timestamp 1670211287
transform 1 0 7392 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_67
timestamp 1670211287
transform 1 0 8624 0 -1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_73
timestamp 1670211287
transform 1 0 9296 0 -1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_78
timestamp 1670211287
transform 1 0 9856 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_84 OpenLane/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1670211287
transform 1 0 10528 0 -1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_100
timestamp 1670211287
transform 1 0 12320 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_104
timestamp 1670211287
transform 1 0 12768 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_108
timestamp 1670211287
transform 1 0 13216 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_110
timestamp 1670211287
transform 1 0 13440 0 -1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_2
timestamp 1670211287
transform 1 0 1344 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_6
timestamp 1670211287
transform 1 0 1792 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_8
timestamp 1670211287
transform 1 0 2016 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_19
timestamp 1670211287
transform 1 0 3248 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_25
timestamp 1670211287
transform 1 0 3920 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_29
timestamp 1670211287
transform 1 0 4368 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_33
timestamp 1670211287
transform 1 0 4816 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_37
timestamp 1670211287
transform 1 0 5264 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_40
timestamp 1670211287
transform 1 0 5600 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_46
timestamp 1670211287
transform 1 0 6272 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_54
timestamp 1670211287
transform 1 0 7168 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_58
timestamp 1670211287
transform 1 0 7616 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_100
timestamp 1670211287
transform 1 0 12320 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_104
timestamp 1670211287
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_108
timestamp 1670211287
transform 1 0 13216 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_110
timestamp 1670211287
transform 1 0 13440 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_2
timestamp 1670211287
transform 1 0 1344 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_6
timestamp 1670211287
transform 1 0 1792 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_12
timestamp 1670211287
transform 1 0 2464 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_16
timestamp 1670211287
transform 1 0 2912 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_22
timestamp 1670211287
transform 1 0 3584 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_38
timestamp 1670211287
transform 1 0 5376 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_46
timestamp 1670211287
transform 1 0 6272 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_49
timestamp 1670211287
transform 1 0 6608 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_59
timestamp 1670211287
transform 1 0 7728 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_67
timestamp 1670211287
transform 1 0 8624 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_73
timestamp 1670211287
transform 1 0 9296 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_81
timestamp 1670211287
transform 1 0 10192 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_89
timestamp 1670211287
transform 1 0 11088 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_97
timestamp 1670211287
transform 1 0 11984 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_105
timestamp 1670211287
transform 1 0 12880 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_109
timestamp 1670211287
transform 1 0 13328 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_2
timestamp 1670211287
transform 1 0 1344 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_34
timestamp 1670211287
transform 1 0 4928 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_37 OpenLane/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1670211287
transform 1 0 5264 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_101
timestamp 1670211287
transform 1 0 12432 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_105
timestamp 1670211287
transform 1 0 12880 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_108
timestamp 1670211287
transform 1 0 13216 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_110
timestamp 1670211287
transform 1 0 13440 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_2
timestamp 1670211287
transform 1 0 1344 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_34
timestamp 1670211287
transform 1 0 4928 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_50
timestamp 1670211287
transform 1 0 6720 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_57
timestamp 1670211287
transform 1 0 7504 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_65
timestamp 1670211287
transform 1 0 8400 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_69
timestamp 1670211287
transform 1 0 8848 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_73
timestamp 1670211287
transform 1 0 9296 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_105
timestamp 1670211287
transform 1 0 12880 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_109
timestamp 1670211287
transform 1 0 13328 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_2
timestamp 1670211287
transform 1 0 1344 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_34
timestamp 1670211287
transform 1 0 4928 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_37
timestamp 1670211287
transform 1 0 5264 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_43
timestamp 1670211287
transform 1 0 5936 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_71
timestamp 1670211287
transform 1 0 9072 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_81
timestamp 1670211287
transform 1 0 10192 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_97
timestamp 1670211287
transform 1 0 11984 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_105
timestamp 1670211287
transform 1 0 12880 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_108
timestamp 1670211287
transform 1 0 13216 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_110
timestamp 1670211287
transform 1 0 13440 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_2
timestamp 1670211287
transform 1 0 1344 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_34
timestamp 1670211287
transform 1 0 4928 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_38
timestamp 1670211287
transform 1 0 5376 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_44
timestamp 1670211287
transform 1 0 6048 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_50
timestamp 1670211287
transform 1 0 6720 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_56
timestamp 1670211287
transform 1 0 7392 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_62
timestamp 1670211287
transform 1 0 8064 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_68
timestamp 1670211287
transform 1 0 8736 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_70
timestamp 1670211287
transform 1 0 8960 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_73
timestamp 1670211287
transform 1 0 9296 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_79
timestamp 1670211287
transform 1 0 9968 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_91
timestamp 1670211287
transform 1 0 11312 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_107
timestamp 1670211287
transform 1 0 13104 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_2
timestamp 1670211287
transform 1 0 1344 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_6
timestamp 1670211287
transform 1 0 1792 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_12
timestamp 1670211287
transform 1 0 2464 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_28
timestamp 1670211287
transform 1 0 4256 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_32
timestamp 1670211287
transform 1 0 4704 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_34
timestamp 1670211287
transform 1 0 4928 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_37
timestamp 1670211287
transform 1 0 5264 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_45
timestamp 1670211287
transform 1 0 6160 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_48
timestamp 1670211287
transform 1 0 6496 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_65
timestamp 1670211287
transform 1 0 8400 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_69
timestamp 1670211287
transform 1 0 8848 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_85
timestamp 1670211287
transform 1 0 10640 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_93
timestamp 1670211287
transform 1 0 11536 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_101
timestamp 1670211287
transform 1 0 12432 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_105
timestamp 1670211287
transform 1 0 12880 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_108
timestamp 1670211287
transform 1 0 13216 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_110
timestamp 1670211287
transform 1 0 13440 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_2
timestamp 1670211287
transform 1 0 1344 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_66
timestamp 1670211287
transform 1 0 8512 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_70
timestamp 1670211287
transform 1 0 8960 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_73
timestamp 1670211287
transform 1 0 9296 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_105
timestamp 1670211287
transform 1 0 12880 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_109
timestamp 1670211287
transform 1 0 13328 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_2
timestamp 1670211287
transform 1 0 1344 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_10
timestamp 1670211287
transform 1 0 2240 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_15
timestamp 1670211287
transform 1 0 2800 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_31
timestamp 1670211287
transform 1 0 4592 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_37
timestamp 1670211287
transform 1 0 5264 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_53
timestamp 1670211287
transform 1 0 7056 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_57
timestamp 1670211287
transform 1 0 7504 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_63
timestamp 1670211287
transform 1 0 8176 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_95
timestamp 1670211287
transform 1 0 11760 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_101
timestamp 1670211287
transform 1 0 12432 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_105
timestamp 1670211287
transform 1 0 12880 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_108
timestamp 1670211287
transform 1 0 13216 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_110
timestamp 1670211287
transform 1 0 13440 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_2
timestamp 1670211287
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_4
timestamp 1670211287
transform 1 0 1568 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_14
timestamp 1670211287
transform 1 0 2688 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_20
timestamp 1670211287
transform 1 0 3360 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_36
timestamp 1670211287
transform 1 0 5152 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_44
timestamp 1670211287
transform 1 0 6048 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_46
timestamp 1670211287
transform 1 0 6272 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_49
timestamp 1670211287
transform 1 0 6608 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_57
timestamp 1670211287
transform 1 0 7504 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_65
timestamp 1670211287
transform 1 0 8400 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_69
timestamp 1670211287
transform 1 0 8848 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_73
timestamp 1670211287
transform 1 0 9296 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_93
timestamp 1670211287
transform 1 0 11536 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_110
timestamp 1670211287
transform 1 0 13440 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_2
timestamp 1670211287
transform 1 0 1344 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_6
timestamp 1670211287
transform 1 0 1792 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_12
timestamp 1670211287
transform 1 0 2464 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_28
timestamp 1670211287
transform 1 0 4256 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_32
timestamp 1670211287
transform 1 0 4704 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_34
timestamp 1670211287
transform 1 0 4928 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_37
timestamp 1670211287
transform 1 0 5264 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_53
timestamp 1670211287
transform 1 0 7056 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_61
timestamp 1670211287
transform 1 0 7952 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_69
timestamp 1670211287
transform 1 0 8848 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_72
timestamp 1670211287
transform 1 0 9184 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_88
timestamp 1670211287
transform 1 0 10976 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_96
timestamp 1670211287
transform 1 0 11872 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_104
timestamp 1670211287
transform 1 0 12768 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_107
timestamp 1670211287
transform 1 0 13104 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_0 OpenLane/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1670211287
transform 1 0 1120 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_1
timestamp 1670211287
transform -1 0 13776 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_2
timestamp 1670211287
transform 1 0 1120 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_3
timestamp 1670211287
transform -1 0 13776 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_4
timestamp 1670211287
transform 1 0 1120 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_5
timestamp 1670211287
transform -1 0 13776 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_6
timestamp 1670211287
transform 1 0 1120 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_7
timestamp 1670211287
transform -1 0 13776 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_8
timestamp 1670211287
transform 1 0 1120 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_9
timestamp 1670211287
transform -1 0 13776 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_10
timestamp 1670211287
transform 1 0 1120 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_11
timestamp 1670211287
transform -1 0 13776 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_12
timestamp 1670211287
transform 1 0 1120 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_13
timestamp 1670211287
transform -1 0 13776 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_14
timestamp 1670211287
transform 1 0 1120 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_15
timestamp 1670211287
transform -1 0 13776 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_16
timestamp 1670211287
transform 1 0 1120 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_17
timestamp 1670211287
transform -1 0 13776 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_18
timestamp 1670211287
transform 1 0 1120 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_19
timestamp 1670211287
transform -1 0 13776 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_20
timestamp 1670211287
transform 1 0 1120 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_21
timestamp 1670211287
transform -1 0 13776 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_22
timestamp 1670211287
transform 1 0 1120 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_23
timestamp 1670211287
transform -1 0 13776 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_24
timestamp 1670211287
transform 1 0 1120 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_25
timestamp 1670211287
transform -1 0 13776 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_26 OpenLane/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1670211287
transform 1 0 5040 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_27
timestamp 1670211287
transform 1 0 8960 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_28
timestamp 1670211287
transform 1 0 12880 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_29
timestamp 1670211287
transform 1 0 9072 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_30
timestamp 1670211287
transform 1 0 5040 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_31
timestamp 1670211287
transform 1 0 12992 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_32
timestamp 1670211287
transform 1 0 9072 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_33
timestamp 1670211287
transform 1 0 5040 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_34
timestamp 1670211287
transform 1 0 12992 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_35
timestamp 1670211287
transform 1 0 9072 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_36
timestamp 1670211287
transform 1 0 5040 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_37
timestamp 1670211287
transform 1 0 12992 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_38
timestamp 1670211287
transform 1 0 9072 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_39
timestamp 1670211287
transform 1 0 5040 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_40
timestamp 1670211287
transform 1 0 12992 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_41
timestamp 1670211287
transform 1 0 9072 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_42
timestamp 1670211287
transform 1 0 5040 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_43
timestamp 1670211287
transform 1 0 12992 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_44
timestamp 1670211287
transform 1 0 9072 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_45
timestamp 1670211287
transform 1 0 5040 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_46
timestamp 1670211287
transform 1 0 8960 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_47
timestamp 1670211287
transform 1 0 12880 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__inv_12  spare_logic_biginv OpenLane/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1670211287
transform -1 0 9072 0 1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  spare_logic_const_one\[0\] OpenLane/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1670211287
transform -1 0 4368 0 1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  spare_logic_const_one\[1\]
timestamp 1670211287
transform -1 0 2464 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  spare_logic_const_one\[2\]
timestamp 1670211287
transform 1 0 12432 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  spare_logic_const_one\[3\]
timestamp 1670211287
transform -1 0 2464 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spare_logic_const_zero\[0\] OpenLane/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1670211287
transform 1 0 7728 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spare_logic_const_zero\[1\]
timestamp 1670211287
transform 1 0 7616 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spare_logic_const_zero\[2\]
timestamp 1670211287
transform -1 0 7168 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spare_logic_const_zero\[3\]
timestamp 1670211287
transform 1 0 7504 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spare_logic_const_zero\[4\]
timestamp 1670211287
transform 1 0 5600 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spare_logic_const_zero\[5\]
timestamp 1670211287
transform -1 0 2800 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spare_logic_const_zero\[6\]
timestamp 1670211287
transform 1 0 8400 0 1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spare_logic_const_zero\[7\]
timestamp 1670211287
transform -1 0 3360 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spare_logic_const_zero\[8\]
timestamp 1670211287
transform -1 0 7728 0 1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spare_logic_const_zero\[9\]
timestamp 1670211287
transform 1 0 3136 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spare_logic_const_zero\[10\]
timestamp 1670211287
transform -1 0 9968 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spare_logic_const_zero\[11\]
timestamp 1670211287
transform -1 0 3920 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spare_logic_const_zero\[12\]
timestamp 1670211287
transform 1 0 11088 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spare_logic_const_zero\[13\]
timestamp 1670211287
transform -1 0 12432 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spare_logic_const_zero\[14\]
timestamp 1670211287
transform 1 0 8288 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spare_logic_const_zero\[15\]
timestamp 1670211287
transform 1 0 11088 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spare_logic_const_zero\[16\]
timestamp 1670211287
transform 1 0 6272 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spare_logic_const_zero\[17\]
timestamp 1670211287
transform -1 0 12768 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spare_logic_const_zero\[18\]
timestamp 1670211287
transform -1 0 7392 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spare_logic_const_zero\[19\]
timestamp 1670211287
transform -1 0 2464 0 1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spare_logic_const_zero\[20\]
timestamp 1670211287
transform -1 0 9856 0 -1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spare_logic_const_zero\[21\]
timestamp 1670211287
transform 1 0 2016 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spare_logic_const_zero\[22\]
timestamp 1670211287
transform 1 0 6048 0 1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spare_logic_const_zero\[23\]
timestamp 1670211287
transform 1 0 5376 0 1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spare_logic_const_zero\[24\]
timestamp 1670211287
transform 1 0 10640 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spare_logic_const_zero\[25\]
timestamp 1670211287
transform 1 0 5824 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spare_logic_const_zero\[26\]
timestamp 1670211287
transform 1 0 10080 0 -1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrsnq_2  spare_logic_flop\[0\] OpenLane/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1670211287
transform 1 0 1568 0 -1 3136
box -86 -86 4678 870
use gf180mcu_fd_sc_mcu7t5v0__dffrsnq_2  spare_logic_flop\[1\]
timestamp 1670211287
transform 1 0 7728 0 1 3136
box -86 -86 4678 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  spare_logic_inv\[0\] OpenLane/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1670211287
transform -1 0 8400 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  spare_logic_inv\[1\]
timestamp 1670211287
transform -1 0 7504 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  spare_logic_inv\[2\]
timestamp 1670211287
transform 1 0 6720 0 -1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  spare_logic_inv\[3\]
timestamp 1670211287
transform -1 0 7504 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  spare_logic_mux\[0\] OpenLane/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1670211287
transform -1 0 13440 0 -1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  spare_logic_mux\[1\]
timestamp 1670211287
transform 1 0 6720 0 1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  spare_logic_nand\[0\] OpenLane/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1670211287
transform -1 0 2688 0 -1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  spare_logic_nand\[1\]
timestamp 1670211287
transform -1 0 8624 0 -1 3136
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  spare_logic_nor\[0\] OpenLane/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1670211287
transform -1 0 3248 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  spare_logic_nor\[1\]
timestamp 1670211287
transform 1 0 10192 0 -1 7840
box -86 -86 1206 870
<< labels >>
flabel metal4 s 4224 1508 4544 11820 0 FreeSans 1280 90 0 0 VDD
port 0 nsew power bidirectional
flabel metal4 s 7414 1508 7734 11820 0 FreeSans 1280 90 0 0 VDD
port 0 nsew power bidirectional
flabel metal4 s 10604 1508 10924 11820 0 FreeSans 1280 90 0 0 VDD
port 0 nsew power bidirectional
flabel metal5 s 1060 4738 13836 5058 0 FreeSans 2304 0 0 0 VDD
port 0 nsew power bidirectional
flabel metal4 s 5819 1508 6139 11820 0 FreeSans 1280 90 0 0 VSS
port 1 nsew ground bidirectional
flabel metal4 s 9009 1508 9329 11820 0 FreeSans 1280 90 0 0 VSS
port 1 nsew ground bidirectional
flabel metal4 s 12199 1508 12519 11820 0 FreeSans 1280 90 0 0 VSS
port 1 nsew ground bidirectional
flabel metal5 s 1060 6096 13836 6416 0 FreeSans 2304 0 0 0 VSS
port 1 nsew ground bidirectional
flabel metal3 s 0 4704 800 4816 0 FreeSans 448 0 0 0 spare_xfq[0]
port 2 nsew signal tristate
flabel metal2 s 13440 0 13552 800 0 FreeSans 448 90 0 0 spare_xfq[1]
port 3 nsew signal tristate
flabel metal2 s 6720 13200 6832 14000 0 FreeSans 448 90 0 0 spare_xi[0]
port 4 nsew signal tristate
flabel metal2 s 5376 0 5488 800 0 FreeSans 448 90 0 0 spare_xi[1]
port 5 nsew signal tristate
flabel metal3 s 14200 2016 15000 2128 0 FreeSans 448 0 0 0 spare_xi[2]
port 6 nsew signal tristate
flabel metal3 s 0 10080 800 10192 0 FreeSans 448 0 0 0 spare_xi[3]
port 7 nsew signal tristate
flabel metal3 s 14200 672 15000 784 0 FreeSans 448 0 0 0 spare_xib
port 8 nsew signal tristate
flabel metal2 s 14784 0 14896 800 0 FreeSans 448 90 0 0 spare_xmx[0]
port 9 nsew signal tristate
flabel metal3 s 14200 10080 15000 10192 0 FreeSans 448 0 0 0 spare_xmx[1]
port 10 nsew signal tristate
flabel metal2 s 0 13200 112 14000 0 FreeSans 448 90 0 0 spare_xna[0]
port 11 nsew signal tristate
flabel metal2 s 8064 0 8176 800 0 FreeSans 448 90 0 0 spare_xna[1]
port 12 nsew signal tristate
flabel metal3 s 0 3360 800 3472 0 FreeSans 448 0 0 0 spare_xno[0]
port 13 nsew signal tristate
flabel metal2 s 10752 0 10864 800 0 FreeSans 448 90 0 0 spare_xno[1]
port 14 nsew signal tristate
flabel metal3 s 14200 11424 15000 11536 0 FreeSans 448 0 0 0 spare_xz[0]
port 15 nsew signal tristate
flabel metal3 s 0 7392 800 7504 0 FreeSans 448 0 0 0 spare_xz[10]
port 16 nsew signal tristate
flabel metal2 s 2688 0 2800 800 0 FreeSans 448 90 0 0 spare_xz[11]
port 17 nsew signal tristate
flabel metal2 s 13440 13200 13552 14000 0 FreeSans 448 90 0 0 spare_xz[12]
port 18 nsew signal tristate
flabel metal2 s 9408 13200 9520 14000 0 FreeSans 448 90 0 0 spare_xz[13]
port 19 nsew signal tristate
flabel metal3 s 14200 7392 15000 7504 0 FreeSans 448 0 0 0 spare_xz[14]
port 20 nsew signal tristate
flabel metal2 s 12096 13200 12208 14000 0 FreeSans 448 90 0 0 spare_xz[15]
port 21 nsew signal tristate
flabel metal3 s 0 2016 800 2128 0 FreeSans 448 0 0 0 spare_xz[16]
port 22 nsew signal tristate
flabel metal3 s 14200 12768 15000 12880 0 FreeSans 448 0 0 0 spare_xz[17]
port 23 nsew signal tristate
flabel metal2 s 2688 13200 2800 14000 0 FreeSans 448 90 0 0 spare_xz[18]
port 24 nsew signal tristate
flabel metal2 s 0 0 112 800 0 FreeSans 448 90 0 0 spare_xz[19]
port 25 nsew signal tristate
flabel metal2 s 8064 13200 8176 14000 0 FreeSans 448 90 0 0 spare_xz[1]
port 26 nsew signal tristate
flabel metal3 s 14200 8736 15000 8848 0 FreeSans 448 0 0 0 spare_xz[20]
port 27 nsew signal tristate
flabel metal2 s 1344 13200 1456 14000 0 FreeSans 448 90 0 0 spare_xz[21]
port 28 nsew signal tristate
flabel metal3 s 0 672 800 784 0 FreeSans 448 0 0 0 spare_xz[22]
port 29 nsew signal tristate
flabel metal2 s 12096 0 12208 800 0 FreeSans 448 90 0 0 spare_xz[23]
port 30 nsew signal tristate
flabel metal2 s 10752 13200 10864 14000 0 FreeSans 448 90 0 0 spare_xz[24]
port 31 nsew signal tristate
flabel metal3 s 14200 3360 15000 3472 0 FreeSans 448 0 0 0 spare_xz[25]
port 32 nsew signal tristate
flabel metal2 s 1344 0 1456 800 0 FreeSans 448 90 0 0 spare_xz[26]
port 33 nsew signal tristate
flabel metal2 s 4032 0 4144 800 0 FreeSans 448 90 0 0 spare_xz[27]
port 34 nsew signal tristate
flabel metal3 s 0 11424 800 11536 0 FreeSans 448 0 0 0 spare_xz[28]
port 35 nsew signal tristate
flabel metal3 s 14200 4704 15000 4816 0 FreeSans 448 0 0 0 spare_xz[29]
port 36 nsew signal tristate
flabel metal2 s 6720 0 6832 800 0 FreeSans 448 90 0 0 spare_xz[2]
port 37 nsew signal tristate
flabel metal3 s 0 8736 800 8848 0 FreeSans 448 0 0 0 spare_xz[30]
port 38 nsew signal tristate
flabel metal2 s 14784 13200 14896 14000 0 FreeSans 448 90 0 0 spare_xz[3]
port 39 nsew signal tristate
flabel metal2 s 4032 13200 4144 14000 0 FreeSans 448 90 0 0 spare_xz[4]
port 40 nsew signal tristate
flabel metal2 s 5376 13200 5488 14000 0 FreeSans 448 90 0 0 spare_xz[5]
port 41 nsew signal tristate
flabel metal2 s 9408 0 9520 800 0 FreeSans 448 90 0 0 spare_xz[6]
port 42 nsew signal tristate
flabel metal3 s 0 6048 800 6160 0 FreeSans 448 0 0 0 spare_xz[7]
port 43 nsew signal tristate
flabel metal3 s 0 12768 800 12880 0 FreeSans 448 0 0 0 spare_xz[8]
port 44 nsew signal tristate
flabel metal3 s 14200 6048 15000 6160 0 FreeSans 448 0 0 0 spare_xz[9]
port 45 nsew signal tristate
rlabel via1 7448 11760 7448 11760 0 VDD
rlabel metal1 7448 10976 7448 10976 0 VSS
rlabel metal3 4704 2856 4704 2856 0 spare_xfq[0]
rlabel metal2 13496 2142 13496 2142 0 spare_xfq[1]
rlabel metal3 7392 10472 7392 10472 0 spare_xi[0]
rlabel metal2 5432 1414 5432 1414 0 spare_xi[1]
rlabel metal2 7224 2576 7224 2576 0 spare_xi[2]
rlabel metal3 910 10136 910 10136 0 spare_xi[3]
rlabel metal3 10808 6776 10808 6776 0 spare_xib
rlabel metal1 14336 10360 14336 10360 0 spare_xmx[0]
rlabel metal2 7000 8372 7000 8372 0 spare_xmx[1]
rlabel metal3 1008 10808 1008 10808 0 spare_xna[0]
rlabel metal2 8120 1694 8120 1694 0 spare_xna[1]
rlabel metal3 1526 3416 1526 3416 0 spare_xno[0]
rlabel metal2 10808 1470 10808 1470 0 spare_xno[1]
rlabel metal2 8232 10528 8232 10528 0 spare_xz[0]
rlabel metal2 9688 7504 9688 7504 0 spare_xz[10]
rlabel metal2 2744 2198 2744 2198 0 spare_xz[11]
rlabel metal3 11200 8008 11200 8008 0 spare_xz[12]
rlabel metal2 12040 10360 12040 10360 0 spare_xz[13]
rlabel metal2 8120 7896 8120 7896 0 spare_xz[14]
rlabel metal2 11368 10976 11368 10976 0 spare_xz[15]
rlabel metal2 6552 7448 6552 7448 0 spare_xz[16]
rlabel metal2 12488 12040 12488 12040 0 spare_xz[17]
rlabel metal3 4480 7672 4480 7672 0 spare_xz[18]
rlabel metal3 1120 1736 1120 1736 0 spare_xz[19]
rlabel metal2 7896 6720 7896 6720 0 spare_xz[1]
rlabel metal3 9016 3528 9016 3528 0 spare_xz[20]
rlabel metal2 2296 4256 2296 4256 0 spare_xz[21]
rlabel metal3 5992 1736 5992 1736 0 spare_xz[22]
rlabel metal2 6552 4144 6552 4144 0 spare_xz[23]
rlabel metal3 11032 4536 11032 4536 0 spare_xz[24]
rlabel metal2 6944 2072 6944 2072 0 spare_xz[25]
rlabel metal2 1400 2254 1400 2254 0 spare_xz[26]
rlabel metal2 4088 1414 4088 1414 0 spare_xz[27]
rlabel metal3 1470 11480 1470 11480 0 spare_xz[28]
rlabel metal2 12712 4480 12712 4480 0 spare_xz[29]
rlabel metal2 6832 2744 6832 2744 0 spare_xz[2]
rlabel metal3 1470 8792 1470 8792 0 spare_xz[30]
rlabel metal2 7336 10920 7336 10920 0 spare_xz[3]
rlabel metal3 6160 6664 6160 6664 0 spare_xz[4]
rlabel metal2 2408 10360 2408 10360 0 spare_xz[5]
rlabel metal3 9072 1736 9072 1736 0 spare_xz[6]
rlabel metal3 2142 6104 2142 6104 0 spare_xz[7]
rlabel metal2 7896 2856 7896 2856 0 spare_xz[8]
rlabel metal2 3416 4760 3416 4760 0 spare_xz[9]
<< properties >>
string FIXED_BBOX 0 0 15000 14000
<< end >>
