magic
tech gf180mcuC
magscale 1 5
timestamp 1654634570
<< metal5 >>
rect 108 648 216 756
rect 72 612 324 648
rect 36 576 324 612
rect 0 540 324 576
rect 0 432 144 540
rect 0 396 252 432
rect 36 360 288 396
rect 72 324 324 360
rect 180 216 324 324
rect 0 180 324 216
rect 0 144 288 180
rect 0 108 252 144
rect 108 0 216 108
<< properties >>
string FIXED_BBOX 0 -216 432 756
<< end >>
