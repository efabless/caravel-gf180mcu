magic
tech gf180mcuD
magscale 1 10
timestamp 1655304105
<< error_p >>
rect -58 309 -47 355
<< nwell >>
rect -378 -586 368 586
<< mvpmos >>
rect -60 -324 50 276
<< mvpdiff >>
rect -148 263 -60 276
rect -148 -311 -135 263
rect -89 -311 -60 263
rect -148 -324 -60 -311
rect 50 263 138 276
rect 50 -311 79 263
rect 125 -311 138 263
rect 50 -324 138 -311
<< mvpdiffc >>
rect -135 -311 -89 263
rect 79 -311 125 263
<< mvnsubdiff >>
rect -292 428 282 500
rect -292 384 -220 428
rect -292 -384 -279 384
rect -233 -384 -220 384
rect 210 384 282 428
rect -292 -428 -220 -384
rect 210 -384 223 384
rect 269 -384 282 384
rect 210 -428 282 -384
rect -292 -441 282 -428
rect -292 -487 -176 -441
rect 166 -487 282 -441
rect -292 -500 282 -487
<< mvnsubdiffcont >>
rect -279 -384 -233 384
rect 223 -384 269 384
rect -176 -487 166 -441
<< polysilicon >>
rect -60 355 50 368
rect -60 309 -47 355
rect 37 309 50 355
rect -60 276 50 309
rect -60 -368 50 -324
<< polycontact >>
rect -47 309 37 355
<< metal1 >>
rect -279 441 269 487
rect -279 384 -233 441
rect 223 384 269 441
rect -58 309 -47 355
rect 37 309 48 355
rect -135 263 -89 274
rect -135 -322 -89 -311
rect 79 263 125 274
rect 79 -322 125 -311
rect -279 -441 -233 -384
rect 223 -441 269 -384
rect -279 -487 -176 -441
rect 166 -487 269 -441
<< properties >>
string FIXED_BBOX -246 -464 246 464
string gencell pmos_6p0
string library gf180mcu
string parameters w 3.0 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.5 wmin 0.3 full_metal 1 compatible {pmos_3p3 pmos_6p0}
<< end >>
