magic
tech gf180mcuC
magscale 1 5
timestamp 1669656465
<< obsm1 >>
rect 672 1538 61320 76257
<< metal2 >>
rect 1960 77600 2016 78000
rect 2800 77600 2856 78000
rect 3640 77600 3696 78000
rect 4480 77600 4536 78000
rect 5320 77600 5376 78000
rect 6160 77600 6216 78000
rect 7000 77600 7056 78000
rect 7840 77600 7896 78000
rect 8680 77600 8736 78000
rect 9520 77600 9576 78000
rect 10360 77600 10416 78000
rect 11200 77600 11256 78000
rect 12040 77600 12096 78000
rect 12880 77600 12936 78000
rect 13720 77600 13776 78000
rect 14560 77600 14616 78000
rect 15400 77600 15456 78000
rect 16240 77600 16296 78000
rect 17080 77600 17136 78000
rect 17920 77600 17976 78000
rect 18760 77600 18816 78000
rect 19600 77600 19656 78000
rect 20440 77600 20496 78000
rect 21280 77600 21336 78000
rect 22120 77600 22176 78000
rect 22960 77600 23016 78000
rect 23800 77600 23856 78000
rect 24640 77600 24696 78000
rect 25480 77600 25536 78000
rect 26320 77600 26376 78000
rect 27160 77600 27216 78000
rect 28000 77600 28056 78000
rect 28840 77600 28896 78000
rect 29680 77600 29736 78000
rect 30520 77600 30576 78000
rect 31360 77600 31416 78000
rect 32200 77600 32256 78000
rect 33040 77600 33096 78000
rect 33880 77600 33936 78000
rect 34720 77600 34776 78000
rect 35560 77600 35616 78000
rect 36400 77600 36456 78000
rect 37240 77600 37296 78000
rect 38080 77600 38136 78000
rect 38920 77600 38976 78000
rect 39760 77600 39816 78000
rect 40600 77600 40656 78000
rect 41440 77600 41496 78000
rect 42280 77600 42336 78000
rect 43120 77600 43176 78000
rect 43960 77600 44016 78000
rect 44800 77600 44856 78000
rect 45640 77600 45696 78000
rect 46480 77600 46536 78000
rect 47320 77600 47376 78000
rect 48160 77600 48216 78000
rect 49000 77600 49056 78000
rect 49840 77600 49896 78000
rect 50680 77600 50736 78000
rect 51520 77600 51576 78000
rect 52360 77600 52416 78000
rect 53200 77600 53256 78000
rect 54040 77600 54096 78000
rect 54880 77600 54936 78000
rect 55720 77600 55776 78000
rect 56560 77600 56616 78000
rect 57400 77600 57456 78000
rect 58240 77600 58296 78000
rect 59080 77600 59136 78000
rect 59920 77600 59976 78000
rect 1064 0 1120 400
rect 1736 0 1792 400
rect 2408 0 2464 400
rect 3080 0 3136 400
rect 3752 0 3808 400
rect 4424 0 4480 400
rect 5096 0 5152 400
rect 5768 0 5824 400
rect 6440 0 6496 400
rect 7112 0 7168 400
rect 7784 0 7840 400
rect 8456 0 8512 400
rect 9128 0 9184 400
rect 9800 0 9856 400
rect 10472 0 10528 400
rect 11144 0 11200 400
rect 11816 0 11872 400
rect 12488 0 12544 400
rect 13160 0 13216 400
rect 13832 0 13888 400
rect 14504 0 14560 400
rect 15176 0 15232 400
rect 15848 0 15904 400
rect 16520 0 16576 400
rect 17192 0 17248 400
rect 17864 0 17920 400
rect 18536 0 18592 400
rect 19208 0 19264 400
rect 19880 0 19936 400
rect 20552 0 20608 400
rect 21224 0 21280 400
rect 21896 0 21952 400
rect 22568 0 22624 400
rect 23240 0 23296 400
rect 23912 0 23968 400
rect 24584 0 24640 400
rect 25256 0 25312 400
rect 25928 0 25984 400
rect 26600 0 26656 400
rect 27272 0 27328 400
rect 27944 0 28000 400
rect 28616 0 28672 400
rect 29288 0 29344 400
rect 29960 0 30016 400
rect 30632 0 30688 400
rect 31304 0 31360 400
rect 31976 0 32032 400
rect 32648 0 32704 400
rect 33320 0 33376 400
rect 33992 0 34048 400
rect 34664 0 34720 400
rect 35336 0 35392 400
rect 36008 0 36064 400
rect 36680 0 36736 400
rect 37352 0 37408 400
rect 38024 0 38080 400
rect 38696 0 38752 400
rect 39368 0 39424 400
rect 40040 0 40096 400
rect 40712 0 40768 400
rect 41384 0 41440 400
rect 42056 0 42112 400
rect 42728 0 42784 400
rect 43400 0 43456 400
rect 44072 0 44128 400
rect 44744 0 44800 400
rect 45416 0 45472 400
rect 46088 0 46144 400
rect 46760 0 46816 400
rect 47432 0 47488 400
rect 48104 0 48160 400
rect 48776 0 48832 400
rect 49448 0 49504 400
rect 50120 0 50176 400
rect 50792 0 50848 400
rect 51464 0 51520 400
rect 52136 0 52192 400
rect 52808 0 52864 400
rect 53480 0 53536 400
rect 54152 0 54208 400
rect 54824 0 54880 400
rect 55496 0 55552 400
rect 56168 0 56224 400
rect 56840 0 56896 400
rect 57512 0 57568 400
rect 58184 0 58240 400
rect 58856 0 58912 400
rect 59528 0 59584 400
rect 60200 0 60256 400
rect 60872 0 60928 400
<< obsm2 >>
rect 406 77570 1930 77600
rect 2046 77570 2770 77600
rect 2886 77570 3610 77600
rect 3726 77570 4450 77600
rect 4566 77570 5290 77600
rect 5406 77570 6130 77600
rect 6246 77570 6970 77600
rect 7086 77570 7810 77600
rect 7926 77570 8650 77600
rect 8766 77570 9490 77600
rect 9606 77570 10330 77600
rect 10446 77570 11170 77600
rect 11286 77570 12010 77600
rect 12126 77570 12850 77600
rect 12966 77570 13690 77600
rect 13806 77570 14530 77600
rect 14646 77570 15370 77600
rect 15486 77570 16210 77600
rect 16326 77570 17050 77600
rect 17166 77570 17890 77600
rect 18006 77570 18730 77600
rect 18846 77570 19570 77600
rect 19686 77570 20410 77600
rect 20526 77570 21250 77600
rect 21366 77570 22090 77600
rect 22206 77570 22930 77600
rect 23046 77570 23770 77600
rect 23886 77570 24610 77600
rect 24726 77570 25450 77600
rect 25566 77570 26290 77600
rect 26406 77570 27130 77600
rect 27246 77570 27970 77600
rect 28086 77570 28810 77600
rect 28926 77570 29650 77600
rect 29766 77570 30490 77600
rect 30606 77570 31330 77600
rect 31446 77570 32170 77600
rect 32286 77570 33010 77600
rect 33126 77570 33850 77600
rect 33966 77570 34690 77600
rect 34806 77570 35530 77600
rect 35646 77570 36370 77600
rect 36486 77570 37210 77600
rect 37326 77570 38050 77600
rect 38166 77570 38890 77600
rect 39006 77570 39730 77600
rect 39846 77570 40570 77600
rect 40686 77570 41410 77600
rect 41526 77570 42250 77600
rect 42366 77570 43090 77600
rect 43206 77570 43930 77600
rect 44046 77570 44770 77600
rect 44886 77570 45610 77600
rect 45726 77570 46450 77600
rect 46566 77570 47290 77600
rect 47406 77570 48130 77600
rect 48246 77570 48970 77600
rect 49086 77570 49810 77600
rect 49926 77570 50650 77600
rect 50766 77570 51490 77600
rect 51606 77570 52330 77600
rect 52446 77570 53170 77600
rect 53286 77570 54010 77600
rect 54126 77570 54850 77600
rect 54966 77570 55690 77600
rect 55806 77570 56530 77600
rect 56646 77570 57370 77600
rect 57486 77570 58210 77600
rect 58326 77570 59050 77600
rect 59166 77570 59890 77600
rect 60006 77570 61530 77600
rect 406 430 61530 77570
rect 406 350 1034 430
rect 1150 350 1706 430
rect 1822 350 2378 430
rect 2494 350 3050 430
rect 3166 350 3722 430
rect 3838 350 4394 430
rect 4510 350 5066 430
rect 5182 350 5738 430
rect 5854 350 6410 430
rect 6526 350 7082 430
rect 7198 350 7754 430
rect 7870 350 8426 430
rect 8542 350 9098 430
rect 9214 350 9770 430
rect 9886 350 10442 430
rect 10558 350 11114 430
rect 11230 350 11786 430
rect 11902 350 12458 430
rect 12574 350 13130 430
rect 13246 350 13802 430
rect 13918 350 14474 430
rect 14590 350 15146 430
rect 15262 350 15818 430
rect 15934 350 16490 430
rect 16606 350 17162 430
rect 17278 350 17834 430
rect 17950 350 18506 430
rect 18622 350 19178 430
rect 19294 350 19850 430
rect 19966 350 20522 430
rect 20638 350 21194 430
rect 21310 350 21866 430
rect 21982 350 22538 430
rect 22654 350 23210 430
rect 23326 350 23882 430
rect 23998 350 24554 430
rect 24670 350 25226 430
rect 25342 350 25898 430
rect 26014 350 26570 430
rect 26686 350 27242 430
rect 27358 350 27914 430
rect 28030 350 28586 430
rect 28702 350 29258 430
rect 29374 350 29930 430
rect 30046 350 30602 430
rect 30718 350 31274 430
rect 31390 350 31946 430
rect 32062 350 32618 430
rect 32734 350 33290 430
rect 33406 350 33962 430
rect 34078 350 34634 430
rect 34750 350 35306 430
rect 35422 350 35978 430
rect 36094 350 36650 430
rect 36766 350 37322 430
rect 37438 350 37994 430
rect 38110 350 38666 430
rect 38782 350 39338 430
rect 39454 350 40010 430
rect 40126 350 40682 430
rect 40798 350 41354 430
rect 41470 350 42026 430
rect 42142 350 42698 430
rect 42814 350 43370 430
rect 43486 350 44042 430
rect 44158 350 44714 430
rect 44830 350 45386 430
rect 45502 350 46058 430
rect 46174 350 46730 430
rect 46846 350 47402 430
rect 47518 350 48074 430
rect 48190 350 48746 430
rect 48862 350 49418 430
rect 49534 350 50090 430
rect 50206 350 50762 430
rect 50878 350 51434 430
rect 51550 350 52106 430
rect 52222 350 52778 430
rect 52894 350 53450 430
rect 53566 350 54122 430
rect 54238 350 54794 430
rect 54910 350 55466 430
rect 55582 350 56138 430
rect 56254 350 56810 430
rect 56926 350 57482 430
rect 57598 350 58154 430
rect 58270 350 58826 430
rect 58942 350 59498 430
rect 59614 350 60170 430
rect 60286 350 60842 430
rect 60958 350 61530 430
<< metal3 >>
rect 61600 76608 62000 76664
rect 0 75600 400 75656
rect 61600 75432 62000 75488
rect 0 74984 400 75040
rect 0 74368 400 74424
rect 61600 74256 62000 74312
rect 0 73752 400 73808
rect 0 73136 400 73192
rect 61600 73080 62000 73136
rect 0 72520 400 72576
rect 0 71904 400 71960
rect 61600 71904 62000 71960
rect 0 71288 400 71344
rect 0 70672 400 70728
rect 61600 70728 62000 70784
rect 0 70056 400 70112
rect 61600 69552 62000 69608
rect 0 69440 400 69496
rect 0 68824 400 68880
rect 61600 68376 62000 68432
rect 0 68208 400 68264
rect 0 67592 400 67648
rect 61600 67200 62000 67256
rect 0 66976 400 67032
rect 0 66360 400 66416
rect 61600 66024 62000 66080
rect 0 65744 400 65800
rect 0 65128 400 65184
rect 61600 64848 62000 64904
rect 0 64512 400 64568
rect 0 63896 400 63952
rect 61600 63672 62000 63728
rect 0 63280 400 63336
rect 0 62664 400 62720
rect 61600 62496 62000 62552
rect 0 62048 400 62104
rect 0 61432 400 61488
rect 61600 61320 62000 61376
rect 0 60816 400 60872
rect 0 60200 400 60256
rect 61600 60144 62000 60200
rect 0 59584 400 59640
rect 0 58968 400 59024
rect 61600 58968 62000 59024
rect 0 58352 400 58408
rect 0 57736 400 57792
rect 61600 57792 62000 57848
rect 0 57120 400 57176
rect 61600 56616 62000 56672
rect 0 56504 400 56560
rect 0 55888 400 55944
rect 61600 55440 62000 55496
rect 0 55272 400 55328
rect 0 54656 400 54712
rect 61600 54264 62000 54320
rect 0 54040 400 54096
rect 0 53424 400 53480
rect 61600 53088 62000 53144
rect 0 52808 400 52864
rect 0 52192 400 52248
rect 61600 51912 62000 51968
rect 0 51576 400 51632
rect 0 50960 400 51016
rect 61600 50736 62000 50792
rect 0 50344 400 50400
rect 0 49728 400 49784
rect 61600 49560 62000 49616
rect 0 49112 400 49168
rect 0 48496 400 48552
rect 61600 48384 62000 48440
rect 0 47880 400 47936
rect 0 47264 400 47320
rect 61600 47208 62000 47264
rect 0 46648 400 46704
rect 0 46032 400 46088
rect 61600 46032 62000 46088
rect 0 45416 400 45472
rect 0 44800 400 44856
rect 61600 44856 62000 44912
rect 0 44184 400 44240
rect 61600 43680 62000 43736
rect 0 43568 400 43624
rect 0 42952 400 43008
rect 61600 42504 62000 42560
rect 0 42336 400 42392
rect 0 41720 400 41776
rect 61600 41328 62000 41384
rect 0 41104 400 41160
rect 0 40488 400 40544
rect 61600 40152 62000 40208
rect 0 39872 400 39928
rect 0 39256 400 39312
rect 61600 38976 62000 39032
rect 0 38640 400 38696
rect 0 38024 400 38080
rect 61600 37800 62000 37856
rect 0 37408 400 37464
rect 0 36792 400 36848
rect 61600 36624 62000 36680
rect 0 36176 400 36232
rect 0 35560 400 35616
rect 61600 35448 62000 35504
rect 0 34944 400 35000
rect 0 34328 400 34384
rect 61600 34272 62000 34328
rect 0 33712 400 33768
rect 0 33096 400 33152
rect 61600 33096 62000 33152
rect 0 32480 400 32536
rect 0 31864 400 31920
rect 61600 31920 62000 31976
rect 0 31248 400 31304
rect 61600 30744 62000 30800
rect 0 30632 400 30688
rect 0 30016 400 30072
rect 61600 29568 62000 29624
rect 0 29400 400 29456
rect 0 28784 400 28840
rect 61600 28392 62000 28448
rect 0 28168 400 28224
rect 0 27552 400 27608
rect 61600 27216 62000 27272
rect 0 26936 400 26992
rect 0 26320 400 26376
rect 61600 26040 62000 26096
rect 0 25704 400 25760
rect 0 25088 400 25144
rect 61600 24864 62000 24920
rect 0 24472 400 24528
rect 0 23856 400 23912
rect 61600 23688 62000 23744
rect 0 23240 400 23296
rect 0 22624 400 22680
rect 61600 22512 62000 22568
rect 0 22008 400 22064
rect 0 21392 400 21448
rect 61600 21336 62000 21392
rect 0 20776 400 20832
rect 0 20160 400 20216
rect 61600 20160 62000 20216
rect 0 19544 400 19600
rect 0 18928 400 18984
rect 61600 18984 62000 19040
rect 0 18312 400 18368
rect 61600 17808 62000 17864
rect 0 17696 400 17752
rect 0 17080 400 17136
rect 61600 16632 62000 16688
rect 0 16464 400 16520
rect 0 15848 400 15904
rect 61600 15456 62000 15512
rect 0 15232 400 15288
rect 0 14616 400 14672
rect 61600 14280 62000 14336
rect 0 14000 400 14056
rect 0 13384 400 13440
rect 61600 13104 62000 13160
rect 0 12768 400 12824
rect 0 12152 400 12208
rect 61600 11928 62000 11984
rect 0 11536 400 11592
rect 0 10920 400 10976
rect 61600 10752 62000 10808
rect 0 10304 400 10360
rect 0 9688 400 9744
rect 61600 9576 62000 9632
rect 0 9072 400 9128
rect 0 8456 400 8512
rect 61600 8400 62000 8456
rect 0 7840 400 7896
rect 0 7224 400 7280
rect 61600 7224 62000 7280
rect 0 6608 400 6664
rect 0 5992 400 6048
rect 61600 6048 62000 6104
rect 0 5376 400 5432
rect 61600 4872 62000 4928
rect 0 4760 400 4816
rect 0 4144 400 4200
rect 61600 3696 62000 3752
rect 0 3528 400 3584
rect 0 2912 400 2968
rect 61600 2520 62000 2576
rect 0 2296 400 2352
rect 61600 1344 62000 1400
<< obsm3 >>
rect 350 76578 61570 76650
rect 350 75686 61642 76578
rect 430 75570 61642 75686
rect 350 75518 61642 75570
rect 350 75402 61570 75518
rect 350 75070 61642 75402
rect 430 74954 61642 75070
rect 350 74454 61642 74954
rect 430 74342 61642 74454
rect 430 74338 61570 74342
rect 350 74226 61570 74338
rect 350 73838 61642 74226
rect 430 73722 61642 73838
rect 350 73222 61642 73722
rect 430 73166 61642 73222
rect 430 73106 61570 73166
rect 350 73050 61570 73106
rect 350 72606 61642 73050
rect 430 72490 61642 72606
rect 350 71990 61642 72490
rect 430 71874 61570 71990
rect 350 71374 61642 71874
rect 430 71258 61642 71374
rect 350 70814 61642 71258
rect 350 70758 61570 70814
rect 430 70698 61570 70758
rect 430 70642 61642 70698
rect 350 70142 61642 70642
rect 430 70026 61642 70142
rect 350 69638 61642 70026
rect 350 69526 61570 69638
rect 430 69522 61570 69526
rect 430 69410 61642 69522
rect 350 68910 61642 69410
rect 430 68794 61642 68910
rect 350 68462 61642 68794
rect 350 68346 61570 68462
rect 350 68294 61642 68346
rect 430 68178 61642 68294
rect 350 67678 61642 68178
rect 430 67562 61642 67678
rect 350 67286 61642 67562
rect 350 67170 61570 67286
rect 350 67062 61642 67170
rect 430 66946 61642 67062
rect 350 66446 61642 66946
rect 430 66330 61642 66446
rect 350 66110 61642 66330
rect 350 65994 61570 66110
rect 350 65830 61642 65994
rect 430 65714 61642 65830
rect 350 65214 61642 65714
rect 430 65098 61642 65214
rect 350 64934 61642 65098
rect 350 64818 61570 64934
rect 350 64598 61642 64818
rect 430 64482 61642 64598
rect 350 63982 61642 64482
rect 430 63866 61642 63982
rect 350 63758 61642 63866
rect 350 63642 61570 63758
rect 350 63366 61642 63642
rect 430 63250 61642 63366
rect 350 62750 61642 63250
rect 430 62634 61642 62750
rect 350 62582 61642 62634
rect 350 62466 61570 62582
rect 350 62134 61642 62466
rect 430 62018 61642 62134
rect 350 61518 61642 62018
rect 430 61406 61642 61518
rect 430 61402 61570 61406
rect 350 61290 61570 61402
rect 350 60902 61642 61290
rect 430 60786 61642 60902
rect 350 60286 61642 60786
rect 430 60230 61642 60286
rect 430 60170 61570 60230
rect 350 60114 61570 60170
rect 350 59670 61642 60114
rect 430 59554 61642 59670
rect 350 59054 61642 59554
rect 430 58938 61570 59054
rect 350 58438 61642 58938
rect 430 58322 61642 58438
rect 350 57878 61642 58322
rect 350 57822 61570 57878
rect 430 57762 61570 57822
rect 430 57706 61642 57762
rect 350 57206 61642 57706
rect 430 57090 61642 57206
rect 350 56702 61642 57090
rect 350 56590 61570 56702
rect 430 56586 61570 56590
rect 430 56474 61642 56586
rect 350 55974 61642 56474
rect 430 55858 61642 55974
rect 350 55526 61642 55858
rect 350 55410 61570 55526
rect 350 55358 61642 55410
rect 430 55242 61642 55358
rect 350 54742 61642 55242
rect 430 54626 61642 54742
rect 350 54350 61642 54626
rect 350 54234 61570 54350
rect 350 54126 61642 54234
rect 430 54010 61642 54126
rect 350 53510 61642 54010
rect 430 53394 61642 53510
rect 350 53174 61642 53394
rect 350 53058 61570 53174
rect 350 52894 61642 53058
rect 430 52778 61642 52894
rect 350 52278 61642 52778
rect 430 52162 61642 52278
rect 350 51998 61642 52162
rect 350 51882 61570 51998
rect 350 51662 61642 51882
rect 430 51546 61642 51662
rect 350 51046 61642 51546
rect 430 50930 61642 51046
rect 350 50822 61642 50930
rect 350 50706 61570 50822
rect 350 50430 61642 50706
rect 430 50314 61642 50430
rect 350 49814 61642 50314
rect 430 49698 61642 49814
rect 350 49646 61642 49698
rect 350 49530 61570 49646
rect 350 49198 61642 49530
rect 430 49082 61642 49198
rect 350 48582 61642 49082
rect 430 48470 61642 48582
rect 430 48466 61570 48470
rect 350 48354 61570 48466
rect 350 47966 61642 48354
rect 430 47850 61642 47966
rect 350 47350 61642 47850
rect 430 47294 61642 47350
rect 430 47234 61570 47294
rect 350 47178 61570 47234
rect 350 46734 61642 47178
rect 430 46618 61642 46734
rect 350 46118 61642 46618
rect 430 46002 61570 46118
rect 350 45502 61642 46002
rect 430 45386 61642 45502
rect 350 44942 61642 45386
rect 350 44886 61570 44942
rect 430 44826 61570 44886
rect 430 44770 61642 44826
rect 350 44270 61642 44770
rect 430 44154 61642 44270
rect 350 43766 61642 44154
rect 350 43654 61570 43766
rect 430 43650 61570 43654
rect 430 43538 61642 43650
rect 350 43038 61642 43538
rect 430 42922 61642 43038
rect 350 42590 61642 42922
rect 350 42474 61570 42590
rect 350 42422 61642 42474
rect 430 42306 61642 42422
rect 350 41806 61642 42306
rect 430 41690 61642 41806
rect 350 41414 61642 41690
rect 350 41298 61570 41414
rect 350 41190 61642 41298
rect 430 41074 61642 41190
rect 350 40574 61642 41074
rect 430 40458 61642 40574
rect 350 40238 61642 40458
rect 350 40122 61570 40238
rect 350 39958 61642 40122
rect 430 39842 61642 39958
rect 350 39342 61642 39842
rect 430 39226 61642 39342
rect 350 39062 61642 39226
rect 350 38946 61570 39062
rect 350 38726 61642 38946
rect 430 38610 61642 38726
rect 350 38110 61642 38610
rect 430 37994 61642 38110
rect 350 37886 61642 37994
rect 350 37770 61570 37886
rect 350 37494 61642 37770
rect 430 37378 61642 37494
rect 350 36878 61642 37378
rect 430 36762 61642 36878
rect 350 36710 61642 36762
rect 350 36594 61570 36710
rect 350 36262 61642 36594
rect 430 36146 61642 36262
rect 350 35646 61642 36146
rect 430 35534 61642 35646
rect 430 35530 61570 35534
rect 350 35418 61570 35530
rect 350 35030 61642 35418
rect 430 34914 61642 35030
rect 350 34414 61642 34914
rect 430 34358 61642 34414
rect 430 34298 61570 34358
rect 350 34242 61570 34298
rect 350 33798 61642 34242
rect 430 33682 61642 33798
rect 350 33182 61642 33682
rect 430 33066 61570 33182
rect 350 32566 61642 33066
rect 430 32450 61642 32566
rect 350 32006 61642 32450
rect 350 31950 61570 32006
rect 430 31890 61570 31950
rect 430 31834 61642 31890
rect 350 31334 61642 31834
rect 430 31218 61642 31334
rect 350 30830 61642 31218
rect 350 30718 61570 30830
rect 430 30714 61570 30718
rect 430 30602 61642 30714
rect 350 30102 61642 30602
rect 430 29986 61642 30102
rect 350 29654 61642 29986
rect 350 29538 61570 29654
rect 350 29486 61642 29538
rect 430 29370 61642 29486
rect 350 28870 61642 29370
rect 430 28754 61642 28870
rect 350 28478 61642 28754
rect 350 28362 61570 28478
rect 350 28254 61642 28362
rect 430 28138 61642 28254
rect 350 27638 61642 28138
rect 430 27522 61642 27638
rect 350 27302 61642 27522
rect 350 27186 61570 27302
rect 350 27022 61642 27186
rect 430 26906 61642 27022
rect 350 26406 61642 26906
rect 430 26290 61642 26406
rect 350 26126 61642 26290
rect 350 26010 61570 26126
rect 350 25790 61642 26010
rect 430 25674 61642 25790
rect 350 25174 61642 25674
rect 430 25058 61642 25174
rect 350 24950 61642 25058
rect 350 24834 61570 24950
rect 350 24558 61642 24834
rect 430 24442 61642 24558
rect 350 23942 61642 24442
rect 430 23826 61642 23942
rect 350 23774 61642 23826
rect 350 23658 61570 23774
rect 350 23326 61642 23658
rect 430 23210 61642 23326
rect 350 22710 61642 23210
rect 430 22598 61642 22710
rect 430 22594 61570 22598
rect 350 22482 61570 22594
rect 350 22094 61642 22482
rect 430 21978 61642 22094
rect 350 21478 61642 21978
rect 430 21422 61642 21478
rect 430 21362 61570 21422
rect 350 21306 61570 21362
rect 350 20862 61642 21306
rect 430 20746 61642 20862
rect 350 20246 61642 20746
rect 430 20130 61570 20246
rect 350 19630 61642 20130
rect 430 19514 61642 19630
rect 350 19070 61642 19514
rect 350 19014 61570 19070
rect 430 18954 61570 19014
rect 430 18898 61642 18954
rect 350 18398 61642 18898
rect 430 18282 61642 18398
rect 350 17894 61642 18282
rect 350 17782 61570 17894
rect 430 17778 61570 17782
rect 430 17666 61642 17778
rect 350 17166 61642 17666
rect 430 17050 61642 17166
rect 350 16718 61642 17050
rect 350 16602 61570 16718
rect 350 16550 61642 16602
rect 430 16434 61642 16550
rect 350 15934 61642 16434
rect 430 15818 61642 15934
rect 350 15542 61642 15818
rect 350 15426 61570 15542
rect 350 15318 61642 15426
rect 430 15202 61642 15318
rect 350 14702 61642 15202
rect 430 14586 61642 14702
rect 350 14366 61642 14586
rect 350 14250 61570 14366
rect 350 14086 61642 14250
rect 430 13970 61642 14086
rect 350 13470 61642 13970
rect 430 13354 61642 13470
rect 350 13190 61642 13354
rect 350 13074 61570 13190
rect 350 12854 61642 13074
rect 430 12738 61642 12854
rect 350 12238 61642 12738
rect 430 12122 61642 12238
rect 350 12014 61642 12122
rect 350 11898 61570 12014
rect 350 11622 61642 11898
rect 430 11506 61642 11622
rect 350 11006 61642 11506
rect 430 10890 61642 11006
rect 350 10838 61642 10890
rect 350 10722 61570 10838
rect 350 10390 61642 10722
rect 430 10274 61642 10390
rect 350 9774 61642 10274
rect 430 9662 61642 9774
rect 430 9658 61570 9662
rect 350 9546 61570 9658
rect 350 9158 61642 9546
rect 430 9042 61642 9158
rect 350 8542 61642 9042
rect 430 8486 61642 8542
rect 430 8426 61570 8486
rect 350 8370 61570 8426
rect 350 7926 61642 8370
rect 430 7810 61642 7926
rect 350 7310 61642 7810
rect 430 7194 61570 7310
rect 350 6694 61642 7194
rect 430 6578 61642 6694
rect 350 6134 61642 6578
rect 350 6078 61570 6134
rect 430 6018 61570 6078
rect 430 5962 61642 6018
rect 350 5462 61642 5962
rect 430 5346 61642 5462
rect 350 4958 61642 5346
rect 350 4846 61570 4958
rect 430 4842 61570 4846
rect 430 4730 61642 4842
rect 350 4230 61642 4730
rect 430 4114 61642 4230
rect 350 3782 61642 4114
rect 350 3666 61570 3782
rect 350 3614 61642 3666
rect 430 3498 61642 3614
rect 350 2998 61642 3498
rect 430 2882 61642 2998
rect 350 2606 61642 2882
rect 350 2490 61570 2606
rect 350 2382 61642 2490
rect 430 2266 61642 2382
rect 350 1430 61642 2266
rect 350 1314 61570 1430
rect 350 126 61642 1314
<< metal4 >>
rect -418 478 -258 77138
rect -88 808 72 76808
rect 2224 478 2384 77138
rect 2554 478 2714 77138
rect 9904 478 10064 77138
rect 10234 478 10394 77138
rect 17584 478 17744 77138
rect 17914 478 18074 77138
rect 25264 478 25424 77138
rect 25594 478 25754 77138
rect 32944 478 33104 77138
rect 33274 478 33434 77138
rect 40624 478 40784 77138
rect 40954 478 41114 77138
rect 48304 478 48464 77138
rect 48634 478 48794 77138
rect 55984 478 56144 77138
rect 56314 478 56474 77138
rect 61920 808 62080 76808
rect 62250 478 62410 77138
<< obsm4 >>
rect 742 448 2194 75871
rect 2414 448 2524 75871
rect 2744 448 9874 75871
rect 10094 448 10204 75871
rect 10424 448 17554 75871
rect 17774 448 17884 75871
rect 18104 448 25234 75871
rect 25454 448 25564 75871
rect 25784 448 32914 75871
rect 33134 448 33244 75871
rect 33464 448 40594 75871
rect 40814 448 40924 75871
rect 41144 448 48274 75871
rect 48494 448 48604 75871
rect 48824 448 55954 75871
rect 56174 448 56284 75871
rect 56504 448 61138 75871
rect 742 9 61138 448
<< metal5 >>
rect -418 76978 62410 77138
rect -88 76648 62080 76808
rect -418 74129 62410 74289
rect -418 71129 62410 71289
rect -418 68129 62410 68289
rect -418 65129 62410 65289
rect -418 62129 62410 62289
rect -418 59129 62410 59289
rect -418 56129 62410 56289
rect -418 53129 62410 53289
rect -418 50129 62410 50289
rect -418 47129 62410 47289
rect -418 44129 62410 44289
rect -418 41129 62410 41289
rect -418 38129 62410 38289
rect -418 35129 62410 35289
rect -418 32129 62410 32289
rect -418 29129 62410 29289
rect -418 26129 62410 26289
rect -418 23129 62410 23289
rect -418 20129 62410 20289
rect -418 17129 62410 17289
rect -418 14129 62410 14289
rect -418 11129 62410 11289
rect -418 8129 62410 8289
rect -418 5129 62410 5289
rect -418 2129 62410 2289
rect -88 808 62080 968
rect -418 478 62410 638
<< obsm5 >>
rect 958 68339 61146 69210
rect 958 65339 61146 68079
rect 958 62339 61146 65079
rect 958 59339 61146 62079
rect 958 56339 61146 59079
rect 958 53339 61146 56079
rect 958 50339 61146 53079
rect 958 47339 61146 50079
rect 958 44339 61146 47079
rect 958 41339 61146 44079
rect 958 38339 61146 41079
rect 958 35339 61146 38079
rect 958 32339 61146 35079
rect 958 29339 61146 32079
rect 958 26339 61146 29079
rect 958 23339 61146 26079
rect 958 20339 61146 23079
rect 958 17339 61146 20079
rect 958 14339 61146 17079
rect 958 11339 61146 14079
rect 958 8339 61146 11079
rect 958 5339 61146 8079
rect 958 2339 61146 5079
rect 958 1018 61146 2079
rect 958 688 61146 758
rect 958 6 61146 428
<< labels >>
rlabel metal4 s -88 808 72 76808 4 VDD
port 1 nsew power bidirectional
rlabel metal5 s -88 808 62080 968 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s -88 76648 62080 76808 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 61920 808 62080 76808 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 2224 478 2384 77138 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 9904 478 10064 77138 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 17584 478 17744 77138 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 25264 478 25424 77138 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 32944 478 33104 77138 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 40624 478 40784 77138 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 48304 478 48464 77138 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 55984 478 56144 77138 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s -418 2129 62410 2289 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s -418 8129 62410 8289 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s -418 14129 62410 14289 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s -418 20129 62410 20289 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s -418 26129 62410 26289 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s -418 32129 62410 32289 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s -418 38129 62410 38289 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s -418 44129 62410 44289 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s -418 50129 62410 50289 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s -418 56129 62410 56289 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s -418 62129 62410 62289 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s -418 68129 62410 68289 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s -418 74129 62410 74289 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s -418 478 -258 77138 4 VSS
port 2 nsew ground bidirectional
rlabel metal5 s -418 478 62410 638 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s -418 76978 62410 77138 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 62250 478 62410 77138 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 2554 478 2714 77138 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 10234 478 10394 77138 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 17914 478 18074 77138 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 25594 478 25754 77138 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 33274 478 33434 77138 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 40954 478 41114 77138 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 48634 478 48794 77138 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 56314 478 56474 77138 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s -418 5129 62410 5289 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s -418 11129 62410 11289 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s -418 17129 62410 17289 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s -418 23129 62410 23289 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s -418 29129 62410 29289 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s -418 35129 62410 35289 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s -418 41129 62410 41289 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s -418 47129 62410 47289 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s -418 53129 62410 53289 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s -418 59129 62410 59289 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s -418 65129 62410 65289 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s -418 71129 62410 71289 6 VSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 2296 400 2352 6 debug_in
port 3 nsew signal output
rlabel metal3 s 0 2912 400 2968 6 debug_mode
port 4 nsew signal input
rlabel metal3 s 0 3528 400 3584 6 debug_oeb
port 5 nsew signal input
rlabel metal3 s 0 4144 400 4200 6 debug_out
port 6 nsew signal input
rlabel metal3 s 0 5376 400 5432 6 irq[0]
port 7 nsew signal output
rlabel metal3 s 0 5992 400 6048 6 irq[1]
port 8 nsew signal output
rlabel metal3 s 0 6608 400 6664 6 irq[2]
port 9 nsew signal output
rlabel metal2 s 39368 0 39424 400 6 mask_rev_in[0]
port 10 nsew signal input
rlabel metal2 s 46088 0 46144 400 6 mask_rev_in[10]
port 11 nsew signal input
rlabel metal2 s 46760 0 46816 400 6 mask_rev_in[11]
port 12 nsew signal input
rlabel metal2 s 47432 0 47488 400 6 mask_rev_in[12]
port 13 nsew signal input
rlabel metal2 s 48104 0 48160 400 6 mask_rev_in[13]
port 14 nsew signal input
rlabel metal2 s 48776 0 48832 400 6 mask_rev_in[14]
port 15 nsew signal input
rlabel metal2 s 49448 0 49504 400 6 mask_rev_in[15]
port 16 nsew signal input
rlabel metal2 s 50120 0 50176 400 6 mask_rev_in[16]
port 17 nsew signal input
rlabel metal2 s 50792 0 50848 400 6 mask_rev_in[17]
port 18 nsew signal input
rlabel metal2 s 51464 0 51520 400 6 mask_rev_in[18]
port 19 nsew signal input
rlabel metal2 s 52136 0 52192 400 6 mask_rev_in[19]
port 20 nsew signal input
rlabel metal2 s 40040 0 40096 400 6 mask_rev_in[1]
port 21 nsew signal input
rlabel metal2 s 52808 0 52864 400 6 mask_rev_in[20]
port 22 nsew signal input
rlabel metal2 s 53480 0 53536 400 6 mask_rev_in[21]
port 23 nsew signal input
rlabel metal2 s 54152 0 54208 400 6 mask_rev_in[22]
port 24 nsew signal input
rlabel metal2 s 54824 0 54880 400 6 mask_rev_in[23]
port 25 nsew signal input
rlabel metal2 s 55496 0 55552 400 6 mask_rev_in[24]
port 26 nsew signal input
rlabel metal2 s 56168 0 56224 400 6 mask_rev_in[25]
port 27 nsew signal input
rlabel metal2 s 56840 0 56896 400 6 mask_rev_in[26]
port 28 nsew signal input
rlabel metal2 s 57512 0 57568 400 6 mask_rev_in[27]
port 29 nsew signal input
rlabel metal2 s 58184 0 58240 400 6 mask_rev_in[28]
port 30 nsew signal input
rlabel metal2 s 58856 0 58912 400 6 mask_rev_in[29]
port 31 nsew signal input
rlabel metal2 s 40712 0 40768 400 6 mask_rev_in[2]
port 32 nsew signal input
rlabel metal2 s 59528 0 59584 400 6 mask_rev_in[30]
port 33 nsew signal input
rlabel metal2 s 60200 0 60256 400 6 mask_rev_in[31]
port 34 nsew signal input
rlabel metal2 s 41384 0 41440 400 6 mask_rev_in[3]
port 35 nsew signal input
rlabel metal2 s 42056 0 42112 400 6 mask_rev_in[4]
port 36 nsew signal input
rlabel metal2 s 42728 0 42784 400 6 mask_rev_in[5]
port 37 nsew signal input
rlabel metal2 s 43400 0 43456 400 6 mask_rev_in[6]
port 38 nsew signal input
rlabel metal2 s 44072 0 44128 400 6 mask_rev_in[7]
port 39 nsew signal input
rlabel metal2 s 44744 0 44800 400 6 mask_rev_in[8]
port 40 nsew signal input
rlabel metal2 s 45416 0 45472 400 6 mask_rev_in[9]
port 41 nsew signal input
rlabel metal3 s 61600 7224 62000 7280 6 mgmt_gpio_in[0]
port 42 nsew signal input
rlabel metal3 s 61600 42504 62000 42560 6 mgmt_gpio_in[10]
port 43 nsew signal input
rlabel metal3 s 61600 46032 62000 46088 6 mgmt_gpio_in[11]
port 44 nsew signal input
rlabel metal3 s 61600 49560 62000 49616 6 mgmt_gpio_in[12]
port 45 nsew signal input
rlabel metal3 s 61600 53088 62000 53144 6 mgmt_gpio_in[13]
port 46 nsew signal input
rlabel metal3 s 61600 56616 62000 56672 6 mgmt_gpio_in[14]
port 47 nsew signal input
rlabel metal3 s 61600 60144 62000 60200 6 mgmt_gpio_in[15]
port 48 nsew signal input
rlabel metal3 s 61600 63672 62000 63728 6 mgmt_gpio_in[16]
port 49 nsew signal input
rlabel metal3 s 61600 67200 62000 67256 6 mgmt_gpio_in[17]
port 50 nsew signal input
rlabel metal3 s 61600 70728 62000 70784 6 mgmt_gpio_in[18]
port 51 nsew signal input
rlabel metal3 s 61600 74256 62000 74312 6 mgmt_gpio_in[19]
port 52 nsew signal input
rlabel metal3 s 61600 10752 62000 10808 6 mgmt_gpio_in[1]
port 53 nsew signal input
rlabel metal3 s 0 42952 400 43008 6 mgmt_gpio_in[20]
port 54 nsew signal input
rlabel metal3 s 0 44800 400 44856 6 mgmt_gpio_in[21]
port 55 nsew signal input
rlabel metal3 s 0 46648 400 46704 6 mgmt_gpio_in[22]
port 56 nsew signal input
rlabel metal3 s 0 48496 400 48552 6 mgmt_gpio_in[23]
port 57 nsew signal input
rlabel metal3 s 0 50344 400 50400 6 mgmt_gpio_in[24]
port 58 nsew signal input
rlabel metal3 s 0 52192 400 52248 6 mgmt_gpio_in[25]
port 59 nsew signal input
rlabel metal3 s 0 54040 400 54096 6 mgmt_gpio_in[26]
port 60 nsew signal input
rlabel metal3 s 0 55888 400 55944 6 mgmt_gpio_in[27]
port 61 nsew signal input
rlabel metal3 s 0 57736 400 57792 6 mgmt_gpio_in[28]
port 62 nsew signal input
rlabel metal3 s 0 59584 400 59640 6 mgmt_gpio_in[29]
port 63 nsew signal input
rlabel metal3 s 61600 14280 62000 14336 6 mgmt_gpio_in[2]
port 64 nsew signal input
rlabel metal3 s 0 61432 400 61488 6 mgmt_gpio_in[30]
port 65 nsew signal input
rlabel metal3 s 0 63280 400 63336 6 mgmt_gpio_in[31]
port 66 nsew signal input
rlabel metal3 s 0 65128 400 65184 6 mgmt_gpio_in[32]
port 67 nsew signal input
rlabel metal3 s 0 66976 400 67032 6 mgmt_gpio_in[33]
port 68 nsew signal input
rlabel metal3 s 0 68824 400 68880 6 mgmt_gpio_in[34]
port 69 nsew signal input
rlabel metal3 s 0 70672 400 70728 6 mgmt_gpio_in[35]
port 70 nsew signal input
rlabel metal3 s 0 72520 400 72576 6 mgmt_gpio_in[36]
port 71 nsew signal input
rlabel metal3 s 0 74368 400 74424 6 mgmt_gpio_in[37]
port 72 nsew signal input
rlabel metal3 s 61600 17808 62000 17864 6 mgmt_gpio_in[3]
port 73 nsew signal input
rlabel metal3 s 61600 21336 62000 21392 6 mgmt_gpio_in[4]
port 74 nsew signal input
rlabel metal3 s 61600 24864 62000 24920 6 mgmt_gpio_in[5]
port 75 nsew signal input
rlabel metal3 s 61600 28392 62000 28448 6 mgmt_gpio_in[6]
port 76 nsew signal input
rlabel metal3 s 61600 31920 62000 31976 6 mgmt_gpio_in[7]
port 77 nsew signal input
rlabel metal3 s 61600 35448 62000 35504 6 mgmt_gpio_in[8]
port 78 nsew signal input
rlabel metal3 s 61600 38976 62000 39032 6 mgmt_gpio_in[9]
port 79 nsew signal input
rlabel metal3 s 61600 8400 62000 8456 6 mgmt_gpio_oeb[0]
port 80 nsew signal output
rlabel metal3 s 61600 43680 62000 43736 6 mgmt_gpio_oeb[10]
port 81 nsew signal output
rlabel metal3 s 61600 47208 62000 47264 6 mgmt_gpio_oeb[11]
port 82 nsew signal output
rlabel metal3 s 61600 50736 62000 50792 6 mgmt_gpio_oeb[12]
port 83 nsew signal output
rlabel metal3 s 61600 54264 62000 54320 6 mgmt_gpio_oeb[13]
port 84 nsew signal output
rlabel metal3 s 61600 57792 62000 57848 6 mgmt_gpio_oeb[14]
port 85 nsew signal output
rlabel metal3 s 61600 61320 62000 61376 6 mgmt_gpio_oeb[15]
port 86 nsew signal output
rlabel metal3 s 61600 64848 62000 64904 6 mgmt_gpio_oeb[16]
port 87 nsew signal output
rlabel metal3 s 61600 68376 62000 68432 6 mgmt_gpio_oeb[17]
port 88 nsew signal output
rlabel metal3 s 61600 71904 62000 71960 6 mgmt_gpio_oeb[18]
port 89 nsew signal output
rlabel metal3 s 61600 75432 62000 75488 6 mgmt_gpio_oeb[19]
port 90 nsew signal output
rlabel metal3 s 61600 11928 62000 11984 6 mgmt_gpio_oeb[1]
port 91 nsew signal output
rlabel metal3 s 0 43568 400 43624 6 mgmt_gpio_oeb[20]
port 92 nsew signal output
rlabel metal3 s 0 45416 400 45472 6 mgmt_gpio_oeb[21]
port 93 nsew signal output
rlabel metal3 s 0 47264 400 47320 6 mgmt_gpio_oeb[22]
port 94 nsew signal output
rlabel metal3 s 0 49112 400 49168 6 mgmt_gpio_oeb[23]
port 95 nsew signal output
rlabel metal3 s 0 50960 400 51016 6 mgmt_gpio_oeb[24]
port 96 nsew signal output
rlabel metal3 s 0 52808 400 52864 6 mgmt_gpio_oeb[25]
port 97 nsew signal output
rlabel metal3 s 0 54656 400 54712 6 mgmt_gpio_oeb[26]
port 98 nsew signal output
rlabel metal3 s 0 56504 400 56560 6 mgmt_gpio_oeb[27]
port 99 nsew signal output
rlabel metal3 s 0 58352 400 58408 6 mgmt_gpio_oeb[28]
port 100 nsew signal output
rlabel metal3 s 0 60200 400 60256 6 mgmt_gpio_oeb[29]
port 101 nsew signal output
rlabel metal3 s 61600 15456 62000 15512 6 mgmt_gpio_oeb[2]
port 102 nsew signal output
rlabel metal3 s 0 62048 400 62104 6 mgmt_gpio_oeb[30]
port 103 nsew signal output
rlabel metal3 s 0 63896 400 63952 6 mgmt_gpio_oeb[31]
port 104 nsew signal output
rlabel metal3 s 0 65744 400 65800 6 mgmt_gpio_oeb[32]
port 105 nsew signal output
rlabel metal3 s 0 67592 400 67648 6 mgmt_gpio_oeb[33]
port 106 nsew signal output
rlabel metal3 s 0 69440 400 69496 6 mgmt_gpio_oeb[34]
port 107 nsew signal output
rlabel metal3 s 0 71288 400 71344 6 mgmt_gpio_oeb[35]
port 108 nsew signal output
rlabel metal3 s 0 73136 400 73192 6 mgmt_gpio_oeb[36]
port 109 nsew signal output
rlabel metal3 s 0 74984 400 75040 6 mgmt_gpio_oeb[37]
port 110 nsew signal output
rlabel metal3 s 61600 18984 62000 19040 6 mgmt_gpio_oeb[3]
port 111 nsew signal output
rlabel metal3 s 61600 22512 62000 22568 6 mgmt_gpio_oeb[4]
port 112 nsew signal output
rlabel metal3 s 61600 26040 62000 26096 6 mgmt_gpio_oeb[5]
port 113 nsew signal output
rlabel metal3 s 61600 29568 62000 29624 6 mgmt_gpio_oeb[6]
port 114 nsew signal output
rlabel metal3 s 61600 33096 62000 33152 6 mgmt_gpio_oeb[7]
port 115 nsew signal output
rlabel metal3 s 61600 36624 62000 36680 6 mgmt_gpio_oeb[8]
port 116 nsew signal output
rlabel metal3 s 61600 40152 62000 40208 6 mgmt_gpio_oeb[9]
port 117 nsew signal output
rlabel metal3 s 61600 9576 62000 9632 6 mgmt_gpio_out[0]
port 118 nsew signal output
rlabel metal3 s 61600 44856 62000 44912 6 mgmt_gpio_out[10]
port 119 nsew signal output
rlabel metal3 s 61600 48384 62000 48440 6 mgmt_gpio_out[11]
port 120 nsew signal output
rlabel metal3 s 61600 51912 62000 51968 6 mgmt_gpio_out[12]
port 121 nsew signal output
rlabel metal3 s 61600 55440 62000 55496 6 mgmt_gpio_out[13]
port 122 nsew signal output
rlabel metal3 s 61600 58968 62000 59024 6 mgmt_gpio_out[14]
port 123 nsew signal output
rlabel metal3 s 61600 62496 62000 62552 6 mgmt_gpio_out[15]
port 124 nsew signal output
rlabel metal3 s 61600 66024 62000 66080 6 mgmt_gpio_out[16]
port 125 nsew signal output
rlabel metal3 s 61600 69552 62000 69608 6 mgmt_gpio_out[17]
port 126 nsew signal output
rlabel metal3 s 61600 73080 62000 73136 6 mgmt_gpio_out[18]
port 127 nsew signal output
rlabel metal3 s 61600 76608 62000 76664 6 mgmt_gpio_out[19]
port 128 nsew signal output
rlabel metal3 s 61600 13104 62000 13160 6 mgmt_gpio_out[1]
port 129 nsew signal output
rlabel metal3 s 0 44184 400 44240 6 mgmt_gpio_out[20]
port 130 nsew signal output
rlabel metal3 s 0 46032 400 46088 6 mgmt_gpio_out[21]
port 131 nsew signal output
rlabel metal3 s 0 47880 400 47936 6 mgmt_gpio_out[22]
port 132 nsew signal output
rlabel metal3 s 0 49728 400 49784 6 mgmt_gpio_out[23]
port 133 nsew signal output
rlabel metal3 s 0 51576 400 51632 6 mgmt_gpio_out[24]
port 134 nsew signal output
rlabel metal3 s 0 53424 400 53480 6 mgmt_gpio_out[25]
port 135 nsew signal output
rlabel metal3 s 0 55272 400 55328 6 mgmt_gpio_out[26]
port 136 nsew signal output
rlabel metal3 s 0 57120 400 57176 6 mgmt_gpio_out[27]
port 137 nsew signal output
rlabel metal3 s 0 58968 400 59024 6 mgmt_gpio_out[28]
port 138 nsew signal output
rlabel metal3 s 0 60816 400 60872 6 mgmt_gpio_out[29]
port 139 nsew signal output
rlabel metal3 s 61600 16632 62000 16688 6 mgmt_gpio_out[2]
port 140 nsew signal output
rlabel metal3 s 0 62664 400 62720 6 mgmt_gpio_out[30]
port 141 nsew signal output
rlabel metal3 s 0 64512 400 64568 6 mgmt_gpio_out[31]
port 142 nsew signal output
rlabel metal3 s 0 66360 400 66416 6 mgmt_gpio_out[32]
port 143 nsew signal output
rlabel metal3 s 0 68208 400 68264 6 mgmt_gpio_out[33]
port 144 nsew signal output
rlabel metal3 s 0 70056 400 70112 6 mgmt_gpio_out[34]
port 145 nsew signal output
rlabel metal3 s 0 71904 400 71960 6 mgmt_gpio_out[35]
port 146 nsew signal output
rlabel metal3 s 0 73752 400 73808 6 mgmt_gpio_out[36]
port 147 nsew signal output
rlabel metal3 s 0 75600 400 75656 6 mgmt_gpio_out[37]
port 148 nsew signal output
rlabel metal3 s 61600 20160 62000 20216 6 mgmt_gpio_out[3]
port 149 nsew signal output
rlabel metal3 s 61600 23688 62000 23744 6 mgmt_gpio_out[4]
port 150 nsew signal output
rlabel metal3 s 61600 27216 62000 27272 6 mgmt_gpio_out[5]
port 151 nsew signal output
rlabel metal3 s 61600 30744 62000 30800 6 mgmt_gpio_out[6]
port 152 nsew signal output
rlabel metal3 s 61600 34272 62000 34328 6 mgmt_gpio_out[7]
port 153 nsew signal output
rlabel metal3 s 61600 37800 62000 37856 6 mgmt_gpio_out[8]
port 154 nsew signal output
rlabel metal3 s 61600 41328 62000 41384 6 mgmt_gpio_out[9]
port 155 nsew signal output
rlabel metal2 s 1736 0 1792 400 6 pad_flash_clk
port 156 nsew signal output
rlabel metal2 s 2408 0 2464 400 6 pad_flash_clk_oe
port 157 nsew signal output
rlabel metal2 s 3080 0 3136 400 6 pad_flash_csb
port 158 nsew signal output
rlabel metal2 s 3752 0 3808 400 6 pad_flash_csb_oe
port 159 nsew signal output
rlabel metal2 s 4424 0 4480 400 6 pad_flash_io0_di
port 160 nsew signal input
rlabel metal2 s 5096 0 5152 400 6 pad_flash_io0_do
port 161 nsew signal output
rlabel metal2 s 5768 0 5824 400 6 pad_flash_io0_ie
port 162 nsew signal output
rlabel metal2 s 6440 0 6496 400 6 pad_flash_io0_oe
port 163 nsew signal output
rlabel metal2 s 7112 0 7168 400 6 pad_flash_io1_di
port 164 nsew signal input
rlabel metal2 s 7784 0 7840 400 6 pad_flash_io1_do
port 165 nsew signal output
rlabel metal2 s 8456 0 8512 400 6 pad_flash_io1_ie
port 166 nsew signal output
rlabel metal2 s 9128 0 9184 400 6 pad_flash_io1_oe
port 167 nsew signal output
rlabel metal2 s 17864 0 17920 400 6 pll90_sel[0]
port 168 nsew signal output
rlabel metal2 s 18536 0 18592 400 6 pll90_sel[1]
port 169 nsew signal output
rlabel metal2 s 19208 0 19264 400 6 pll90_sel[2]
port 170 nsew signal output
rlabel metal2 s 37352 0 37408 400 6 pll_bypass
port 171 nsew signal output
rlabel metal2 s 11816 0 11872 400 6 pll_dco_ena
port 172 nsew signal output
rlabel metal2 s 12488 0 12544 400 6 pll_div[0]
port 173 nsew signal output
rlabel metal2 s 13160 0 13216 400 6 pll_div[1]
port 174 nsew signal output
rlabel metal2 s 13832 0 13888 400 6 pll_div[2]
port 175 nsew signal output
rlabel metal2 s 14504 0 14560 400 6 pll_div[3]
port 176 nsew signal output
rlabel metal2 s 15176 0 15232 400 6 pll_div[4]
port 177 nsew signal output
rlabel metal2 s 11144 0 11200 400 6 pll_ena
port 178 nsew signal output
rlabel metal2 s 15848 0 15904 400 6 pll_sel[0]
port 179 nsew signal output
rlabel metal2 s 16520 0 16576 400 6 pll_sel[1]
port 180 nsew signal output
rlabel metal2 s 17192 0 17248 400 6 pll_sel[2]
port 181 nsew signal output
rlabel metal2 s 19880 0 19936 400 6 pll_trim[0]
port 182 nsew signal output
rlabel metal2 s 26600 0 26656 400 6 pll_trim[10]
port 183 nsew signal output
rlabel metal2 s 27272 0 27328 400 6 pll_trim[11]
port 184 nsew signal output
rlabel metal2 s 27944 0 28000 400 6 pll_trim[12]
port 185 nsew signal output
rlabel metal2 s 28616 0 28672 400 6 pll_trim[13]
port 186 nsew signal output
rlabel metal2 s 29288 0 29344 400 6 pll_trim[14]
port 187 nsew signal output
rlabel metal2 s 29960 0 30016 400 6 pll_trim[15]
port 188 nsew signal output
rlabel metal2 s 30632 0 30688 400 6 pll_trim[16]
port 189 nsew signal output
rlabel metal2 s 31304 0 31360 400 6 pll_trim[17]
port 190 nsew signal output
rlabel metal2 s 31976 0 32032 400 6 pll_trim[18]
port 191 nsew signal output
rlabel metal2 s 32648 0 32704 400 6 pll_trim[19]
port 192 nsew signal output
rlabel metal2 s 20552 0 20608 400 6 pll_trim[1]
port 193 nsew signal output
rlabel metal2 s 33320 0 33376 400 6 pll_trim[20]
port 194 nsew signal output
rlabel metal2 s 33992 0 34048 400 6 pll_trim[21]
port 195 nsew signal output
rlabel metal2 s 34664 0 34720 400 6 pll_trim[22]
port 196 nsew signal output
rlabel metal2 s 35336 0 35392 400 6 pll_trim[23]
port 197 nsew signal output
rlabel metal2 s 36008 0 36064 400 6 pll_trim[24]
port 198 nsew signal output
rlabel metal2 s 36680 0 36736 400 6 pll_trim[25]
port 199 nsew signal output
rlabel metal2 s 21224 0 21280 400 6 pll_trim[2]
port 200 nsew signal output
rlabel metal2 s 21896 0 21952 400 6 pll_trim[3]
port 201 nsew signal output
rlabel metal2 s 22568 0 22624 400 6 pll_trim[4]
port 202 nsew signal output
rlabel metal2 s 23240 0 23296 400 6 pll_trim[5]
port 203 nsew signal output
rlabel metal2 s 23912 0 23968 400 6 pll_trim[6]
port 204 nsew signal output
rlabel metal2 s 24584 0 24640 400 6 pll_trim[7]
port 205 nsew signal output
rlabel metal2 s 25256 0 25312 400 6 pll_trim[8]
port 206 nsew signal output
rlabel metal2 s 25928 0 25984 400 6 pll_trim[9]
port 207 nsew signal output
rlabel metal2 s 9800 0 9856 400 6 porb
port 208 nsew signal input
rlabel metal2 s 60872 0 60928 400 6 pwr_ctrl_out
port 209 nsew signal output
rlabel metal3 s 0 11536 400 11592 6 qspi_enabled
port 210 nsew signal input
rlabel metal2 s 10472 0 10528 400 6 reset
port 211 nsew signal output
rlabel metal3 s 0 10920 400 10976 6 ser_rx
port 212 nsew signal output
rlabel metal3 s 0 10304 400 10360 6 ser_tx
port 213 nsew signal input
rlabel metal3 s 61600 1344 62000 1400 6 serial_clock
port 214 nsew signal output
rlabel metal3 s 61600 4872 62000 4928 6 serial_data_1
port 215 nsew signal output
rlabel metal3 s 61600 6048 62000 6104 6 serial_data_2
port 216 nsew signal output
rlabel metal3 s 61600 3696 62000 3752 6 serial_load
port 217 nsew signal output
rlabel metal3 s 61600 2520 62000 2576 6 serial_resetn
port 218 nsew signal output
rlabel metal3 s 0 9072 400 9128 6 spi_csb
port 219 nsew signal input
rlabel metal3 s 0 12768 400 12824 6 spi_enabled
port 220 nsew signal input
rlabel metal3 s 0 8456 400 8512 6 spi_sck
port 221 nsew signal input
rlabel metal3 s 0 9688 400 9744 6 spi_sdi
port 222 nsew signal output
rlabel metal3 s 0 7840 400 7896 6 spi_sdo
port 223 nsew signal input
rlabel metal3 s 0 7224 400 7280 6 spi_sdoenb
port 224 nsew signal input
rlabel metal3 s 0 34328 400 34384 6 spimemio_flash_clk
port 225 nsew signal input
rlabel metal3 s 0 34944 400 35000 6 spimemio_flash_csb
port 226 nsew signal input
rlabel metal3 s 0 35560 400 35616 6 spimemio_flash_io0_di
port 227 nsew signal output
rlabel metal3 s 0 36176 400 36232 6 spimemio_flash_io0_do
port 228 nsew signal input
rlabel metal3 s 0 36792 400 36848 6 spimemio_flash_io0_oeb
port 229 nsew signal input
rlabel metal3 s 0 37408 400 37464 6 spimemio_flash_io1_di
port 230 nsew signal output
rlabel metal3 s 0 38024 400 38080 6 spimemio_flash_io1_do
port 231 nsew signal input
rlabel metal3 s 0 38640 400 38696 6 spimemio_flash_io1_oeb
port 232 nsew signal input
rlabel metal3 s 0 39256 400 39312 6 spimemio_flash_io2_di
port 233 nsew signal output
rlabel metal3 s 0 39872 400 39928 6 spimemio_flash_io2_do
port 234 nsew signal input
rlabel metal3 s 0 40488 400 40544 6 spimemio_flash_io2_oeb
port 235 nsew signal input
rlabel metal3 s 0 41104 400 41160 6 spimemio_flash_io3_di
port 236 nsew signal output
rlabel metal3 s 0 41720 400 41776 6 spimemio_flash_io3_do
port 237 nsew signal input
rlabel metal3 s 0 42336 400 42392 6 spimemio_flash_io3_oeb
port 238 nsew signal input
rlabel metal3 s 0 4760 400 4816 6 trap
port 239 nsew signal input
rlabel metal3 s 0 12152 400 12208 6 uart_enabled
port 240 nsew signal input
rlabel metal2 s 1064 0 1120 400 6 user_clock
port 241 nsew signal input
rlabel metal3 s 0 13384 400 13440 6 wb_ack_o
port 242 nsew signal output
rlabel metal2 s 1960 77600 2016 78000 6 wb_adr_i[0]
port 243 nsew signal input
rlabel metal2 s 10360 77600 10416 78000 6 wb_adr_i[10]
port 244 nsew signal input
rlabel metal2 s 11200 77600 11256 78000 6 wb_adr_i[11]
port 245 nsew signal input
rlabel metal2 s 12040 77600 12096 78000 6 wb_adr_i[12]
port 246 nsew signal input
rlabel metal2 s 12880 77600 12936 78000 6 wb_adr_i[13]
port 247 nsew signal input
rlabel metal2 s 13720 77600 13776 78000 6 wb_adr_i[14]
port 248 nsew signal input
rlabel metal2 s 14560 77600 14616 78000 6 wb_adr_i[15]
port 249 nsew signal input
rlabel metal2 s 15400 77600 15456 78000 6 wb_adr_i[16]
port 250 nsew signal input
rlabel metal2 s 16240 77600 16296 78000 6 wb_adr_i[17]
port 251 nsew signal input
rlabel metal2 s 17080 77600 17136 78000 6 wb_adr_i[18]
port 252 nsew signal input
rlabel metal2 s 17920 77600 17976 78000 6 wb_adr_i[19]
port 253 nsew signal input
rlabel metal2 s 2800 77600 2856 78000 6 wb_adr_i[1]
port 254 nsew signal input
rlabel metal2 s 18760 77600 18816 78000 6 wb_adr_i[20]
port 255 nsew signal input
rlabel metal2 s 19600 77600 19656 78000 6 wb_adr_i[21]
port 256 nsew signal input
rlabel metal2 s 20440 77600 20496 78000 6 wb_adr_i[22]
port 257 nsew signal input
rlabel metal2 s 21280 77600 21336 78000 6 wb_adr_i[23]
port 258 nsew signal input
rlabel metal2 s 22120 77600 22176 78000 6 wb_adr_i[24]
port 259 nsew signal input
rlabel metal2 s 22960 77600 23016 78000 6 wb_adr_i[25]
port 260 nsew signal input
rlabel metal2 s 23800 77600 23856 78000 6 wb_adr_i[26]
port 261 nsew signal input
rlabel metal2 s 24640 77600 24696 78000 6 wb_adr_i[27]
port 262 nsew signal input
rlabel metal2 s 25480 77600 25536 78000 6 wb_adr_i[28]
port 263 nsew signal input
rlabel metal2 s 26320 77600 26376 78000 6 wb_adr_i[29]
port 264 nsew signal input
rlabel metal2 s 3640 77600 3696 78000 6 wb_adr_i[2]
port 265 nsew signal input
rlabel metal2 s 27160 77600 27216 78000 6 wb_adr_i[30]
port 266 nsew signal input
rlabel metal2 s 28000 77600 28056 78000 6 wb_adr_i[31]
port 267 nsew signal input
rlabel metal2 s 4480 77600 4536 78000 6 wb_adr_i[3]
port 268 nsew signal input
rlabel metal2 s 5320 77600 5376 78000 6 wb_adr_i[4]
port 269 nsew signal input
rlabel metal2 s 6160 77600 6216 78000 6 wb_adr_i[5]
port 270 nsew signal input
rlabel metal2 s 7000 77600 7056 78000 6 wb_adr_i[6]
port 271 nsew signal input
rlabel metal2 s 7840 77600 7896 78000 6 wb_adr_i[7]
port 272 nsew signal input
rlabel metal2 s 8680 77600 8736 78000 6 wb_adr_i[8]
port 273 nsew signal input
rlabel metal2 s 9520 77600 9576 78000 6 wb_adr_i[9]
port 274 nsew signal input
rlabel metal2 s 38024 0 38080 400 6 wb_clk_i
port 275 nsew signal input
rlabel metal2 s 59920 77600 59976 78000 6 wb_cyc_i
port 276 nsew signal input
rlabel metal2 s 28840 77600 28896 78000 6 wb_dat_i[0]
port 277 nsew signal input
rlabel metal2 s 37240 77600 37296 78000 6 wb_dat_i[10]
port 278 nsew signal input
rlabel metal2 s 38080 77600 38136 78000 6 wb_dat_i[11]
port 279 nsew signal input
rlabel metal2 s 38920 77600 38976 78000 6 wb_dat_i[12]
port 280 nsew signal input
rlabel metal2 s 39760 77600 39816 78000 6 wb_dat_i[13]
port 281 nsew signal input
rlabel metal2 s 40600 77600 40656 78000 6 wb_dat_i[14]
port 282 nsew signal input
rlabel metal2 s 41440 77600 41496 78000 6 wb_dat_i[15]
port 283 nsew signal input
rlabel metal2 s 42280 77600 42336 78000 6 wb_dat_i[16]
port 284 nsew signal input
rlabel metal2 s 43120 77600 43176 78000 6 wb_dat_i[17]
port 285 nsew signal input
rlabel metal2 s 43960 77600 44016 78000 6 wb_dat_i[18]
port 286 nsew signal input
rlabel metal2 s 44800 77600 44856 78000 6 wb_dat_i[19]
port 287 nsew signal input
rlabel metal2 s 29680 77600 29736 78000 6 wb_dat_i[1]
port 288 nsew signal input
rlabel metal2 s 45640 77600 45696 78000 6 wb_dat_i[20]
port 289 nsew signal input
rlabel metal2 s 46480 77600 46536 78000 6 wb_dat_i[21]
port 290 nsew signal input
rlabel metal2 s 47320 77600 47376 78000 6 wb_dat_i[22]
port 291 nsew signal input
rlabel metal2 s 48160 77600 48216 78000 6 wb_dat_i[23]
port 292 nsew signal input
rlabel metal2 s 49000 77600 49056 78000 6 wb_dat_i[24]
port 293 nsew signal input
rlabel metal2 s 49840 77600 49896 78000 6 wb_dat_i[25]
port 294 nsew signal input
rlabel metal2 s 50680 77600 50736 78000 6 wb_dat_i[26]
port 295 nsew signal input
rlabel metal2 s 51520 77600 51576 78000 6 wb_dat_i[27]
port 296 nsew signal input
rlabel metal2 s 52360 77600 52416 78000 6 wb_dat_i[28]
port 297 nsew signal input
rlabel metal2 s 53200 77600 53256 78000 6 wb_dat_i[29]
port 298 nsew signal input
rlabel metal2 s 30520 77600 30576 78000 6 wb_dat_i[2]
port 299 nsew signal input
rlabel metal2 s 54040 77600 54096 78000 6 wb_dat_i[30]
port 300 nsew signal input
rlabel metal2 s 54880 77600 54936 78000 6 wb_dat_i[31]
port 301 nsew signal input
rlabel metal2 s 31360 77600 31416 78000 6 wb_dat_i[3]
port 302 nsew signal input
rlabel metal2 s 32200 77600 32256 78000 6 wb_dat_i[4]
port 303 nsew signal input
rlabel metal2 s 33040 77600 33096 78000 6 wb_dat_i[5]
port 304 nsew signal input
rlabel metal2 s 33880 77600 33936 78000 6 wb_dat_i[6]
port 305 nsew signal input
rlabel metal2 s 34720 77600 34776 78000 6 wb_dat_i[7]
port 306 nsew signal input
rlabel metal2 s 35560 77600 35616 78000 6 wb_dat_i[8]
port 307 nsew signal input
rlabel metal2 s 36400 77600 36456 78000 6 wb_dat_i[9]
port 308 nsew signal input
rlabel metal3 s 0 14616 400 14672 6 wb_dat_o[0]
port 309 nsew signal output
rlabel metal3 s 0 20776 400 20832 6 wb_dat_o[10]
port 310 nsew signal output
rlabel metal3 s 0 21392 400 21448 6 wb_dat_o[11]
port 311 nsew signal output
rlabel metal3 s 0 22008 400 22064 6 wb_dat_o[12]
port 312 nsew signal output
rlabel metal3 s 0 22624 400 22680 6 wb_dat_o[13]
port 313 nsew signal output
rlabel metal3 s 0 23240 400 23296 6 wb_dat_o[14]
port 314 nsew signal output
rlabel metal3 s 0 23856 400 23912 6 wb_dat_o[15]
port 315 nsew signal output
rlabel metal3 s 0 24472 400 24528 6 wb_dat_o[16]
port 316 nsew signal output
rlabel metal3 s 0 25088 400 25144 6 wb_dat_o[17]
port 317 nsew signal output
rlabel metal3 s 0 25704 400 25760 6 wb_dat_o[18]
port 318 nsew signal output
rlabel metal3 s 0 26320 400 26376 6 wb_dat_o[19]
port 319 nsew signal output
rlabel metal3 s 0 15232 400 15288 6 wb_dat_o[1]
port 320 nsew signal output
rlabel metal3 s 0 26936 400 26992 6 wb_dat_o[20]
port 321 nsew signal output
rlabel metal3 s 0 27552 400 27608 6 wb_dat_o[21]
port 322 nsew signal output
rlabel metal3 s 0 28168 400 28224 6 wb_dat_o[22]
port 323 nsew signal output
rlabel metal3 s 0 28784 400 28840 6 wb_dat_o[23]
port 324 nsew signal output
rlabel metal3 s 0 29400 400 29456 6 wb_dat_o[24]
port 325 nsew signal output
rlabel metal3 s 0 30016 400 30072 6 wb_dat_o[25]
port 326 nsew signal output
rlabel metal3 s 0 30632 400 30688 6 wb_dat_o[26]
port 327 nsew signal output
rlabel metal3 s 0 31248 400 31304 6 wb_dat_o[27]
port 328 nsew signal output
rlabel metal3 s 0 31864 400 31920 6 wb_dat_o[28]
port 329 nsew signal output
rlabel metal3 s 0 32480 400 32536 6 wb_dat_o[29]
port 330 nsew signal output
rlabel metal3 s 0 15848 400 15904 6 wb_dat_o[2]
port 331 nsew signal output
rlabel metal3 s 0 33096 400 33152 6 wb_dat_o[30]
port 332 nsew signal output
rlabel metal3 s 0 33712 400 33768 6 wb_dat_o[31]
port 333 nsew signal output
rlabel metal3 s 0 16464 400 16520 6 wb_dat_o[3]
port 334 nsew signal output
rlabel metal3 s 0 17080 400 17136 6 wb_dat_o[4]
port 335 nsew signal output
rlabel metal3 s 0 17696 400 17752 6 wb_dat_o[5]
port 336 nsew signal output
rlabel metal3 s 0 18312 400 18368 6 wb_dat_o[6]
port 337 nsew signal output
rlabel metal3 s 0 18928 400 18984 6 wb_dat_o[7]
port 338 nsew signal output
rlabel metal3 s 0 19544 400 19600 6 wb_dat_o[8]
port 339 nsew signal output
rlabel metal3 s 0 20160 400 20216 6 wb_dat_o[9]
port 340 nsew signal output
rlabel metal2 s 38696 0 38752 400 6 wb_rstn_i
port 341 nsew signal input
rlabel metal2 s 55720 77600 55776 78000 6 wb_sel_i[0]
port 342 nsew signal input
rlabel metal2 s 56560 77600 56616 78000 6 wb_sel_i[1]
port 343 nsew signal input
rlabel metal2 s 57400 77600 57456 78000 6 wb_sel_i[2]
port 344 nsew signal input
rlabel metal2 s 58240 77600 58296 78000 6 wb_sel_i[3]
port 345 nsew signal input
rlabel metal3 s 0 14000 400 14056 6 wb_stb_i
port 346 nsew signal input
rlabel metal2 s 59080 77600 59136 78000 6 wb_we_i
port 347 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 62000 78000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 12152444
string GDS_FILE /home/hosni/GF180/PnR_2/caravel-gf180mcu/openlane/housekeeping/runs/RUN_2022.11.28_17.23.38/results/signoff/housekeeping.magic.gds
string GDS_START 457500
<< end >>

