/* Gate level verilog for user_id_programming */

module user_id_programming(VDD, VSS, mask_rev);
   input VDD;
   input VSS;
   output [31:0] mask_rev;
   wire \user_proj_id_nc[0] ;
   wire \user_proj_id_nc[1] ;
   wire \user_proj_id_nc[2] ;
   wire \user_proj_id_nc[3] ;
   wire \user_proj_id_nc[4] ;
   wire \user_proj_id_nc[5] ;
   wire \user_proj_id_nc[6] ;
   wire \user_proj_id_nc[7] ;
   wire \user_proj_id_nc[8] ;
   wire \user_proj_id_nc[9] ;
   wire \user_proj_id_nc[10] ;
   wire \user_proj_id_nc[11] ;
   wire \user_proj_id_nc[12] ;
   wire \user_proj_id_nc[13] ;
   wire \user_proj_id_nc[14] ;
   wire \user_proj_id_nc[15] ;
   wire \user_proj_id_nc[16] ;
   wire \user_proj_id_nc[17] ;
   wire \user_proj_id_nc[18] ;
   wire \user_proj_id_nc[19] ;
   wire \user_proj_id_nc[20] ;
   wire \user_proj_id_nc[21] ;
   wire \user_proj_id_nc[22] ;
   wire \user_proj_id_nc[23] ;
   wire \user_proj_id_nc[24] ;
   wire \user_proj_id_nc[25] ;
   wire \user_proj_id_nc[26] ;
   wire \user_proj_id_nc[27] ;
   wire \user_proj_id_nc[28] ;
   wire \user_proj_id_nc[29] ;
   wire \user_proj_id_nc[30] ;
   wire \user_proj_id_nc[31] ;

   /* 4 endcaps */
   gf180mcu_fd_sc_mcu7t5v0__endcap ENDCAP_0 (.VDD(VDD), .VSS(VSS));
   gf180mcu_fd_sc_mcu7t5v0__endcap ENDCAP_1 (.VDD(VDD), .VSS(VSS));
   gf180mcu_fd_sc_mcu7t5v0__endcap ENDCAP_2 (.VDD(VDD), .VSS(VSS));
   gf180mcu_fd_sc_mcu7t5v0__endcap ENDCAP_3 (.VDD(VDD), .VSS(VSS));

   /* 14 fillties */
   gf180mcu_fd_sc_mcu7t5v0__filltie FILLTIE_0 (.VDD(VDD), .VSS(VSS));
   gf180mcu_fd_sc_mcu7t5v0__filltie FILLTIE_1 (.VDD(VDD), .VSS(VSS));
   gf180mcu_fd_sc_mcu7t5v0__filltie FILLTIE_2 (.VDD(VDD), .VSS(VSS));
   gf180mcu_fd_sc_mcu7t5v0__filltie FILLTIE_3 (.VDD(VDD), .VSS(VSS));
   gf180mcu_fd_sc_mcu7t5v0__filltie FILLTIE_4 (.VDD(VDD), .VSS(VSS));
   gf180mcu_fd_sc_mcu7t5v0__filltie FILLTIE_5 (.VDD(VDD), .VSS(VSS));
   gf180mcu_fd_sc_mcu7t5v0__filltie FILLTIE_6 (.VDD(VDD), .VSS(VSS));
   gf180mcu_fd_sc_mcu7t5v0__filltie FILLTIE_7 (.VDD(VDD), .VSS(VSS));
   gf180mcu_fd_sc_mcu7t5v0__filltie FILLTIE_8 (.VDD(VDD), .VSS(VSS));
   gf180mcu_fd_sc_mcu7t5v0__filltie FILLTIE_9 (.VDD(VDD), .VSS(VSS));
   gf180mcu_fd_sc_mcu7t5v0__filltie FILLTIE_10 (.VDD(VDD), .VSS(VSS));
   gf180mcu_fd_sc_mcu7t5v0__filltie FILLTIE_11 (.VDD(VDD), .VSS(VSS));
   gf180mcu_fd_sc_mcu7t5v0__filltie FILLTIE_12 (.VDD(VDD), .VSS(VSS));
   gf180mcu_fd_sc_mcu7t5v0__filltie FILLTIE_13 (.VDD(VDD), .VSS(VSS));

   /* 24 fillcap_4s */
   gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLCAP_4_0 (.VDD(VDD),
		.VSS(VSS), .VPW(VSS), .VNW(VDD));
   gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLCAP_4_1 (.VDD(VDD),
		.VSS(VSS), .VPW(VSS), .VNW(VDD));
   gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLCAP_4_2 (.VDD(VDD),
		.VSS(VSS), .VPW(VSS), .VNW(VDD));
   gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLCAP_4_3 (.VDD(VDD),
		.VSS(VSS), .VPW(VSS), .VNW(VDD));
   gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLCAP_4_4 (.VDD(VDD),
		.VSS(VSS), .VPW(VSS), .VNW(VDD));
   gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLCAP_4_5 (.VDD(VDD),
		.VSS(VSS), .VPW(VSS), .VNW(VDD));
   gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLCAP_4_6 (.VDD(VDD),
		.VSS(VSS), .VPW(VSS), .VNW(VDD));
   gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLCAP_4_7 (.VDD(VDD),
		.VSS(VSS), .VPW(VSS), .VNW(VDD));
   gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLCAP_4_8 (.VDD(VDD),
		.VSS(VSS), .VPW(VSS), .VNW(VDD));
   gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLCAP_4_9 (.VDD(VDD),
		.VSS(VSS), .VPW(VSS), .VNW(VDD));
   gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLCAP_4_10 (.VDD(VDD),
		.VSS(VSS), .VPW(VSS), .VNW(VDD));
   gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLCAP_4_11 (.VDD(VDD),
		.VSS(VSS), .VPW(VSS), .VNW(VDD));
   gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLCAP_4_12 (.VDD(VDD),
		.VSS(VSS), .VPW(VSS), .VNW(VDD));
   gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLCAP_4_13 (.VDD(VDD),
		.VSS(VSS), .VPW(VSS), .VNW(VDD));
   gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLCAP_4_14 (.VDD(VDD),
		.VSS(VSS), .VPW(VSS), .VNW(VDD));
   gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLCAP_4_15 (.VDD(VDD),
		.VSS(VSS), .VPW(VSS), .VNW(VDD));
   gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLCAP_4_16 (.VDD(VDD),
		.VSS(VSS), .VPW(VSS), .VNW(VDD));
   gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLCAP_4_17 (.VDD(VDD),
		.VSS(VSS), .VPW(VSS), .VNW(VDD));
   gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLCAP_4_18 (.VDD(VDD),
		.VSS(VSS), .VPW(VSS), .VNW(VDD));
   gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLCAP_4_19 (.VDD(VDD),
		.VSS(VSS), .VPW(VSS), .VNW(VDD));
   gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLCAP_4_20 (.VDD(VDD),
		.VSS(VSS), .VPW(VSS), .VNW(VDD));
   gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLCAP_4_21 (.VDD(VDD),
		.VSS(VSS), .VPW(VSS), .VNW(VDD));
   gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLCAP_4_22 (.VDD(VDD),
		.VSS(VSS), .VPW(VSS), .VNW(VDD));
   gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLCAP_4_23 (.VDD(VDD),
		.VSS(VSS), .VPW(VSS), .VNW(VDD));

   /* 32 tiehs */
   gf180mcu_fd_sc_mcu7t5v0__tieh \mask_rev_value_one[0]  (
	.VDD(VDD), .VSS(VSS), .VPW(VSS), .VNW(VDD),
	.Z(\user_proj_id_nc[0] )
   );
   gf180mcu_fd_sc_mcu7t5v0__tieh \mask_rev_value_one[1]  (
	.VDD(VDD), .VSS(VSS), .VPW(VSS), .VNW(VDD),
	.Z(\user_proj_id_nc[1] )
   );
   gf180mcu_fd_sc_mcu7t5v0__tieh \mask_rev_value_one[2]  (
	.VDD(VDD), .VSS(VSS), .VPW(VSS), .VNW(VDD),
	.Z(\user_proj_id_nc[2] )
   );
   gf180mcu_fd_sc_mcu7t5v0__tieh \mask_rev_value_one[3]  (
	.VDD(VDD), .VSS(VSS), .VPW(VSS), .VNW(VDD),
	.Z(\user_proj_id_nc[3] )
   );
   gf180mcu_fd_sc_mcu7t5v0__tieh \mask_rev_value_one[4]  (
	.VDD(VDD), .VSS(VSS), .VPW(VSS), .VNW(VDD),
	.Z(\user_proj_id_nc[4] )
   );
   gf180mcu_fd_sc_mcu7t5v0__tieh \mask_rev_value_one[5]  (
	.VDD(VDD), .VSS(VSS), .VPW(VSS), .VNW(VDD),
	.Z(\user_proj_id_nc[5] )
   );
   gf180mcu_fd_sc_mcu7t5v0__tieh \mask_rev_value_one[6]  (
	.VDD(VDD), .VSS(VSS), .VPW(VSS), .VNW(VDD),
	.Z(\user_proj_id_nc[6] )
   );
   gf180mcu_fd_sc_mcu7t5v0__tieh \mask_rev_value_one[7]  (
	.VDD(VDD), .VSS(VSS), .VPW(VSS), .VNW(VDD),
	.Z(\user_proj_id_nc[7] )
   );
   gf180mcu_fd_sc_mcu7t5v0__tieh \mask_rev_value_one[8]  (
	.VDD(VDD), .VSS(VSS), .VPW(VSS), .VNW(VDD),
	.Z(\user_proj_id_nc[8] )
   );
   gf180mcu_fd_sc_mcu7t5v0__tieh \mask_rev_value_one[9]  (
	.VDD(VDD), .VSS(VSS), .VPW(VSS), .VNW(VDD),
	.Z(\user_proj_id_nc[9] )
   );
   gf180mcu_fd_sc_mcu7t5v0__tieh \mask_rev_value_one[10]  (
	.VDD(VDD), .VSS(VSS), .VPW(VSS), .VNW(VDD),
	.Z(\user_proj_id_nc[10] )
   );
   gf180mcu_fd_sc_mcu7t5v0__tieh \mask_rev_value_one[11]  (
	.VDD(VDD), .VSS(VSS), .VPW(VSS), .VNW(VDD),
	.Z(\user_proj_id_nc[11] )
   );
   gf180mcu_fd_sc_mcu7t5v0__tieh \mask_rev_value_one[12]  (
	.VDD(VDD), .VSS(VSS), .VPW(VSS), .VNW(VDD),
	.Z(\user_proj_id_nc[12] )
   );
   gf180mcu_fd_sc_mcu7t5v0__tieh \mask_rev_value_one[13]  (
	.VDD(VDD), .VSS(VSS), .VPW(VSS), .VNW(VDD),
	.Z(\user_proj_id_nc[13] )
   );
   gf180mcu_fd_sc_mcu7t5v0__tieh \mask_rev_value_one[14]  (
	.VDD(VDD), .VSS(VSS), .VPW(VSS), .VNW(VDD),
	.Z(\user_proj_id_nc[14] )
   );
   gf180mcu_fd_sc_mcu7t5v0__tieh \mask_rev_value_one[15]  (
	.VDD(VDD), .VSS(VSS), .VPW(VSS), .VNW(VDD),
	.Z(\user_proj_id_nc[15] )
   );
   gf180mcu_fd_sc_mcu7t5v0__tieh \mask_rev_value_one[16]  (
	.VDD(VDD), .VSS(VSS), .VPW(VSS), .VNW(VDD),
	.Z(\user_proj_id_nc[16] )
   );
   gf180mcu_fd_sc_mcu7t5v0__tieh \mask_rev_value_one[17]  (
	.VDD(VDD), .VSS(VSS), .VPW(VSS), .VNW(VDD),
	.Z(\user_proj_id_nc[17] )
   );
   gf180mcu_fd_sc_mcu7t5v0__tieh \mask_rev_value_one[18]  (
	.VDD(VDD), .VSS(VSS), .VPW(VSS), .VNW(VDD),
	.Z(\user_proj_id_nc[18] )
   );
   gf180mcu_fd_sc_mcu7t5v0__tieh \mask_rev_value_one[19]  (
	.VDD(VDD), .VSS(VSS), .VPW(VSS), .VNW(VDD),
	.Z(\user_proj_id_nc[19] )
   );
   gf180mcu_fd_sc_mcu7t5v0__tieh \mask_rev_value_one[20]  (
	.VDD(VDD), .VSS(VSS), .VPW(VSS), .VNW(VDD),
	.Z(\user_proj_id_nc[20] )
   );
   gf180mcu_fd_sc_mcu7t5v0__tieh \mask_rev_value_one[21]  (
	.VDD(VDD), .VSS(VSS), .VPW(VSS), .VNW(VDD),
	.Z(\user_proj_id_nc[21] )
   );
   gf180mcu_fd_sc_mcu7t5v0__tieh \mask_rev_value_one[22]  (
	.VDD(VDD), .VSS(VSS), .VPW(VSS), .VNW(VDD),
	.Z(\user_proj_id_nc[22] )
   );
   gf180mcu_fd_sc_mcu7t5v0__tieh \mask_rev_value_one[23]  (
	.VDD(VDD), .VSS(VSS), .VPW(VSS), .VNW(VDD),
	.Z(\user_proj_id_nc[23] )
   );
   gf180mcu_fd_sc_mcu7t5v0__tieh \mask_rev_value_one[24]  (
	.VDD(VDD), .VSS(VSS), .VPW(VSS), .VNW(VDD),
	.Z(\user_proj_id_nc[24] )
   );
   gf180mcu_fd_sc_mcu7t5v0__tieh \mask_rev_value_one[25]  (
	.VDD(VDD), .VSS(VSS), .VPW(VSS), .VNW(VDD),
	.Z(\user_proj_id_nc[25] )
   );
   gf180mcu_fd_sc_mcu7t5v0__tieh \mask_rev_value_one[26]  (
	.VDD(VDD), .VSS(VSS), .VPW(VSS), .VNW(VDD),
	.Z(\user_proj_id_nc[26] )
   );
   gf180mcu_fd_sc_mcu7t5v0__tieh \mask_rev_value_one[27]  (
	.VDD(VDD), .VSS(VSS), .VPW(VSS), .VNW(VDD),
	.Z(\user_proj_id_nc[27] )
   );
   gf180mcu_fd_sc_mcu7t5v0__tieh \mask_rev_value_one[28]  (
	.VDD(VDD), .VSS(VSS), .VPW(VSS), .VNW(VDD),
	.Z(\user_proj_id_nc[28] )
   );
   gf180mcu_fd_sc_mcu7t5v0__tieh \mask_rev_value_one[29]  (
	.VDD(VDD), .VSS(VSS), .VPW(VSS), .VNW(VDD),
	.Z(\user_proj_id_nc[29] )
   );
   gf180mcu_fd_sc_mcu7t5v0__tieh \mask_rev_value_one[30]  (
	.VDD(VDD), .VSS(VSS), .VPW(VSS), .VNW(VDD),
	.Z(\user_proj_id_nc[30] )
   );
   gf180mcu_fd_sc_mcu7t5v0__tieh \mask_rev_value_one[31]  (
	.VDD(VDD), .VSS(VSS), .VPW(VSS), .VNW(VDD),
	.Z(\user_proj_id_nc[31] )
   );

   /* 32 tiels */
   gf180mcu_fd_sc_mcu7t5v0__tiel \mask_rev_value_zero[0]  (
	.VDD(VDD), .VSS(VSS), .VPW(VSS), .VNW(VDD),
	.ZN(mask_rev[0] )
   );
   gf180mcu_fd_sc_mcu7t5v0__tiel \mask_rev_value_zero[1]  (
	.VDD(VDD), .VSS(VSS), .VPW(VSS), .VNW(VDD),
	.ZN(mask_rev[1] )
   );
   gf180mcu_fd_sc_mcu7t5v0__tiel \mask_rev_value_zero[2]  (
	.VDD(VDD), .VSS(VSS), .VPW(VSS), .VNW(VDD),
	.ZN(mask_rev[2] )
   );
   gf180mcu_fd_sc_mcu7t5v0__tiel \mask_rev_value_zero[3]  (
	.VDD(VDD), .VSS(VSS), .VPW(VSS), .VNW(VDD),
	.ZN(mask_rev[3] )
   );
   gf180mcu_fd_sc_mcu7t5v0__tiel \mask_rev_value_zero[4]  (
	.VDD(VDD), .VSS(VSS), .VPW(VSS), .VNW(VDD),
	.ZN(mask_rev[4] )
   );
   gf180mcu_fd_sc_mcu7t5v0__tiel \mask_rev_value_zero[5]  (
	.VDD(VDD), .VSS(VSS), .VPW(VSS), .VNW(VDD),
	.ZN(mask_rev[5] )
   );
   gf180mcu_fd_sc_mcu7t5v0__tiel \mask_rev_value_zero[6]  (
	.VDD(VDD), .VSS(VSS), .VPW(VSS), .VNW(VDD),
	.ZN(mask_rev[6] )
   );
   gf180mcu_fd_sc_mcu7t5v0__tiel \mask_rev_value_zero[7]  (
	.VDD(VDD), .VSS(VSS), .VPW(VSS), .VNW(VDD),
	.ZN(mask_rev[7] )
   );
   gf180mcu_fd_sc_mcu7t5v0__tiel \mask_rev_value_zero[8]  (
	.VDD(VDD), .VSS(VSS), .VPW(VSS), .VNW(VDD),
	.ZN(mask_rev[8] )
   );
   gf180mcu_fd_sc_mcu7t5v0__tiel \mask_rev_value_zero[9]  (
	.VDD(VDD), .VSS(VSS), .VPW(VSS), .VNW(VDD),
	.ZN(mask_rev[9] )
   );
   gf180mcu_fd_sc_mcu7t5v0__tiel \mask_rev_value_zero[10]  (
	.VDD(VDD), .VSS(VSS), .VPW(VSS), .VNW(VDD),
	.ZN(mask_rev[10] )
   );
   gf180mcu_fd_sc_mcu7t5v0__tiel \mask_rev_value_zero[11]  (
	.VDD(VDD), .VSS(VSS), .VPW(VSS), .VNW(VDD),
	.ZN(mask_rev[11] )
   );
   gf180mcu_fd_sc_mcu7t5v0__tiel \mask_rev_value_zero[12]  (
	.VDD(VDD), .VSS(VSS), .VPW(VSS), .VNW(VDD),
	.ZN(mask_rev[12] )
   );
   gf180mcu_fd_sc_mcu7t5v0__tiel \mask_rev_value_zero[13]  (
	.VDD(VDD), .VSS(VSS), .VPW(VSS), .VNW(VDD),
	.ZN(mask_rev[13] )
   );
   gf180mcu_fd_sc_mcu7t5v0__tiel \mask_rev_value_zero[14]  (
	.VDD(VDD), .VSS(VSS), .VPW(VSS), .VNW(VDD),
	.ZN(mask_rev[14] )
   );
   gf180mcu_fd_sc_mcu7t5v0__tiel \mask_rev_value_zero[15]  (
	.VDD(VDD), .VSS(VSS), .VPW(VSS), .VNW(VDD),
	.ZN(mask_rev[15] )
   );
   gf180mcu_fd_sc_mcu7t5v0__tiel \mask_rev_value_zero[16]  (
	.VDD(VDD), .VSS(VSS), .VPW(VSS), .VNW(VDD),
	.ZN(mask_rev[16] )
   );
   gf180mcu_fd_sc_mcu7t5v0__tiel \mask_rev_value_zero[17]  (
	.VDD(VDD), .VSS(VSS), .VPW(VSS), .VNW(VDD),
	.ZN(mask_rev[17] )
   );
   gf180mcu_fd_sc_mcu7t5v0__tiel \mask_rev_value_zero[18]  (
	.VDD(VDD), .VSS(VSS), .VPW(VSS), .VNW(VDD),
	.ZN(mask_rev[18] )
   );
   gf180mcu_fd_sc_mcu7t5v0__tiel \mask_rev_value_zero[19]  (
	.VDD(VDD), .VSS(VSS), .VPW(VSS), .VNW(VDD),
	.ZN(mask_rev[19] )
   );
   gf180mcu_fd_sc_mcu7t5v0__tiel \mask_rev_value_zero[20]  (
	.VDD(VDD), .VSS(VSS), .VPW(VSS), .VNW(VDD),
	.ZN(mask_rev[20] )
   );
   gf180mcu_fd_sc_mcu7t5v0__tiel \mask_rev_value_zero[21]  (
	.VDD(VDD), .VSS(VSS), .VPW(VSS), .VNW(VDD),
	.ZN(mask_rev[21] )
   );
   gf180mcu_fd_sc_mcu7t5v0__tiel \mask_rev_value_zero[22]  (
	.VDD(VDD), .VSS(VSS), .VPW(VSS), .VNW(VDD),
	.ZN(mask_rev[22] )
   );
   gf180mcu_fd_sc_mcu7t5v0__tiel \mask_rev_value_zero[23]  (
	.VDD(VDD), .VSS(VSS), .VPW(VSS), .VNW(VDD),
	.ZN(mask_rev[23] )
   );
   gf180mcu_fd_sc_mcu7t5v0__tiel \mask_rev_value_zero[24]  (
	.VDD(VDD), .VSS(VSS), .VPW(VSS), .VNW(VDD),
	.ZN(mask_rev[24] )
   );
   gf180mcu_fd_sc_mcu7t5v0__tiel \mask_rev_value_zero[25]  (
	.VDD(VDD), .VSS(VSS), .VPW(VSS), .VNW(VDD),
	.ZN(mask_rev[25] )
   );
   gf180mcu_fd_sc_mcu7t5v0__tiel \mask_rev_value_zero[26]  (
	.VDD(VDD), .VSS(VSS), .VPW(VSS), .VNW(VDD),
	.ZN(mask_rev[26] )
   );
   gf180mcu_fd_sc_mcu7t5v0__tiel \mask_rev_value_zero[27]  (
	.VDD(VDD), .VSS(VSS), .VPW(VSS), .VNW(VDD),
	.ZN(mask_rev[27] )
   );
   gf180mcu_fd_sc_mcu7t5v0__tiel \mask_rev_value_zero[28]  (
	.VDD(VDD), .VSS(VSS), .VPW(VSS), .VNW(VDD),
	.ZN(mask_rev[28] )
   );
   gf180mcu_fd_sc_mcu7t5v0__tiel \mask_rev_value_zero[29]  (
	.VDD(VDD), .VSS(VSS), .VPW(VSS), .VNW(VDD),
	.ZN(mask_rev[29] )
   );
   gf180mcu_fd_sc_mcu7t5v0__tiel \mask_rev_value_zero[30]  (
	.VDD(VDD), .VSS(VSS), .VPW(VSS), .VNW(VDD),
	.ZN(mask_rev[30] )
   );
   gf180mcu_fd_sc_mcu7t5v0__tiel \mask_rev_value_zero[31]  (
	.VDD(VDD), .VSS(VSS), .VPW(VSS), .VNW(VDD),
	.ZN(mask_rev[31] )
   );
endmodule
