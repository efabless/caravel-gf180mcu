magic
tech gf180mcuC
magscale 1 10
timestamp 1670447911
<< fillblock >>
rect 0 0 41440 10810
use alpha_0  alphaX_0 hexdigits
timestamp 1654634570
transform 1 0 36895 0 1 890
box 0 0 3888 9072
use alpha_0  alphaX_1
timestamp 1654634570
transform 1 0 31710 0 1 890
box 0 0 3888 9072
use alpha_0  alphaX_2
timestamp 1654634570
transform 1 0 26585 0 1 890
box 0 0 3888 9072
use alpha_0  alphaX_3
timestamp 1654634570
transform 1 0 21460 0 1 890
box 0 0 3888 9072
use alpha_0  alphaX_4
timestamp 1654634570
transform 1 0 16335 0 1 890
box 0 0 3888 9072
use alpha_0  alphaX_5
timestamp 1654634570
transform 1 0 11210 0 1 890
box 0 0 3888 9072
use alpha_0  alphaX_6
timestamp 1654634570
transform 1 0 6085 0 1 890
box 0 0 3888 9072
use alpha_0  alphaX_7
timestamp 1654634570
transform 1 0 960 0 1 890
box 0 0 3888 9072
<< end >>
