* NGSPICE file created from spare_logic_block.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tieh abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tieh Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrsnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrsnq_2 D RN SETN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_12 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_12 I ZN VDD VSS
.ends

.subckt spare_logic_block VDD VSS spare_xfq[0] spare_xfq[1] spare_xi[0] spare_xi[1]
+ spare_xi[2] spare_xi[3] spare_xib spare_xmx[0] spare_xmx[1] spare_xna[0] spare_xna[1]
+ spare_xno[0] spare_xno[1] spare_xz[0] spare_xz[10] spare_xz[11] spare_xz[12] spare_xz[13]
+ spare_xz[14] spare_xz[15] spare_xz[16] spare_xz[17] spare_xz[18] spare_xz[19] spare_xz[1]
+ spare_xz[20] spare_xz[21] spare_xz[22] spare_xz[23] spare_xz[24] spare_xz[25] spare_xz[26]
+ spare_xz[27] spare_xz[28] spare_xz[29] spare_xz[2] spare_xz[30] spare_xz[3] spare_xz[4]
+ spare_xz[5] spare_xz[6] spare_xz[7] spare_xz[8] spare_xz[9]
XFILLER_3_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xspare_logic_const_one\[1\] spare_xz[28] VDD VSS gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_9_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xspare_logic_const_zero\[12\] spare_xz[12] VDD VSS gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_3_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_12_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xspare_logic_nor\[0\] spare_xz[9] spare_xz[11] spare_xno[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_2_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_12_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xspare_logic_const_zero\[6\] spare_xz[6] VDD VSS gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_11_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xspare_logic_const_zero\[10\] spare_xz[10] VDD VSS gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xspare_logic_const_zero\[4\] spare_xz[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_2_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_1_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xspare_logic_const_zero\[26\] spare_xz[26] VDD VSS gf180mcu_fd_sc_mcu7t5v0__tiel
XPHY_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xspare_logic_const_zero\[19\] spare_xz[19] VDD VSS gf180mcu_fd_sc_mcu7t5v0__tiel
Xspare_logic_const_zero\[2\] spare_xz[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_10_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xspare_logic_flop\[0\] spare_xz[19] spare_xz[25] spare_xz[23] spare_xz[21] spare_xfq[0]
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrsnq_2
Xspare_logic_mux\[1\] spare_xz[14] spare_xz[16] spare_xz[18] spare_xmx[1] VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_5_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_2_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xspare_logic_const_zero\[24\] spare_xz[24] VDD VSS gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_4_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xspare_logic_const_zero\[17\] spare_xz[17] VDD VSS gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_7_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_5 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xspare_logic_inv\[3\] spare_xz[3] spare_xi[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_8_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xspare_logic_const_zero\[0\] spare_xz[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_10_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_5_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xspare_logic_const_zero\[22\] spare_xz[22] VDD VSS gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_10_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_4_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xspare_logic_const_zero\[15\] spare_xz[15] VDD VSS gf180mcu_fd_sc_mcu7t5v0__tiel
Xspare_logic_inv\[1\] spare_xz[1] spare_xi[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_10_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_4_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xspare_logic_const_zero\[9\] spare_xz[9] VDD VSS gf180mcu_fd_sc_mcu7t5v0__tiel
Xspare_logic_nand\[1\] spare_xz[6] spare_xz[8] spare_xna[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_5_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xspare_logic_const_zero\[20\] spare_xz[20] VDD VSS gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_4_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xspare_logic_const_one\[2\] spare_xz[29] VDD VSS gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_7_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xspare_logic_const_zero\[13\] spare_xz[13] VDD VSS gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xspare_logic_nor\[1\] spare_xz[10] spare_xz[12] spare_xno[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_2_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_71 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xspare_logic_const_zero\[7\] spare_xz[7] VDD VSS gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_4_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_12_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xspare_logic_const_one\[0\] spare_xz[27] VDD VSS gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_4_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xspare_logic_const_zero\[11\] spare_xz[11] VDD VSS gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xspare_logic_biginv spare_xz[4] spare_xib VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_12
XFILLER_2_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xspare_logic_const_zero\[5\] spare_xz[5] VDD VSS gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_5_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xspare_logic_const_zero\[3\] spare_xz[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_11_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_2_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xspare_logic_flop\[1\] spare_xz[20] spare_xz[26] spare_xz[24] spare_xz[22] spare_xfq[1]
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrsnq_2
XFILLER_5_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xspare_logic_const_zero\[25\] spare_xz[25] VDD VSS gf180mcu_fd_sc_mcu7t5v0__tiel
XPHY_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_2_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xspare_logic_const_zero\[18\] spare_xz[18] VDD VSS gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_11_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xspare_logic_const_zero\[1\] spare_xz[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_8_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xspare_logic_mux\[0\] spare_xz[13] spare_xz[15] spare_xz[17] spare_xmx[0] VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xspare_logic_const_zero\[23\] spare_xz[23] VDD VSS gf180mcu_fd_sc_mcu7t5v0__tiel
XPHY_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xspare_logic_const_zero\[16\] spare_xz[16] VDD VSS gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_6_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xspare_logic_inv\[2\] spare_xz[2] spare_xi[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_3_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xspare_logic_const_zero\[21\] spare_xz[21] VDD VSS gf180mcu_fd_sc_mcu7t5v0__tiel
Xspare_logic_const_one\[3\] spare_xz[30] VDD VSS gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_6_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xspare_logic_const_zero\[14\] spare_xz[14] VDD VSS gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_12_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_12_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xspare_logic_inv\[0\] spare_xz[0] spare_xi[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_10_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xspare_logic_const_zero\[8\] spare_xz[8] VDD VSS gf180mcu_fd_sc_mcu7t5v0__tiel
Xspare_logic_nand\[0\] spare_xz[5] spare_xz[7] spare_xna[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_3_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_12_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
.ends

