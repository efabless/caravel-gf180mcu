magic
tech gf180mcuC
magscale 1 5
timestamp 1654634570
<< metal5 >>
rect 0 432 108 756
rect 216 432 324 540
rect 0 360 324 432
rect 0 324 288 360
rect 0 216 216 324
rect 0 180 288 216
rect 0 108 324 180
rect 0 0 108 108
rect 216 0 324 108
<< properties >>
string FIXED_BBOX 0 -216 432 756
<< end >>
