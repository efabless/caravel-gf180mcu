magic
tech gf180mcuD
magscale 1 10
timestamp 1655304105
<< pwell >>
rect -12578 -2920 12578 2920
<< mvpsubdiff >>
rect -12492 2821 12492 2834
rect -12492 2775 -12345 2821
rect 12356 2775 12492 2821
rect -12492 2762 12492 2775
rect -12492 2718 -12420 2762
rect -12492 -2718 -12479 2718
rect -12433 -2718 -12420 2718
rect 12420 2718 12492 2762
rect -12492 -2762 -12420 -2718
rect 12420 -2718 12433 2718
rect 12479 -2718 12492 2718
rect 12420 -2762 12492 -2718
rect -12492 -2775 12492 -2762
rect -12492 -2821 -12372 -2775
rect 12329 -2821 12492 -2775
rect -12492 -2834 12492 -2821
<< mvpsubdiffcont >>
rect -12345 2775 12356 2821
rect -12479 -2718 -12433 2718
rect 12433 -2718 12479 2718
rect -12372 -2821 12329 -2775
<< polysilicon >>
rect -12280 2609 -12080 2622
rect -12280 2563 -12267 2609
rect -12093 2563 -12080 2609
rect -12280 2500 -12080 2563
rect -12280 -2563 -12080 -2500
rect -12280 -2609 -12267 -2563
rect -12093 -2609 -12080 -2563
rect -12280 -2622 -12080 -2609
rect -12000 2609 -11800 2622
rect -12000 2563 -11987 2609
rect -11813 2563 -11800 2609
rect -12000 2500 -11800 2563
rect -12000 -2563 -11800 -2500
rect -12000 -2609 -11987 -2563
rect -11813 -2609 -11800 -2563
rect -12000 -2622 -11800 -2609
rect -11720 2609 -11520 2622
rect -11720 2563 -11707 2609
rect -11533 2563 -11520 2609
rect -11720 2500 -11520 2563
rect -11720 -2563 -11520 -2500
rect -11720 -2609 -11707 -2563
rect -11533 -2609 -11520 -2563
rect -11720 -2622 -11520 -2609
rect -11440 2609 -11240 2622
rect -11440 2563 -11427 2609
rect -11253 2563 -11240 2609
rect -11440 2500 -11240 2563
rect -11440 -2563 -11240 -2500
rect -11440 -2609 -11427 -2563
rect -11253 -2609 -11240 -2563
rect -11440 -2622 -11240 -2609
rect -11160 2609 -10960 2622
rect -11160 2563 -11147 2609
rect -10973 2563 -10960 2609
rect -11160 2500 -10960 2563
rect -11160 -2563 -10960 -2500
rect -11160 -2609 -11147 -2563
rect -10973 -2609 -10960 -2563
rect -11160 -2622 -10960 -2609
rect -10880 2609 -10680 2622
rect -10880 2563 -10867 2609
rect -10693 2563 -10680 2609
rect -10880 2500 -10680 2563
rect -10880 -2563 -10680 -2500
rect -10880 -2609 -10867 -2563
rect -10693 -2609 -10680 -2563
rect -10880 -2622 -10680 -2609
rect -10600 2609 -10400 2622
rect -10600 2563 -10587 2609
rect -10413 2563 -10400 2609
rect -10600 2500 -10400 2563
rect -10600 -2563 -10400 -2500
rect -10600 -2609 -10587 -2563
rect -10413 -2609 -10400 -2563
rect -10600 -2622 -10400 -2609
rect -10320 2609 -10120 2622
rect -10320 2563 -10307 2609
rect -10133 2563 -10120 2609
rect -10320 2500 -10120 2563
rect -10320 -2563 -10120 -2500
rect -10320 -2609 -10307 -2563
rect -10133 -2609 -10120 -2563
rect -10320 -2622 -10120 -2609
rect -10040 2609 -9840 2622
rect -10040 2563 -10027 2609
rect -9853 2563 -9840 2609
rect -10040 2500 -9840 2563
rect -10040 -2563 -9840 -2500
rect -10040 -2609 -10027 -2563
rect -9853 -2609 -9840 -2563
rect -10040 -2622 -9840 -2609
rect -9760 2609 -9560 2622
rect -9760 2563 -9747 2609
rect -9573 2563 -9560 2609
rect -9760 2500 -9560 2563
rect -9760 -2563 -9560 -2500
rect -9760 -2609 -9747 -2563
rect -9573 -2609 -9560 -2563
rect -9760 -2622 -9560 -2609
rect -9480 2609 -9280 2622
rect -9480 2563 -9467 2609
rect -9293 2563 -9280 2609
rect -9480 2500 -9280 2563
rect -9480 -2563 -9280 -2500
rect -9480 -2609 -9467 -2563
rect -9293 -2609 -9280 -2563
rect -9480 -2622 -9280 -2609
rect -9200 2609 -9000 2622
rect -9200 2563 -9187 2609
rect -9013 2563 -9000 2609
rect -9200 2500 -9000 2563
rect -9200 -2563 -9000 -2500
rect -9200 -2609 -9187 -2563
rect -9013 -2609 -9000 -2563
rect -9200 -2622 -9000 -2609
rect -8920 2609 -8720 2622
rect -8920 2563 -8907 2609
rect -8733 2563 -8720 2609
rect -8920 2500 -8720 2563
rect -8920 -2563 -8720 -2500
rect -8920 -2609 -8907 -2563
rect -8733 -2609 -8720 -2563
rect -8920 -2622 -8720 -2609
rect -8640 2609 -8440 2622
rect -8640 2563 -8627 2609
rect -8453 2563 -8440 2609
rect -8640 2500 -8440 2563
rect -8640 -2563 -8440 -2500
rect -8640 -2609 -8627 -2563
rect -8453 -2609 -8440 -2563
rect -8640 -2622 -8440 -2609
rect -8360 2609 -8160 2622
rect -8360 2563 -8347 2609
rect -8173 2563 -8160 2609
rect -8360 2500 -8160 2563
rect -8360 -2563 -8160 -2500
rect -8360 -2609 -8347 -2563
rect -8173 -2609 -8160 -2563
rect -8360 -2622 -8160 -2609
rect -8080 2609 -7880 2622
rect -8080 2563 -8067 2609
rect -7893 2563 -7880 2609
rect -8080 2500 -7880 2563
rect -8080 -2563 -7880 -2500
rect -8080 -2609 -8067 -2563
rect -7893 -2609 -7880 -2563
rect -8080 -2622 -7880 -2609
rect -7800 2609 -7600 2622
rect -7800 2563 -7787 2609
rect -7613 2563 -7600 2609
rect -7800 2500 -7600 2563
rect -7800 -2563 -7600 -2500
rect -7800 -2609 -7787 -2563
rect -7613 -2609 -7600 -2563
rect -7800 -2622 -7600 -2609
rect -7520 2609 -7320 2622
rect -7520 2563 -7507 2609
rect -7333 2563 -7320 2609
rect -7520 2500 -7320 2563
rect -7520 -2563 -7320 -2500
rect -7520 -2609 -7507 -2563
rect -7333 -2609 -7320 -2563
rect -7520 -2622 -7320 -2609
rect -7240 2609 -7040 2622
rect -7240 2563 -7227 2609
rect -7053 2563 -7040 2609
rect -7240 2500 -7040 2563
rect -7240 -2563 -7040 -2500
rect -7240 -2609 -7227 -2563
rect -7053 -2609 -7040 -2563
rect -7240 -2622 -7040 -2609
rect -6960 2609 -6760 2622
rect -6960 2563 -6947 2609
rect -6773 2563 -6760 2609
rect -6960 2500 -6760 2563
rect -6960 -2563 -6760 -2500
rect -6960 -2609 -6947 -2563
rect -6773 -2609 -6760 -2563
rect -6960 -2622 -6760 -2609
rect -6680 2609 -6480 2622
rect -6680 2563 -6667 2609
rect -6493 2563 -6480 2609
rect -6680 2500 -6480 2563
rect -6680 -2563 -6480 -2500
rect -6680 -2609 -6667 -2563
rect -6493 -2609 -6480 -2563
rect -6680 -2622 -6480 -2609
rect -6400 2609 -6200 2622
rect -6400 2563 -6387 2609
rect -6213 2563 -6200 2609
rect -6400 2500 -6200 2563
rect -6400 -2563 -6200 -2500
rect -6400 -2609 -6387 -2563
rect -6213 -2609 -6200 -2563
rect -6400 -2622 -6200 -2609
rect -6120 2609 -5920 2622
rect -6120 2563 -6107 2609
rect -5933 2563 -5920 2609
rect -6120 2500 -5920 2563
rect -6120 -2563 -5920 -2500
rect -6120 -2609 -6107 -2563
rect -5933 -2609 -5920 -2563
rect -6120 -2622 -5920 -2609
rect -5840 2609 -5640 2622
rect -5840 2563 -5827 2609
rect -5653 2563 -5640 2609
rect -5840 2500 -5640 2563
rect -5840 -2563 -5640 -2500
rect -5840 -2609 -5827 -2563
rect -5653 -2609 -5640 -2563
rect -5840 -2622 -5640 -2609
rect -5560 2609 -5360 2622
rect -5560 2563 -5547 2609
rect -5373 2563 -5360 2609
rect -5560 2500 -5360 2563
rect -5560 -2563 -5360 -2500
rect -5560 -2609 -5547 -2563
rect -5373 -2609 -5360 -2563
rect -5560 -2622 -5360 -2609
rect -5280 2609 -5080 2622
rect -5280 2563 -5267 2609
rect -5093 2563 -5080 2609
rect -5280 2500 -5080 2563
rect -5280 -2563 -5080 -2500
rect -5280 -2609 -5267 -2563
rect -5093 -2609 -5080 -2563
rect -5280 -2622 -5080 -2609
rect -5000 2609 -4800 2622
rect -5000 2563 -4987 2609
rect -4813 2563 -4800 2609
rect -5000 2500 -4800 2563
rect -5000 -2563 -4800 -2500
rect -5000 -2609 -4987 -2563
rect -4813 -2609 -4800 -2563
rect -5000 -2622 -4800 -2609
rect -4720 2609 -4520 2622
rect -4720 2563 -4707 2609
rect -4533 2563 -4520 2609
rect -4720 2500 -4520 2563
rect -4720 -2563 -4520 -2500
rect -4720 -2609 -4707 -2563
rect -4533 -2609 -4520 -2563
rect -4720 -2622 -4520 -2609
rect -4440 2609 -4240 2622
rect -4440 2563 -4427 2609
rect -4253 2563 -4240 2609
rect -4440 2500 -4240 2563
rect -4440 -2563 -4240 -2500
rect -4440 -2609 -4427 -2563
rect -4253 -2609 -4240 -2563
rect -4440 -2622 -4240 -2609
rect -4160 2609 -3960 2622
rect -4160 2563 -4147 2609
rect -3973 2563 -3960 2609
rect -4160 2500 -3960 2563
rect -4160 -2563 -3960 -2500
rect -4160 -2609 -4147 -2563
rect -3973 -2609 -3960 -2563
rect -4160 -2622 -3960 -2609
rect -3880 2609 -3680 2622
rect -3880 2563 -3867 2609
rect -3693 2563 -3680 2609
rect -3880 2500 -3680 2563
rect -3880 -2563 -3680 -2500
rect -3880 -2609 -3867 -2563
rect -3693 -2609 -3680 -2563
rect -3880 -2622 -3680 -2609
rect -3600 2609 -3400 2622
rect -3600 2563 -3587 2609
rect -3413 2563 -3400 2609
rect -3600 2500 -3400 2563
rect -3600 -2563 -3400 -2500
rect -3600 -2609 -3587 -2563
rect -3413 -2609 -3400 -2563
rect -3600 -2622 -3400 -2609
rect -3320 2609 -3120 2622
rect -3320 2563 -3307 2609
rect -3133 2563 -3120 2609
rect -3320 2500 -3120 2563
rect -3320 -2563 -3120 -2500
rect -3320 -2609 -3307 -2563
rect -3133 -2609 -3120 -2563
rect -3320 -2622 -3120 -2609
rect -3040 2609 -2840 2622
rect -3040 2563 -3027 2609
rect -2853 2563 -2840 2609
rect -3040 2500 -2840 2563
rect -3040 -2563 -2840 -2500
rect -3040 -2609 -3027 -2563
rect -2853 -2609 -2840 -2563
rect -3040 -2622 -2840 -2609
rect -2760 2609 -2560 2622
rect -2760 2563 -2747 2609
rect -2573 2563 -2560 2609
rect -2760 2500 -2560 2563
rect -2760 -2563 -2560 -2500
rect -2760 -2609 -2747 -2563
rect -2573 -2609 -2560 -2563
rect -2760 -2622 -2560 -2609
rect -2480 2609 -2280 2622
rect -2480 2563 -2467 2609
rect -2293 2563 -2280 2609
rect -2480 2500 -2280 2563
rect -2480 -2563 -2280 -2500
rect -2480 -2609 -2467 -2563
rect -2293 -2609 -2280 -2563
rect -2480 -2622 -2280 -2609
rect -2200 2609 -2000 2622
rect -2200 2563 -2187 2609
rect -2013 2563 -2000 2609
rect -2200 2500 -2000 2563
rect -2200 -2563 -2000 -2500
rect -2200 -2609 -2187 -2563
rect -2013 -2609 -2000 -2563
rect -2200 -2622 -2000 -2609
rect -1920 2609 -1720 2622
rect -1920 2563 -1907 2609
rect -1733 2563 -1720 2609
rect -1920 2500 -1720 2563
rect -1920 -2563 -1720 -2500
rect -1920 -2609 -1907 -2563
rect -1733 -2609 -1720 -2563
rect -1920 -2622 -1720 -2609
rect -1640 2609 -1440 2622
rect -1640 2563 -1627 2609
rect -1453 2563 -1440 2609
rect -1640 2500 -1440 2563
rect -1640 -2563 -1440 -2500
rect -1640 -2609 -1627 -2563
rect -1453 -2609 -1440 -2563
rect -1640 -2622 -1440 -2609
rect -1360 2609 -1160 2622
rect -1360 2563 -1347 2609
rect -1173 2563 -1160 2609
rect -1360 2500 -1160 2563
rect -1360 -2563 -1160 -2500
rect -1360 -2609 -1347 -2563
rect -1173 -2609 -1160 -2563
rect -1360 -2622 -1160 -2609
rect -1080 2609 -880 2622
rect -1080 2563 -1067 2609
rect -893 2563 -880 2609
rect -1080 2500 -880 2563
rect -1080 -2563 -880 -2500
rect -1080 -2609 -1067 -2563
rect -893 -2609 -880 -2563
rect -1080 -2622 -880 -2609
rect -800 2609 -600 2622
rect -800 2563 -787 2609
rect -613 2563 -600 2609
rect -800 2500 -600 2563
rect -800 -2563 -600 -2500
rect -800 -2609 -787 -2563
rect -613 -2609 -600 -2563
rect -800 -2622 -600 -2609
rect -520 2609 -320 2622
rect -520 2563 -507 2609
rect -333 2563 -320 2609
rect -520 2500 -320 2563
rect -520 -2563 -320 -2500
rect -520 -2609 -507 -2563
rect -333 -2609 -320 -2563
rect -520 -2622 -320 -2609
rect -240 2609 -40 2622
rect -240 2563 -227 2609
rect -53 2563 -40 2609
rect -240 2500 -40 2563
rect -240 -2563 -40 -2500
rect -240 -2609 -227 -2563
rect -53 -2609 -40 -2563
rect -240 -2622 -40 -2609
rect 40 2609 240 2622
rect 40 2563 53 2609
rect 227 2563 240 2609
rect 40 2500 240 2563
rect 40 -2563 240 -2500
rect 40 -2609 53 -2563
rect 227 -2609 240 -2563
rect 40 -2622 240 -2609
rect 320 2609 520 2622
rect 320 2563 333 2609
rect 507 2563 520 2609
rect 320 2500 520 2563
rect 320 -2563 520 -2500
rect 320 -2609 333 -2563
rect 507 -2609 520 -2563
rect 320 -2622 520 -2609
rect 600 2609 800 2622
rect 600 2563 613 2609
rect 787 2563 800 2609
rect 600 2500 800 2563
rect 600 -2563 800 -2500
rect 600 -2609 613 -2563
rect 787 -2609 800 -2563
rect 600 -2622 800 -2609
rect 880 2609 1080 2622
rect 880 2563 893 2609
rect 1067 2563 1080 2609
rect 880 2500 1080 2563
rect 880 -2563 1080 -2500
rect 880 -2609 893 -2563
rect 1067 -2609 1080 -2563
rect 880 -2622 1080 -2609
rect 1160 2609 1360 2622
rect 1160 2563 1173 2609
rect 1347 2563 1360 2609
rect 1160 2500 1360 2563
rect 1160 -2563 1360 -2500
rect 1160 -2609 1173 -2563
rect 1347 -2609 1360 -2563
rect 1160 -2622 1360 -2609
rect 1440 2609 1640 2622
rect 1440 2563 1453 2609
rect 1627 2563 1640 2609
rect 1440 2500 1640 2563
rect 1440 -2563 1640 -2500
rect 1440 -2609 1453 -2563
rect 1627 -2609 1640 -2563
rect 1440 -2622 1640 -2609
rect 1720 2609 1920 2622
rect 1720 2563 1733 2609
rect 1907 2563 1920 2609
rect 1720 2500 1920 2563
rect 1720 -2563 1920 -2500
rect 1720 -2609 1733 -2563
rect 1907 -2609 1920 -2563
rect 1720 -2622 1920 -2609
rect 2000 2609 2200 2622
rect 2000 2563 2013 2609
rect 2187 2563 2200 2609
rect 2000 2500 2200 2563
rect 2000 -2563 2200 -2500
rect 2000 -2609 2013 -2563
rect 2187 -2609 2200 -2563
rect 2000 -2622 2200 -2609
rect 2280 2609 2480 2622
rect 2280 2563 2293 2609
rect 2467 2563 2480 2609
rect 2280 2500 2480 2563
rect 2280 -2563 2480 -2500
rect 2280 -2609 2293 -2563
rect 2467 -2609 2480 -2563
rect 2280 -2622 2480 -2609
rect 2560 2609 2760 2622
rect 2560 2563 2573 2609
rect 2747 2563 2760 2609
rect 2560 2500 2760 2563
rect 2560 -2563 2760 -2500
rect 2560 -2609 2573 -2563
rect 2747 -2609 2760 -2563
rect 2560 -2622 2760 -2609
rect 2840 2609 3040 2622
rect 2840 2563 2853 2609
rect 3027 2563 3040 2609
rect 2840 2500 3040 2563
rect 2840 -2563 3040 -2500
rect 2840 -2609 2853 -2563
rect 3027 -2609 3040 -2563
rect 2840 -2622 3040 -2609
rect 3120 2609 3320 2622
rect 3120 2563 3133 2609
rect 3307 2563 3320 2609
rect 3120 2500 3320 2563
rect 3120 -2563 3320 -2500
rect 3120 -2609 3133 -2563
rect 3307 -2609 3320 -2563
rect 3120 -2622 3320 -2609
rect 3400 2609 3600 2622
rect 3400 2563 3413 2609
rect 3587 2563 3600 2609
rect 3400 2500 3600 2563
rect 3400 -2563 3600 -2500
rect 3400 -2609 3413 -2563
rect 3587 -2609 3600 -2563
rect 3400 -2622 3600 -2609
rect 3680 2609 3880 2622
rect 3680 2563 3693 2609
rect 3867 2563 3880 2609
rect 3680 2500 3880 2563
rect 3680 -2563 3880 -2500
rect 3680 -2609 3693 -2563
rect 3867 -2609 3880 -2563
rect 3680 -2622 3880 -2609
rect 3960 2609 4160 2622
rect 3960 2563 3973 2609
rect 4147 2563 4160 2609
rect 3960 2500 4160 2563
rect 3960 -2563 4160 -2500
rect 3960 -2609 3973 -2563
rect 4147 -2609 4160 -2563
rect 3960 -2622 4160 -2609
rect 4240 2609 4440 2622
rect 4240 2563 4253 2609
rect 4427 2563 4440 2609
rect 4240 2500 4440 2563
rect 4240 -2563 4440 -2500
rect 4240 -2609 4253 -2563
rect 4427 -2609 4440 -2563
rect 4240 -2622 4440 -2609
rect 4520 2609 4720 2622
rect 4520 2563 4533 2609
rect 4707 2563 4720 2609
rect 4520 2500 4720 2563
rect 4520 -2563 4720 -2500
rect 4520 -2609 4533 -2563
rect 4707 -2609 4720 -2563
rect 4520 -2622 4720 -2609
rect 4800 2609 5000 2622
rect 4800 2563 4813 2609
rect 4987 2563 5000 2609
rect 4800 2500 5000 2563
rect 4800 -2563 5000 -2500
rect 4800 -2609 4813 -2563
rect 4987 -2609 5000 -2563
rect 4800 -2622 5000 -2609
rect 5080 2609 5280 2622
rect 5080 2563 5093 2609
rect 5267 2563 5280 2609
rect 5080 2500 5280 2563
rect 5080 -2563 5280 -2500
rect 5080 -2609 5093 -2563
rect 5267 -2609 5280 -2563
rect 5080 -2622 5280 -2609
rect 5360 2609 5560 2622
rect 5360 2563 5373 2609
rect 5547 2563 5560 2609
rect 5360 2500 5560 2563
rect 5360 -2563 5560 -2500
rect 5360 -2609 5373 -2563
rect 5547 -2609 5560 -2563
rect 5360 -2622 5560 -2609
rect 5640 2609 5840 2622
rect 5640 2563 5653 2609
rect 5827 2563 5840 2609
rect 5640 2500 5840 2563
rect 5640 -2563 5840 -2500
rect 5640 -2609 5653 -2563
rect 5827 -2609 5840 -2563
rect 5640 -2622 5840 -2609
rect 5920 2609 6120 2622
rect 5920 2563 5933 2609
rect 6107 2563 6120 2609
rect 5920 2500 6120 2563
rect 5920 -2563 6120 -2500
rect 5920 -2609 5933 -2563
rect 6107 -2609 6120 -2563
rect 5920 -2622 6120 -2609
rect 6200 2609 6400 2622
rect 6200 2563 6213 2609
rect 6387 2563 6400 2609
rect 6200 2500 6400 2563
rect 6200 -2563 6400 -2500
rect 6200 -2609 6213 -2563
rect 6387 -2609 6400 -2563
rect 6200 -2622 6400 -2609
rect 6480 2609 6680 2622
rect 6480 2563 6493 2609
rect 6667 2563 6680 2609
rect 6480 2500 6680 2563
rect 6480 -2563 6680 -2500
rect 6480 -2609 6493 -2563
rect 6667 -2609 6680 -2563
rect 6480 -2622 6680 -2609
rect 6760 2609 6960 2622
rect 6760 2563 6773 2609
rect 6947 2563 6960 2609
rect 6760 2500 6960 2563
rect 6760 -2563 6960 -2500
rect 6760 -2609 6773 -2563
rect 6947 -2609 6960 -2563
rect 6760 -2622 6960 -2609
rect 7040 2609 7240 2622
rect 7040 2563 7053 2609
rect 7227 2563 7240 2609
rect 7040 2500 7240 2563
rect 7040 -2563 7240 -2500
rect 7040 -2609 7053 -2563
rect 7227 -2609 7240 -2563
rect 7040 -2622 7240 -2609
rect 7320 2609 7520 2622
rect 7320 2563 7333 2609
rect 7507 2563 7520 2609
rect 7320 2500 7520 2563
rect 7320 -2563 7520 -2500
rect 7320 -2609 7333 -2563
rect 7507 -2609 7520 -2563
rect 7320 -2622 7520 -2609
rect 7600 2609 7800 2622
rect 7600 2563 7613 2609
rect 7787 2563 7800 2609
rect 7600 2500 7800 2563
rect 7600 -2563 7800 -2500
rect 7600 -2609 7613 -2563
rect 7787 -2609 7800 -2563
rect 7600 -2622 7800 -2609
rect 7880 2609 8080 2622
rect 7880 2563 7893 2609
rect 8067 2563 8080 2609
rect 7880 2500 8080 2563
rect 7880 -2563 8080 -2500
rect 7880 -2609 7893 -2563
rect 8067 -2609 8080 -2563
rect 7880 -2622 8080 -2609
rect 8160 2609 8360 2622
rect 8160 2563 8173 2609
rect 8347 2563 8360 2609
rect 8160 2500 8360 2563
rect 8160 -2563 8360 -2500
rect 8160 -2609 8173 -2563
rect 8347 -2609 8360 -2563
rect 8160 -2622 8360 -2609
rect 8440 2609 8640 2622
rect 8440 2563 8453 2609
rect 8627 2563 8640 2609
rect 8440 2500 8640 2563
rect 8440 -2563 8640 -2500
rect 8440 -2609 8453 -2563
rect 8627 -2609 8640 -2563
rect 8440 -2622 8640 -2609
rect 8720 2609 8920 2622
rect 8720 2563 8733 2609
rect 8907 2563 8920 2609
rect 8720 2500 8920 2563
rect 8720 -2563 8920 -2500
rect 8720 -2609 8733 -2563
rect 8907 -2609 8920 -2563
rect 8720 -2622 8920 -2609
rect 9000 2609 9200 2622
rect 9000 2563 9013 2609
rect 9187 2563 9200 2609
rect 9000 2500 9200 2563
rect 9000 -2563 9200 -2500
rect 9000 -2609 9013 -2563
rect 9187 -2609 9200 -2563
rect 9000 -2622 9200 -2609
rect 9280 2609 9480 2622
rect 9280 2563 9293 2609
rect 9467 2563 9480 2609
rect 9280 2500 9480 2563
rect 9280 -2563 9480 -2500
rect 9280 -2609 9293 -2563
rect 9467 -2609 9480 -2563
rect 9280 -2622 9480 -2609
rect 9560 2609 9760 2622
rect 9560 2563 9573 2609
rect 9747 2563 9760 2609
rect 9560 2500 9760 2563
rect 9560 -2563 9760 -2500
rect 9560 -2609 9573 -2563
rect 9747 -2609 9760 -2563
rect 9560 -2622 9760 -2609
rect 9840 2609 10040 2622
rect 9840 2563 9853 2609
rect 10027 2563 10040 2609
rect 9840 2500 10040 2563
rect 9840 -2563 10040 -2500
rect 9840 -2609 9853 -2563
rect 10027 -2609 10040 -2563
rect 9840 -2622 10040 -2609
rect 10120 2609 10320 2622
rect 10120 2563 10133 2609
rect 10307 2563 10320 2609
rect 10120 2500 10320 2563
rect 10120 -2563 10320 -2500
rect 10120 -2609 10133 -2563
rect 10307 -2609 10320 -2563
rect 10120 -2622 10320 -2609
rect 10400 2609 10600 2622
rect 10400 2563 10413 2609
rect 10587 2563 10600 2609
rect 10400 2500 10600 2563
rect 10400 -2563 10600 -2500
rect 10400 -2609 10413 -2563
rect 10587 -2609 10600 -2563
rect 10400 -2622 10600 -2609
rect 10680 2609 10880 2622
rect 10680 2563 10693 2609
rect 10867 2563 10880 2609
rect 10680 2500 10880 2563
rect 10680 -2563 10880 -2500
rect 10680 -2609 10693 -2563
rect 10867 -2609 10880 -2563
rect 10680 -2622 10880 -2609
rect 10960 2609 11160 2622
rect 10960 2563 10973 2609
rect 11147 2563 11160 2609
rect 10960 2500 11160 2563
rect 10960 -2563 11160 -2500
rect 10960 -2609 10973 -2563
rect 11147 -2609 11160 -2563
rect 10960 -2622 11160 -2609
rect 11240 2609 11440 2622
rect 11240 2563 11253 2609
rect 11427 2563 11440 2609
rect 11240 2500 11440 2563
rect 11240 -2563 11440 -2500
rect 11240 -2609 11253 -2563
rect 11427 -2609 11440 -2563
rect 11240 -2622 11440 -2609
rect 11520 2609 11720 2622
rect 11520 2563 11533 2609
rect 11707 2563 11720 2609
rect 11520 2500 11720 2563
rect 11520 -2563 11720 -2500
rect 11520 -2609 11533 -2563
rect 11707 -2609 11720 -2563
rect 11520 -2622 11720 -2609
rect 11800 2609 12000 2622
rect 11800 2563 11813 2609
rect 11987 2563 12000 2609
rect 11800 2500 12000 2563
rect 11800 -2563 12000 -2500
rect 11800 -2609 11813 -2563
rect 11987 -2609 12000 -2563
rect 11800 -2622 12000 -2609
rect 12080 2609 12280 2622
rect 12080 2563 12093 2609
rect 12267 2563 12280 2609
rect 12080 2500 12280 2563
rect 12080 -2563 12280 -2500
rect 12080 -2609 12093 -2563
rect 12267 -2609 12280 -2563
rect 12080 -2622 12280 -2609
<< polycontact >>
rect -12267 2563 -12093 2609
rect -12267 -2609 -12093 -2563
rect -11987 2563 -11813 2609
rect -11987 -2609 -11813 -2563
rect -11707 2563 -11533 2609
rect -11707 -2609 -11533 -2563
rect -11427 2563 -11253 2609
rect -11427 -2609 -11253 -2563
rect -11147 2563 -10973 2609
rect -11147 -2609 -10973 -2563
rect -10867 2563 -10693 2609
rect -10867 -2609 -10693 -2563
rect -10587 2563 -10413 2609
rect -10587 -2609 -10413 -2563
rect -10307 2563 -10133 2609
rect -10307 -2609 -10133 -2563
rect -10027 2563 -9853 2609
rect -10027 -2609 -9853 -2563
rect -9747 2563 -9573 2609
rect -9747 -2609 -9573 -2563
rect -9467 2563 -9293 2609
rect -9467 -2609 -9293 -2563
rect -9187 2563 -9013 2609
rect -9187 -2609 -9013 -2563
rect -8907 2563 -8733 2609
rect -8907 -2609 -8733 -2563
rect -8627 2563 -8453 2609
rect -8627 -2609 -8453 -2563
rect -8347 2563 -8173 2609
rect -8347 -2609 -8173 -2563
rect -8067 2563 -7893 2609
rect -8067 -2609 -7893 -2563
rect -7787 2563 -7613 2609
rect -7787 -2609 -7613 -2563
rect -7507 2563 -7333 2609
rect -7507 -2609 -7333 -2563
rect -7227 2563 -7053 2609
rect -7227 -2609 -7053 -2563
rect -6947 2563 -6773 2609
rect -6947 -2609 -6773 -2563
rect -6667 2563 -6493 2609
rect -6667 -2609 -6493 -2563
rect -6387 2563 -6213 2609
rect -6387 -2609 -6213 -2563
rect -6107 2563 -5933 2609
rect -6107 -2609 -5933 -2563
rect -5827 2563 -5653 2609
rect -5827 -2609 -5653 -2563
rect -5547 2563 -5373 2609
rect -5547 -2609 -5373 -2563
rect -5267 2563 -5093 2609
rect -5267 -2609 -5093 -2563
rect -4987 2563 -4813 2609
rect -4987 -2609 -4813 -2563
rect -4707 2563 -4533 2609
rect -4707 -2609 -4533 -2563
rect -4427 2563 -4253 2609
rect -4427 -2609 -4253 -2563
rect -4147 2563 -3973 2609
rect -4147 -2609 -3973 -2563
rect -3867 2563 -3693 2609
rect -3867 -2609 -3693 -2563
rect -3587 2563 -3413 2609
rect -3587 -2609 -3413 -2563
rect -3307 2563 -3133 2609
rect -3307 -2609 -3133 -2563
rect -3027 2563 -2853 2609
rect -3027 -2609 -2853 -2563
rect -2747 2563 -2573 2609
rect -2747 -2609 -2573 -2563
rect -2467 2563 -2293 2609
rect -2467 -2609 -2293 -2563
rect -2187 2563 -2013 2609
rect -2187 -2609 -2013 -2563
rect -1907 2563 -1733 2609
rect -1907 -2609 -1733 -2563
rect -1627 2563 -1453 2609
rect -1627 -2609 -1453 -2563
rect -1347 2563 -1173 2609
rect -1347 -2609 -1173 -2563
rect -1067 2563 -893 2609
rect -1067 -2609 -893 -2563
rect -787 2563 -613 2609
rect -787 -2609 -613 -2563
rect -507 2563 -333 2609
rect -507 -2609 -333 -2563
rect -227 2563 -53 2609
rect -227 -2609 -53 -2563
rect 53 2563 227 2609
rect 53 -2609 227 -2563
rect 333 2563 507 2609
rect 333 -2609 507 -2563
rect 613 2563 787 2609
rect 613 -2609 787 -2563
rect 893 2563 1067 2609
rect 893 -2609 1067 -2563
rect 1173 2563 1347 2609
rect 1173 -2609 1347 -2563
rect 1453 2563 1627 2609
rect 1453 -2609 1627 -2563
rect 1733 2563 1907 2609
rect 1733 -2609 1907 -2563
rect 2013 2563 2187 2609
rect 2013 -2609 2187 -2563
rect 2293 2563 2467 2609
rect 2293 -2609 2467 -2563
rect 2573 2563 2747 2609
rect 2573 -2609 2747 -2563
rect 2853 2563 3027 2609
rect 2853 -2609 3027 -2563
rect 3133 2563 3307 2609
rect 3133 -2609 3307 -2563
rect 3413 2563 3587 2609
rect 3413 -2609 3587 -2563
rect 3693 2563 3867 2609
rect 3693 -2609 3867 -2563
rect 3973 2563 4147 2609
rect 3973 -2609 4147 -2563
rect 4253 2563 4427 2609
rect 4253 -2609 4427 -2563
rect 4533 2563 4707 2609
rect 4533 -2609 4707 -2563
rect 4813 2563 4987 2609
rect 4813 -2609 4987 -2563
rect 5093 2563 5267 2609
rect 5093 -2609 5267 -2563
rect 5373 2563 5547 2609
rect 5373 -2609 5547 -2563
rect 5653 2563 5827 2609
rect 5653 -2609 5827 -2563
rect 5933 2563 6107 2609
rect 5933 -2609 6107 -2563
rect 6213 2563 6387 2609
rect 6213 -2609 6387 -2563
rect 6493 2563 6667 2609
rect 6493 -2609 6667 -2563
rect 6773 2563 6947 2609
rect 6773 -2609 6947 -2563
rect 7053 2563 7227 2609
rect 7053 -2609 7227 -2563
rect 7333 2563 7507 2609
rect 7333 -2609 7507 -2563
rect 7613 2563 7787 2609
rect 7613 -2609 7787 -2563
rect 7893 2563 8067 2609
rect 7893 -2609 8067 -2563
rect 8173 2563 8347 2609
rect 8173 -2609 8347 -2563
rect 8453 2563 8627 2609
rect 8453 -2609 8627 -2563
rect 8733 2563 8907 2609
rect 8733 -2609 8907 -2563
rect 9013 2563 9187 2609
rect 9013 -2609 9187 -2563
rect 9293 2563 9467 2609
rect 9293 -2609 9467 -2563
rect 9573 2563 9747 2609
rect 9573 -2609 9747 -2563
rect 9853 2563 10027 2609
rect 9853 -2609 10027 -2563
rect 10133 2563 10307 2609
rect 10133 -2609 10307 -2563
rect 10413 2563 10587 2609
rect 10413 -2609 10587 -2563
rect 10693 2563 10867 2609
rect 10693 -2609 10867 -2563
rect 10973 2563 11147 2609
rect 10973 -2609 11147 -2563
rect 11253 2563 11427 2609
rect 11253 -2609 11427 -2563
rect 11533 2563 11707 2609
rect 11533 -2609 11707 -2563
rect 11813 2563 11987 2609
rect 11813 -2609 11987 -2563
rect 12093 2563 12267 2609
rect 12093 -2609 12267 -2563
<< mvnhighres >>
rect -12280 -2500 -12080 2500
rect -12000 -2500 -11800 2500
rect -11720 -2500 -11520 2500
rect -11440 -2500 -11240 2500
rect -11160 -2500 -10960 2500
rect -10880 -2500 -10680 2500
rect -10600 -2500 -10400 2500
rect -10320 -2500 -10120 2500
rect -10040 -2500 -9840 2500
rect -9760 -2500 -9560 2500
rect -9480 -2500 -9280 2500
rect -9200 -2500 -9000 2500
rect -8920 -2500 -8720 2500
rect -8640 -2500 -8440 2500
rect -8360 -2500 -8160 2500
rect -8080 -2500 -7880 2500
rect -7800 -2500 -7600 2500
rect -7520 -2500 -7320 2500
rect -7240 -2500 -7040 2500
rect -6960 -2500 -6760 2500
rect -6680 -2500 -6480 2500
rect -6400 -2500 -6200 2500
rect -6120 -2500 -5920 2500
rect -5840 -2500 -5640 2500
rect -5560 -2500 -5360 2500
rect -5280 -2500 -5080 2500
rect -5000 -2500 -4800 2500
rect -4720 -2500 -4520 2500
rect -4440 -2500 -4240 2500
rect -4160 -2500 -3960 2500
rect -3880 -2500 -3680 2500
rect -3600 -2500 -3400 2500
rect -3320 -2500 -3120 2500
rect -3040 -2500 -2840 2500
rect -2760 -2500 -2560 2500
rect -2480 -2500 -2280 2500
rect -2200 -2500 -2000 2500
rect -1920 -2500 -1720 2500
rect -1640 -2500 -1440 2500
rect -1360 -2500 -1160 2500
rect -1080 -2500 -880 2500
rect -800 -2500 -600 2500
rect -520 -2500 -320 2500
rect -240 -2500 -40 2500
rect 40 -2500 240 2500
rect 320 -2500 520 2500
rect 600 -2500 800 2500
rect 880 -2500 1080 2500
rect 1160 -2500 1360 2500
rect 1440 -2500 1640 2500
rect 1720 -2500 1920 2500
rect 2000 -2500 2200 2500
rect 2280 -2500 2480 2500
rect 2560 -2500 2760 2500
rect 2840 -2500 3040 2500
rect 3120 -2500 3320 2500
rect 3400 -2500 3600 2500
rect 3680 -2500 3880 2500
rect 3960 -2500 4160 2500
rect 4240 -2500 4440 2500
rect 4520 -2500 4720 2500
rect 4800 -2500 5000 2500
rect 5080 -2500 5280 2500
rect 5360 -2500 5560 2500
rect 5640 -2500 5840 2500
rect 5920 -2500 6120 2500
rect 6200 -2500 6400 2500
rect 6480 -2500 6680 2500
rect 6760 -2500 6960 2500
rect 7040 -2500 7240 2500
rect 7320 -2500 7520 2500
rect 7600 -2500 7800 2500
rect 7880 -2500 8080 2500
rect 8160 -2500 8360 2500
rect 8440 -2500 8640 2500
rect 8720 -2500 8920 2500
rect 9000 -2500 9200 2500
rect 9280 -2500 9480 2500
rect 9560 -2500 9760 2500
rect 9840 -2500 10040 2500
rect 10120 -2500 10320 2500
rect 10400 -2500 10600 2500
rect 10680 -2500 10880 2500
rect 10960 -2500 11160 2500
rect 11240 -2500 11440 2500
rect 11520 -2500 11720 2500
rect 11800 -2500 12000 2500
rect 12080 -2500 12280 2500
<< metal1 >>
rect -12479 2775 -12345 2821
rect 12356 2775 12479 2821
rect -12479 2718 -12433 2775
rect 12433 2718 12479 2775
rect -12278 2563 -12267 2609
rect -12093 2563 -12082 2609
rect -11998 2563 -11987 2609
rect -11813 2563 -11802 2609
rect -11718 2563 -11707 2609
rect -11533 2563 -11522 2609
rect -11438 2563 -11427 2609
rect -11253 2563 -11242 2609
rect -11158 2563 -11147 2609
rect -10973 2563 -10962 2609
rect -10878 2563 -10867 2609
rect -10693 2563 -10682 2609
rect -10598 2563 -10587 2609
rect -10413 2563 -10402 2609
rect -10318 2563 -10307 2609
rect -10133 2563 -10122 2609
rect -10038 2563 -10027 2609
rect -9853 2563 -9842 2609
rect -9758 2563 -9747 2609
rect -9573 2563 -9562 2609
rect -9478 2563 -9467 2609
rect -9293 2563 -9282 2609
rect -9198 2563 -9187 2609
rect -9013 2563 -9002 2609
rect -8918 2563 -8907 2609
rect -8733 2563 -8722 2609
rect -8638 2563 -8627 2609
rect -8453 2563 -8442 2609
rect -8358 2563 -8347 2609
rect -8173 2563 -8162 2609
rect -8078 2563 -8067 2609
rect -7893 2563 -7882 2609
rect -7798 2563 -7787 2609
rect -7613 2563 -7602 2609
rect -7518 2563 -7507 2609
rect -7333 2563 -7322 2609
rect -7238 2563 -7227 2609
rect -7053 2563 -7042 2609
rect -6958 2563 -6947 2609
rect -6773 2563 -6762 2609
rect -6678 2563 -6667 2609
rect -6493 2563 -6482 2609
rect -6398 2563 -6387 2609
rect -6213 2563 -6202 2609
rect -6118 2563 -6107 2609
rect -5933 2563 -5922 2609
rect -5838 2563 -5827 2609
rect -5653 2563 -5642 2609
rect -5558 2563 -5547 2609
rect -5373 2563 -5362 2609
rect -5278 2563 -5267 2609
rect -5093 2563 -5082 2609
rect -4998 2563 -4987 2609
rect -4813 2563 -4802 2609
rect -4718 2563 -4707 2609
rect -4533 2563 -4522 2609
rect -4438 2563 -4427 2609
rect -4253 2563 -4242 2609
rect -4158 2563 -4147 2609
rect -3973 2563 -3962 2609
rect -3878 2563 -3867 2609
rect -3693 2563 -3682 2609
rect -3598 2563 -3587 2609
rect -3413 2563 -3402 2609
rect -3318 2563 -3307 2609
rect -3133 2563 -3122 2609
rect -3038 2563 -3027 2609
rect -2853 2563 -2842 2609
rect -2758 2563 -2747 2609
rect -2573 2563 -2562 2609
rect -2478 2563 -2467 2609
rect -2293 2563 -2282 2609
rect -2198 2563 -2187 2609
rect -2013 2563 -2002 2609
rect -1918 2563 -1907 2609
rect -1733 2563 -1722 2609
rect -1638 2563 -1627 2609
rect -1453 2563 -1442 2609
rect -1358 2563 -1347 2609
rect -1173 2563 -1162 2609
rect -1078 2563 -1067 2609
rect -893 2563 -882 2609
rect -798 2563 -787 2609
rect -613 2563 -602 2609
rect -518 2563 -507 2609
rect -333 2563 -322 2609
rect -238 2563 -227 2609
rect -53 2563 -42 2609
rect 42 2563 53 2609
rect 227 2563 238 2609
rect 322 2563 333 2609
rect 507 2563 518 2609
rect 602 2563 613 2609
rect 787 2563 798 2609
rect 882 2563 893 2609
rect 1067 2563 1078 2609
rect 1162 2563 1173 2609
rect 1347 2563 1358 2609
rect 1442 2563 1453 2609
rect 1627 2563 1638 2609
rect 1722 2563 1733 2609
rect 1907 2563 1918 2609
rect 2002 2563 2013 2609
rect 2187 2563 2198 2609
rect 2282 2563 2293 2609
rect 2467 2563 2478 2609
rect 2562 2563 2573 2609
rect 2747 2563 2758 2609
rect 2842 2563 2853 2609
rect 3027 2563 3038 2609
rect 3122 2563 3133 2609
rect 3307 2563 3318 2609
rect 3402 2563 3413 2609
rect 3587 2563 3598 2609
rect 3682 2563 3693 2609
rect 3867 2563 3878 2609
rect 3962 2563 3973 2609
rect 4147 2563 4158 2609
rect 4242 2563 4253 2609
rect 4427 2563 4438 2609
rect 4522 2563 4533 2609
rect 4707 2563 4718 2609
rect 4802 2563 4813 2609
rect 4987 2563 4998 2609
rect 5082 2563 5093 2609
rect 5267 2563 5278 2609
rect 5362 2563 5373 2609
rect 5547 2563 5558 2609
rect 5642 2563 5653 2609
rect 5827 2563 5838 2609
rect 5922 2563 5933 2609
rect 6107 2563 6118 2609
rect 6202 2563 6213 2609
rect 6387 2563 6398 2609
rect 6482 2563 6493 2609
rect 6667 2563 6678 2609
rect 6762 2563 6773 2609
rect 6947 2563 6958 2609
rect 7042 2563 7053 2609
rect 7227 2563 7238 2609
rect 7322 2563 7333 2609
rect 7507 2563 7518 2609
rect 7602 2563 7613 2609
rect 7787 2563 7798 2609
rect 7882 2563 7893 2609
rect 8067 2563 8078 2609
rect 8162 2563 8173 2609
rect 8347 2563 8358 2609
rect 8442 2563 8453 2609
rect 8627 2563 8638 2609
rect 8722 2563 8733 2609
rect 8907 2563 8918 2609
rect 9002 2563 9013 2609
rect 9187 2563 9198 2609
rect 9282 2563 9293 2609
rect 9467 2563 9478 2609
rect 9562 2563 9573 2609
rect 9747 2563 9758 2609
rect 9842 2563 9853 2609
rect 10027 2563 10038 2609
rect 10122 2563 10133 2609
rect 10307 2563 10318 2609
rect 10402 2563 10413 2609
rect 10587 2563 10598 2609
rect 10682 2563 10693 2609
rect 10867 2563 10878 2609
rect 10962 2563 10973 2609
rect 11147 2563 11158 2609
rect 11242 2563 11253 2609
rect 11427 2563 11438 2609
rect 11522 2563 11533 2609
rect 11707 2563 11718 2609
rect 11802 2563 11813 2609
rect 11987 2563 11998 2609
rect 12082 2563 12093 2609
rect 12267 2563 12278 2609
rect -12278 -2609 -12267 -2563
rect -12093 -2609 -12082 -2563
rect -11998 -2609 -11987 -2563
rect -11813 -2609 -11802 -2563
rect -11718 -2609 -11707 -2563
rect -11533 -2609 -11522 -2563
rect -11438 -2609 -11427 -2563
rect -11253 -2609 -11242 -2563
rect -11158 -2609 -11147 -2563
rect -10973 -2609 -10962 -2563
rect -10878 -2609 -10867 -2563
rect -10693 -2609 -10682 -2563
rect -10598 -2609 -10587 -2563
rect -10413 -2609 -10402 -2563
rect -10318 -2609 -10307 -2563
rect -10133 -2609 -10122 -2563
rect -10038 -2609 -10027 -2563
rect -9853 -2609 -9842 -2563
rect -9758 -2609 -9747 -2563
rect -9573 -2609 -9562 -2563
rect -9478 -2609 -9467 -2563
rect -9293 -2609 -9282 -2563
rect -9198 -2609 -9187 -2563
rect -9013 -2609 -9002 -2563
rect -8918 -2609 -8907 -2563
rect -8733 -2609 -8722 -2563
rect -8638 -2609 -8627 -2563
rect -8453 -2609 -8442 -2563
rect -8358 -2609 -8347 -2563
rect -8173 -2609 -8162 -2563
rect -8078 -2609 -8067 -2563
rect -7893 -2609 -7882 -2563
rect -7798 -2609 -7787 -2563
rect -7613 -2609 -7602 -2563
rect -7518 -2609 -7507 -2563
rect -7333 -2609 -7322 -2563
rect -7238 -2609 -7227 -2563
rect -7053 -2609 -7042 -2563
rect -6958 -2609 -6947 -2563
rect -6773 -2609 -6762 -2563
rect -6678 -2609 -6667 -2563
rect -6493 -2609 -6482 -2563
rect -6398 -2609 -6387 -2563
rect -6213 -2609 -6202 -2563
rect -6118 -2609 -6107 -2563
rect -5933 -2609 -5922 -2563
rect -5838 -2609 -5827 -2563
rect -5653 -2609 -5642 -2563
rect -5558 -2609 -5547 -2563
rect -5373 -2609 -5362 -2563
rect -5278 -2609 -5267 -2563
rect -5093 -2609 -5082 -2563
rect -4998 -2609 -4987 -2563
rect -4813 -2609 -4802 -2563
rect -4718 -2609 -4707 -2563
rect -4533 -2609 -4522 -2563
rect -4438 -2609 -4427 -2563
rect -4253 -2609 -4242 -2563
rect -4158 -2609 -4147 -2563
rect -3973 -2609 -3962 -2563
rect -3878 -2609 -3867 -2563
rect -3693 -2609 -3682 -2563
rect -3598 -2609 -3587 -2563
rect -3413 -2609 -3402 -2563
rect -3318 -2609 -3307 -2563
rect -3133 -2609 -3122 -2563
rect -3038 -2609 -3027 -2563
rect -2853 -2609 -2842 -2563
rect -2758 -2609 -2747 -2563
rect -2573 -2609 -2562 -2563
rect -2478 -2609 -2467 -2563
rect -2293 -2609 -2282 -2563
rect -2198 -2609 -2187 -2563
rect -2013 -2609 -2002 -2563
rect -1918 -2609 -1907 -2563
rect -1733 -2609 -1722 -2563
rect -1638 -2609 -1627 -2563
rect -1453 -2609 -1442 -2563
rect -1358 -2609 -1347 -2563
rect -1173 -2609 -1162 -2563
rect -1078 -2609 -1067 -2563
rect -893 -2609 -882 -2563
rect -798 -2609 -787 -2563
rect -613 -2609 -602 -2563
rect -518 -2609 -507 -2563
rect -333 -2609 -322 -2563
rect -238 -2609 -227 -2563
rect -53 -2609 -42 -2563
rect 42 -2609 53 -2563
rect 227 -2609 238 -2563
rect 322 -2609 333 -2563
rect 507 -2609 518 -2563
rect 602 -2609 613 -2563
rect 787 -2609 798 -2563
rect 882 -2609 893 -2563
rect 1067 -2609 1078 -2563
rect 1162 -2609 1173 -2563
rect 1347 -2609 1358 -2563
rect 1442 -2609 1453 -2563
rect 1627 -2609 1638 -2563
rect 1722 -2609 1733 -2563
rect 1907 -2609 1918 -2563
rect 2002 -2609 2013 -2563
rect 2187 -2609 2198 -2563
rect 2282 -2609 2293 -2563
rect 2467 -2609 2478 -2563
rect 2562 -2609 2573 -2563
rect 2747 -2609 2758 -2563
rect 2842 -2609 2853 -2563
rect 3027 -2609 3038 -2563
rect 3122 -2609 3133 -2563
rect 3307 -2609 3318 -2563
rect 3402 -2609 3413 -2563
rect 3587 -2609 3598 -2563
rect 3682 -2609 3693 -2563
rect 3867 -2609 3878 -2563
rect 3962 -2609 3973 -2563
rect 4147 -2609 4158 -2563
rect 4242 -2609 4253 -2563
rect 4427 -2609 4438 -2563
rect 4522 -2609 4533 -2563
rect 4707 -2609 4718 -2563
rect 4802 -2609 4813 -2563
rect 4987 -2609 4998 -2563
rect 5082 -2609 5093 -2563
rect 5267 -2609 5278 -2563
rect 5362 -2609 5373 -2563
rect 5547 -2609 5558 -2563
rect 5642 -2609 5653 -2563
rect 5827 -2609 5838 -2563
rect 5922 -2609 5933 -2563
rect 6107 -2609 6118 -2563
rect 6202 -2609 6213 -2563
rect 6387 -2609 6398 -2563
rect 6482 -2609 6493 -2563
rect 6667 -2609 6678 -2563
rect 6762 -2609 6773 -2563
rect 6947 -2609 6958 -2563
rect 7042 -2609 7053 -2563
rect 7227 -2609 7238 -2563
rect 7322 -2609 7333 -2563
rect 7507 -2609 7518 -2563
rect 7602 -2609 7613 -2563
rect 7787 -2609 7798 -2563
rect 7882 -2609 7893 -2563
rect 8067 -2609 8078 -2563
rect 8162 -2609 8173 -2563
rect 8347 -2609 8358 -2563
rect 8442 -2609 8453 -2563
rect 8627 -2609 8638 -2563
rect 8722 -2609 8733 -2563
rect 8907 -2609 8918 -2563
rect 9002 -2609 9013 -2563
rect 9187 -2609 9198 -2563
rect 9282 -2609 9293 -2563
rect 9467 -2609 9478 -2563
rect 9562 -2609 9573 -2563
rect 9747 -2609 9758 -2563
rect 9842 -2609 9853 -2563
rect 10027 -2609 10038 -2563
rect 10122 -2609 10133 -2563
rect 10307 -2609 10318 -2563
rect 10402 -2609 10413 -2563
rect 10587 -2609 10598 -2563
rect 10682 -2609 10693 -2563
rect 10867 -2609 10878 -2563
rect 10962 -2609 10973 -2563
rect 11147 -2609 11158 -2563
rect 11242 -2609 11253 -2563
rect 11427 -2609 11438 -2563
rect 11522 -2609 11533 -2563
rect 11707 -2609 11718 -2563
rect 11802 -2609 11813 -2563
rect 11987 -2609 11998 -2563
rect 12082 -2609 12093 -2563
rect 12267 -2609 12278 -2563
rect -12479 -2775 -12433 -2718
rect 12433 -2775 12479 -2718
rect -12479 -2821 -12372 -2775
rect 12329 -2821 12479 -2775
<< properties >>
string FIXED_BBOX -12404 -2784 12404 2784
string gencell ppolyf_u_1k_6p0
string library gf180mcu
string parameters w 1.000 l 25.000 m 1 nx 88 wmin 1.000 lmin 1.000 rho 1000 val 25.0k dummy 0 dw 0.0 term 0.0 sterm 0.0 caplen 0.4 snake 0 glc 1 grc 1 gtc 0 gbc 0 roverlap 0 endcov 100 full_metal 1 compatible {ppolyf_u_1k ppolyf_u_1k_6p0}
<< end >>
