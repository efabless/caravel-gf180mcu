magic
tech gf180mcuC
magscale 1 10
timestamp 1654981632
<< metal1 >>
rect 11610 14870 11622 14922
rect 11674 14919 11686 14922
rect 11674 14873 38662 14919
rect 11674 14870 11686 14873
rect 38616 14807 38662 14873
rect 63242 14870 63254 14922
rect 63306 14919 63318 14922
rect 63306 14873 71815 14919
rect 63306 14870 63318 14873
rect 68394 14807 68406 14810
rect 38616 14761 68406 14807
rect 68394 14758 68406 14761
rect 68458 14758 68470 14810
rect 71769 14807 71815 14873
rect 73322 14870 73334 14922
rect 73386 14919 73398 14922
rect 79482 14919 79494 14922
rect 73386 14873 79494 14919
rect 73386 14870 73398 14873
rect 79482 14870 79494 14873
rect 79546 14870 79558 14922
rect 80714 14870 80726 14922
rect 80778 14919 80790 14922
rect 80778 14873 103175 14919
rect 80778 14870 80790 14873
rect 103129 14807 103175 14873
rect 103226 14870 103238 14922
rect 103290 14919 103302 14922
rect 103290 14873 104183 14919
rect 103290 14870 103302 14873
rect 104010 14807 104022 14810
rect 71769 14761 102839 14807
rect 103129 14761 104022 14807
rect 9482 14646 9494 14698
rect 9546 14695 9558 14698
rect 63130 14695 63142 14698
rect 9546 14649 63142 14695
rect 9546 14646 9558 14649
rect 63130 14646 63142 14649
rect 63194 14646 63206 14698
rect 64026 14646 64038 14698
rect 64090 14695 64102 14698
rect 73322 14695 73334 14698
rect 64090 14649 73334 14695
rect 64090 14646 64102 14649
rect 73322 14646 73334 14649
rect 73386 14646 73398 14698
rect 73546 14646 73558 14698
rect 73610 14695 73622 14698
rect 78698 14695 78710 14698
rect 73610 14649 78710 14695
rect 73610 14646 73622 14649
rect 78698 14646 78710 14649
rect 78762 14646 78774 14698
rect 79258 14695 79270 14698
rect 78825 14649 79270 14695
rect 10042 14534 10054 14586
rect 10106 14583 10118 14586
rect 78825 14583 78871 14649
rect 79258 14646 79270 14649
rect 79322 14646 79334 14698
rect 79930 14695 79942 14698
rect 79385 14649 79942 14695
rect 79385 14583 79431 14649
rect 79930 14646 79942 14649
rect 79994 14646 80006 14698
rect 80154 14646 80166 14698
rect 80218 14695 80230 14698
rect 80714 14695 80726 14698
rect 80218 14649 80726 14695
rect 80218 14646 80230 14649
rect 80714 14646 80726 14649
rect 80778 14646 80790 14698
rect 80938 14646 80950 14698
rect 81002 14695 81014 14698
rect 82842 14695 82854 14698
rect 81002 14649 82854 14695
rect 81002 14646 81014 14649
rect 82842 14646 82854 14649
rect 82906 14646 82918 14698
rect 83066 14646 83078 14698
rect 83130 14695 83142 14698
rect 84410 14695 84422 14698
rect 83130 14649 84422 14695
rect 83130 14646 83142 14649
rect 84410 14646 84422 14649
rect 84474 14646 84486 14698
rect 84970 14646 84982 14698
rect 85034 14695 85046 14698
rect 90794 14695 90806 14698
rect 85034 14649 90806 14695
rect 85034 14646 85046 14649
rect 90794 14646 90806 14649
rect 90858 14646 90870 14698
rect 91018 14646 91030 14698
rect 91082 14695 91094 14698
rect 102666 14695 102678 14698
rect 91082 14649 102678 14695
rect 91082 14646 91094 14649
rect 102666 14646 102678 14649
rect 102730 14646 102742 14698
rect 102793 14695 102839 14761
rect 104010 14758 104022 14761
rect 104074 14758 104086 14810
rect 104137 14807 104183 14873
rect 104794 14870 104806 14922
rect 104858 14919 104870 14922
rect 104858 14873 120982 14919
rect 104858 14870 104870 14873
rect 104137 14761 115831 14807
rect 115658 14695 115670 14698
rect 102793 14649 115670 14695
rect 115658 14646 115670 14649
rect 115722 14646 115734 14698
rect 10106 14537 78871 14583
rect 78937 14537 79431 14583
rect 10106 14534 10118 14537
rect 51034 14422 51046 14474
rect 51098 14471 51110 14474
rect 74890 14471 74902 14474
rect 51098 14425 74902 14471
rect 51098 14422 51110 14425
rect 74890 14422 74902 14425
rect 74954 14422 74966 14474
rect 75562 14422 75574 14474
rect 75626 14471 75638 14474
rect 78937 14471 78983 14537
rect 79482 14534 79494 14586
rect 79546 14583 79558 14586
rect 81498 14583 81510 14586
rect 79546 14537 81510 14583
rect 79546 14534 79558 14537
rect 81498 14534 81510 14537
rect 81562 14534 81574 14586
rect 103898 14583 103910 14586
rect 81625 14537 103910 14583
rect 75626 14425 78983 14471
rect 75626 14422 75638 14425
rect 79370 14422 79382 14474
rect 79434 14471 79446 14474
rect 81625 14471 81671 14537
rect 103898 14534 103910 14537
rect 103962 14534 103974 14586
rect 104682 14534 104694 14586
rect 104746 14583 104758 14586
rect 113418 14583 113430 14586
rect 104746 14537 113430 14583
rect 104746 14534 104758 14537
rect 113418 14534 113430 14537
rect 113482 14534 113494 14586
rect 113545 14537 115159 14583
rect 79434 14425 81671 14471
rect 83193 14425 91751 14471
rect 79434 14422 79446 14425
rect 8474 14310 8486 14362
rect 8538 14359 8550 14362
rect 8538 14313 80887 14359
rect 8538 14310 8550 14313
rect 53050 14198 53062 14250
rect 53114 14247 53126 14250
rect 73546 14247 73558 14250
rect 53114 14201 73558 14247
rect 53114 14198 53126 14201
rect 73546 14198 73558 14201
rect 73610 14198 73622 14250
rect 80714 14247 80726 14250
rect 73785 14201 80726 14247
rect 1866 14086 1878 14138
rect 1930 14135 1942 14138
rect 57530 14135 57542 14138
rect 1930 14089 57542 14135
rect 1930 14086 1942 14089
rect 57530 14086 57542 14089
rect 57594 14086 57606 14138
rect 61674 14086 61686 14138
rect 61738 14135 61750 14138
rect 64138 14135 64150 14138
rect 61738 14089 64150 14135
rect 61738 14086 61750 14089
rect 64138 14086 64150 14089
rect 64202 14086 64214 14138
rect 65930 14086 65942 14138
rect 65994 14135 66006 14138
rect 73785 14135 73831 14201
rect 80714 14198 80726 14201
rect 80778 14198 80790 14250
rect 80841 14247 80887 14313
rect 80938 14310 80950 14362
rect 81002 14359 81014 14362
rect 83066 14359 83078 14362
rect 81002 14313 83078 14359
rect 81002 14310 81014 14313
rect 83066 14310 83078 14313
rect 83130 14310 83142 14362
rect 83193 14247 83239 14425
rect 84522 14310 84534 14362
rect 84586 14359 84598 14362
rect 91578 14359 91590 14362
rect 84586 14313 91590 14359
rect 84586 14310 84598 14313
rect 91578 14310 91590 14313
rect 91642 14310 91654 14362
rect 91705 14359 91751 14425
rect 98298 14422 98310 14474
rect 98362 14471 98374 14474
rect 98362 14425 102335 14471
rect 98362 14422 98374 14425
rect 101994 14359 102006 14362
rect 91705 14313 102006 14359
rect 101994 14310 102006 14313
rect 102058 14310 102070 14362
rect 88218 14247 88230 14250
rect 80841 14201 83239 14247
rect 83305 14201 88230 14247
rect 65994 14089 73831 14135
rect 65994 14086 66006 14089
rect 73994 14086 74006 14138
rect 74058 14135 74070 14138
rect 75562 14135 75574 14138
rect 74058 14089 75574 14135
rect 74058 14086 74070 14089
rect 75562 14086 75574 14089
rect 75626 14086 75638 14138
rect 76906 14086 76918 14138
rect 76970 14135 76982 14138
rect 77354 14135 77366 14138
rect 76970 14089 77366 14135
rect 76970 14086 76982 14089
rect 77354 14086 77366 14089
rect 77418 14086 77430 14138
rect 77578 14086 77590 14138
rect 77642 14135 77654 14138
rect 78026 14135 78038 14138
rect 77642 14089 78038 14135
rect 77642 14086 77654 14089
rect 78026 14086 78038 14089
rect 78090 14086 78102 14138
rect 78362 14086 78374 14138
rect 78426 14135 78438 14138
rect 78810 14135 78822 14138
rect 78426 14089 78822 14135
rect 78426 14086 78438 14089
rect 78810 14086 78822 14089
rect 78874 14086 78886 14138
rect 79034 14086 79046 14138
rect 79098 14135 79110 14138
rect 79098 14089 79991 14135
rect 79098 14086 79110 14089
rect 45434 13974 45446 14026
rect 45498 14023 45510 14026
rect 64026 14023 64038 14026
rect 45498 13977 64038 14023
rect 45498 13974 45510 13977
rect 64026 13974 64038 13977
rect 64090 13974 64102 14026
rect 64474 13974 64486 14026
rect 64538 14023 64550 14026
rect 70410 14023 70422 14026
rect 64538 13977 70422 14023
rect 64538 13974 64550 13977
rect 70410 13974 70422 13977
rect 70474 13974 70486 14026
rect 71642 13974 71654 14026
rect 71706 14023 71718 14026
rect 74666 14023 74678 14026
rect 71706 13977 74678 14023
rect 71706 13974 71718 13977
rect 74666 13974 74678 13977
rect 74730 13974 74742 14026
rect 75002 13974 75014 14026
rect 75066 14023 75078 14026
rect 79945 14023 79991 14089
rect 80490 14086 80502 14138
rect 80554 14135 80566 14138
rect 81722 14135 81734 14138
rect 80554 14089 81734 14135
rect 80554 14086 80566 14089
rect 81722 14086 81734 14089
rect 81786 14086 81798 14138
rect 82170 14086 82182 14138
rect 82234 14135 82246 14138
rect 83305 14135 83351 14201
rect 88218 14198 88230 14201
rect 88282 14198 88294 14250
rect 88666 14198 88678 14250
rect 88730 14247 88742 14250
rect 100986 14247 100998 14250
rect 88730 14201 100998 14247
rect 88730 14198 88742 14201
rect 100986 14198 100998 14201
rect 101050 14198 101062 14250
rect 102289 14247 102335 14425
rect 102554 14422 102566 14474
rect 102618 14471 102630 14474
rect 113545 14471 113591 14537
rect 114874 14471 114886 14474
rect 102618 14425 113591 14471
rect 113657 14425 114886 14471
rect 102618 14422 102630 14425
rect 102442 14310 102454 14362
rect 102506 14359 102518 14362
rect 102506 14313 102839 14359
rect 102506 14310 102518 14313
rect 102666 14247 102678 14250
rect 102289 14201 102678 14247
rect 102666 14198 102678 14201
rect 102730 14198 102742 14250
rect 102793 14247 102839 14313
rect 104234 14310 104246 14362
rect 104298 14359 104310 14362
rect 113657 14359 113703 14425
rect 114874 14422 114886 14425
rect 114938 14422 114950 14474
rect 114986 14359 114998 14362
rect 104298 14313 113703 14359
rect 113769 14313 114998 14359
rect 104298 14310 104310 14313
rect 113769 14247 113815 14313
rect 114986 14310 114998 14313
rect 115050 14310 115062 14362
rect 115113 14359 115159 14537
rect 115785 14471 115831 14761
rect 115882 14758 115894 14810
rect 115946 14807 115958 14810
rect 120250 14807 120262 14810
rect 115946 14761 120262 14807
rect 115946 14758 115958 14761
rect 120250 14758 120262 14761
rect 120314 14758 120326 14810
rect 120936 14807 120982 14873
rect 121034 14870 121046 14922
rect 121098 14919 121110 14922
rect 127418 14919 127430 14922
rect 121098 14873 127430 14919
rect 121098 14870 121110 14873
rect 127418 14870 127430 14873
rect 127482 14870 127494 14922
rect 131114 14870 131126 14922
rect 131178 14919 131190 14922
rect 148586 14919 148598 14922
rect 131178 14873 148598 14919
rect 131178 14870 131190 14873
rect 148586 14870 148598 14873
rect 148650 14870 148662 14922
rect 121482 14807 121494 14810
rect 120936 14761 121494 14807
rect 121482 14758 121494 14761
rect 121546 14758 121558 14810
rect 122490 14758 122502 14810
rect 122554 14807 122566 14810
rect 151498 14807 151510 14810
rect 122554 14761 151510 14807
rect 122554 14758 122566 14761
rect 151498 14758 151510 14761
rect 151562 14758 151574 14810
rect 116330 14646 116342 14698
rect 116394 14695 116406 14698
rect 148362 14695 148374 14698
rect 116394 14649 148374 14695
rect 116394 14646 116406 14649
rect 148362 14646 148374 14649
rect 148426 14646 148438 14698
rect 116554 14534 116566 14586
rect 116618 14583 116630 14586
rect 116618 14537 137111 14583
rect 116618 14534 116630 14537
rect 116666 14471 116678 14474
rect 115785 14425 116678 14471
rect 116666 14422 116678 14425
rect 116730 14422 116742 14474
rect 117114 14422 117126 14474
rect 117178 14471 117190 14474
rect 137065 14471 137111 14537
rect 138954 14534 138966 14586
rect 139018 14583 139030 14586
rect 167514 14583 167526 14586
rect 139018 14537 167526 14583
rect 139018 14534 139030 14537
rect 167514 14534 167526 14537
rect 167578 14534 167590 14586
rect 149818 14471 149830 14474
rect 117178 14425 136999 14471
rect 137065 14425 149830 14471
rect 117178 14422 117190 14425
rect 115113 14313 118743 14359
rect 118697 14250 118743 14313
rect 118794 14310 118806 14362
rect 118858 14359 118870 14362
rect 120698 14359 120710 14362
rect 118858 14313 120710 14359
rect 118858 14310 118870 14313
rect 120698 14310 120710 14313
rect 120762 14310 120774 14362
rect 121594 14310 121606 14362
rect 121658 14359 121670 14362
rect 136266 14359 136278 14362
rect 121658 14313 136278 14359
rect 121658 14310 121670 14313
rect 136266 14310 136278 14313
rect 136330 14310 136342 14362
rect 136953 14359 136999 14425
rect 149818 14422 149830 14425
rect 149882 14422 149894 14474
rect 141082 14359 141094 14362
rect 136953 14313 141094 14359
rect 141082 14310 141094 14313
rect 141146 14310 141158 14362
rect 147914 14310 147926 14362
rect 147978 14359 147990 14362
rect 147978 14313 191542 14359
rect 147978 14310 147990 14313
rect 102793 14201 113815 14247
rect 114202 14198 114214 14250
rect 114266 14247 114278 14250
rect 116330 14247 116342 14250
rect 114266 14201 116342 14247
rect 114266 14198 114278 14201
rect 116330 14198 116342 14201
rect 116394 14198 116406 14250
rect 116457 14201 117511 14247
rect 83738 14135 83750 14138
rect 82234 14089 83351 14135
rect 83417 14089 83750 14135
rect 82234 14086 82246 14089
rect 80826 14023 80838 14026
rect 75066 13977 79879 14023
rect 79945 13977 80838 14023
rect 75066 13974 75078 13977
rect 43642 13862 43654 13914
rect 43706 13911 43718 13914
rect 75114 13911 75126 13914
rect 43706 13865 75126 13911
rect 43706 13862 43718 13865
rect 75114 13862 75126 13865
rect 75178 13862 75190 13914
rect 79833 13911 79879 13977
rect 80826 13974 80838 13977
rect 80890 13974 80902 14026
rect 81050 13974 81062 14026
rect 81114 14023 81126 14026
rect 83417 14023 83463 14089
rect 83738 14086 83750 14089
rect 83802 14086 83814 14138
rect 84298 14086 84310 14138
rect 84362 14135 84374 14138
rect 91018 14135 91030 14138
rect 84362 14089 91030 14135
rect 84362 14086 84374 14089
rect 91018 14086 91030 14089
rect 91082 14086 91094 14138
rect 92698 14135 92710 14138
rect 91145 14089 92710 14135
rect 81114 13977 83463 14023
rect 81114 13974 81126 13977
rect 83514 13974 83526 14026
rect 83578 14023 83590 14026
rect 87210 14023 87222 14026
rect 83578 13977 87222 14023
rect 83578 13974 83590 13977
rect 87210 13974 87222 13977
rect 87274 13974 87286 14026
rect 88218 13974 88230 14026
rect 88282 14023 88294 14026
rect 90010 14023 90022 14026
rect 88282 13977 90022 14023
rect 88282 13974 88294 13977
rect 90010 13974 90022 13977
rect 90074 13974 90086 14026
rect 91145 14023 91191 14089
rect 92698 14086 92710 14089
rect 92762 14086 92774 14138
rect 92922 14086 92934 14138
rect 92986 14135 92998 14138
rect 97514 14135 97526 14138
rect 92986 14089 97526 14135
rect 92986 14086 92998 14089
rect 97514 14086 97526 14089
rect 97578 14086 97590 14138
rect 98074 14086 98086 14138
rect 98138 14135 98150 14138
rect 99194 14135 99206 14138
rect 98138 14089 99206 14135
rect 98138 14086 98150 14089
rect 99194 14086 99206 14089
rect 99258 14086 99270 14138
rect 99418 14086 99430 14138
rect 99482 14135 99494 14138
rect 116457 14135 116503 14201
rect 99482 14089 116503 14135
rect 99482 14086 99494 14089
rect 116666 14086 116678 14138
rect 116730 14135 116742 14138
rect 117338 14135 117350 14138
rect 116730 14089 117350 14135
rect 116730 14086 116742 14089
rect 117338 14086 117350 14089
rect 117402 14086 117414 14138
rect 117465 14135 117511 14201
rect 118682 14198 118694 14250
rect 118746 14198 118758 14250
rect 148698 14247 148710 14250
rect 118809 14201 148710 14247
rect 118809 14135 118855 14201
rect 148698 14198 148710 14201
rect 148762 14198 148774 14250
rect 149258 14198 149270 14250
rect 149322 14247 149334 14250
rect 149322 14201 179782 14247
rect 149322 14198 149334 14201
rect 117465 14089 118855 14135
rect 119242 14086 119254 14138
rect 119306 14135 119318 14138
rect 149370 14135 149382 14138
rect 119306 14089 149382 14135
rect 119306 14086 119318 14089
rect 149370 14086 149382 14089
rect 149434 14086 149446 14138
rect 176362 14135 176374 14138
rect 156216 14089 176374 14135
rect 90585 13977 91191 14023
rect 90585 13911 90631 13977
rect 91578 13974 91590 14026
rect 91642 14023 91654 14026
rect 102554 14023 102566 14026
rect 91642 13977 102566 14023
rect 91642 13974 91654 13977
rect 102554 13974 102566 13977
rect 102618 13974 102630 14026
rect 103898 13974 103910 14026
rect 103962 14023 103974 14026
rect 111178 14023 111190 14026
rect 103962 13977 111190 14023
rect 103962 13974 103974 13977
rect 111178 13974 111190 13977
rect 111242 13974 111254 14026
rect 111962 13974 111974 14026
rect 112026 14023 112038 14026
rect 112970 14023 112982 14026
rect 112026 13977 112982 14023
rect 112026 13974 112038 13977
rect 112970 13974 112982 13977
rect 113034 13974 113046 14026
rect 113418 13974 113430 14026
rect 113482 14023 113494 14026
rect 114202 14023 114214 14026
rect 113482 13977 114214 14023
rect 113482 13974 113494 13977
rect 114202 13974 114214 13977
rect 114266 13974 114278 14026
rect 114986 13974 114998 14026
rect 115050 14023 115062 14026
rect 120026 14023 120038 14026
rect 115050 13977 120038 14023
rect 115050 13974 115062 13977
rect 120026 13974 120038 13977
rect 120090 13974 120102 14026
rect 134138 14023 134150 14026
rect 120936 13977 134150 14023
rect 117114 13911 117126 13914
rect 75577 13865 79767 13911
rect 79833 13865 90631 13911
rect 90696 13865 117126 13911
rect 47562 13750 47574 13802
rect 47626 13799 47638 13802
rect 75450 13799 75462 13802
rect 47626 13753 75462 13799
rect 47626 13750 47638 13753
rect 75450 13750 75462 13753
rect 75514 13750 75526 13802
rect 6794 13638 6806 13690
rect 6858 13687 6870 13690
rect 55738 13687 55750 13690
rect 6858 13641 55750 13687
rect 6858 13638 6870 13641
rect 55738 13638 55750 13641
rect 55802 13638 55814 13690
rect 58202 13638 58214 13690
rect 58266 13687 58278 13690
rect 75577 13687 75623 13865
rect 75674 13750 75686 13802
rect 75738 13799 75750 13802
rect 79594 13799 79606 13802
rect 75738 13753 79606 13799
rect 75738 13750 75750 13753
rect 79594 13750 79606 13753
rect 79658 13750 79670 13802
rect 79721 13799 79767 13865
rect 82506 13799 82518 13802
rect 79721 13753 82518 13799
rect 82506 13750 82518 13753
rect 82570 13750 82582 13802
rect 82730 13799 82742 13802
rect 82633 13753 82742 13799
rect 58266 13641 75623 13687
rect 58266 13638 58278 13641
rect 75786 13638 75798 13690
rect 75850 13687 75862 13690
rect 82058 13687 82070 13690
rect 75850 13641 82070 13687
rect 75850 13638 75862 13641
rect 82058 13638 82070 13641
rect 82122 13638 82134 13690
rect 82185 13641 82342 13687
rect 54394 13526 54406 13578
rect 54458 13575 54470 13578
rect 82185 13575 82231 13641
rect 54458 13529 82231 13575
rect 82296 13575 82342 13641
rect 82394 13638 82406 13690
rect 82458 13687 82470 13690
rect 82633 13687 82679 13753
rect 82730 13750 82742 13753
rect 82794 13750 82806 13802
rect 82954 13750 82966 13802
rect 83018 13799 83030 13802
rect 84298 13799 84310 13802
rect 83018 13753 84310 13799
rect 83018 13750 83030 13753
rect 84298 13750 84310 13753
rect 84362 13750 84374 13802
rect 84522 13750 84534 13802
rect 84586 13799 84598 13802
rect 90696 13799 90742 13865
rect 117114 13862 117126 13865
rect 117178 13862 117190 13914
rect 117338 13862 117350 13914
rect 117402 13911 117414 13914
rect 119914 13911 119926 13914
rect 117402 13865 119926 13911
rect 117402 13862 117414 13865
rect 119914 13862 119926 13865
rect 119978 13862 119990 13914
rect 120936 13911 120982 13977
rect 134138 13974 134150 13977
rect 134202 13974 134214 14026
rect 138506 13974 138518 14026
rect 138570 14023 138582 14026
rect 156216 14023 156262 14089
rect 176362 14086 176374 14089
rect 176426 14086 176438 14138
rect 138570 13977 156262 14023
rect 179736 14023 179782 14201
rect 191496 14135 191542 14313
rect 196410 14135 196422 14138
rect 191496 14089 196422 14135
rect 196410 14086 196422 14089
rect 196474 14086 196486 14138
rect 197194 14023 197206 14026
rect 179736 13977 197206 14023
rect 138570 13974 138582 13977
rect 197194 13974 197206 13977
rect 197258 13974 197270 14026
rect 120041 13865 120982 13911
rect 84586 13753 90742 13799
rect 90809 13753 100711 13799
rect 84586 13750 84598 13753
rect 90809 13687 90855 13753
rect 100538 13687 100550 13690
rect 82458 13641 82679 13687
rect 82745 13641 90855 13687
rect 90921 13641 100550 13687
rect 82458 13638 82470 13641
rect 82745 13575 82791 13641
rect 82296 13529 82791 13575
rect 54458 13526 54470 13529
rect 82842 13526 82854 13578
rect 82906 13575 82918 13578
rect 90122 13575 90134 13578
rect 82906 13529 90134 13575
rect 82906 13526 82918 13529
rect 90122 13526 90134 13529
rect 90186 13526 90198 13578
rect 90346 13526 90358 13578
rect 90410 13575 90422 13578
rect 90921 13575 90967 13641
rect 100538 13638 100550 13641
rect 100602 13638 100614 13690
rect 100665 13687 100711 13753
rect 100986 13750 100998 13802
rect 101050 13799 101062 13802
rect 101322 13799 101334 13802
rect 101050 13753 101334 13799
rect 101050 13750 101062 13753
rect 101322 13750 101334 13753
rect 101386 13750 101398 13802
rect 101770 13750 101782 13802
rect 101834 13799 101846 13802
rect 102106 13799 102118 13802
rect 101834 13753 102118 13799
rect 101834 13750 101846 13753
rect 102106 13750 102118 13753
rect 102170 13750 102182 13802
rect 103129 13753 103287 13799
rect 102442 13687 102454 13690
rect 100665 13641 102454 13687
rect 102442 13638 102454 13641
rect 102506 13638 102518 13690
rect 103129 13687 103175 13753
rect 102961 13641 103175 13687
rect 103241 13687 103287 13753
rect 104570 13750 104582 13802
rect 104634 13799 104646 13802
rect 119354 13799 119366 13802
rect 104634 13753 119366 13799
rect 104634 13750 104646 13753
rect 119354 13750 119366 13753
rect 119418 13750 119430 13802
rect 119578 13750 119590 13802
rect 119642 13799 119654 13802
rect 120041 13799 120087 13865
rect 121034 13862 121046 13914
rect 121098 13911 121110 13914
rect 122490 13911 122502 13914
rect 121098 13865 122502 13911
rect 121098 13862 121110 13865
rect 122490 13862 122502 13865
rect 122554 13862 122566 13914
rect 122938 13862 122950 13914
rect 123002 13911 123014 13914
rect 125962 13911 125974 13914
rect 123002 13865 125974 13911
rect 123002 13862 123014 13865
rect 125962 13862 125974 13865
rect 126026 13862 126038 13914
rect 126186 13862 126198 13914
rect 126250 13911 126262 13914
rect 134250 13911 134262 13914
rect 126250 13865 134262 13911
rect 126250 13862 126262 13865
rect 134250 13862 134262 13865
rect 134314 13862 134326 13914
rect 134698 13862 134710 13914
rect 134762 13911 134774 13914
rect 142874 13911 142886 13914
rect 134762 13865 142886 13911
rect 134762 13862 134774 13865
rect 142874 13862 142886 13865
rect 142938 13862 142950 13914
rect 143210 13862 143222 13914
rect 143274 13911 143286 13914
rect 212762 13911 212774 13914
rect 143274 13865 212774 13911
rect 143274 13862 143286 13865
rect 212762 13862 212774 13865
rect 212826 13862 212838 13914
rect 119642 13753 120087 13799
rect 119642 13750 119654 13753
rect 120250 13750 120262 13802
rect 120314 13799 120326 13802
rect 120314 13753 146743 13799
rect 120314 13750 120326 13753
rect 103241 13641 103399 13687
rect 90410 13529 90967 13575
rect 90410 13526 90422 13529
rect 91018 13526 91030 13578
rect 91082 13575 91094 13578
rect 102961 13575 103007 13641
rect 91082 13529 103007 13575
rect 103353 13575 103399 13641
rect 103450 13638 103462 13690
rect 103514 13687 103526 13690
rect 118458 13687 118470 13690
rect 103514 13641 118470 13687
rect 103514 13638 103526 13641
rect 118458 13638 118470 13641
rect 118522 13638 118534 13690
rect 118682 13638 118694 13690
rect 118746 13687 118758 13690
rect 118746 13641 144502 13687
rect 118746 13638 118758 13641
rect 116218 13575 116230 13578
rect 103353 13529 116230 13575
rect 91082 13526 91094 13529
rect 116218 13526 116230 13529
rect 116282 13526 116294 13578
rect 116442 13526 116454 13578
rect 116506 13575 116518 13578
rect 138506 13575 138518 13578
rect 116506 13529 138518 13575
rect 116506 13526 116518 13529
rect 138506 13526 138518 13529
rect 138570 13526 138582 13578
rect 139066 13575 139078 13578
rect 138633 13529 139078 13575
rect 53834 13414 53846 13466
rect 53898 13463 53910 13466
rect 75786 13463 75798 13466
rect 53898 13417 75798 13463
rect 53898 13414 53910 13417
rect 75786 13414 75798 13417
rect 75850 13414 75862 13466
rect 76010 13414 76022 13466
rect 76074 13463 76086 13466
rect 76074 13417 82455 13463
rect 76074 13414 76086 13417
rect 49802 13302 49814 13354
rect 49866 13351 49878 13354
rect 49866 13305 82342 13351
rect 49866 13302 49878 13305
rect 55962 13190 55974 13242
rect 56026 13239 56038 13242
rect 56026 13193 68007 13239
rect 56026 13190 56038 13193
rect 74 13078 86 13130
rect 138 13127 150 13130
rect 67498 13127 67510 13130
rect 138 13081 67510 13127
rect 138 13078 150 13081
rect 67498 13078 67510 13081
rect 67562 13078 67574 13130
rect 41066 12966 41078 13018
rect 41130 13015 41142 13018
rect 67834 13015 67846 13018
rect 41130 12969 67846 13015
rect 41130 12966 41142 12969
rect 67834 12966 67846 12969
rect 67898 12966 67910 13018
rect 67961 13015 68007 13193
rect 68394 13190 68406 13242
rect 68458 13239 68470 13242
rect 79034 13239 79046 13242
rect 68458 13193 79046 13239
rect 68458 13190 68470 13193
rect 79034 13190 79046 13193
rect 79098 13190 79110 13242
rect 79594 13190 79606 13242
rect 79658 13239 79670 13242
rect 80826 13239 80838 13242
rect 79658 13193 80838 13239
rect 79658 13190 79670 13193
rect 80826 13190 80838 13193
rect 80890 13190 80902 13242
rect 81162 13190 81174 13242
rect 81226 13239 81238 13242
rect 81722 13239 81734 13242
rect 81226 13193 81734 13239
rect 81226 13190 81238 13193
rect 81722 13190 81734 13193
rect 81786 13190 81798 13242
rect 68058 13078 68070 13130
rect 68122 13127 68134 13130
rect 80714 13127 80726 13130
rect 68122 13081 80726 13127
rect 68122 13078 68134 13081
rect 80714 13078 80726 13081
rect 80778 13078 80790 13130
rect 82170 13127 82182 13130
rect 80841 13081 82182 13127
rect 73770 13015 73782 13018
rect 67961 12969 73782 13015
rect 73770 12966 73782 12969
rect 73834 12966 73846 13018
rect 74442 13015 74454 13018
rect 73896 12969 74454 13015
rect 43194 12854 43206 12906
rect 43258 12903 43270 12906
rect 68058 12903 68070 12906
rect 43258 12857 68070 12903
rect 43258 12854 43270 12857
rect 68058 12854 68070 12857
rect 68122 12854 68134 12906
rect 69962 12854 69974 12906
rect 70026 12903 70038 12906
rect 73896 12903 73942 12969
rect 74442 12966 74454 12969
rect 74506 12966 74518 13018
rect 75114 12966 75126 13018
rect 75178 13015 75190 13018
rect 78698 13015 78710 13018
rect 75178 12969 78710 13015
rect 75178 12966 75190 12969
rect 78698 12966 78710 12969
rect 78762 12966 78774 13018
rect 78922 12966 78934 13018
rect 78986 13015 78998 13018
rect 80841 13015 80887 13081
rect 82170 13078 82182 13081
rect 82234 13078 82246 13130
rect 82296 13015 82342 13305
rect 82409 13127 82455 13417
rect 83178 13414 83190 13466
rect 83242 13463 83254 13466
rect 90234 13463 90246 13466
rect 83242 13417 90246 13463
rect 83242 13414 83254 13417
rect 90234 13414 90246 13417
rect 90298 13414 90310 13466
rect 90794 13414 90806 13466
rect 90858 13463 90870 13466
rect 103338 13463 103350 13466
rect 90858 13417 103350 13463
rect 90858 13414 90870 13417
rect 103338 13414 103350 13417
rect 103402 13414 103414 13466
rect 104122 13414 104134 13466
rect 104186 13463 104198 13466
rect 138633 13463 138679 13529
rect 139066 13526 139078 13529
rect 139130 13526 139142 13578
rect 139514 13526 139526 13578
rect 139578 13575 139590 13578
rect 143210 13575 143222 13578
rect 139578 13529 143222 13575
rect 139578 13526 139590 13529
rect 143210 13526 143222 13529
rect 143274 13526 143286 13578
rect 104186 13417 138679 13463
rect 104186 13414 104198 13417
rect 138730 13414 138742 13466
rect 138794 13463 138806 13466
rect 140634 13463 140646 13466
rect 138794 13417 140646 13463
rect 138794 13414 138806 13417
rect 140634 13414 140646 13417
rect 140698 13414 140710 13466
rect 144456 13463 144502 13641
rect 146697 13575 146743 13753
rect 149146 13750 149158 13802
rect 149210 13799 149222 13802
rect 153178 13799 153190 13802
rect 149210 13753 153190 13799
rect 149210 13750 149222 13753
rect 153178 13750 153190 13753
rect 153242 13750 153254 13802
rect 159226 13750 159238 13802
rect 159290 13799 159302 13802
rect 178266 13799 178278 13802
rect 159290 13753 178278 13799
rect 159290 13750 159302 13753
rect 178266 13750 178278 13753
rect 178330 13750 178342 13802
rect 149370 13638 149382 13690
rect 149434 13687 149446 13690
rect 210410 13687 210422 13690
rect 149434 13641 210422 13687
rect 149434 13638 149446 13641
rect 210410 13638 210422 13641
rect 210474 13638 210486 13690
rect 146697 13529 156262 13575
rect 148362 13463 148374 13466
rect 144456 13417 148374 13463
rect 148362 13414 148374 13417
rect 148426 13414 148438 13466
rect 156216 13463 156262 13529
rect 161242 13526 161254 13578
rect 161306 13575 161318 13578
rect 182522 13575 182534 13578
rect 161306 13529 182534 13575
rect 161306 13526 161318 13529
rect 182522 13526 182534 13529
rect 182586 13526 182598 13578
rect 184538 13463 184550 13466
rect 156216 13417 184550 13463
rect 184538 13414 184550 13417
rect 184602 13414 184614 13466
rect 82730 13302 82742 13354
rect 82794 13351 82806 13354
rect 84186 13351 84198 13354
rect 82794 13305 84198 13351
rect 82794 13302 82806 13305
rect 84186 13302 84198 13305
rect 84250 13302 84262 13354
rect 84410 13302 84422 13354
rect 84474 13351 84486 13354
rect 84474 13305 114823 13351
rect 84474 13302 84486 13305
rect 103226 13239 103238 13242
rect 82633 13193 103238 13239
rect 82633 13127 82679 13193
rect 103226 13190 103238 13193
rect 103290 13190 103302 13242
rect 114650 13239 114662 13242
rect 103353 13193 114662 13239
rect 82409 13081 82679 13127
rect 82730 13078 82742 13130
rect 82794 13127 82806 13130
rect 101098 13127 101110 13130
rect 82794 13081 101110 13127
rect 82794 13078 82806 13081
rect 101098 13078 101110 13081
rect 101162 13078 101174 13130
rect 102554 13078 102566 13130
rect 102618 13127 102630 13130
rect 103353 13127 103399 13193
rect 114650 13190 114662 13193
rect 114714 13190 114726 13242
rect 114777 13239 114823 13305
rect 115210 13302 115222 13354
rect 115274 13351 115286 13354
rect 149146 13351 149158 13354
rect 115274 13305 149158 13351
rect 115274 13302 115286 13305
rect 149146 13302 149158 13305
rect 149210 13302 149222 13354
rect 149370 13302 149382 13354
rect 149434 13351 149446 13354
rect 211642 13351 211654 13354
rect 149434 13305 211654 13351
rect 149434 13302 149446 13305
rect 211642 13302 211654 13305
rect 211706 13302 211718 13354
rect 138954 13239 138966 13242
rect 114777 13193 138966 13239
rect 138954 13190 138966 13193
rect 139018 13190 139030 13242
rect 144442 13190 144454 13242
rect 144506 13239 144518 13242
rect 149482 13239 149494 13242
rect 144506 13193 149494 13239
rect 144506 13190 144518 13193
rect 149482 13190 149494 13193
rect 149546 13190 149558 13242
rect 151050 13190 151062 13242
rect 151114 13239 151126 13242
rect 155306 13239 155318 13242
rect 151114 13193 155318 13239
rect 151114 13190 151126 13193
rect 155306 13190 155318 13193
rect 155370 13190 155382 13242
rect 165050 13190 165062 13242
rect 165114 13239 165126 13242
rect 173674 13239 173686 13242
rect 165114 13193 173686 13239
rect 165114 13190 165126 13193
rect 173674 13190 173686 13193
rect 173738 13190 173750 13242
rect 102618 13081 103399 13127
rect 102618 13078 102630 13081
rect 103450 13078 103462 13130
rect 103514 13127 103526 13130
rect 120586 13127 120598 13130
rect 103514 13081 120598 13127
rect 103514 13078 103526 13081
rect 120586 13078 120598 13081
rect 120650 13078 120662 13130
rect 120810 13078 120822 13130
rect 120874 13127 120886 13130
rect 126186 13127 126198 13130
rect 120874 13081 126198 13127
rect 120874 13078 120886 13081
rect 126186 13078 126198 13081
rect 126250 13078 126262 13130
rect 126746 13078 126758 13130
rect 126810 13127 126822 13130
rect 142650 13127 142662 13130
rect 126810 13081 142662 13127
rect 126810 13078 126822 13081
rect 142650 13078 142662 13081
rect 142714 13078 142726 13130
rect 149258 13078 149270 13130
rect 149322 13127 149334 13130
rect 185882 13127 185894 13130
rect 149322 13081 185894 13127
rect 149322 13078 149334 13081
rect 185882 13078 185894 13081
rect 185946 13078 185958 13130
rect 99418 13015 99430 13018
rect 78986 12969 80887 13015
rect 81737 12969 82119 13015
rect 82296 12969 99430 13015
rect 78986 12966 78998 12969
rect 70026 12857 73942 12903
rect 70026 12854 70038 12857
rect 73994 12854 74006 12906
rect 74058 12903 74070 12906
rect 77354 12903 77366 12906
rect 74058 12857 77366 12903
rect 74058 12854 74070 12857
rect 77354 12854 77366 12857
rect 77418 12854 77430 12906
rect 77802 12854 77814 12906
rect 77866 12903 77878 12906
rect 81737 12903 81783 12969
rect 77866 12857 81783 12903
rect 77866 12854 77878 12857
rect 81946 12854 81958 12906
rect 82010 12854 82022 12906
rect 82073 12903 82119 12969
rect 99418 12966 99430 12969
rect 99482 12966 99494 13018
rect 102778 13015 102790 13018
rect 99545 12969 102790 13015
rect 88442 12903 88454 12906
rect 82073 12857 88454 12903
rect 88442 12854 88454 12857
rect 88506 12854 88518 12906
rect 88666 12854 88678 12906
rect 88730 12903 88742 12906
rect 89450 12903 89462 12906
rect 88730 12857 89462 12903
rect 88730 12854 88742 12857
rect 89450 12854 89462 12857
rect 89514 12854 89526 12906
rect 89786 12854 89798 12906
rect 89850 12903 89862 12906
rect 99545 12903 99591 12969
rect 102778 12966 102790 12969
rect 102842 12966 102854 13018
rect 103002 12966 103014 13018
rect 103066 13015 103078 13018
rect 103786 13015 103798 13018
rect 103066 12969 103798 13015
rect 103066 12966 103078 12969
rect 103786 12966 103798 12969
rect 103850 12966 103862 13018
rect 104010 12966 104022 13018
rect 104074 13015 104086 13018
rect 117226 13015 117238 13018
rect 104074 12969 117238 13015
rect 104074 12966 104086 12969
rect 117226 12966 117238 12969
rect 117290 12966 117302 13018
rect 117450 12966 117462 13018
rect 117514 13015 117526 13018
rect 122266 13015 122278 13018
rect 117514 12969 122278 13015
rect 117514 12966 117526 12969
rect 122266 12966 122278 12969
rect 122330 12966 122342 13018
rect 122490 12966 122502 13018
rect 122554 13015 122566 13018
rect 138170 13015 138182 13018
rect 122554 12969 138182 13015
rect 122554 12966 122566 12969
rect 138170 12966 138182 12969
rect 138234 12966 138246 13018
rect 138394 12966 138406 13018
rect 138458 13015 138470 13018
rect 142314 13015 142326 13018
rect 138458 12969 142326 13015
rect 138458 12966 138470 12969
rect 142314 12966 142326 12969
rect 142378 12966 142390 13018
rect 148586 12966 148598 13018
rect 148650 13015 148662 13018
rect 186554 13015 186566 13018
rect 148650 12969 186566 13015
rect 148650 12966 148662 12969
rect 186554 12966 186566 12969
rect 186618 12966 186630 13018
rect 89850 12857 99591 12903
rect 89850 12854 89862 12857
rect 99642 12854 99654 12906
rect 99706 12903 99718 12906
rect 102330 12903 102342 12906
rect 99706 12857 102342 12903
rect 99706 12854 99718 12857
rect 102330 12854 102342 12857
rect 102394 12854 102406 12906
rect 102554 12854 102566 12906
rect 102618 12903 102630 12906
rect 102890 12903 102902 12906
rect 102618 12857 102902 12903
rect 102618 12854 102630 12857
rect 102890 12854 102902 12857
rect 102954 12854 102966 12906
rect 104794 12903 104806 12906
rect 103017 12857 104806 12903
rect 5338 12742 5350 12794
rect 5402 12791 5414 12794
rect 56970 12791 56982 12794
rect 5402 12745 56982 12791
rect 5402 12742 5414 12745
rect 56970 12742 56982 12745
rect 57034 12742 57046 12794
rect 58538 12742 58550 12794
rect 58602 12791 58614 12794
rect 81961 12791 82007 12854
rect 58602 12745 82007 12791
rect 58602 12742 58614 12745
rect 82394 12742 82406 12794
rect 82458 12791 82470 12794
rect 103017 12791 103063 12857
rect 104794 12854 104806 12857
rect 104858 12854 104870 12906
rect 109162 12854 109174 12906
rect 109226 12903 109238 12906
rect 109834 12903 109846 12906
rect 109226 12857 109846 12903
rect 109226 12854 109238 12857
rect 109834 12854 109846 12857
rect 109898 12854 109910 12906
rect 110842 12854 110854 12906
rect 110906 12903 110918 12906
rect 114426 12903 114438 12906
rect 110906 12857 114438 12903
rect 110906 12854 110918 12857
rect 114426 12854 114438 12857
rect 114490 12854 114502 12906
rect 114650 12854 114662 12906
rect 114714 12903 114726 12906
rect 121594 12903 121606 12906
rect 114714 12857 121606 12903
rect 114714 12854 114726 12857
rect 121594 12854 121606 12857
rect 121658 12854 121670 12906
rect 125850 12854 125862 12906
rect 125914 12903 125926 12906
rect 126746 12903 126758 12906
rect 125914 12857 126758 12903
rect 125914 12854 125926 12857
rect 126746 12854 126758 12857
rect 126810 12854 126822 12906
rect 127418 12854 127430 12906
rect 127482 12903 127494 12906
rect 149034 12903 149046 12906
rect 127482 12857 149046 12903
rect 127482 12854 127494 12857
rect 149034 12854 149046 12857
rect 149098 12854 149110 12906
rect 149258 12854 149270 12906
rect 149322 12903 149334 12906
rect 188458 12903 188470 12906
rect 149322 12857 188470 12903
rect 149322 12854 149334 12857
rect 188458 12854 188470 12857
rect 188522 12854 188534 12906
rect 82458 12745 103063 12791
rect 82458 12742 82470 12745
rect 103114 12742 103126 12794
rect 103178 12791 103190 12794
rect 114538 12791 114550 12794
rect 103178 12745 114550 12791
rect 103178 12742 103190 12745
rect 114538 12742 114550 12745
rect 114602 12742 114614 12794
rect 114721 12745 115159 12791
rect 29418 12630 29430 12682
rect 29482 12679 29494 12682
rect 71754 12679 71766 12682
rect 29482 12633 71766 12679
rect 29482 12630 29494 12633
rect 71754 12630 71766 12633
rect 71818 12630 71830 12682
rect 71978 12630 71990 12682
rect 72042 12679 72054 12682
rect 76794 12679 76806 12682
rect 72042 12633 76806 12679
rect 72042 12630 72054 12633
rect 76794 12630 76806 12633
rect 76858 12630 76870 12682
rect 77369 12633 78647 12679
rect 56410 12518 56422 12570
rect 56474 12567 56486 12570
rect 77369 12567 77415 12633
rect 78601 12567 78647 12633
rect 78698 12630 78710 12682
rect 78762 12679 78774 12682
rect 80602 12679 80614 12682
rect 78762 12633 80614 12679
rect 78762 12630 78774 12633
rect 80602 12630 80614 12633
rect 80666 12630 80678 12682
rect 80826 12630 80838 12682
rect 80890 12679 80902 12682
rect 80890 12633 81335 12679
rect 80890 12630 80902 12633
rect 81289 12567 81335 12633
rect 81386 12630 81398 12682
rect 81450 12679 81462 12682
rect 84522 12679 84534 12682
rect 81450 12633 84534 12679
rect 81450 12630 81462 12633
rect 84522 12630 84534 12633
rect 84586 12630 84598 12682
rect 84858 12630 84870 12682
rect 84922 12679 84934 12682
rect 102666 12679 102678 12682
rect 84922 12633 102678 12679
rect 84922 12630 84934 12633
rect 102666 12630 102678 12633
rect 102730 12630 102742 12682
rect 103562 12679 103574 12682
rect 102793 12633 103574 12679
rect 82282 12567 82294 12570
rect 56474 12521 77415 12567
rect 77481 12521 78087 12567
rect 78601 12521 81223 12567
rect 81289 12521 82294 12567
rect 56474 12518 56486 12521
rect 51930 12406 51942 12458
rect 51994 12455 52006 12458
rect 77481 12455 77527 12521
rect 77914 12455 77926 12458
rect 51994 12409 77527 12455
rect 77593 12409 77926 12455
rect 51994 12406 52006 12409
rect 54170 12294 54182 12346
rect 54234 12343 54246 12346
rect 75226 12343 75238 12346
rect 54234 12297 75238 12343
rect 54234 12294 54246 12297
rect 75226 12294 75238 12297
rect 75290 12294 75302 12346
rect 77593 12343 77639 12409
rect 77914 12406 77926 12409
rect 77978 12406 77990 12458
rect 78041 12455 78087 12521
rect 79930 12455 79942 12458
rect 78041 12409 79942 12455
rect 79930 12406 79942 12409
rect 79994 12406 80006 12458
rect 80602 12406 80614 12458
rect 80666 12455 80678 12458
rect 81050 12455 81062 12458
rect 80666 12409 81062 12455
rect 80666 12406 80678 12409
rect 81050 12406 81062 12409
rect 81114 12406 81126 12458
rect 81177 12455 81223 12521
rect 82282 12518 82294 12521
rect 82346 12518 82358 12570
rect 83066 12518 83078 12570
rect 83130 12567 83142 12570
rect 87882 12567 87894 12570
rect 83130 12521 87894 12567
rect 83130 12518 83142 12521
rect 87882 12518 87894 12521
rect 87946 12518 87958 12570
rect 102793 12567 102839 12633
rect 103562 12630 103574 12633
rect 103626 12630 103638 12682
rect 114721 12679 114767 12745
rect 103689 12633 114767 12679
rect 89913 12521 102839 12567
rect 81177 12409 81335 12455
rect 76361 12297 77639 12343
rect 4666 12182 4678 12234
rect 4730 12231 4742 12234
rect 64474 12231 64486 12234
rect 4730 12185 64486 12231
rect 4730 12182 4742 12185
rect 64474 12182 64486 12185
rect 64538 12182 64550 12234
rect 67722 12182 67734 12234
rect 67786 12231 67798 12234
rect 69626 12231 69638 12234
rect 67786 12185 69638 12231
rect 67786 12182 67798 12185
rect 69626 12182 69638 12185
rect 69690 12182 69702 12234
rect 69850 12182 69862 12234
rect 69914 12231 69926 12234
rect 76361 12231 76407 12297
rect 78250 12294 78262 12346
rect 78314 12343 78326 12346
rect 78314 12297 78535 12343
rect 78314 12294 78326 12297
rect 69914 12185 76407 12231
rect 69914 12182 69926 12185
rect 76682 12182 76694 12234
rect 76746 12231 76758 12234
rect 78362 12231 78374 12234
rect 76746 12185 78374 12231
rect 76746 12182 76758 12185
rect 78362 12182 78374 12185
rect 78426 12182 78438 12234
rect 78489 12231 78535 12297
rect 78586 12294 78598 12346
rect 78650 12343 78662 12346
rect 80266 12343 80278 12346
rect 78650 12297 80278 12343
rect 78650 12294 78662 12297
rect 80266 12294 80278 12297
rect 80330 12294 80342 12346
rect 81289 12343 81335 12409
rect 81722 12406 81734 12458
rect 81786 12455 81798 12458
rect 89786 12455 89798 12458
rect 81786 12409 89798 12455
rect 81786 12406 81798 12409
rect 89786 12406 89798 12409
rect 89850 12406 89862 12458
rect 89913 12343 89959 12521
rect 102890 12518 102902 12570
rect 102954 12567 102966 12570
rect 103689 12567 103735 12633
rect 114986 12630 114998 12682
rect 115050 12630 115062 12682
rect 115113 12679 115159 12745
rect 115546 12742 115558 12794
rect 115610 12791 115622 12794
rect 142650 12791 142662 12794
rect 115610 12745 142662 12791
rect 115610 12742 115622 12745
rect 142650 12742 142662 12745
rect 142714 12742 142726 12794
rect 142874 12742 142886 12794
rect 142938 12791 142950 12794
rect 188570 12791 188582 12794
rect 142938 12745 188582 12791
rect 142938 12742 142950 12745
rect 188570 12742 188582 12745
rect 188634 12742 188646 12794
rect 138394 12679 138406 12682
rect 115113 12633 138406 12679
rect 138394 12630 138406 12633
rect 138458 12630 138470 12682
rect 139066 12630 139078 12682
rect 139130 12679 139142 12682
rect 189802 12679 189814 12682
rect 139130 12633 189814 12679
rect 139130 12630 139142 12633
rect 189802 12630 189814 12633
rect 189866 12630 189878 12682
rect 102954 12521 103735 12567
rect 102954 12518 102966 12521
rect 104122 12518 104134 12570
rect 104186 12567 104198 12570
rect 114874 12567 114886 12570
rect 104186 12521 114886 12567
rect 104186 12518 104198 12521
rect 114874 12518 114886 12521
rect 114938 12518 114950 12570
rect 115001 12567 115047 12630
rect 116554 12567 116566 12570
rect 115001 12521 116566 12567
rect 116554 12518 116566 12521
rect 116618 12518 116630 12570
rect 119578 12567 119590 12570
rect 116681 12521 119590 12567
rect 116681 12455 116727 12521
rect 119578 12518 119590 12521
rect 119642 12518 119654 12570
rect 119914 12518 119926 12570
rect 119978 12567 119990 12570
rect 120810 12567 120822 12570
rect 119978 12521 120822 12567
rect 119978 12518 119990 12521
rect 120810 12518 120822 12521
rect 120874 12518 120886 12570
rect 120936 12521 145287 12567
rect 81289 12297 89959 12343
rect 90025 12409 116727 12455
rect 78489 12185 80327 12231
rect 20682 12070 20694 12122
rect 20746 12119 20758 12122
rect 63690 12119 63702 12122
rect 20746 12073 63702 12119
rect 20746 12070 20758 12073
rect 63690 12070 63702 12073
rect 63754 12070 63766 12122
rect 65146 12070 65158 12122
rect 65210 12119 65222 12122
rect 80281 12119 80327 12185
rect 80714 12182 80726 12234
rect 80778 12231 80790 12234
rect 81946 12231 81958 12234
rect 80778 12185 81958 12231
rect 80778 12182 80790 12185
rect 81946 12182 81958 12185
rect 82010 12182 82022 12234
rect 90025 12231 90071 12409
rect 116778 12406 116790 12458
rect 116842 12455 116854 12458
rect 118458 12455 118470 12458
rect 116842 12409 118470 12455
rect 116842 12406 116854 12409
rect 118458 12406 118470 12409
rect 118522 12406 118534 12458
rect 118682 12406 118694 12458
rect 118746 12455 118758 12458
rect 120936 12455 120982 12521
rect 118746 12409 120982 12455
rect 118746 12406 118758 12409
rect 121034 12406 121046 12458
rect 121098 12455 121110 12458
rect 145114 12455 145126 12458
rect 121098 12409 145126 12455
rect 121098 12406 121110 12409
rect 145114 12406 145126 12409
rect 145178 12406 145190 12458
rect 90234 12294 90246 12346
rect 90298 12343 90310 12346
rect 103338 12343 103350 12346
rect 90298 12297 103350 12343
rect 90298 12294 90310 12297
rect 103338 12294 103350 12297
rect 103402 12294 103414 12346
rect 103674 12294 103686 12346
rect 103738 12343 103750 12346
rect 145241 12343 145287 12521
rect 148698 12518 148710 12570
rect 148762 12567 148774 12570
rect 149258 12567 149270 12570
rect 148762 12521 149270 12567
rect 148762 12518 148774 12521
rect 149258 12518 149270 12521
rect 149322 12518 149334 12570
rect 152842 12518 152854 12570
rect 152906 12567 152918 12570
rect 196298 12567 196310 12570
rect 152906 12521 196310 12567
rect 152906 12518 152918 12521
rect 196298 12518 196310 12521
rect 196362 12518 196374 12570
rect 145338 12406 145350 12458
rect 145402 12455 145414 12458
rect 150378 12455 150390 12458
rect 145402 12409 150390 12455
rect 145402 12406 145414 12409
rect 150378 12406 150390 12409
rect 150442 12406 150454 12458
rect 162810 12406 162822 12458
rect 162874 12455 162886 12458
rect 209290 12455 209302 12458
rect 162874 12409 209302 12455
rect 162874 12406 162886 12409
rect 209290 12406 209302 12409
rect 209354 12406 209366 12458
rect 193050 12343 193062 12346
rect 103738 12297 145175 12343
rect 145241 12297 193062 12343
rect 103738 12294 103750 12297
rect 82185 12185 90071 12231
rect 80826 12119 80838 12122
rect 65210 12073 80215 12119
rect 80281 12073 80838 12119
rect 65210 12070 65222 12073
rect 43530 11958 43542 12010
rect 43594 12007 43606 12010
rect 58314 12007 58326 12010
rect 43594 11961 58326 12007
rect 43594 11958 43606 11961
rect 58314 11958 58326 11961
rect 58378 11958 58390 12010
rect 61226 11958 61238 12010
rect 61290 12007 61302 12010
rect 68282 12007 68294 12010
rect 61290 11961 68294 12007
rect 61290 11958 61302 11961
rect 68282 11958 68294 11961
rect 68346 11958 68358 12010
rect 69514 11958 69526 12010
rect 69578 12007 69590 12010
rect 69578 11961 77751 12007
rect 69578 11958 69590 11961
rect 55178 11846 55190 11898
rect 55242 11895 55254 11898
rect 67834 11895 67846 11898
rect 55242 11849 67846 11895
rect 55242 11846 55254 11849
rect 67834 11846 67846 11849
rect 67898 11846 67910 11898
rect 73210 11895 73222 11898
rect 67961 11849 73222 11895
rect 33786 11734 33798 11786
rect 33850 11783 33862 11786
rect 57082 11783 57094 11786
rect 33850 11737 57094 11783
rect 33850 11734 33862 11737
rect 57082 11734 57094 11737
rect 57146 11734 57158 11786
rect 65706 11783 65718 11786
rect 58776 11737 65718 11783
rect 56970 11622 56982 11674
rect 57034 11671 57046 11674
rect 58776 11671 58822 11737
rect 65706 11734 65718 11737
rect 65770 11734 65782 11786
rect 67961 11671 68007 11849
rect 73210 11846 73222 11849
rect 73274 11846 73286 11898
rect 74106 11895 74118 11898
rect 73337 11849 74118 11895
rect 68058 11734 68070 11786
rect 68122 11783 68134 11786
rect 73337 11783 73383 11849
rect 74106 11846 74118 11849
rect 74170 11846 74182 11898
rect 74666 11846 74678 11898
rect 74730 11895 74742 11898
rect 77578 11895 77590 11898
rect 74730 11849 77590 11895
rect 74730 11846 74742 11849
rect 77578 11846 77590 11849
rect 77642 11846 77654 11898
rect 77705 11895 77751 11961
rect 77802 11958 77814 12010
rect 77866 12007 77878 12010
rect 79594 12007 79606 12010
rect 77866 11961 79606 12007
rect 77866 11958 77878 11961
rect 79594 11958 79606 11961
rect 79658 11958 79670 12010
rect 80169 12007 80215 12073
rect 80826 12070 80838 12073
rect 80890 12070 80902 12122
rect 82058 12119 82070 12122
rect 80953 12073 82070 12119
rect 80169 11961 80327 12007
rect 80281 11898 80327 11961
rect 80602 11958 80614 12010
rect 80666 12007 80678 12010
rect 80953 12007 80999 12073
rect 82058 12070 82070 12073
rect 82122 12070 82134 12122
rect 80666 11961 80999 12007
rect 80666 11958 80678 11961
rect 81050 11958 81062 12010
rect 81114 12007 81126 12010
rect 81946 12007 81958 12010
rect 81114 11961 81958 12007
rect 81114 11958 81126 11961
rect 81946 11958 81958 11961
rect 82010 11958 82022 12010
rect 82185 12007 82231 12185
rect 90122 12182 90134 12234
rect 90186 12231 90198 12234
rect 98186 12231 98198 12234
rect 90186 12185 98198 12231
rect 90186 12182 90198 12185
rect 98186 12182 98198 12185
rect 98250 12182 98262 12234
rect 98522 12182 98534 12234
rect 98586 12231 98598 12234
rect 103226 12231 103238 12234
rect 98586 12185 103238 12231
rect 98586 12182 98598 12185
rect 103226 12182 103238 12185
rect 103290 12182 103302 12234
rect 103450 12182 103462 12234
rect 103514 12231 103526 12234
rect 115210 12231 115222 12234
rect 103514 12185 115222 12231
rect 103514 12182 103526 12185
rect 115210 12182 115222 12185
rect 115274 12182 115286 12234
rect 116666 12182 116678 12234
rect 116730 12231 116742 12234
rect 117002 12231 117014 12234
rect 116730 12185 117014 12231
rect 116730 12182 116742 12185
rect 117002 12182 117014 12185
rect 117066 12182 117078 12234
rect 117226 12182 117238 12234
rect 117290 12231 117302 12234
rect 144442 12231 144454 12234
rect 117290 12185 144454 12231
rect 117290 12182 117302 12185
rect 144442 12182 144454 12185
rect 144506 12182 144518 12234
rect 145129 12231 145175 12297
rect 193050 12294 193062 12297
rect 193114 12294 193126 12346
rect 148586 12231 148598 12234
rect 145129 12185 148598 12231
rect 148586 12182 148598 12185
rect 148650 12182 148662 12234
rect 158778 12182 158790 12234
rect 158842 12231 158854 12234
rect 175914 12231 175926 12234
rect 158842 12185 175926 12231
rect 158842 12182 158854 12185
rect 175914 12182 175926 12185
rect 175978 12182 175990 12234
rect 82730 12070 82742 12122
rect 82794 12119 82806 12122
rect 83290 12119 83302 12122
rect 82794 12073 83302 12119
rect 82794 12070 82806 12073
rect 83290 12070 83302 12073
rect 83354 12070 83366 12122
rect 83738 12070 83750 12122
rect 83802 12119 83814 12122
rect 91354 12119 91366 12122
rect 83802 12073 91366 12119
rect 83802 12070 83814 12073
rect 91354 12070 91366 12073
rect 91418 12070 91430 12122
rect 102890 12119 102902 12122
rect 91481 12073 102902 12119
rect 82073 11961 82231 12007
rect 77705 11849 80103 11895
rect 68122 11737 73383 11783
rect 68122 11734 68134 11737
rect 73546 11734 73558 11786
rect 73610 11783 73622 11786
rect 80057 11783 80103 11849
rect 80266 11846 80278 11898
rect 80330 11846 80342 11898
rect 81274 11895 81286 11898
rect 80393 11849 81286 11895
rect 80393 11783 80439 11849
rect 81274 11846 81286 11849
rect 81338 11846 81350 11898
rect 81834 11846 81846 11898
rect 81898 11895 81910 11898
rect 82073 11895 82119 11961
rect 82506 11958 82518 12010
rect 82570 12007 82582 12010
rect 91481 12007 91527 12073
rect 102890 12070 102902 12073
rect 102954 12070 102966 12122
rect 103114 12070 103126 12122
rect 103178 12119 103190 12122
rect 114538 12119 114550 12122
rect 103178 12073 114550 12119
rect 103178 12070 103190 12073
rect 114538 12070 114550 12073
rect 114602 12070 114614 12122
rect 114762 12070 114774 12122
rect 114826 12119 114838 12122
rect 115658 12119 115670 12122
rect 114826 12073 115670 12119
rect 114826 12070 114838 12073
rect 115658 12070 115670 12073
rect 115722 12070 115734 12122
rect 115882 12070 115894 12122
rect 115946 12119 115958 12122
rect 122490 12119 122502 12122
rect 115946 12073 122502 12119
rect 115946 12070 115958 12073
rect 122490 12070 122502 12073
rect 122554 12070 122566 12122
rect 122714 12070 122726 12122
rect 122778 12119 122790 12122
rect 131114 12119 131126 12122
rect 122778 12073 131126 12119
rect 122778 12070 122790 12073
rect 131114 12070 131126 12073
rect 131178 12070 131190 12122
rect 136266 12070 136278 12122
rect 136330 12119 136342 12122
rect 136330 12073 139127 12119
rect 136330 12070 136342 12073
rect 117450 12007 117462 12010
rect 82570 11961 91527 12007
rect 91593 11961 117462 12007
rect 82570 11958 82582 11961
rect 81898 11849 82119 11895
rect 81898 11846 81910 11849
rect 82394 11846 82406 11898
rect 82458 11895 82470 11898
rect 91593 11895 91639 11961
rect 117450 11958 117462 11961
rect 117514 11958 117526 12010
rect 138842 12007 138854 12010
rect 117577 11961 138854 12007
rect 82458 11849 91639 11895
rect 82458 11846 82470 11849
rect 91690 11846 91702 11898
rect 91754 11895 91766 11898
rect 97738 11895 97750 11898
rect 91754 11849 97750 11895
rect 91754 11846 91766 11849
rect 97738 11846 97750 11849
rect 97802 11846 97814 11898
rect 98298 11846 98310 11898
rect 98362 11895 98374 11898
rect 99194 11895 99206 11898
rect 98362 11849 99206 11895
rect 98362 11846 98374 11849
rect 99194 11846 99206 11849
rect 99258 11846 99270 11898
rect 99321 11849 100935 11895
rect 73610 11737 79767 11783
rect 80057 11737 80439 11783
rect 73610 11734 73622 11737
rect 57034 11625 58822 11671
rect 58889 11625 68007 11671
rect 57034 11622 57046 11625
rect 51034 11510 51046 11562
rect 51098 11559 51110 11562
rect 58889 11559 58935 11625
rect 68170 11622 68182 11674
rect 68234 11671 68246 11674
rect 79594 11671 79606 11674
rect 68234 11625 79606 11671
rect 68234 11622 68246 11625
rect 79594 11622 79606 11625
rect 79658 11622 79670 11674
rect 79721 11671 79767 11737
rect 80490 11734 80502 11786
rect 80554 11783 80566 11786
rect 92922 11783 92934 11786
rect 80554 11737 92934 11783
rect 80554 11734 80566 11737
rect 92922 11734 92934 11737
rect 92986 11734 92998 11786
rect 93146 11734 93158 11786
rect 93210 11783 93222 11786
rect 99321 11783 99367 11849
rect 100426 11783 100438 11786
rect 93210 11737 99367 11783
rect 99433 11737 100438 11783
rect 93210 11734 93222 11737
rect 79721 11625 80327 11671
rect 51098 11513 58935 11559
rect 51098 11510 51110 11513
rect 64026 11510 64038 11562
rect 64090 11559 64102 11562
rect 80154 11559 80166 11562
rect 64090 11513 80166 11559
rect 64090 11510 64102 11513
rect 80154 11510 80166 11513
rect 80218 11510 80230 11562
rect 80281 11559 80327 11625
rect 80378 11622 80390 11674
rect 80442 11671 80454 11674
rect 81386 11671 81398 11674
rect 80442 11625 81398 11671
rect 80442 11622 80454 11625
rect 81386 11622 81398 11625
rect 81450 11622 81462 11674
rect 81722 11622 81734 11674
rect 81786 11671 81798 11674
rect 99433 11671 99479 11737
rect 100426 11734 100438 11737
rect 100490 11734 100502 11786
rect 100889 11783 100935 11849
rect 100986 11846 100998 11898
rect 101050 11895 101062 11898
rect 102554 11895 102566 11898
rect 101050 11849 102566 11895
rect 101050 11846 101062 11849
rect 102554 11846 102566 11849
rect 102618 11846 102630 11898
rect 103002 11846 103014 11898
rect 103066 11895 103078 11898
rect 103066 11849 103847 11895
rect 103066 11846 103078 11849
rect 102218 11783 102230 11786
rect 100889 11737 102230 11783
rect 102218 11734 102230 11737
rect 102282 11734 102294 11786
rect 102442 11734 102454 11786
rect 102506 11783 102518 11786
rect 103674 11783 103686 11786
rect 102506 11737 103686 11783
rect 102506 11734 102518 11737
rect 103674 11734 103686 11737
rect 103738 11734 103750 11786
rect 103801 11783 103847 11849
rect 104010 11846 104022 11898
rect 104074 11895 104086 11898
rect 108714 11895 108726 11898
rect 104074 11849 108726 11895
rect 104074 11846 104086 11849
rect 108714 11846 108726 11849
rect 108778 11846 108790 11898
rect 108938 11846 108950 11898
rect 109002 11895 109014 11898
rect 110954 11895 110966 11898
rect 109002 11849 110966 11895
rect 109002 11846 109014 11849
rect 110954 11846 110966 11849
rect 111018 11846 111030 11898
rect 111178 11846 111190 11898
rect 111242 11895 111254 11898
rect 117577 11895 117623 11961
rect 138842 11958 138854 11961
rect 138906 11958 138918 12010
rect 139081 12007 139127 12073
rect 139178 12070 139190 12122
rect 139242 12119 139254 12122
rect 144218 12119 144230 12122
rect 139242 12073 144230 12119
rect 139242 12070 139254 12073
rect 144218 12070 144230 12073
rect 144282 12070 144294 12122
rect 159562 12070 159574 12122
rect 159626 12119 159638 12122
rect 159626 12073 168022 12119
rect 159626 12070 159638 12073
rect 139738 12007 139750 12010
rect 139081 11961 139750 12007
rect 139738 11958 139750 11961
rect 139802 11958 139814 12010
rect 141082 11958 141094 12010
rect 141146 12007 141158 12010
rect 162362 12007 162374 12010
rect 141146 11961 162374 12007
rect 141146 11958 141158 11961
rect 162362 11958 162374 11961
rect 162426 11958 162438 12010
rect 167976 12007 168022 12073
rect 170986 12070 170998 12122
rect 171050 12119 171062 12122
rect 192042 12119 192054 12122
rect 171050 12073 192054 12119
rect 171050 12070 171062 12073
rect 192042 12070 192054 12073
rect 192106 12070 192118 12122
rect 213658 12007 213670 12010
rect 167976 11961 213670 12007
rect 213658 11958 213670 11961
rect 213722 11958 213734 12010
rect 111242 11849 117623 11895
rect 111242 11846 111254 11849
rect 118234 11846 118246 11898
rect 118298 11846 118310 11898
rect 118458 11846 118470 11898
rect 118522 11895 118534 11898
rect 118522 11849 126023 11895
rect 118522 11846 118534 11849
rect 104570 11783 104582 11786
rect 103801 11737 104582 11783
rect 104570 11734 104582 11737
rect 104634 11734 104646 11786
rect 105802 11734 105814 11786
rect 105866 11783 105878 11786
rect 114986 11783 114998 11786
rect 105866 11737 114998 11783
rect 105866 11734 105878 11737
rect 114986 11734 114998 11737
rect 115050 11734 115062 11786
rect 115210 11734 115222 11786
rect 115274 11783 115286 11786
rect 118249 11783 118295 11846
rect 115274 11737 118295 11783
rect 115274 11734 115286 11737
rect 119242 11734 119254 11786
rect 119306 11783 119318 11786
rect 120362 11783 120374 11786
rect 119306 11737 120374 11783
rect 119306 11734 119318 11737
rect 120362 11734 120374 11737
rect 120426 11734 120438 11786
rect 120586 11734 120598 11786
rect 120650 11783 120662 11786
rect 125850 11783 125862 11786
rect 120650 11737 125862 11783
rect 120650 11734 120662 11737
rect 125850 11734 125862 11737
rect 125914 11734 125926 11786
rect 125977 11783 126023 11849
rect 126074 11846 126086 11898
rect 126138 11895 126150 11898
rect 148138 11895 148150 11898
rect 126138 11849 148150 11895
rect 126138 11846 126150 11849
rect 148138 11846 148150 11849
rect 148202 11846 148214 11898
rect 148922 11846 148934 11898
rect 148986 11895 148998 11898
rect 151498 11895 151510 11898
rect 148986 11849 151510 11895
rect 148986 11846 148998 11849
rect 151498 11846 151510 11849
rect 151562 11846 151574 11898
rect 154858 11846 154870 11898
rect 154922 11895 154934 11898
rect 170650 11895 170662 11898
rect 154922 11849 170662 11895
rect 154922 11846 154934 11849
rect 170650 11846 170662 11849
rect 170714 11895 170726 11898
rect 192378 11895 192390 11898
rect 170714 11849 192390 11895
rect 170714 11846 170726 11849
rect 192378 11846 192390 11849
rect 192442 11846 192454 11898
rect 141082 11783 141094 11786
rect 125977 11737 141094 11783
rect 141082 11734 141094 11737
rect 141146 11734 141158 11786
rect 164602 11734 164614 11786
rect 164666 11783 164678 11786
rect 191706 11783 191718 11786
rect 164666 11737 191718 11783
rect 164666 11734 164678 11737
rect 191706 11734 191718 11737
rect 191770 11734 191782 11786
rect 100986 11671 100998 11674
rect 81786 11625 99479 11671
rect 99545 11625 100998 11671
rect 81786 11622 81798 11625
rect 82058 11559 82070 11562
rect 80281 11513 82070 11559
rect 82058 11510 82070 11513
rect 82122 11510 82134 11562
rect 82745 11513 83575 11559
rect 50586 11398 50598 11450
rect 50650 11447 50662 11450
rect 66938 11447 66950 11450
rect 50650 11401 66950 11447
rect 50650 11398 50662 11401
rect 66938 11398 66950 11401
rect 67002 11398 67014 11450
rect 67610 11398 67622 11450
rect 67674 11447 67686 11450
rect 69066 11447 69078 11450
rect 67674 11401 69078 11447
rect 67674 11398 67686 11401
rect 69066 11398 69078 11401
rect 69130 11398 69142 11450
rect 69402 11398 69414 11450
rect 69466 11447 69478 11450
rect 71866 11447 71878 11450
rect 69466 11401 71878 11447
rect 69466 11398 69478 11401
rect 71866 11398 71878 11401
rect 71930 11398 71942 11450
rect 72090 11398 72102 11450
rect 72154 11447 72166 11450
rect 82745 11447 82791 11513
rect 72154 11401 82791 11447
rect 72154 11398 72166 11401
rect 82842 11398 82854 11450
rect 82906 11447 82918 11450
rect 83402 11447 83414 11450
rect 82906 11401 83414 11447
rect 82906 11398 82918 11401
rect 83402 11398 83414 11401
rect 83466 11398 83478 11450
rect 83529 11447 83575 11513
rect 83962 11510 83974 11562
rect 84026 11559 84038 11562
rect 90570 11559 90582 11562
rect 84026 11513 90582 11559
rect 84026 11510 84038 11513
rect 90570 11510 90582 11513
rect 90634 11510 90646 11562
rect 90794 11510 90806 11562
rect 90858 11559 90870 11562
rect 91914 11559 91926 11562
rect 90858 11513 91926 11559
rect 90858 11510 90870 11513
rect 91914 11510 91926 11513
rect 91978 11510 91990 11562
rect 92922 11510 92934 11562
rect 92986 11559 92998 11562
rect 94714 11559 94726 11562
rect 92986 11513 94726 11559
rect 92986 11510 92998 11513
rect 94714 11510 94726 11513
rect 94778 11510 94790 11562
rect 94938 11510 94950 11562
rect 95002 11559 95014 11562
rect 98074 11559 98086 11562
rect 95002 11513 98086 11559
rect 95002 11510 95014 11513
rect 98074 11510 98086 11513
rect 98138 11510 98150 11562
rect 99545 11559 99591 11625
rect 100986 11622 100998 11625
rect 101050 11622 101062 11674
rect 101546 11622 101558 11674
rect 101610 11671 101622 11674
rect 109274 11671 109286 11674
rect 101610 11625 109286 11671
rect 101610 11622 101622 11625
rect 109274 11622 109286 11625
rect 109338 11622 109350 11674
rect 109722 11622 109734 11674
rect 109786 11671 109798 11674
rect 127754 11671 127766 11674
rect 109786 11625 127766 11671
rect 109786 11622 109798 11625
rect 127754 11622 127766 11625
rect 127818 11622 127830 11674
rect 134026 11622 134038 11674
rect 134090 11671 134102 11674
rect 138282 11671 138294 11674
rect 134090 11625 138294 11671
rect 134090 11622 134102 11625
rect 138282 11622 138294 11625
rect 138346 11622 138358 11674
rect 138506 11622 138518 11674
rect 138570 11671 138582 11674
rect 151274 11671 151286 11674
rect 138570 11625 151286 11671
rect 138570 11622 138582 11625
rect 151274 11622 151286 11625
rect 151338 11622 151350 11674
rect 98201 11513 99591 11559
rect 98201 11447 98247 11513
rect 99642 11510 99654 11562
rect 99706 11559 99718 11562
rect 112074 11559 112086 11562
rect 99706 11513 112086 11559
rect 99706 11510 99718 11513
rect 112074 11510 112086 11513
rect 112138 11510 112150 11562
rect 119018 11559 119030 11562
rect 113769 11513 117623 11559
rect 83529 11401 98247 11447
rect 98298 11398 98310 11450
rect 98362 11447 98374 11450
rect 103338 11447 103350 11450
rect 98362 11401 103350 11447
rect 98362 11398 98374 11401
rect 103338 11398 103350 11401
rect 103402 11398 103414 11450
rect 103562 11398 103574 11450
rect 103626 11447 103638 11450
rect 108042 11447 108054 11450
rect 103626 11401 108054 11447
rect 103626 11398 103638 11401
rect 108042 11398 108054 11401
rect 108106 11398 108118 11450
rect 113642 11447 113654 11450
rect 108169 11401 113654 11447
rect 49018 11286 49030 11338
rect 49082 11335 49094 11338
rect 61786 11335 61798 11338
rect 49082 11289 61798 11335
rect 49082 11286 49094 11289
rect 61786 11286 61798 11289
rect 61850 11286 61862 11338
rect 62346 11286 62358 11338
rect 62410 11335 62422 11338
rect 108169 11335 108215 11401
rect 113642 11398 113654 11401
rect 113706 11398 113718 11450
rect 62410 11289 108215 11335
rect 62410 11286 62422 11289
rect 109274 11286 109286 11338
rect 109338 11335 109350 11338
rect 113769 11335 113815 11513
rect 113866 11398 113878 11450
rect 113930 11447 113942 11450
rect 117226 11447 117238 11450
rect 113930 11401 117238 11447
rect 113930 11398 113942 11401
rect 117226 11398 117238 11401
rect 117290 11398 117302 11450
rect 117450 11398 117462 11450
rect 117514 11398 117526 11450
rect 109338 11289 113815 11335
rect 109338 11286 109350 11289
rect 114090 11286 114102 11338
rect 114154 11335 114166 11338
rect 116442 11335 116454 11338
rect 114154 11289 116454 11335
rect 114154 11286 114166 11289
rect 116442 11286 116454 11289
rect 116506 11286 116518 11338
rect 16314 11174 16326 11226
rect 16378 11223 16390 11226
rect 79146 11223 79158 11226
rect 16378 11177 79158 11223
rect 16378 11174 16390 11177
rect 79146 11174 79158 11177
rect 79210 11174 79222 11226
rect 79482 11174 79494 11226
rect 79546 11223 79558 11226
rect 80602 11223 80614 11226
rect 79546 11177 80614 11223
rect 79546 11174 79558 11177
rect 80602 11174 80614 11177
rect 80666 11174 80678 11226
rect 80826 11174 80838 11226
rect 80890 11223 80902 11226
rect 82506 11223 82518 11226
rect 80890 11177 82518 11223
rect 80890 11174 80902 11177
rect 82506 11174 82518 11177
rect 82570 11174 82582 11226
rect 82730 11174 82742 11226
rect 82794 11223 82806 11226
rect 86426 11223 86438 11226
rect 82794 11177 86438 11223
rect 82794 11174 82806 11177
rect 86426 11174 86438 11177
rect 86490 11174 86502 11226
rect 86650 11174 86662 11226
rect 86714 11223 86726 11226
rect 88778 11223 88790 11226
rect 86714 11177 88790 11223
rect 86714 11174 86726 11177
rect 88778 11174 88790 11177
rect 88842 11174 88854 11226
rect 89002 11174 89014 11226
rect 89066 11223 89078 11226
rect 117465 11223 117511 11398
rect 89066 11177 117511 11223
rect 117577 11223 117623 11513
rect 117689 11513 119030 11559
rect 117689 11338 117735 11513
rect 119018 11510 119030 11513
rect 119082 11510 119094 11562
rect 119578 11510 119590 11562
rect 119642 11559 119654 11562
rect 126298 11559 126310 11562
rect 119642 11513 126310 11559
rect 119642 11510 119654 11513
rect 126298 11510 126310 11513
rect 126362 11510 126374 11562
rect 126522 11510 126534 11562
rect 126586 11559 126598 11562
rect 126586 11513 135655 11559
rect 126586 11510 126598 11513
rect 117786 11398 117798 11450
rect 117850 11447 117862 11450
rect 124394 11447 124406 11450
rect 117850 11401 124406 11447
rect 117850 11398 117862 11401
rect 124394 11398 124406 11401
rect 124458 11398 124470 11450
rect 129210 11398 129222 11450
rect 129274 11447 129286 11450
rect 135370 11447 135382 11450
rect 129274 11401 135382 11447
rect 129274 11398 129286 11401
rect 135370 11398 135382 11401
rect 135434 11398 135446 11450
rect 135609 11447 135655 11513
rect 135706 11510 135718 11562
rect 135770 11559 135782 11562
rect 147466 11559 147478 11562
rect 135770 11513 147478 11559
rect 135770 11510 135782 11513
rect 147466 11510 147478 11513
rect 147530 11510 147542 11562
rect 138618 11447 138630 11450
rect 135609 11401 138630 11447
rect 138618 11398 138630 11401
rect 138682 11398 138694 11450
rect 150042 11398 150054 11450
rect 150106 11447 150118 11450
rect 153514 11447 153526 11450
rect 150106 11401 153526 11447
rect 150106 11398 150118 11401
rect 153514 11398 153526 11401
rect 153578 11398 153590 11450
rect 117674 11286 117686 11338
rect 117738 11286 117750 11338
rect 117898 11286 117910 11338
rect 117962 11335 117974 11338
rect 121034 11335 121046 11338
rect 117962 11289 121046 11335
rect 117962 11286 117974 11289
rect 121034 11286 121046 11289
rect 121098 11286 121110 11338
rect 121818 11286 121830 11338
rect 121882 11335 121894 11338
rect 136602 11335 136614 11338
rect 121882 11289 136614 11335
rect 121882 11286 121894 11289
rect 136602 11286 136614 11289
rect 136666 11286 136678 11338
rect 151162 11335 151174 11338
rect 137065 11289 151174 11335
rect 118346 11223 118358 11226
rect 117577 11177 118358 11223
rect 89066 11174 89078 11177
rect 118346 11174 118358 11177
rect 118410 11174 118422 11226
rect 118570 11174 118582 11226
rect 118634 11223 118646 11226
rect 124954 11223 124966 11226
rect 118634 11177 124966 11223
rect 118634 11174 118646 11177
rect 124954 11174 124966 11177
rect 125018 11174 125030 11226
rect 127754 11174 127766 11226
rect 127818 11223 127830 11226
rect 137065 11223 137111 11289
rect 151162 11286 151174 11289
rect 151226 11286 151238 11338
rect 127818 11177 137111 11223
rect 127818 11174 127830 11177
rect 138058 11174 138070 11226
rect 138122 11223 138134 11226
rect 138954 11223 138966 11226
rect 138122 11177 138966 11223
rect 138122 11174 138134 11177
rect 138954 11174 138966 11177
rect 139018 11174 139030 11226
rect 139514 11174 139526 11226
rect 139578 11223 139590 11226
rect 139578 11177 141031 11223
rect 139578 11174 139590 11177
rect 53386 11062 53398 11114
rect 53450 11111 53462 11114
rect 129994 11111 130006 11114
rect 53450 11065 130006 11111
rect 53450 11062 53462 11065
rect 129994 11062 130006 11065
rect 130058 11062 130070 11114
rect 130442 11062 130454 11114
rect 130506 11111 130518 11114
rect 132906 11111 132918 11114
rect 130506 11065 132918 11111
rect 130506 11062 130518 11065
rect 132906 11062 132918 11065
rect 132970 11062 132982 11114
rect 133578 11062 133590 11114
rect 133642 11111 133654 11114
rect 135146 11111 135158 11114
rect 133642 11065 135158 11111
rect 133642 11062 133654 11065
rect 135146 11062 135158 11065
rect 135210 11062 135222 11114
rect 135370 11062 135382 11114
rect 135434 11111 135446 11114
rect 140858 11111 140870 11114
rect 135434 11065 140870 11111
rect 135434 11062 135446 11065
rect 140858 11062 140870 11065
rect 140922 11062 140934 11114
rect 140985 11111 141031 11177
rect 143322 11174 143334 11226
rect 143386 11223 143398 11226
rect 146010 11223 146022 11226
rect 143386 11177 146022 11223
rect 143386 11174 143398 11177
rect 146010 11174 146022 11177
rect 146074 11174 146086 11226
rect 150378 11111 150390 11114
rect 140985 11065 150390 11111
rect 150378 11062 150390 11065
rect 150442 11062 150454 11114
rect 166618 11062 166630 11114
rect 166682 11111 166694 11114
rect 206378 11111 206390 11114
rect 166682 11065 206390 11111
rect 166682 11062 166694 11065
rect 206378 11062 206390 11065
rect 206442 11062 206454 11114
rect 6458 10950 6470 11002
rect 6522 10999 6534 11002
rect 83626 10999 83638 11002
rect 6522 10953 83638 10999
rect 6522 10950 6534 10953
rect 83626 10950 83638 10953
rect 83690 10950 83702 11002
rect 84298 10950 84310 11002
rect 84362 10999 84374 11002
rect 85082 10999 85094 11002
rect 84362 10953 85094 10999
rect 84362 10950 84374 10953
rect 85082 10950 85094 10953
rect 85146 10950 85158 11002
rect 85306 10950 85318 11002
rect 85370 10999 85382 11002
rect 89562 10999 89574 11002
rect 85370 10953 89574 10999
rect 85370 10950 85382 10953
rect 89562 10950 89574 10953
rect 89626 10950 89638 11002
rect 90010 10950 90022 11002
rect 90074 10999 90086 11002
rect 98746 10999 98758 11002
rect 90074 10953 98758 10999
rect 90074 10950 90086 10953
rect 98746 10950 98758 10953
rect 98810 10950 98822 11002
rect 98970 10950 98982 11002
rect 99034 10999 99046 11002
rect 103002 10999 103014 11002
rect 99034 10953 103014 10999
rect 99034 10950 99046 10953
rect 103002 10950 103014 10953
rect 103066 10950 103078 11002
rect 103338 10950 103350 11002
rect 103402 10999 103414 11002
rect 135706 10999 135718 11002
rect 103402 10953 135718 10999
rect 103402 10950 103414 10953
rect 135706 10950 135718 10953
rect 135770 10950 135782 11002
rect 135930 10950 135942 11002
rect 135994 10999 136006 11002
rect 150266 10999 150278 11002
rect 135994 10953 150278 10999
rect 135994 10950 136006 10953
rect 150266 10950 150278 10953
rect 150330 10950 150342 11002
rect 151050 10950 151062 11002
rect 151114 10999 151126 11002
rect 190026 10999 190038 11002
rect 151114 10953 190038 10999
rect 151114 10950 151126 10953
rect 190026 10950 190038 10953
rect 190090 10950 190102 11002
rect 21802 10838 21814 10890
rect 21866 10887 21878 10890
rect 125514 10887 125526 10890
rect 21866 10841 125526 10887
rect 21866 10838 21878 10841
rect 125514 10838 125526 10841
rect 125578 10838 125590 10890
rect 125738 10838 125750 10890
rect 125802 10887 125814 10890
rect 138506 10887 138518 10890
rect 125802 10841 138518 10887
rect 125802 10838 125814 10841
rect 138506 10838 138518 10841
rect 138570 10838 138582 10890
rect 138954 10838 138966 10890
rect 139018 10887 139030 10890
rect 139018 10841 144502 10887
rect 139018 10838 139030 10841
rect 41290 10726 41302 10778
rect 41354 10775 41366 10778
rect 60778 10775 60790 10778
rect 41354 10729 60790 10775
rect 41354 10726 41366 10729
rect 60778 10726 60790 10729
rect 60842 10726 60854 10778
rect 61002 10726 61014 10778
rect 61066 10775 61078 10778
rect 65258 10775 65270 10778
rect 61066 10729 65270 10775
rect 61066 10726 61078 10729
rect 65258 10726 65270 10729
rect 65322 10726 65334 10778
rect 65482 10726 65494 10778
rect 65546 10775 65558 10778
rect 69290 10775 69302 10778
rect 65546 10729 69302 10775
rect 65546 10726 65558 10729
rect 69290 10726 69302 10729
rect 69354 10726 69366 10778
rect 71306 10726 71318 10778
rect 71370 10775 71382 10778
rect 73434 10775 73446 10778
rect 71370 10729 73446 10775
rect 71370 10726 71382 10729
rect 73434 10726 73446 10729
rect 73498 10726 73510 10778
rect 73770 10726 73782 10778
rect 73834 10775 73846 10778
rect 125626 10775 125638 10778
rect 73834 10729 125638 10775
rect 73834 10726 73846 10729
rect 125626 10726 125638 10729
rect 125690 10726 125702 10778
rect 125850 10726 125862 10778
rect 125914 10775 125926 10778
rect 134810 10775 134822 10778
rect 125914 10729 134822 10775
rect 125914 10726 125926 10729
rect 134810 10726 134822 10729
rect 134874 10726 134886 10778
rect 136378 10726 136390 10778
rect 136442 10775 136454 10778
rect 143546 10775 143558 10778
rect 136442 10729 143558 10775
rect 136442 10726 136454 10729
rect 143546 10726 143558 10729
rect 143610 10726 143622 10778
rect 144456 10775 144502 10841
rect 151386 10838 151398 10890
rect 151450 10887 151462 10890
rect 194506 10887 194518 10890
rect 151450 10841 194518 10887
rect 151450 10838 151462 10841
rect 194506 10838 194518 10841
rect 194570 10838 194582 10890
rect 187786 10775 187798 10778
rect 144456 10729 187798 10775
rect 187786 10726 187798 10729
rect 187850 10726 187862 10778
rect 54282 10614 54294 10666
rect 54346 10663 54358 10666
rect 109722 10663 109734 10666
rect 54346 10617 109734 10663
rect 54346 10614 54358 10617
rect 109722 10614 109734 10617
rect 109786 10614 109798 10666
rect 109946 10614 109958 10666
rect 110010 10663 110022 10666
rect 114202 10663 114214 10666
rect 110010 10617 114214 10663
rect 110010 10614 110022 10617
rect 114202 10614 114214 10617
rect 114266 10614 114278 10666
rect 114426 10614 114438 10666
rect 114490 10663 114502 10666
rect 117338 10663 117350 10666
rect 114490 10617 117350 10663
rect 114490 10614 114502 10617
rect 117338 10614 117350 10617
rect 117402 10614 117414 10666
rect 117674 10614 117686 10666
rect 117738 10663 117750 10666
rect 120474 10663 120486 10666
rect 117738 10617 120486 10663
rect 117738 10614 117750 10617
rect 120474 10614 120486 10617
rect 120538 10614 120550 10666
rect 121594 10614 121606 10666
rect 121658 10663 121670 10666
rect 129098 10663 129110 10666
rect 121658 10617 129110 10663
rect 121658 10614 121670 10617
rect 129098 10614 129110 10617
rect 129162 10614 129174 10666
rect 130890 10614 130902 10666
rect 130954 10663 130966 10666
rect 181066 10663 181078 10666
rect 130954 10617 134535 10663
rect 130954 10614 130966 10617
rect 50026 10502 50038 10554
rect 50090 10551 50102 10554
rect 133914 10551 133926 10554
rect 50090 10505 133926 10551
rect 50090 10502 50102 10505
rect 133914 10502 133926 10505
rect 133978 10502 133990 10554
rect 21578 10390 21590 10442
rect 21642 10439 21654 10442
rect 83738 10439 83750 10442
rect 21642 10393 83750 10439
rect 21642 10390 21654 10393
rect 83738 10390 83750 10393
rect 83802 10390 83814 10442
rect 83962 10390 83974 10442
rect 84026 10439 84038 10442
rect 89338 10439 89350 10442
rect 84026 10393 89350 10439
rect 84026 10390 84038 10393
rect 89338 10390 89350 10393
rect 89402 10390 89414 10442
rect 89562 10390 89574 10442
rect 89626 10439 89638 10442
rect 134250 10439 134262 10442
rect 89626 10393 134262 10439
rect 89626 10390 89638 10393
rect 134250 10390 134262 10393
rect 134314 10390 134326 10442
rect 134489 10439 134535 10617
rect 134825 10617 181078 10663
rect 134825 10439 134871 10617
rect 181066 10614 181078 10617
rect 181130 10614 181142 10666
rect 186554 10614 186566 10666
rect 186618 10663 186630 10666
rect 200890 10663 200902 10666
rect 186618 10617 200902 10663
rect 186618 10614 186630 10617
rect 200890 10614 200902 10617
rect 200954 10614 200966 10666
rect 137722 10502 137734 10554
rect 137786 10551 137798 10554
rect 194954 10551 194966 10554
rect 137786 10505 194966 10551
rect 137786 10502 137798 10505
rect 194954 10502 194966 10505
rect 195018 10502 195030 10554
rect 134489 10393 134871 10439
rect 136826 10390 136838 10442
rect 136890 10439 136902 10442
rect 143322 10439 143334 10442
rect 136890 10393 143334 10439
rect 136890 10390 136902 10393
rect 143322 10390 143334 10393
rect 143386 10390 143398 10442
rect 143546 10390 143558 10442
rect 143610 10439 143622 10442
rect 211418 10439 211430 10442
rect 143610 10393 211430 10439
rect 143610 10390 143622 10393
rect 211418 10390 211430 10393
rect 211482 10390 211494 10442
rect 1344 10218 218624 10252
rect 1344 10166 28378 10218
rect 28430 10166 28482 10218
rect 28534 10166 28586 10218
rect 28638 10166 82706 10218
rect 82758 10166 82810 10218
rect 82862 10166 82914 10218
rect 82966 10166 137034 10218
rect 137086 10166 137138 10218
rect 137190 10166 137242 10218
rect 137294 10166 191362 10218
rect 191414 10166 191466 10218
rect 191518 10166 191570 10218
rect 191622 10166 218624 10218
rect 1344 10132 218624 10166
rect 78362 10047 78374 10050
rect 9830 9994 9882 10006
rect 9830 9930 9882 9942
rect 10726 9994 10778 10006
rect 10726 9930 10778 9942
rect 11622 9994 11674 10006
rect 11622 9930 11674 9942
rect 45558 9994 45610 10006
rect 76582 9994 76634 10006
rect 54506 9942 54518 9994
rect 54570 9942 54582 9994
rect 45558 9930 45610 9942
rect 76582 9930 76634 9942
rect 77590 9994 77642 10006
rect 77590 9930 77642 9942
rect 78321 9998 78374 10047
rect 78426 9998 78438 10050
rect 42590 9882 42642 9894
rect 42590 9818 42642 9830
rect 43486 9882 43538 9894
rect 43486 9818 43538 9830
rect 47966 9882 48018 9894
rect 47966 9818 48018 9830
rect 48862 9882 48914 9894
rect 48862 9818 48914 9830
rect 50542 9882 50594 9894
rect 50542 9818 50594 9830
rect 52782 9882 52834 9894
rect 52782 9818 52834 9830
rect 70926 9882 70978 9894
rect 8318 9770 8370 9782
rect 53566 9770 53618 9782
rect 55178 9774 55190 9826
rect 55242 9774 55254 9826
rect 55402 9774 55414 9826
rect 55466 9774 55478 9826
rect 70926 9818 70978 9830
rect 11050 9718 11062 9770
rect 11114 9718 11126 9770
rect 8318 9706 8370 9718
rect 53566 9706 53618 9718
rect 56590 9770 56642 9782
rect 56590 9706 56642 9718
rect 8878 9658 8930 9670
rect 8878 9594 8930 9606
rect 10166 9658 10218 9670
rect 10166 9594 10218 9606
rect 11958 9658 12010 9670
rect 11958 9594 12010 9606
rect 12574 9658 12626 9670
rect 12574 9594 12626 9606
rect 22542 9658 22594 9670
rect 22542 9594 22594 9606
rect 25230 9658 25282 9670
rect 25230 9594 25282 9606
rect 43934 9658 43986 9670
rect 43934 9594 43986 9606
rect 45222 9658 45274 9670
rect 45222 9594 45274 9606
rect 46062 9658 46114 9670
rect 46062 9594 46114 9606
rect 46510 9658 46562 9670
rect 46510 9594 46562 9606
rect 47070 9658 47122 9670
rect 47070 9594 47122 9606
rect 57038 9658 57090 9670
rect 57038 9594 57090 9606
rect 57374 9658 57426 9670
rect 57374 9594 57426 9606
rect 58046 9658 58098 9670
rect 58046 9594 58098 9606
rect 76246 9658 76298 9670
rect 76246 9594 76298 9606
rect 77254 9658 77306 9670
rect 78321 9658 78367 9998
rect 79270 9994 79322 10006
rect 79270 9930 79322 9942
rect 80950 9994 81002 10006
rect 80950 9930 81002 9942
rect 81846 9994 81898 10006
rect 81846 9930 81898 9942
rect 86774 9994 86826 10006
rect 86774 9930 86826 9942
rect 104022 9994 104074 10006
rect 104022 9930 104074 9942
rect 109958 9994 110010 10006
rect 109958 9930 110010 9942
rect 111862 9994 111914 10006
rect 111862 9930 111914 9942
rect 115782 9994 115834 10006
rect 115782 9930 115834 9942
rect 121382 9994 121434 10006
rect 121382 9930 121434 9942
rect 129222 9994 129274 10006
rect 129222 9930 129274 9942
rect 131574 9994 131626 10006
rect 137398 9994 137450 10006
rect 132570 9942 132582 9994
rect 132634 9942 132646 9994
rect 135482 9942 135494 9994
rect 135546 9942 135558 9994
rect 131574 9930 131626 9942
rect 137398 9930 137450 9942
rect 139302 9994 139354 10006
rect 139302 9930 139354 9942
rect 143222 9994 143274 10006
rect 143222 9930 143274 9942
rect 144118 9994 144170 10006
rect 144118 9930 144170 9942
rect 147142 9994 147194 10006
rect 147142 9930 147194 9942
rect 151062 9994 151114 10006
rect 151062 9930 151114 9942
rect 154982 9994 155034 10006
rect 154982 9930 155034 9942
rect 165622 9994 165674 10006
rect 165622 9930 165674 9942
rect 172454 9994 172506 10006
rect 172454 9930 172506 9942
rect 176934 9994 176986 10006
rect 176934 9930 176986 9942
rect 180070 9994 180122 10006
rect 183990 9994 184042 10006
rect 182522 9942 182534 9994
rect 182586 9942 182598 9994
rect 180070 9930 180122 9942
rect 183990 9930 184042 9942
rect 187910 9994 187962 10006
rect 187910 9930 187962 9942
rect 191830 9994 191882 10006
rect 109062 9882 109114 9894
rect 109062 9818 109114 9830
rect 114718 9882 114770 9894
rect 114718 9818 114770 9830
rect 137790 9882 137842 9894
rect 80110 9770 80162 9782
rect 83134 9770 83186 9782
rect 78922 9718 78934 9770
rect 78986 9718 78998 9770
rect 80602 9718 80614 9770
rect 80666 9718 80678 9770
rect 82394 9718 82406 9770
rect 82458 9718 82470 9770
rect 80110 9706 80162 9718
rect 83134 9706 83186 9718
rect 102958 9770 103010 9782
rect 120542 9770 120594 9782
rect 132010 9774 132022 9826
rect 132074 9774 132086 9826
rect 133466 9774 133478 9826
rect 133530 9774 133542 9826
rect 134922 9774 134934 9826
rect 134986 9774 134998 9826
rect 137790 9818 137842 9830
rect 141710 9882 141762 9894
rect 139738 9774 139750 9826
rect 139802 9774 139814 9826
rect 141710 9818 141762 9830
rect 144510 9882 144562 9894
rect 144510 9818 144562 9830
rect 147534 9882 147586 9894
rect 147534 9818 147586 9830
rect 147982 9882 148034 9894
rect 147982 9818 148034 9830
rect 148430 9882 148482 9894
rect 148430 9818 148482 9830
rect 149774 9882 149826 9894
rect 149774 9818 149826 9830
rect 151454 9882 151506 9894
rect 151454 9818 151506 9830
rect 153022 9882 153074 9894
rect 153022 9818 153074 9830
rect 155374 9882 155426 9894
rect 155374 9818 155426 9830
rect 161422 9882 161474 9894
rect 144958 9770 145010 9782
rect 156314 9774 156326 9826
rect 156378 9774 156390 9826
rect 157770 9774 157782 9826
rect 157834 9774 157846 9826
rect 159338 9774 159350 9826
rect 159402 9774 159414 9826
rect 160794 9774 160806 9826
rect 160858 9774 160870 9826
rect 161422 9818 161474 9830
rect 164334 9882 164386 9894
rect 162362 9774 162374 9826
rect 162426 9774 162438 9826
rect 164334 9818 164386 9830
rect 168702 9882 168754 9894
rect 166618 9774 166630 9826
rect 166682 9774 166694 9826
rect 168702 9818 168754 9830
rect 173294 9882 173346 9894
rect 188750 9882 188802 9894
rect 191370 9886 191382 9938
rect 191434 9886 191446 9938
rect 191830 9930 191882 9942
rect 193734 9994 193786 10006
rect 193734 9930 193786 9942
rect 195078 9994 195130 10006
rect 195078 9930 195130 9942
rect 195974 9994 196026 10006
rect 195974 9930 196026 9942
rect 196422 9994 196474 10006
rect 196422 9930 196474 9942
rect 198102 9994 198154 10006
rect 198102 9930 198154 9942
rect 199446 9994 199498 10006
rect 199446 9930 199498 9942
rect 202022 9994 202074 10006
rect 202022 9930 202074 9942
rect 204822 9994 204874 10006
rect 204822 9930 204874 9942
rect 206166 9994 206218 10006
rect 206166 9930 206218 9942
rect 211878 9994 211930 10006
rect 171210 9774 171222 9826
rect 171274 9774 171286 9826
rect 173294 9818 173346 9830
rect 181134 9826 181186 9838
rect 185054 9826 185106 9838
rect 174190 9770 174242 9782
rect 174794 9774 174806 9826
rect 174858 9774 174870 9826
rect 179610 9774 179622 9826
rect 179674 9774 179686 9826
rect 182746 9774 182758 9826
rect 182810 9774 182822 9826
rect 185882 9774 185894 9826
rect 185946 9774 185958 9826
rect 188750 9818 188802 9830
rect 198494 9882 198546 9894
rect 189802 9774 189814 9826
rect 189866 9774 189878 9826
rect 198494 9818 198546 9830
rect 200398 9882 200450 9894
rect 200398 9818 200450 9830
rect 200734 9882 200786 9894
rect 200734 9818 200786 9830
rect 202414 9882 202466 9894
rect 202414 9818 202466 9830
rect 203310 9882 203362 9894
rect 208170 9886 208182 9938
rect 208234 9886 208246 9938
rect 211878 9930 211930 9942
rect 213782 9994 213834 10006
rect 213782 9930 213834 9942
rect 203310 9818 203362 9830
rect 208058 9774 208070 9826
rect 208122 9774 208134 9826
rect 210970 9774 210982 9826
rect 211034 9774 211046 9826
rect 103674 9718 103686 9770
rect 103738 9718 103750 9770
rect 108714 9718 108726 9770
rect 108778 9718 108790 9770
rect 111514 9718 111526 9770
rect 111578 9718 111590 9770
rect 115434 9718 115446 9770
rect 115498 9718 115510 9770
rect 121034 9718 121046 9770
rect 121098 9718 121110 9770
rect 129994 9718 130006 9770
rect 130058 9718 130070 9770
rect 131226 9718 131238 9770
rect 131290 9718 131302 9770
rect 137050 9718 137062 9770
rect 137114 9718 137126 9770
rect 142874 9718 142886 9770
rect 142938 9718 142950 9770
rect 146794 9718 146806 9770
rect 146858 9718 146870 9770
rect 150714 9718 150726 9770
rect 150778 9718 150790 9770
rect 154634 9718 154646 9770
rect 154698 9718 154710 9770
rect 165274 9718 165286 9770
rect 165338 9718 165350 9770
rect 172778 9718 172790 9770
rect 172842 9718 172854 9770
rect 177258 9718 177270 9770
rect 177322 9718 177334 9770
rect 180394 9718 180406 9770
rect 180458 9718 180470 9770
rect 181134 9762 181186 9774
rect 185054 9762 185106 9774
rect 217310 9770 217362 9782
rect 192154 9718 192166 9770
rect 192218 9718 192230 9770
rect 194730 9718 194742 9770
rect 194794 9718 194806 9770
rect 204474 9718 204486 9770
rect 204538 9718 204550 9770
rect 102958 9706 103010 9718
rect 120542 9706 120594 9718
rect 78250 9606 78262 9658
rect 78314 9609 78367 9658
rect 78430 9658 78482 9670
rect 78314 9606 78326 9609
rect 77254 9594 77306 9606
rect 78430 9594 78482 9606
rect 81510 9658 81562 9670
rect 81510 9594 81562 9606
rect 82742 9658 82794 9670
rect 82742 9594 82794 9606
rect 83918 9658 83970 9670
rect 83918 9594 83970 9606
rect 85934 9658 85986 9670
rect 85934 9594 85986 9606
rect 86438 9658 86490 9670
rect 86438 9594 86490 9606
rect 96014 9658 96066 9670
rect 96014 9594 96066 9606
rect 98926 9658 98978 9670
rect 98926 9594 98978 9606
rect 99710 9658 99762 9670
rect 99710 9594 99762 9606
rect 100046 9658 100098 9670
rect 100046 9594 100098 9606
rect 106878 9658 106930 9670
rect 106878 9594 106930 9606
rect 107830 9658 107882 9670
rect 107830 9594 107882 9606
rect 108166 9658 108218 9670
rect 108166 9594 108218 9606
rect 109622 9658 109674 9670
rect 109622 9594 109674 9606
rect 110798 9658 110850 9670
rect 110798 9594 110850 9606
rect 128382 9658 128434 9670
rect 128382 9594 128434 9606
rect 128886 9658 128938 9670
rect 128886 9594 128938 9606
rect 130342 9658 130394 9670
rect 130342 9594 130394 9606
rect 134094 9658 134146 9670
rect 135930 9662 135942 9714
rect 135994 9662 136006 9714
rect 134094 9594 134146 9606
rect 138966 9658 139018 9670
rect 140746 9662 140758 9714
rect 140810 9662 140822 9714
rect 144958 9706 145010 9718
rect 138966 9594 139018 9606
rect 143782 9658 143834 9670
rect 140970 9550 140982 9602
rect 141034 9550 141046 9602
rect 143782 9594 143834 9606
rect 145518 9658 145570 9670
rect 145518 9594 145570 9606
rect 145966 9658 146018 9670
rect 145966 9594 146018 9606
rect 148878 9658 148930 9670
rect 148878 9594 148930 9606
rect 149438 9658 149490 9670
rect 149438 9594 149490 9606
rect 152238 9658 152290 9670
rect 152238 9594 152290 9606
rect 152686 9658 152738 9670
rect 152686 9594 152738 9606
rect 153582 9658 153634 9670
rect 153582 9594 153634 9606
rect 158566 9658 158618 9670
rect 156314 9550 156326 9602
rect 156378 9550 156390 9602
rect 158566 9594 158618 9606
rect 158902 9658 158954 9670
rect 163706 9662 163718 9714
rect 163770 9662 163782 9714
rect 166730 9662 166742 9714
rect 166794 9662 166806 9714
rect 158902 9594 158954 9606
rect 169150 9658 169202 9670
rect 171658 9662 171670 9714
rect 171722 9662 171734 9714
rect 174190 9706 174242 9718
rect 175130 9662 175142 9714
rect 175194 9662 175206 9714
rect 178266 9662 178278 9714
rect 178330 9662 178342 9714
rect 160570 9550 160582 9602
rect 160634 9550 160646 9602
rect 163594 9550 163606 9602
rect 163658 9550 163670 9602
rect 169150 9594 169202 9606
rect 181022 9658 181074 9670
rect 182074 9662 182086 9714
rect 182138 9662 182150 9714
rect 170314 9550 170326 9602
rect 170378 9550 170390 9602
rect 178154 9550 178166 9602
rect 178218 9550 178230 9602
rect 181022 9594 181074 9606
rect 184326 9658 184378 9670
rect 184326 9594 184378 9606
rect 184942 9658 184994 9670
rect 185994 9662 186006 9714
rect 186058 9662 186070 9714
rect 184942 9594 184994 9606
rect 188246 9658 188298 9670
rect 189914 9662 189926 9714
rect 189978 9662 189990 9714
rect 187338 9550 187350 9602
rect 187402 9550 187414 9602
rect 188246 9594 188298 9606
rect 192782 9658 192834 9670
rect 192782 9594 192834 9606
rect 194070 9658 194122 9670
rect 194070 9594 194122 9606
rect 195638 9658 195690 9670
rect 195638 9594 195690 9606
rect 196758 9658 196810 9670
rect 196758 9594 196810 9606
rect 197766 9658 197818 9670
rect 197766 9594 197818 9606
rect 199110 9658 199162 9670
rect 199110 9594 199162 9606
rect 199950 9658 200002 9670
rect 199950 9594 200002 9606
rect 201686 9658 201738 9670
rect 201686 9594 201738 9606
rect 202862 9658 202914 9670
rect 202862 9594 202914 9606
rect 203870 9658 203922 9670
rect 203870 9594 203922 9606
rect 205830 9658 205882 9670
rect 210746 9662 210758 9714
rect 210810 9662 210822 9714
rect 217310 9706 217362 9718
rect 205830 9594 205882 9606
rect 211542 9658 211594 9670
rect 209514 9550 209526 9602
rect 209578 9550 209590 9602
rect 211542 9594 211594 9606
rect 212270 9658 212322 9670
rect 212270 9594 212322 9606
rect 213446 9658 213498 9670
rect 213446 9594 213498 9606
rect 214174 9658 214226 9670
rect 214174 9594 214226 9606
rect 214622 9658 214674 9670
rect 214622 9594 214674 9606
rect 215070 9658 215122 9670
rect 215070 9594 215122 9606
rect 215518 9658 215570 9670
rect 215518 9594 215570 9606
rect 215966 9658 216018 9670
rect 215966 9594 216018 9606
rect 216414 9658 216466 9670
rect 216414 9594 216466 9606
rect 1344 9434 218624 9468
rect 1344 9382 55542 9434
rect 55594 9382 55646 9434
rect 55698 9382 55750 9434
rect 55802 9382 109870 9434
rect 109922 9382 109974 9434
rect 110026 9382 110078 9434
rect 110130 9382 164198 9434
rect 164250 9382 164302 9434
rect 164354 9382 164406 9434
rect 164458 9382 218624 9434
rect 1344 9348 218624 9382
rect 9718 9210 9770 9222
rect 9718 9146 9770 9158
rect 10614 9210 10666 9222
rect 10614 9146 10666 9158
rect 15598 9210 15650 9222
rect 15598 9146 15650 9158
rect 17782 9210 17834 9222
rect 17782 9146 17834 9158
rect 18118 9210 18170 9222
rect 18118 9146 18170 9158
rect 18510 9210 18562 9222
rect 18510 9146 18562 9158
rect 19910 9210 19962 9222
rect 19910 9146 19962 9158
rect 20246 9210 20298 9222
rect 20246 9146 20298 9158
rect 20638 9210 20690 9222
rect 20638 9146 20690 9158
rect 22262 9210 22314 9222
rect 22262 9146 22314 9158
rect 25958 9210 26010 9222
rect 25958 9146 26010 9158
rect 41974 9210 42026 9222
rect 41974 9146 42026 9158
rect 42310 9210 42362 9222
rect 42310 9146 42362 9158
rect 43206 9210 43258 9222
rect 43206 9146 43258 9158
rect 44046 9210 44098 9222
rect 44046 9146 44098 9158
rect 44550 9210 44602 9222
rect 44550 9146 44602 9158
rect 44886 9210 44938 9222
rect 44886 9146 44938 9158
rect 45390 9210 45442 9222
rect 45390 9146 45442 9158
rect 47350 9210 47402 9222
rect 47350 9146 47402 9158
rect 47686 9210 47738 9222
rect 47686 9146 47738 9158
rect 48582 9210 48634 9222
rect 48582 9146 48634 9158
rect 49926 9210 49978 9222
rect 49926 9146 49978 9158
rect 50262 9210 50314 9222
rect 50262 9146 50314 9158
rect 50822 9210 50874 9222
rect 50822 9146 50874 9158
rect 51158 9210 51210 9222
rect 51158 9146 51210 9158
rect 51550 9210 51602 9222
rect 51550 9146 51602 9158
rect 52166 9210 52218 9222
rect 52166 9146 52218 9158
rect 52502 9210 52554 9222
rect 52502 9146 52554 9158
rect 57766 9210 57818 9222
rect 57766 9146 57818 9158
rect 61238 9210 61290 9222
rect 61238 9146 61290 9158
rect 61574 9210 61626 9222
rect 61574 9146 61626 9158
rect 61966 9210 62018 9222
rect 61966 9146 62018 9158
rect 70198 9210 70250 9222
rect 70198 9146 70250 9158
rect 74118 9210 74170 9222
rect 74118 9146 74170 9158
rect 74454 9210 74506 9222
rect 74454 9146 74506 9158
rect 76750 9210 76802 9222
rect 76750 9146 76802 9158
rect 78654 9210 78706 9222
rect 78654 9146 78706 9158
rect 79606 9210 79658 9222
rect 79606 9146 79658 9158
rect 80502 9210 80554 9222
rect 80502 9146 80554 9158
rect 82518 9210 82570 9222
rect 86494 9210 86546 9222
rect 82518 9146 82570 9158
rect 86046 9154 86098 9166
rect 8990 9098 9042 9110
rect 46846 9098 46898 9110
rect 58382 9098 58434 9110
rect 10042 9046 10054 9098
rect 10106 9046 10118 9098
rect 10938 9046 10950 9098
rect 11002 9046 11014 9098
rect 8990 9034 9042 9046
rect 15094 9042 15146 9054
rect 21914 9046 21926 9098
rect 21978 9046 21990 9098
rect 25610 9046 25622 9098
rect 25674 9046 25686 9098
rect 42858 9046 42870 9098
rect 42922 9046 42934 9098
rect 45882 9046 45894 9098
rect 45946 9046 45958 9098
rect 48234 9046 48246 9098
rect 48298 9046 48310 9098
rect 14074 8990 14086 9042
rect 14138 8990 14150 9042
rect 15094 8978 15146 8990
rect 16046 8986 16098 8998
rect 23370 8990 23382 9042
rect 23434 8990 23446 9042
rect 46846 9034 46898 9046
rect 16046 8922 16098 8934
rect 26350 8986 26402 8998
rect 23034 8878 23046 8930
rect 23098 8878 23110 8930
rect 26350 8922 26402 8934
rect 36990 8986 37042 8998
rect 36990 8922 37042 8934
rect 38110 8986 38162 8998
rect 38110 8922 38162 8934
rect 41470 8986 41522 8998
rect 41470 8922 41522 8934
rect 49310 8986 49362 8998
rect 54842 8990 54854 9042
rect 54906 8990 54918 9042
rect 56410 9001 56422 9053
rect 56474 9001 56486 9053
rect 57418 9046 57430 9098
rect 57482 9046 57494 9098
rect 58382 9034 58434 9046
rect 58830 9098 58882 9110
rect 71262 9098 71314 9110
rect 86494 9146 86546 9158
rect 87726 9210 87778 9222
rect 87726 9146 87778 9158
rect 90694 9210 90746 9222
rect 90694 9146 90746 9158
rect 92206 9210 92258 9222
rect 92206 9146 92258 9158
rect 92822 9210 92874 9222
rect 92822 9146 92874 9158
rect 93158 9210 93210 9222
rect 93158 9146 93210 9158
rect 94894 9210 94946 9222
rect 97738 9214 97750 9266
rect 97802 9214 97814 9266
rect 94894 9146 94946 9158
rect 99766 9210 99818 9222
rect 99082 9102 99094 9154
rect 99146 9102 99158 9154
rect 99766 9146 99818 9158
rect 104302 9210 104354 9222
rect 104302 9146 104354 9158
rect 105142 9210 105194 9222
rect 105142 9146 105194 9158
rect 108334 9210 108386 9222
rect 108334 9146 108386 9158
rect 118414 9210 118466 9222
rect 129614 9210 129666 9222
rect 118414 9146 118466 9158
rect 118526 9154 118578 9166
rect 129614 9146 129666 9158
rect 130846 9210 130898 9222
rect 130846 9146 130898 9158
rect 131406 9210 131458 9222
rect 131406 9146 131458 9158
rect 141318 9210 141370 9222
rect 141318 9146 141370 9158
rect 141710 9210 141762 9222
rect 141710 9146 141762 9158
rect 146974 9210 147026 9222
rect 146974 9146 147026 9158
rect 159182 9210 159234 9222
rect 153066 9102 153078 9154
rect 153130 9102 153142 9154
rect 159182 9146 159234 9158
rect 159630 9210 159682 9222
rect 159630 9146 159682 9158
rect 161310 9210 161362 9222
rect 161310 9146 161362 9158
rect 166462 9210 166514 9222
rect 172566 9210 172618 9222
rect 166462 9146 166514 9158
rect 167918 9154 167970 9166
rect 62794 9046 62806 9098
rect 62858 9046 62870 9098
rect 69850 9046 69862 9098
rect 69914 9046 69926 9098
rect 79258 9046 79270 9098
rect 79322 9046 79334 9098
rect 80154 9046 80166 9098
rect 80218 9046 80230 9098
rect 81274 9046 81286 9098
rect 81338 9046 81350 9098
rect 82170 9046 82182 9098
rect 82234 9046 82246 9098
rect 86046 9090 86098 9102
rect 58830 9034 58882 9046
rect 71262 9034 71314 9046
rect 88398 9042 88450 9054
rect 90346 9046 90358 9098
rect 90410 9046 90422 9098
rect 49310 8922 49362 8934
rect 59390 8986 59442 8998
rect 59390 8922 59442 8934
rect 63534 8986 63586 8998
rect 63534 8922 63586 8934
rect 65326 8986 65378 8998
rect 65326 8922 65378 8934
rect 68686 8986 68738 8998
rect 68686 8922 68738 8934
rect 70590 8986 70642 8998
rect 70590 8922 70642 8934
rect 72046 8986 72098 8998
rect 72046 8922 72098 8934
rect 73278 8986 73330 8998
rect 73278 8922 73330 8934
rect 74846 8986 74898 8998
rect 74846 8922 74898 8934
rect 77758 8986 77810 8998
rect 77758 8922 77810 8934
rect 78206 8986 78258 8998
rect 83066 8990 83078 9042
rect 83130 8990 83142 9042
rect 78206 8922 78258 8934
rect 83806 8986 83858 8998
rect 83806 8922 83858 8934
rect 84254 8986 84306 8998
rect 84254 8922 84306 8934
rect 84702 8986 84754 8998
rect 84702 8922 84754 8934
rect 87054 8986 87106 8998
rect 91310 9042 91362 9054
rect 95946 9046 95958 9098
rect 96010 9046 96022 9098
rect 118526 9090 118578 9102
rect 161758 9098 161810 9110
rect 100830 9042 100882 9054
rect 140970 9046 140982 9098
rect 141034 9046 141046 9098
rect 160862 9042 160914 9054
rect 88398 8978 88450 8990
rect 89070 8986 89122 8998
rect 87054 8922 87106 8934
rect 89070 8922 89122 8934
rect 89742 8986 89794 8998
rect 91310 8978 91362 8990
rect 91758 8986 91810 8998
rect 89742 8922 89794 8934
rect 91758 8922 91810 8934
rect 95342 8986 95394 8998
rect 98970 8990 98982 9042
rect 99034 8990 99046 9042
rect 100830 8978 100882 8990
rect 101278 8986 101330 8998
rect 95342 8922 95394 8934
rect 101278 8922 101330 8934
rect 109230 8986 109282 8998
rect 109230 8922 109282 8934
rect 118974 8986 119026 8998
rect 118974 8922 119026 8934
rect 124798 8986 124850 8998
rect 131786 8990 131798 9042
rect 131850 8990 131862 9042
rect 133242 8990 133254 9042
rect 133306 8990 133318 9042
rect 134250 8990 134262 9042
rect 134314 8990 134326 9042
rect 135258 8990 135270 9042
rect 135322 8990 135334 9042
rect 124798 8922 124850 8934
rect 135774 8986 135826 8998
rect 137610 8990 137622 9042
rect 137674 8990 137686 9042
rect 138282 8990 138294 9042
rect 138346 8990 138358 9042
rect 138842 8990 138854 9042
rect 138906 8990 138918 9042
rect 140298 8990 140310 9042
rect 140362 8990 140374 9042
rect 142314 8990 142326 9042
rect 142378 8990 142390 9042
rect 143770 8990 143782 9042
rect 143834 8990 143846 9042
rect 145114 8990 145126 9042
rect 145178 8990 145190 9042
rect 146458 8990 146470 9042
rect 146522 8990 146534 9042
rect 46230 8874 46282 8886
rect 13066 8822 13078 8874
rect 13130 8822 13142 8874
rect 46230 8810 46282 8822
rect 53286 8874 53338 8886
rect 53286 8810 53338 8822
rect 58270 8874 58322 8886
rect 58270 8810 58322 8822
rect 63142 8874 63194 8886
rect 63142 8810 63194 8822
rect 81622 8874 81674 8886
rect 81622 8810 81674 8822
rect 83414 8874 83466 8886
rect 83414 8810 83466 8822
rect 85934 8874 85986 8886
rect 85934 8810 85986 8822
rect 88286 8874 88338 8886
rect 88286 8810 88338 8822
rect 91198 8874 91250 8886
rect 91198 8810 91250 8822
rect 96294 8874 96346 8886
rect 96294 8810 96346 8822
rect 100102 8874 100154 8886
rect 100102 8810 100154 8822
rect 100718 8874 100770 8886
rect 100718 8810 100770 8822
rect 105478 8874 105530 8886
rect 133130 8878 133142 8930
rect 133194 8878 133206 8930
rect 135370 8878 135382 8930
rect 135434 8878 135446 8930
rect 135774 8922 135826 8934
rect 147422 8986 147474 8998
rect 148138 8990 148150 9042
rect 148202 8990 148214 9042
rect 149482 8990 149494 9042
rect 149546 8990 149558 9042
rect 150490 8990 150502 9042
rect 150554 8990 150566 9042
rect 151834 8990 151846 9042
rect 151898 8990 151910 9042
rect 152954 8990 152966 9042
rect 153018 8990 153030 9042
rect 155194 8990 155206 9042
rect 155258 8990 155270 9042
rect 156314 8990 156326 9042
rect 156378 8990 156390 9042
rect 157210 8990 157222 9042
rect 157274 8990 157286 9042
rect 158666 8990 158678 9042
rect 158730 8990 158742 9042
rect 172566 9146 172618 9158
rect 175478 9210 175530 9222
rect 175478 9146 175530 9158
rect 176598 9210 176650 9222
rect 181850 9214 181862 9266
rect 181914 9214 181926 9266
rect 176598 9146 176650 9158
rect 190598 9210 190650 9222
rect 167918 9090 167970 9102
rect 170830 9098 170882 9110
rect 161758 9034 161810 9046
rect 166070 9042 166122 9054
rect 164378 8990 164390 9042
rect 164442 8990 164454 9042
rect 160862 8978 160914 8990
rect 166070 8978 166122 8990
rect 166910 8986 166962 8998
rect 168858 8990 168870 9042
rect 168922 8990 168934 9042
rect 170090 8990 170102 9042
rect 170154 8990 170166 9042
rect 170830 9034 170882 9046
rect 170942 9098 170994 9110
rect 182746 9102 182758 9154
rect 182810 9102 182822 9154
rect 185098 9102 185110 9154
rect 185162 9102 185174 9154
rect 186666 9102 186678 9154
rect 186730 9102 186742 9154
rect 188682 9102 188694 9154
rect 188746 9102 188758 9154
rect 190598 9146 190650 9158
rect 190934 9210 190986 9222
rect 190934 9146 190986 9158
rect 191438 9210 191490 9222
rect 191438 9146 191490 9158
rect 194518 9210 194570 9222
rect 192826 9102 192838 9154
rect 192890 9102 192902 9154
rect 194518 9146 194570 9158
rect 195414 9210 195466 9222
rect 195414 9146 195466 9158
rect 196310 9210 196362 9222
rect 196310 9146 196362 9158
rect 197206 9210 197258 9222
rect 197206 9146 197258 9158
rect 198046 9210 198098 9222
rect 198046 9146 198098 9158
rect 198494 9210 198546 9222
rect 198494 9146 198546 9158
rect 199390 9210 199442 9222
rect 199390 9146 199442 9158
rect 200398 9210 200450 9222
rect 200398 9146 200450 9158
rect 200846 9210 200898 9222
rect 200846 9146 200898 9158
rect 201294 9210 201346 9222
rect 201294 9146 201346 9158
rect 202190 9210 202242 9222
rect 202190 9146 202242 9158
rect 203254 9210 203306 9222
rect 203254 9146 203306 9158
rect 212774 9210 212826 9222
rect 207498 9102 207510 9154
rect 207562 9102 207574 9154
rect 209850 9102 209862 9154
rect 209914 9102 209926 9154
rect 211082 9102 211094 9154
rect 211146 9102 211158 9154
rect 212774 9146 212826 9158
rect 213110 9210 213162 9222
rect 213110 9146 213162 9158
rect 214846 9210 214898 9222
rect 214846 9146 214898 9158
rect 216750 9210 216802 9222
rect 216750 9146 216802 9158
rect 216302 9098 216354 9110
rect 170942 9034 170994 9046
rect 173338 8990 173350 9042
rect 173402 8990 173414 9042
rect 175030 9038 175082 9050
rect 175802 9046 175814 9098
rect 175866 9046 175878 9098
rect 176922 9046 176934 9098
rect 176986 9046 176998 9098
rect 140410 8878 140422 8930
rect 140474 8878 140486 8930
rect 143882 8878 143894 8930
rect 143946 8878 143958 8930
rect 147422 8922 147474 8934
rect 179610 8990 179622 9042
rect 179674 8990 179686 9042
rect 181302 9038 181354 9050
rect 194842 9046 194854 9098
rect 194906 9046 194918 9098
rect 195738 9046 195750 9098
rect 195802 9046 195814 9098
rect 196634 9046 196646 9098
rect 196698 9046 196710 9098
rect 197530 9046 197542 9098
rect 197594 9046 197606 9098
rect 202906 9046 202918 9098
rect 202970 9046 202982 9098
rect 175030 8974 175082 8986
rect 182970 8990 182982 9042
rect 183034 8990 183046 9042
rect 181302 8974 181354 8986
rect 183710 8986 183762 8998
rect 184538 8990 184550 9042
rect 184602 8990 184614 9042
rect 186554 8990 186566 9042
rect 186618 8990 186630 9042
rect 188570 8990 188582 9042
rect 188634 8990 188646 9042
rect 193050 8990 193062 9042
rect 193114 8990 193126 9042
rect 154410 8878 154422 8930
rect 154474 8878 154486 8930
rect 166910 8922 166962 8934
rect 183710 8922 183762 8934
rect 198942 8986 198994 8998
rect 160750 8874 160802 8886
rect 137386 8822 137398 8874
rect 137450 8822 137462 8874
rect 145562 8822 145574 8874
rect 145626 8822 145638 8874
rect 148586 8822 148598 8874
rect 148650 8822 148662 8874
rect 150938 8822 150950 8874
rect 151002 8822 151014 8874
rect 155418 8822 155430 8874
rect 155482 8822 155494 8874
rect 157770 8822 157782 8874
rect 157834 8822 157846 8874
rect 105478 8810 105530 8822
rect 160750 8810 160802 8822
rect 162822 8874 162874 8886
rect 162822 8810 162874 8822
rect 167806 8874 167858 8886
rect 186106 8878 186118 8930
rect 186170 8878 186182 8930
rect 187898 8878 187910 8930
rect 187962 8878 187974 8930
rect 192714 8878 192726 8930
rect 192778 8878 192790 8930
rect 198942 8922 198994 8934
rect 201742 8986 201794 8998
rect 204026 8990 204038 9042
rect 204090 8990 204102 9042
rect 206490 8990 206502 9042
rect 206554 8990 206566 9042
rect 209514 8990 209526 9042
rect 209578 8990 209590 9042
rect 211418 8990 211430 9042
rect 211482 8990 211494 9042
rect 216302 9034 216354 9046
rect 201742 8922 201794 8934
rect 213502 8986 213554 8998
rect 204138 8878 204150 8930
rect 204202 8878 204214 8930
rect 211978 8878 211990 8930
rect 212042 8878 212054 8930
rect 213502 8922 213554 8934
rect 213950 8986 214002 8998
rect 213950 8922 214002 8934
rect 214398 8986 214450 8998
rect 214398 8922 214450 8934
rect 215294 8986 215346 8998
rect 215294 8922 215346 8934
rect 169194 8822 169206 8874
rect 169258 8822 169270 8874
rect 179274 8822 179286 8874
rect 179338 8822 179350 8874
rect 189130 8822 189142 8874
rect 189194 8822 189206 8874
rect 206714 8822 206726 8874
rect 206778 8822 206790 8874
rect 167806 8810 167858 8822
rect 1344 8650 218624 8684
rect 1344 8598 28378 8650
rect 28430 8598 28482 8650
rect 28534 8598 28586 8650
rect 28638 8598 82706 8650
rect 82758 8598 82810 8650
rect 82862 8598 82914 8650
rect 82966 8598 137034 8650
rect 137086 8598 137138 8650
rect 137190 8598 137242 8650
rect 137294 8598 191362 8650
rect 191414 8598 191466 8650
rect 191518 8598 191570 8650
rect 191622 8598 218624 8650
rect 1344 8564 218624 8598
rect 21814 8426 21866 8438
rect 71766 8426 71818 8438
rect 16314 8374 16326 8426
rect 16378 8374 16390 8426
rect 56410 8374 56422 8426
rect 56474 8374 56486 8426
rect 70186 8374 70198 8426
rect 70250 8374 70262 8426
rect 21814 8362 21866 8374
rect 71766 8362 71818 8374
rect 87726 8426 87778 8438
rect 87726 8362 87778 8374
rect 90414 8426 90466 8438
rect 171334 8426 171386 8438
rect 186566 8426 186618 8438
rect 98298 8374 98310 8426
rect 98362 8374 98374 8426
rect 118906 8374 118918 8426
rect 118970 8374 118982 8426
rect 139514 8374 139526 8426
rect 139578 8374 139590 8426
rect 145674 8374 145686 8426
rect 145738 8374 145750 8426
rect 149258 8374 149270 8426
rect 149322 8374 149334 8426
rect 153962 8374 153974 8426
rect 154026 8374 154038 8426
rect 158890 8374 158902 8426
rect 158954 8374 158966 8426
rect 179050 8374 179062 8426
rect 179114 8374 179126 8426
rect 181514 8374 181526 8426
rect 181578 8374 181590 8426
rect 183530 8374 183542 8426
rect 183594 8374 183606 8426
rect 185546 8374 185558 8426
rect 185610 8374 185622 8426
rect 90414 8362 90466 8374
rect 10278 8314 10330 8326
rect 13582 8314 13634 8326
rect 10278 8250 10330 8262
rect 12854 8262 12906 8274
rect 11610 8206 11622 8258
rect 11674 8206 11686 8258
rect 26966 8314 27018 8326
rect 13582 8250 13634 8262
rect 18342 8258 18394 8270
rect 25062 8258 25114 8270
rect 12854 8198 12906 8210
rect 16650 8206 16662 8258
rect 16714 8206 16726 8258
rect 23370 8206 23382 8258
rect 23434 8206 23446 8258
rect 26966 8250 27018 8262
rect 29878 8314 29930 8326
rect 29878 8250 29930 8262
rect 31894 8314 31946 8326
rect 31894 8250 31946 8262
rect 34358 8314 34410 8326
rect 34358 8250 34410 8262
rect 35254 8314 35306 8326
rect 35254 8250 35306 8262
rect 36710 8314 36762 8326
rect 36710 8250 36762 8262
rect 37830 8314 37882 8326
rect 37830 8250 37882 8262
rect 39062 8314 39114 8326
rect 39062 8250 39114 8262
rect 39958 8314 40010 8326
rect 39958 8250 40010 8262
rect 41078 8314 41130 8326
rect 41078 8250 41130 8262
rect 41974 8314 42026 8326
rect 41974 8250 42026 8262
rect 42870 8314 42922 8326
rect 42870 8250 42922 8262
rect 43766 8314 43818 8326
rect 43766 8250 43818 8262
rect 44662 8314 44714 8326
rect 44662 8250 44714 8262
rect 45894 8314 45946 8326
rect 45894 8250 45946 8262
rect 46790 8314 46842 8326
rect 46790 8250 46842 8262
rect 47686 8314 47738 8326
rect 47686 8250 47738 8262
rect 48582 8314 48634 8326
rect 48582 8250 48634 8262
rect 50038 8314 50090 8326
rect 54406 8314 54458 8326
rect 50038 8250 50090 8262
rect 52614 8258 52666 8270
rect 51594 8206 51606 8258
rect 51658 8206 51670 8258
rect 59334 8314 59386 8326
rect 54406 8250 54458 8262
rect 58438 8258 58490 8270
rect 56746 8206 56758 8258
rect 56810 8206 56822 8258
rect 59334 8250 59386 8262
rect 62358 8314 62410 8326
rect 66558 8314 66610 8326
rect 62358 8250 62410 8262
rect 64934 8262 64986 8274
rect 63242 8206 63254 8258
rect 63306 8206 63318 8258
rect 66558 8250 66610 8262
rect 67398 8314 67450 8326
rect 73782 8314 73834 8326
rect 67398 8250 67450 8262
rect 68462 8258 68514 8270
rect 77982 8314 78034 8326
rect 18342 8194 18394 8206
rect 25062 8194 25114 8206
rect 26618 8150 26630 8202
rect 26682 8150 26694 8202
rect 29530 8150 29542 8202
rect 29594 8150 29606 8202
rect 31546 8150 31558 8202
rect 31610 8150 31622 8202
rect 34906 8150 34918 8202
rect 34970 8150 34982 8202
rect 45546 8150 45558 8202
rect 45610 8150 45622 8202
rect 48234 8150 48246 8202
rect 48298 8150 48310 8202
rect 52614 8194 52666 8206
rect 58438 8194 58490 8206
rect 58986 8150 58998 8202
rect 59050 8150 59062 8202
rect 64934 8198 64986 8210
rect 66054 8202 66106 8214
rect 59950 8146 60002 8158
rect 65706 8150 65718 8202
rect 65770 8150 65782 8202
rect 70746 8206 70758 8258
rect 70810 8206 70822 8258
rect 73782 8250 73834 8262
rect 76470 8258 76522 8270
rect 74778 8206 74790 8258
rect 74842 8206 74854 8258
rect 89910 8314 89962 8326
rect 93930 8318 93942 8370
rect 93994 8318 94006 8370
rect 101658 8318 101670 8370
rect 101722 8318 101734 8370
rect 171334 8362 171386 8374
rect 186566 8362 186618 8374
rect 199670 8426 199722 8438
rect 199670 8362 199722 8374
rect 77982 8250 78034 8262
rect 84422 8258 84474 8270
rect 83290 8206 83302 8258
rect 83354 8206 83366 8258
rect 68462 8194 68514 8206
rect 71418 8150 71430 8202
rect 71482 8150 71494 8202
rect 76470 8194 76522 8206
rect 84422 8194 84474 8206
rect 88510 8258 88562 8270
rect 107886 8314 107938 8326
rect 89910 8250 89962 8262
rect 100326 8262 100378 8274
rect 13918 8090 13970 8102
rect 13918 8026 13970 8038
rect 18734 8090 18786 8102
rect 18734 8026 18786 8038
rect 19182 8090 19234 8102
rect 19182 8026 19234 8038
rect 25454 8090 25506 8102
rect 25454 8026 25506 8038
rect 25902 8090 25954 8102
rect 25902 8026 25954 8038
rect 27470 8090 27522 8102
rect 27470 8026 27522 8038
rect 30382 8090 30434 8102
rect 30382 8026 30434 8038
rect 32398 8090 32450 8102
rect 32398 8026 32450 8038
rect 34022 8090 34074 8102
rect 34022 8026 34074 8038
rect 35758 8090 35810 8102
rect 35758 8026 35810 8038
rect 36374 8090 36426 8102
rect 36374 8026 36426 8038
rect 37494 8090 37546 8102
rect 37494 8026 37546 8038
rect 38726 8090 38778 8102
rect 38726 8026 38778 8038
rect 39622 8090 39674 8102
rect 39622 8026 39674 8038
rect 40742 8090 40794 8102
rect 40742 8026 40794 8038
rect 41638 8090 41690 8102
rect 41638 8026 41690 8038
rect 42534 8090 42586 8102
rect 42534 8026 42586 8038
rect 43430 8090 43482 8102
rect 43430 8026 43482 8038
rect 44326 8090 44378 8102
rect 44326 8026 44378 8038
rect 46454 8090 46506 8102
rect 46454 8026 46506 8038
rect 47350 8090 47402 8102
rect 47350 8026 47402 8038
rect 53566 8090 53618 8102
rect 53566 8026 53618 8038
rect 54070 8090 54122 8102
rect 54070 8026 54122 8038
rect 59838 8090 59890 8102
rect 66054 8138 66106 8150
rect 79438 8146 79490 8158
rect 59950 8082 60002 8094
rect 60510 8090 60562 8102
rect 59838 8026 59890 8038
rect 60510 8026 60562 8038
rect 67062 8090 67114 8102
rect 67062 8026 67114 8038
rect 67902 8090 67954 8102
rect 67902 8026 67954 8038
rect 68350 8090 68402 8102
rect 70634 8094 70646 8146
rect 70698 8094 70710 8146
rect 68350 8026 68402 8038
rect 72382 8090 72434 8102
rect 72382 8026 72434 8038
rect 78318 8090 78370 8102
rect 78318 8026 78370 8038
rect 78878 8090 78930 8102
rect 78878 8026 78930 8038
rect 79326 8090 79378 8102
rect 85822 8146 85874 8158
rect 86538 8150 86550 8202
rect 86602 8150 86614 8202
rect 88510 8194 88562 8206
rect 91198 8202 91250 8214
rect 79438 8082 79490 8094
rect 80054 8090 80106 8102
rect 79326 8026 79378 8038
rect 80054 8026 80106 8038
rect 80390 8090 80442 8102
rect 80390 8026 80442 8038
rect 81958 8090 82010 8102
rect 81958 8026 82010 8038
rect 85262 8090 85314 8102
rect 85262 8026 85314 8038
rect 85710 8090 85762 8102
rect 87838 8146 87890 8158
rect 85822 8082 85874 8094
rect 86886 8090 86938 8102
rect 85710 8026 85762 8038
rect 90526 8146 90578 8158
rect 87838 8082 87890 8094
rect 88398 8090 88450 8102
rect 86886 8026 86938 8038
rect 88398 8026 88450 8038
rect 89070 8090 89122 8102
rect 89070 8026 89122 8038
rect 89574 8090 89626 8102
rect 91198 8138 91250 8150
rect 91646 8202 91698 8214
rect 94826 8206 94838 8258
rect 94890 8206 94902 8258
rect 98634 8206 98646 8258
rect 98698 8206 98710 8258
rect 132078 8314 132130 8326
rect 100326 8198 100378 8210
rect 102554 8206 102566 8258
rect 102618 8206 102630 8258
rect 107886 8250 107938 8262
rect 110462 8258 110514 8270
rect 117002 8225 117014 8277
rect 117066 8225 117078 8277
rect 110462 8194 110514 8206
rect 116174 8202 116226 8214
rect 117898 8206 117910 8258
rect 117962 8206 117974 8258
rect 125066 8225 125078 8277
rect 125130 8225 125142 8277
rect 130510 8258 130562 8270
rect 125962 8206 125974 8258
rect 126026 8206 126038 8258
rect 132078 8250 132130 8262
rect 133590 8314 133642 8326
rect 133590 8250 133642 8262
rect 133982 8314 134034 8326
rect 133982 8250 134034 8262
rect 147086 8314 147138 8326
rect 91646 8138 91698 8150
rect 130510 8194 130562 8206
rect 130958 8202 131010 8214
rect 90526 8082 90578 8094
rect 91086 8090 91138 8102
rect 95386 8094 95398 8146
rect 95450 8094 95462 8146
rect 89574 8026 89626 8038
rect 91086 8026 91138 8038
rect 96238 8090 96290 8102
rect 103002 8094 103014 8146
rect 103066 8094 103078 8146
rect 116174 8138 116226 8150
rect 123342 8146 123394 8158
rect 96238 8026 96290 8038
rect 103630 8090 103682 8102
rect 103630 8026 103682 8038
rect 104078 8090 104130 8102
rect 104078 8026 104130 8038
rect 104526 8090 104578 8102
rect 104526 8026 104578 8038
rect 107550 8090 107602 8102
rect 107550 8026 107602 8038
rect 110350 8090 110402 8102
rect 110350 8026 110402 8038
rect 110910 8090 110962 8102
rect 110910 8026 110962 8038
rect 121662 8090 121714 8102
rect 121662 8026 121714 8038
rect 123230 8090 123282 8102
rect 133242 8150 133254 8202
rect 133306 8150 133318 8202
rect 134586 8195 134598 8247
rect 134650 8195 134662 8247
rect 135482 8206 135494 8258
rect 135546 8206 135558 8258
rect 139178 8206 139190 8258
rect 139242 8206 139254 8258
rect 143322 8206 143334 8258
rect 143386 8206 143398 8258
rect 144218 8195 144230 8247
rect 144282 8195 144294 8247
rect 145114 8206 145126 8258
rect 145178 8206 145190 8258
rect 146570 8206 146582 8258
rect 146634 8206 146646 8258
rect 147086 8250 147138 8262
rect 147534 8314 147586 8326
rect 147534 8250 147586 8262
rect 151118 8314 151170 8326
rect 190486 8314 190538 8326
rect 148698 8206 148710 8258
rect 148762 8206 148774 8258
rect 151118 8250 151170 8262
rect 151902 8258 151954 8270
rect 155990 8258 156042 8270
rect 160918 8258 160970 8270
rect 163886 8258 163938 8270
rect 170774 8258 170826 8270
rect 177606 8258 177658 8270
rect 187630 8258 187682 8270
rect 200398 8314 200450 8326
rect 150670 8202 150722 8214
rect 154298 8206 154310 8258
rect 154362 8206 154374 8258
rect 159226 8206 159238 8258
rect 159290 8206 159302 8258
rect 161466 8206 161478 8258
rect 161530 8206 161542 8258
rect 164714 8206 164726 8258
rect 164778 8206 164790 8258
rect 166954 8206 166966 8258
rect 167018 8206 167030 8258
rect 175914 8206 175926 8258
rect 175978 8206 175990 8258
rect 179162 8206 179174 8258
rect 179226 8206 179238 8258
rect 181178 8206 181190 8258
rect 181242 8206 181254 8258
rect 182858 8206 182870 8258
rect 182922 8206 182934 8258
rect 186106 8206 186118 8258
rect 186170 8206 186182 8258
rect 151902 8194 151954 8206
rect 155990 8194 156042 8206
rect 160918 8194 160970 8206
rect 163886 8194 163938 8206
rect 170774 8194 170826 8206
rect 177606 8194 177658 8206
rect 187518 8202 187570 8214
rect 130958 8138 131010 8150
rect 123342 8082 123394 8094
rect 123790 8090 123842 8102
rect 129054 8090 129106 8102
rect 123230 8026 123282 8038
rect 127530 8038 127542 8090
rect 127594 8038 127606 8090
rect 123790 8026 123842 8038
rect 129054 8026 129106 8038
rect 130398 8090 130450 8102
rect 130398 8026 130450 8038
rect 131630 8090 131682 8102
rect 138954 8094 138966 8146
rect 139018 8094 139030 8146
rect 141878 8090 141930 8102
rect 137274 8038 137286 8090
rect 137338 8038 137350 8090
rect 131630 8026 131682 8038
rect 141878 8026 141930 8038
rect 147982 8090 148034 8102
rect 150042 8094 150054 8146
rect 150106 8094 150118 8146
rect 150670 8138 150722 8150
rect 188458 8206 188470 8258
rect 188522 8206 188534 8258
rect 190486 8250 190538 8262
rect 196422 8258 196474 8270
rect 187630 8194 187682 8206
rect 192266 8195 192278 8247
rect 192330 8195 192342 8247
rect 193610 8206 193622 8258
rect 193674 8206 193686 8258
rect 197530 8206 197542 8258
rect 197594 8206 197606 8258
rect 200398 8250 200450 8262
rect 201406 8314 201458 8326
rect 201406 8250 201458 8262
rect 204318 8314 204370 8326
rect 204318 8250 204370 8262
rect 205942 8314 205994 8326
rect 209850 8318 209862 8370
rect 209914 8318 209926 8370
rect 211262 8314 211314 8326
rect 205942 8250 205994 8262
rect 208630 8258 208682 8270
rect 196422 8194 196474 8206
rect 202190 8202 202242 8214
rect 206938 8206 206950 8258
rect 207002 8206 207014 8258
rect 209178 8206 209190 8258
rect 209242 8206 209254 8258
rect 211262 8250 211314 8262
rect 215070 8314 215122 8326
rect 215070 8250 215122 8262
rect 215518 8314 215570 8326
rect 215518 8250 215570 8262
rect 147982 8026 148034 8038
rect 151790 8090 151842 8102
rect 151790 8026 151842 8038
rect 156606 8090 156658 8102
rect 162362 8094 162374 8146
rect 162426 8094 162438 8146
rect 156606 8026 156658 8038
rect 163774 8090 163826 8102
rect 166058 8094 166070 8146
rect 166122 8094 166134 8146
rect 167402 8094 167414 8146
rect 167466 8094 167478 8146
rect 169306 8094 169318 8146
rect 169370 8094 169382 8146
rect 163774 8026 163826 8038
rect 171670 8090 171722 8102
rect 171670 8026 171722 8038
rect 172566 8090 172618 8102
rect 172566 8026 172618 8038
rect 172902 8090 172954 8102
rect 172902 8026 172954 8038
rect 173406 8090 173458 8102
rect 179386 8094 179398 8146
rect 179450 8094 179462 8146
rect 180954 8094 180966 8146
rect 181018 8094 181030 8146
rect 182970 8094 182982 8146
rect 183034 8094 183046 8146
rect 185882 8094 185894 8146
rect 185946 8094 185958 8146
rect 187518 8138 187570 8150
rect 208630 8194 208682 8206
rect 214510 8202 214562 8214
rect 186902 8090 186954 8102
rect 188682 8094 188694 8146
rect 188746 8094 188758 8146
rect 202190 8138 202242 8150
rect 214510 8138 214562 8150
rect 175018 8038 175030 8090
rect 175082 8038 175094 8090
rect 173406 8026 173458 8038
rect 186902 8026 186954 8038
rect 190822 8090 190874 8102
rect 189354 7982 189366 8034
rect 189418 7982 189430 8034
rect 190822 8026 190874 8038
rect 191326 8090 191378 8102
rect 191326 8026 191378 8038
rect 194630 8090 194682 8102
rect 194630 8026 194682 8038
rect 200846 8090 200898 8102
rect 200846 8026 200898 8038
rect 201742 8090 201794 8102
rect 201742 8026 201794 8038
rect 202638 8090 202690 8102
rect 202638 8026 202690 8038
rect 203086 8090 203138 8102
rect 203086 8026 203138 8038
rect 203646 8090 203698 8102
rect 203646 8026 203698 8038
rect 212270 8090 212322 8102
rect 212270 8026 212322 8038
rect 212718 8090 212770 8102
rect 212718 8026 212770 8038
rect 213166 8090 213218 8102
rect 213166 8026 213218 8038
rect 213614 8090 213666 8102
rect 213614 8026 213666 8038
rect 214062 8090 214114 8102
rect 214062 8026 214114 8038
rect 215854 8090 215906 8102
rect 215854 8026 215906 8038
rect 216302 8090 216354 8102
rect 216302 8026 216354 8038
rect 1344 7866 218624 7900
rect 1344 7814 55542 7866
rect 55594 7814 55646 7866
rect 55698 7814 55750 7866
rect 55802 7814 109870 7866
rect 109922 7814 109974 7866
rect 110026 7814 110078 7866
rect 110130 7814 164198 7866
rect 164250 7814 164302 7866
rect 164354 7814 164406 7866
rect 164458 7814 218624 7866
rect 1344 7780 218624 7814
rect 6470 7642 6522 7654
rect 6470 7578 6522 7590
rect 9550 7642 9602 7654
rect 9550 7578 9602 7590
rect 21590 7642 21642 7654
rect 40798 7642 40850 7654
rect 26842 7590 26854 7642
rect 26906 7590 26918 7642
rect 21590 7578 21642 7590
rect 40798 7578 40850 7590
rect 42198 7642 42250 7654
rect 42198 7578 42250 7590
rect 43094 7642 43146 7654
rect 43094 7578 43146 7590
rect 46230 7642 46282 7654
rect 46230 7578 46282 7590
rect 49814 7642 49866 7654
rect 50698 7646 50710 7698
rect 50762 7646 50774 7698
rect 49814 7578 49866 7590
rect 59502 7642 59554 7654
rect 51930 7534 51942 7586
rect 51994 7534 52006 7586
rect 58650 7534 58662 7586
rect 58714 7534 58726 7586
rect 59502 7578 59554 7590
rect 63422 7642 63474 7654
rect 62906 7534 62918 7586
rect 62970 7534 62982 7586
rect 63422 7578 63474 7590
rect 63870 7642 63922 7654
rect 63870 7578 63922 7590
rect 79438 7642 79490 7654
rect 66714 7534 66726 7586
rect 66778 7534 66790 7586
rect 74666 7534 74678 7586
rect 74730 7534 74742 7586
rect 78362 7534 78374 7586
rect 78426 7534 78438 7586
rect 79438 7578 79490 7590
rect 88510 7642 88562 7654
rect 115950 7642 116002 7654
rect 118794 7646 118806 7698
rect 118858 7646 118870 7698
rect 95610 7590 95622 7642
rect 95674 7590 95686 7642
rect 84858 7534 84870 7586
rect 84922 7534 84934 7586
rect 87210 7534 87222 7586
rect 87274 7534 87286 7586
rect 88510 7578 88562 7590
rect 90346 7534 90358 7586
rect 90410 7534 90422 7586
rect 104122 7534 104134 7586
rect 104186 7534 104198 7586
rect 107146 7534 107158 7586
rect 107210 7534 107222 7586
rect 115434 7534 115446 7586
rect 115498 7534 115510 7586
rect 115950 7578 116002 7590
rect 120878 7642 120930 7654
rect 117786 7534 117798 7586
rect 117850 7534 117862 7586
rect 119914 7534 119926 7586
rect 119978 7534 119990 7586
rect 120878 7578 120930 7590
rect 126702 7642 126754 7654
rect 127262 7642 127314 7654
rect 126702 7578 126754 7590
rect 126814 7586 126866 7598
rect 127262 7578 127314 7590
rect 135214 7642 135266 7654
rect 133578 7534 133590 7586
rect 133642 7534 133654 7586
rect 135214 7578 135266 7590
rect 135998 7642 136050 7654
rect 135998 7578 136050 7590
rect 142830 7642 142882 7654
rect 139962 7534 139974 7586
rect 140026 7534 140038 7586
rect 142830 7578 142882 7590
rect 143726 7642 143778 7654
rect 143726 7578 143778 7590
rect 145294 7642 145346 7654
rect 145294 7578 145346 7590
rect 150446 7642 150498 7654
rect 150446 7578 150498 7590
rect 151006 7642 151058 7654
rect 151006 7578 151058 7590
rect 151342 7642 151394 7654
rect 151342 7578 151394 7590
rect 151790 7642 151842 7654
rect 151790 7578 151842 7590
rect 157166 7642 157218 7654
rect 8934 7474 8986 7486
rect 7914 7422 7926 7474
rect 7978 7422 7990 7474
rect 8934 7410 8986 7422
rect 10334 7418 10386 7430
rect 12730 7422 12742 7474
rect 12794 7422 12806 7474
rect 15866 7422 15878 7474
rect 15930 7422 15942 7474
rect 16886 7470 16938 7482
rect 16886 7406 16938 7418
rect 17614 7418 17666 7430
rect 10334 7354 10386 7366
rect 11386 7310 11398 7362
rect 11450 7310 11462 7362
rect 17614 7354 17666 7366
rect 18062 7418 18114 7430
rect 18062 7354 18114 7366
rect 18622 7418 18674 7430
rect 18622 7354 18674 7366
rect 19182 7418 19234 7430
rect 23034 7422 23046 7474
rect 23098 7422 23110 7474
rect 24054 7470 24106 7482
rect 24054 7406 24106 7418
rect 24558 7418 24610 7430
rect 19182 7354 19234 7366
rect 24558 7354 24610 7366
rect 25566 7418 25618 7430
rect 28186 7422 28198 7474
rect 28250 7422 28262 7474
rect 29654 7470 29706 7482
rect 41850 7478 41862 7530
rect 41914 7478 41926 7530
rect 42746 7478 42758 7530
rect 42810 7478 42822 7530
rect 43642 7478 43654 7530
rect 43706 7478 43718 7530
rect 49466 7478 49478 7530
rect 49530 7478 49542 7530
rect 56646 7474 56698 7486
rect 72550 7474 72602 7486
rect 79550 7474 79602 7486
rect 80154 7478 80166 7530
rect 80218 7478 80230 7530
rect 126814 7522 126866 7534
rect 149998 7530 150050 7542
rect 152954 7534 152966 7586
rect 153018 7534 153030 7586
rect 156090 7534 156102 7586
rect 156154 7534 156166 7586
rect 157166 7578 157218 7590
rect 166966 7642 167018 7654
rect 174918 7642 174970 7654
rect 169418 7590 169430 7642
rect 169482 7590 169494 7642
rect 166966 7578 167018 7590
rect 174918 7578 174970 7590
rect 177718 7642 177770 7654
rect 183710 7642 183762 7654
rect 184762 7646 184774 7698
rect 184826 7646 184838 7698
rect 177718 7578 177770 7590
rect 180798 7586 180850 7598
rect 175758 7530 175810 7542
rect 29654 7406 29706 7418
rect 30158 7418 30210 7430
rect 25566 7354 25618 7366
rect 30158 7354 30210 7366
rect 30606 7418 30658 7430
rect 30606 7354 30658 7366
rect 34526 7418 34578 7430
rect 37818 7422 37830 7474
rect 37882 7422 37894 7474
rect 38714 7403 38726 7455
rect 38778 7403 38790 7455
rect 39230 7418 39282 7430
rect 34526 7354 34578 7366
rect 39230 7354 39282 7366
rect 39790 7418 39842 7430
rect 39790 7354 39842 7366
rect 40126 7418 40178 7430
rect 40126 7354 40178 7366
rect 44606 7418 44658 7430
rect 47674 7422 47686 7474
rect 47738 7422 47750 7474
rect 48570 7403 48582 7455
rect 48634 7403 48646 7455
rect 52154 7422 52166 7474
rect 52218 7422 52230 7474
rect 52670 7418 52722 7430
rect 54954 7422 54966 7474
rect 55018 7422 55030 7474
rect 58986 7422 58998 7474
rect 59050 7422 59062 7474
rect 44606 7354 44658 7366
rect 56646 7410 56698 7422
rect 60174 7418 60226 7430
rect 63018 7422 63030 7474
rect 63082 7422 63094 7474
rect 66378 7422 66390 7474
rect 66442 7422 66454 7474
rect 52670 7354 52722 7366
rect 43990 7306 44042 7318
rect 14858 7254 14870 7306
rect 14922 7254 14934 7306
rect 36810 7254 36822 7306
rect 36874 7254 36886 7306
rect 43990 7242 44042 7254
rect 53398 7306 53450 7318
rect 57418 7310 57430 7362
rect 57482 7310 57494 7362
rect 60174 7354 60226 7366
rect 67230 7418 67282 7430
rect 67230 7354 67282 7366
rect 68126 7418 68178 7430
rect 68126 7354 68178 7366
rect 68574 7418 68626 7430
rect 70858 7422 70870 7474
rect 70922 7422 70934 7474
rect 74554 7422 74566 7474
rect 74618 7422 74630 7474
rect 72550 7410 72602 7422
rect 75182 7418 75234 7430
rect 68574 7354 68626 7366
rect 75182 7354 75234 7366
rect 75630 7418 75682 7430
rect 75630 7354 75682 7366
rect 76078 7418 76130 7430
rect 78026 7422 78038 7474
rect 78090 7422 78102 7474
rect 76078 7354 76130 7366
rect 78878 7418 78930 7430
rect 81274 7422 81286 7474
rect 81338 7422 81350 7474
rect 81834 7422 81846 7474
rect 81898 7422 81910 7474
rect 84970 7422 84982 7474
rect 85034 7422 85046 7474
rect 79550 7410 79602 7422
rect 85374 7418 85426 7430
rect 87434 7422 87446 7474
rect 87498 7422 87510 7474
rect 78878 7354 78930 7366
rect 80502 7306 80554 7318
rect 81162 7310 81174 7362
rect 81226 7310 81238 7362
rect 85374 7354 85426 7366
rect 87950 7418 88002 7430
rect 90570 7422 90582 7474
rect 90634 7422 90646 7474
rect 92822 7470 92874 7482
rect 85978 7310 85990 7362
rect 86042 7310 86054 7362
rect 87950 7354 88002 7366
rect 91086 7418 91138 7430
rect 89114 7310 89126 7362
rect 89178 7310 89190 7362
rect 91086 7354 91138 7366
rect 91534 7418 91586 7430
rect 91534 7354 91586 7366
rect 92430 7418 92482 7430
rect 93818 7422 93830 7474
rect 93882 7422 93894 7474
rect 98086 7470 98138 7482
rect 92822 7406 92874 7418
rect 97694 7418 97746 7430
rect 92430 7354 92482 7366
rect 99082 7422 99094 7474
rect 99146 7422 99158 7474
rect 98086 7406 98138 7418
rect 100662 7418 100714 7430
rect 104234 7422 104246 7474
rect 104298 7422 104310 7474
rect 97694 7354 97746 7366
rect 100662 7354 100714 7366
rect 104974 7418 105026 7430
rect 107258 7422 107270 7474
rect 107322 7422 107334 7474
rect 107818 7403 107830 7455
rect 107882 7403 107894 7455
rect 108714 7422 108726 7474
rect 108778 7422 108790 7474
rect 115546 7422 115558 7474
rect 115610 7422 115622 7474
rect 118122 7422 118134 7474
rect 118186 7422 118198 7474
rect 120250 7422 120262 7474
rect 120314 7422 120326 7474
rect 121930 7433 121942 7485
rect 121994 7433 122006 7485
rect 136110 7474 136162 7486
rect 143614 7474 143666 7486
rect 121326 7418 121378 7430
rect 122826 7422 122838 7474
rect 122890 7422 122902 7474
rect 102778 7310 102790 7362
rect 102842 7310 102854 7362
rect 104974 7354 105026 7366
rect 105690 7310 105702 7362
rect 105754 7310 105766 7362
rect 110966 7306 111018 7318
rect 113978 7310 113990 7362
rect 114042 7310 114054 7362
rect 117002 7310 117014 7362
rect 117066 7310 117078 7362
rect 121326 7354 121378 7366
rect 128270 7418 128322 7430
rect 129378 7422 129390 7474
rect 129442 7422 129454 7474
rect 130218 7422 130230 7474
rect 130282 7422 130294 7474
rect 133354 7422 133366 7474
rect 133418 7422 133430 7474
rect 136938 7422 136950 7474
rect 137002 7422 137014 7474
rect 138282 7422 138294 7474
rect 138346 7422 138358 7474
rect 140298 7422 140310 7474
rect 140362 7422 140374 7474
rect 140970 7422 140982 7474
rect 141034 7422 141046 7474
rect 142426 7422 142438 7474
rect 142490 7422 142502 7474
rect 136110 7410 136162 7422
rect 143614 7410 143666 7422
rect 144734 7418 144786 7430
rect 147914 7422 147926 7474
rect 147978 7422 147990 7474
rect 149606 7470 149658 7482
rect 128270 7354 128322 7366
rect 149998 7466 150050 7478
rect 164278 7474 164330 7486
rect 167290 7478 167302 7530
rect 167354 7478 167366 7530
rect 172230 7474 172282 7486
rect 153402 7422 153414 7474
rect 153466 7422 153478 7474
rect 155530 7422 155542 7474
rect 155594 7422 155606 7474
rect 149606 7406 149658 7418
rect 156718 7418 156770 7430
rect 144734 7354 144786 7366
rect 156718 7354 156770 7366
rect 157614 7418 157666 7430
rect 159450 7422 159462 7474
rect 159514 7422 159526 7474
rect 162586 7422 162598 7474
rect 162650 7422 162662 7474
rect 164826 7422 164838 7474
rect 164890 7422 164902 7474
rect 164278 7410 164330 7422
rect 167806 7418 167858 7430
rect 170650 7422 170662 7474
rect 170714 7422 170726 7474
rect 157614 7354 157666 7366
rect 172230 7410 172282 7422
rect 174358 7474 174410 7486
rect 175242 7478 175254 7530
rect 175306 7478 175318 7530
rect 190598 7642 190650 7654
rect 183710 7578 183762 7590
rect 183822 7586 183874 7598
rect 180798 7522 180850 7534
rect 189914 7534 189926 7586
rect 189978 7534 189990 7586
rect 190598 7578 190650 7590
rect 190934 7642 190986 7654
rect 192446 7642 192498 7654
rect 190934 7578 190986 7590
rect 191774 7586 191826 7598
rect 192446 7578 192498 7590
rect 192894 7642 192946 7654
rect 192894 7578 192946 7590
rect 193790 7642 193842 7654
rect 195134 7642 195186 7654
rect 193790 7578 193842 7590
rect 193902 7586 193954 7598
rect 183822 7522 183874 7534
rect 191774 7522 191826 7534
rect 193902 7522 193954 7534
rect 195022 7586 195074 7598
rect 195134 7578 195186 7590
rect 195582 7642 195634 7654
rect 195582 7578 195634 7590
rect 196030 7642 196082 7654
rect 196030 7578 196082 7590
rect 196926 7642 196978 7654
rect 196926 7578 196978 7590
rect 197374 7642 197426 7654
rect 197374 7578 197426 7590
rect 198270 7642 198322 7654
rect 198270 7578 198322 7590
rect 198718 7642 198770 7654
rect 198718 7578 198770 7590
rect 203086 7642 203138 7654
rect 203086 7578 203138 7590
rect 210870 7642 210922 7654
rect 195022 7522 195074 7534
rect 199614 7530 199666 7542
rect 209626 7534 209638 7586
rect 209690 7534 209702 7586
rect 210870 7578 210922 7590
rect 211710 7642 211762 7654
rect 211710 7578 211762 7590
rect 212158 7642 212210 7654
rect 212158 7578 212210 7590
rect 212606 7642 212658 7654
rect 212606 7578 212658 7590
rect 213054 7642 213106 7654
rect 213054 7578 213106 7590
rect 215294 7642 215346 7654
rect 215294 7578 215346 7590
rect 213950 7530 214002 7542
rect 175758 7466 175810 7478
rect 178490 7422 178502 7474
rect 178554 7422 178566 7474
rect 180182 7470 180234 7482
rect 174358 7410 174410 7422
rect 182970 7422 182982 7474
rect 183034 7422 183046 7474
rect 184650 7422 184662 7474
rect 184714 7422 184726 7474
rect 185770 7422 185782 7474
rect 185834 7422 185846 7474
rect 186666 7422 186678 7474
rect 186730 7422 186742 7474
rect 188010 7422 188022 7474
rect 188074 7422 188086 7474
rect 189690 7422 189702 7474
rect 189754 7422 189766 7474
rect 199614 7466 199666 7478
rect 180182 7406 180234 7418
rect 194350 7418 194402 7430
rect 132470 7306 132522 7318
rect 158442 7310 158454 7362
rect 158506 7310 158518 7362
rect 161030 7306 161082 7318
rect 166170 7310 166182 7362
rect 166234 7310 166246 7362
rect 167806 7354 167858 7366
rect 173114 7310 173126 7362
rect 173178 7310 173190 7362
rect 62458 7254 62470 7306
rect 62522 7254 62534 7306
rect 66266 7254 66278 7306
rect 66330 7254 66342 7306
rect 70522 7254 70534 7306
rect 70586 7254 70598 7306
rect 74218 7254 74230 7306
rect 74282 7254 74294 7306
rect 77914 7254 77926 7306
rect 77978 7254 77990 7306
rect 84410 7254 84422 7306
rect 84474 7254 84486 7306
rect 123834 7254 123846 7306
rect 123898 7254 123910 7306
rect 133802 7254 133814 7306
rect 133866 7254 133878 7306
rect 137386 7254 137398 7306
rect 137450 7254 137462 7306
rect 139850 7254 139862 7306
rect 139914 7254 139926 7306
rect 141866 7254 141878 7306
rect 141930 7254 141942 7306
rect 147578 7254 147590 7306
rect 147642 7254 147654 7306
rect 153738 7254 153750 7306
rect 153802 7254 153814 7306
rect 155306 7254 155318 7306
rect 155370 7254 155382 7306
rect 53398 7242 53450 7254
rect 80502 7242 80554 7254
rect 110966 7242 111018 7254
rect 132470 7242 132522 7254
rect 161030 7242 161082 7254
rect 180686 7306 180738 7318
rect 181626 7310 181638 7362
rect 181690 7310 181702 7362
rect 186554 7310 186566 7362
rect 186618 7310 186630 7362
rect 194350 7354 194402 7366
rect 196478 7418 196530 7430
rect 196478 7354 196530 7366
rect 197822 7418 197874 7430
rect 197822 7354 197874 7366
rect 199166 7418 199218 7430
rect 200554 7422 200566 7474
rect 200618 7422 200630 7474
rect 199166 7354 199218 7366
rect 202638 7418 202690 7430
rect 191662 7306 191714 7318
rect 201562 7310 201574 7362
rect 201626 7310 201638 7362
rect 202638 7354 202690 7366
rect 203534 7418 203586 7430
rect 206042 7422 206054 7474
rect 206106 7422 206118 7474
rect 207734 7470 207786 7482
rect 210522 7478 210534 7530
rect 210586 7478 210598 7530
rect 209850 7422 209862 7474
rect 209914 7422 209926 7474
rect 213950 7466 214002 7478
rect 207734 7406 207786 7418
rect 211262 7418 211314 7430
rect 203534 7354 203586 7366
rect 189578 7254 189590 7306
rect 189642 7254 189654 7306
rect 180686 7242 180738 7254
rect 191662 7242 191714 7254
rect 204486 7306 204538 7318
rect 208394 7310 208406 7362
rect 208458 7310 208470 7362
rect 211262 7354 211314 7366
rect 213502 7418 213554 7430
rect 213502 7354 213554 7366
rect 214398 7418 214450 7430
rect 214398 7354 214450 7366
rect 214846 7418 214898 7430
rect 214846 7354 214898 7366
rect 204486 7242 204538 7254
rect 1344 7082 218624 7116
rect 1344 7030 28378 7082
rect 28430 7030 28482 7082
rect 28534 7030 28586 7082
rect 28638 7030 82706 7082
rect 82758 7030 82810 7082
rect 82862 7030 82914 7082
rect 82966 7030 137034 7082
rect 137086 7030 137138 7082
rect 137190 7030 137242 7082
rect 137294 7030 191362 7082
rect 191414 7030 191466 7082
rect 191518 7030 191570 7082
rect 191622 7030 218624 7082
rect 1344 6996 218624 7030
rect 58046 6858 58098 6870
rect 69358 6858 69410 6870
rect 187126 6858 187178 6870
rect 210702 6858 210754 6870
rect 10826 6806 10838 6858
rect 10890 6806 10902 6858
rect 16202 6806 16214 6858
rect 16266 6806 16278 6858
rect 32666 6806 32678 6858
rect 32730 6806 32742 6858
rect 41402 6806 41414 6858
rect 41466 6806 41478 6858
rect 48346 6806 48358 6858
rect 48410 6806 48422 6858
rect 63802 6806 63814 6858
rect 63866 6806 63878 6858
rect 72202 6806 72214 6858
rect 72266 6806 72278 6858
rect 105466 6806 105478 6858
rect 105530 6855 105542 6858
rect 105690 6855 105702 6858
rect 105530 6809 105702 6855
rect 105530 6806 105542 6809
rect 105690 6806 105702 6809
rect 105754 6806 105766 6858
rect 127978 6806 127990 6858
rect 128042 6806 128054 6858
rect 137834 6806 137846 6858
rect 137898 6806 137910 6858
rect 141754 6806 141766 6858
rect 141818 6806 141830 6858
rect 145786 6806 145798 6858
rect 145850 6806 145862 6858
rect 152170 6806 152182 6858
rect 152234 6806 152246 6858
rect 157322 6806 157334 6858
rect 157386 6806 157398 6858
rect 174122 6806 174134 6858
rect 174186 6806 174198 6858
rect 182634 6806 182646 6858
rect 182698 6806 182710 6858
rect 200554 6806 200566 6858
rect 200618 6806 200630 6858
rect 58046 6794 58098 6806
rect 69358 6794 69410 6806
rect 43934 6746 43986 6758
rect 12854 6690 12906 6702
rect 18230 6690 18282 6702
rect 34694 6690 34746 6702
rect 11498 6638 11510 6690
rect 11562 6638 11574 6690
rect 12854 6626 12906 6638
rect 13582 6634 13634 6646
rect 16650 6638 16662 6690
rect 16714 6638 16726 6690
rect 20682 6638 20694 6690
rect 20746 6638 20758 6690
rect 24378 6638 24390 6690
rect 24442 6638 24454 6690
rect 27738 6638 27750 6690
rect 27802 6638 27814 6690
rect 18230 6626 18282 6638
rect 28702 6634 28754 6646
rect 13582 6570 13634 6582
rect 8766 6522 8818 6534
rect 8766 6458 8818 6470
rect 14030 6522 14082 6534
rect 19338 6526 19350 6578
rect 19402 6526 19414 6578
rect 14030 6458 14082 6470
rect 21534 6522 21586 6534
rect 23034 6526 23046 6578
rect 23098 6526 23110 6578
rect 21534 6458 21586 6470
rect 25006 6522 25058 6534
rect 26394 6526 26406 6578
rect 26458 6526 26470 6578
rect 28702 6570 28754 6582
rect 30606 6634 30658 6646
rect 33450 6638 33462 6690
rect 33514 6638 33526 6690
rect 41850 6638 41862 6690
rect 41914 6638 41926 6690
rect 43934 6682 43986 6694
rect 47406 6746 47458 6758
rect 47406 6682 47458 6694
rect 49870 6746 49922 6758
rect 50990 6746 51042 6758
rect 34694 6626 34746 6638
rect 43306 6627 43318 6679
rect 43370 6627 43382 6679
rect 49018 6638 49030 6690
rect 49082 6638 49094 6690
rect 49870 6682 49922 6694
rect 50542 6690 50594 6702
rect 50990 6682 51042 6694
rect 51774 6746 51826 6758
rect 51774 6682 51826 6694
rect 54294 6746 54346 6758
rect 66558 6746 66610 6758
rect 54294 6682 54346 6694
rect 65830 6694 65882 6706
rect 55178 6638 55190 6690
rect 55242 6638 55254 6690
rect 50542 6626 50594 6638
rect 56746 6627 56758 6679
rect 56810 6627 56822 6679
rect 58606 6634 58658 6646
rect 30606 6570 30658 6582
rect 57486 6578 57538 6590
rect 25006 6458 25058 6470
rect 28366 6522 28418 6534
rect 28366 6458 28418 6470
rect 35086 6522 35138 6534
rect 35086 6458 35138 6470
rect 35534 6522 35586 6534
rect 35534 6458 35586 6470
rect 39006 6522 39058 6534
rect 39006 6458 39058 6470
rect 44382 6522 44434 6534
rect 48346 6526 48358 6578
rect 48410 6526 48422 6578
rect 44382 6458 44434 6470
rect 50430 6522 50482 6534
rect 50430 6458 50482 6470
rect 52110 6522 52162 6534
rect 52110 6458 52162 6470
rect 52558 6522 52610 6534
rect 52558 6458 52610 6470
rect 57374 6522 57426 6534
rect 57486 6514 57538 6526
rect 58158 6578 58210 6590
rect 58606 6570 58658 6582
rect 59390 6634 59442 6646
rect 64138 6638 64150 6690
rect 64202 6638 64214 6690
rect 66558 6682 66610 6694
rect 67902 6746 67954 6758
rect 67902 6682 67954 6694
rect 70030 6746 70082 6758
rect 76302 6746 76354 6758
rect 70030 6682 70082 6694
rect 70142 6690 70194 6702
rect 74230 6690 74282 6702
rect 65830 6630 65882 6642
rect 72538 6638 72550 6690
rect 72602 6638 72614 6690
rect 70142 6626 70194 6638
rect 74230 6626 74282 6638
rect 75070 6690 75122 6702
rect 75854 6690 75906 6702
rect 75070 6626 75122 6638
rect 75182 6634 75234 6646
rect 59390 6570 59442 6582
rect 68462 6578 68514 6590
rect 58158 6514 58210 6526
rect 59950 6522 60002 6534
rect 57374 6458 57426 6470
rect 59950 6458 60002 6470
rect 61742 6522 61794 6534
rect 61742 6458 61794 6470
rect 67006 6522 67058 6534
rect 67006 6458 67058 6470
rect 67454 6522 67506 6534
rect 67454 6458 67506 6470
rect 68350 6522 68402 6534
rect 68462 6514 68514 6526
rect 69470 6578 69522 6590
rect 78318 6746 78370 6758
rect 76302 6682 76354 6694
rect 77198 6690 77250 6702
rect 75854 6626 75906 6638
rect 81510 6746 81562 6758
rect 78318 6682 78370 6694
rect 78822 6690 78874 6702
rect 83470 6746 83522 6758
rect 77198 6626 77250 6638
rect 79818 6638 79830 6690
rect 79882 6638 79894 6690
rect 81510 6682 81562 6694
rect 82910 6690 82962 6702
rect 83470 6682 83522 6694
rect 84030 6746 84082 6758
rect 91758 6746 91810 6758
rect 98746 6750 98758 6802
rect 98810 6750 98822 6802
rect 84030 6682 84082 6694
rect 86662 6690 86714 6702
rect 90750 6690 90802 6702
rect 78822 6626 78874 6638
rect 82910 6626 82962 6638
rect 87658 6638 87670 6690
rect 87722 6638 87734 6690
rect 113262 6746 113314 6758
rect 91758 6682 91810 6694
rect 102118 6690 102170 6702
rect 86662 6626 86714 6638
rect 90750 6626 90802 6638
rect 90862 6634 90914 6646
rect 97402 6638 97414 6690
rect 97466 6638 97478 6690
rect 100314 6638 100326 6690
rect 100378 6638 100390 6690
rect 103114 6638 103126 6690
rect 103178 6638 103190 6690
rect 110506 6638 110518 6690
rect 110570 6638 110582 6690
rect 112746 6638 112758 6690
rect 112810 6638 112822 6690
rect 113262 6682 113314 6694
rect 115950 6746 116002 6758
rect 121034 6750 121046 6802
rect 121098 6750 121110 6802
rect 124842 6750 124854 6802
rect 124906 6750 124918 6802
rect 129322 6750 129334 6802
rect 129386 6750 129398 6802
rect 132794 6750 132806 6802
rect 132858 6750 132870 6802
rect 134810 6750 134822 6802
rect 134874 6750 134886 6802
rect 115950 6682 116002 6694
rect 138798 6746 138850 6758
rect 142762 6750 142774 6802
rect 142826 6750 142838 6802
rect 148698 6750 148710 6802
rect 148762 6750 148774 6802
rect 170202 6750 170214 6802
rect 170266 6750 170278 6802
rect 177146 6750 177158 6802
rect 177210 6750 177222 6802
rect 180462 6746 180514 6758
rect 185098 6750 185110 6802
rect 185162 6750 185174 6802
rect 187126 6794 187178 6806
rect 188458 6750 188470 6802
rect 188522 6750 188534 6802
rect 210702 6794 210754 6806
rect 75182 6570 75234 6582
rect 85150 6578 85202 6590
rect 69470 6514 69522 6526
rect 75742 6522 75794 6534
rect 68350 6458 68402 6470
rect 75742 6458 75794 6470
rect 77310 6522 77362 6534
rect 77310 6458 77362 6470
rect 77982 6522 78034 6534
rect 77982 6458 78034 6470
rect 83022 6522 83074 6534
rect 83022 6458 83074 6470
rect 84478 6522 84530 6534
rect 102118 6626 102170 6638
rect 118414 6634 118466 6646
rect 122602 6638 122614 6690
rect 122666 6638 122678 6690
rect 126410 6638 126422 6690
rect 126474 6638 126486 6690
rect 128538 6638 128550 6690
rect 128602 6638 128614 6690
rect 130890 6638 130902 6690
rect 130954 6638 130966 6690
rect 90862 6570 90914 6582
rect 85150 6514 85202 6526
rect 85262 6522 85314 6534
rect 84478 6458 84530 6470
rect 85262 6458 85314 6470
rect 85822 6522 85874 6534
rect 85822 6458 85874 6470
rect 86158 6522 86210 6534
rect 91422 6522 91474 6534
rect 97290 6526 97302 6578
rect 97354 6526 97366 6578
rect 89450 6470 89462 6522
rect 89514 6470 89526 6522
rect 86158 6458 86210 6470
rect 91422 6458 91474 6470
rect 97918 6522 97970 6534
rect 95946 6414 95958 6466
rect 96010 6414 96022 6466
rect 97918 6458 97970 6470
rect 98366 6522 98418 6534
rect 100202 6526 100214 6578
rect 100266 6526 100278 6578
rect 98366 6458 98418 6470
rect 101054 6522 101106 6534
rect 101054 6458 101106 6470
rect 101614 6522 101666 6534
rect 107662 6522 107714 6534
rect 110394 6526 110406 6578
rect 110458 6526 110470 6578
rect 112298 6526 112310 6578
rect 112362 6526 112374 6578
rect 118414 6570 118466 6582
rect 131406 6634 131458 6646
rect 134362 6638 134374 6690
rect 134426 6638 134438 6690
rect 135818 6638 135830 6690
rect 135882 6638 135894 6690
rect 136938 6638 136950 6690
rect 137002 6638 137014 6690
rect 137162 6638 137174 6690
rect 137226 6638 137238 6690
rect 138798 6682 138850 6694
rect 104906 6470 104918 6522
rect 104970 6470 104982 6522
rect 101614 6458 101666 6470
rect 107662 6458 107714 6470
rect 113710 6522 113762 6534
rect 109274 6414 109286 6466
rect 109338 6414 109350 6466
rect 111290 6414 111302 6466
rect 111354 6414 111366 6466
rect 113710 6458 113762 6470
rect 118750 6522 118802 6534
rect 122490 6526 122502 6578
rect 122554 6526 122566 6578
rect 118750 6458 118802 6470
rect 123118 6522 123170 6534
rect 123118 6458 123170 6470
rect 123566 6522 123618 6534
rect 126298 6526 126310 6578
rect 126362 6526 126374 6578
rect 128426 6526 128438 6578
rect 128490 6526 128502 6578
rect 130778 6526 130790 6578
rect 130842 6526 130854 6578
rect 131406 6570 131458 6582
rect 139694 6634 139746 6646
rect 142314 6638 142326 6690
rect 142378 6638 142390 6690
rect 144330 6638 144342 6690
rect 144394 6638 144406 6690
rect 146346 6638 146358 6690
rect 146410 6638 146422 6690
rect 150266 6638 150278 6690
rect 150330 6638 150342 6690
rect 123566 6458 123618 6470
rect 131854 6522 131906 6534
rect 133802 6526 133814 6578
rect 133866 6526 133878 6578
rect 135370 6526 135382 6578
rect 135434 6526 135446 6578
rect 139694 6570 139746 6582
rect 150782 6634 150834 6646
rect 151722 6638 151734 6690
rect 151786 6638 151798 6690
rect 153066 6638 153078 6690
rect 153130 6638 153142 6690
rect 131854 6458 131906 6470
rect 139246 6522 139298 6534
rect 140970 6526 140982 6578
rect 141034 6526 141046 6578
rect 142986 6526 142998 6578
rect 143050 6526 143062 6578
rect 145338 6526 145350 6578
rect 145402 6526 145414 6578
rect 139246 6458 139298 6470
rect 146750 6522 146802 6534
rect 146750 6458 146802 6470
rect 147198 6522 147250 6534
rect 147198 6458 147250 6470
rect 147646 6522 147698 6534
rect 149258 6526 149270 6578
rect 149322 6526 149334 6578
rect 150782 6570 150834 6582
rect 153694 6634 153746 6646
rect 155978 6638 155990 6690
rect 156042 6638 156054 6690
rect 156762 6638 156774 6690
rect 156826 6638 156838 6690
rect 158218 6638 158230 6690
rect 158282 6638 158294 6690
rect 159338 6638 159350 6690
rect 159402 6638 159414 6690
rect 161130 6638 161142 6690
rect 161194 6638 161206 6690
rect 153694 6570 153746 6582
rect 163326 6634 163378 6646
rect 167626 6638 167638 6690
rect 167690 6638 167702 6690
rect 169194 6657 169206 6709
rect 169258 6657 169270 6709
rect 176150 6690 176202 6702
rect 193118 6746 193170 6758
rect 171210 6638 171222 6690
rect 171274 6638 171286 6690
rect 174458 6638 174470 6690
rect 174522 6638 174534 6690
rect 177930 6638 177942 6690
rect 177994 6638 178006 6690
rect 180462 6682 180514 6694
rect 190654 6690 190706 6702
rect 176150 6626 176202 6638
rect 178838 6634 178890 6646
rect 147646 6458 147698 6470
rect 151118 6522 151170 6534
rect 155418 6526 155430 6578
rect 155482 6526 155494 6578
rect 159002 6526 159014 6578
rect 159066 6526 159078 6578
rect 162474 6526 162486 6578
rect 162538 6526 162550 6578
rect 163326 6570 163378 6582
rect 178838 6570 178890 6582
rect 179678 6634 179730 6646
rect 182970 6638 182982 6690
rect 183034 6638 183046 6690
rect 184482 6638 184494 6690
rect 184546 6638 184558 6690
rect 185658 6638 185670 6690
rect 185722 6638 185734 6690
rect 189466 6638 189478 6690
rect 189530 6638 189542 6690
rect 193118 6682 193170 6694
rect 195694 6746 195746 6758
rect 195694 6682 195746 6694
rect 196814 6746 196866 6758
rect 205270 6746 205322 6758
rect 196814 6682 196866 6694
rect 202582 6690 202634 6702
rect 190654 6626 190706 6638
rect 191774 6634 191826 6646
rect 179678 6570 179730 6582
rect 191326 6578 191378 6590
rect 151118 6458 151170 6470
rect 163662 6522 163714 6534
rect 154522 6414 154534 6466
rect 154586 6414 154598 6466
rect 163662 6458 163714 6470
rect 164558 6522 164610 6534
rect 164558 6458 164610 6470
rect 165006 6522 165058 6534
rect 165006 6458 165058 6470
rect 166854 6522 166906 6534
rect 166854 6458 166906 6470
rect 179174 6522 179226 6534
rect 186330 6526 186342 6578
rect 186394 6526 186406 6578
rect 179174 6458 179226 6470
rect 187462 6522 187514 6534
rect 188682 6526 188694 6578
rect 188746 6526 188758 6578
rect 187462 6458 187514 6470
rect 190542 6522 190594 6534
rect 190542 6458 190594 6470
rect 191214 6522 191266 6534
rect 196366 6634 196418 6646
rect 191774 6570 191826 6582
rect 194350 6578 194402 6590
rect 191326 6514 191378 6526
rect 192222 6522 192274 6534
rect 191214 6458 191266 6470
rect 192222 6458 192274 6470
rect 192670 6522 192722 6534
rect 192670 6458 192722 6470
rect 193566 6522 193618 6534
rect 193566 6458 193618 6470
rect 194238 6522 194290 6534
rect 196366 6570 196418 6582
rect 197262 6634 197314 6646
rect 200890 6638 200902 6690
rect 200954 6638 200966 6690
rect 205270 6682 205322 6694
rect 207958 6690 208010 6702
rect 202582 6626 202634 6638
rect 203086 6634 203138 6646
rect 206490 6638 206502 6690
rect 206554 6638 206566 6690
rect 209850 6638 209862 6690
rect 209914 6638 209926 6690
rect 197262 6570 197314 6582
rect 207958 6626 208010 6638
rect 214510 6634 214562 6646
rect 203086 6570 203138 6582
rect 203198 6578 203250 6590
rect 210814 6578 210866 6590
rect 194350 6514 194402 6526
rect 194798 6522 194850 6534
rect 194238 6458 194290 6470
rect 194798 6458 194850 6470
rect 195246 6522 195298 6534
rect 195246 6458 195298 6470
rect 197710 6522 197762 6534
rect 197710 6458 197762 6470
rect 198158 6522 198210 6534
rect 203198 6514 203250 6526
rect 203646 6522 203698 6534
rect 209738 6526 209750 6578
rect 209802 6526 209814 6578
rect 198158 6458 198210 6470
rect 210814 6514 210866 6526
rect 211374 6578 211426 6590
rect 214510 6570 214562 6582
rect 211374 6514 211426 6526
rect 211486 6522 211538 6534
rect 203646 6458 203698 6470
rect 211486 6458 211538 6470
rect 212270 6522 212322 6534
rect 212270 6458 212322 6470
rect 212718 6522 212770 6534
rect 212718 6458 212770 6470
rect 213166 6522 213218 6534
rect 213166 6458 213218 6470
rect 213614 6522 213666 6534
rect 213614 6458 213666 6470
rect 214062 6522 214114 6534
rect 214062 6458 214114 6470
rect 214958 6522 215010 6534
rect 214958 6458 215010 6470
rect 215406 6522 215458 6534
rect 215406 6458 215458 6470
rect 1344 6298 218624 6332
rect 1344 6246 55542 6298
rect 55594 6246 55646 6298
rect 55698 6246 55750 6298
rect 55802 6246 109870 6298
rect 109922 6246 109974 6298
rect 110026 6246 110078 6298
rect 110130 6246 164198 6298
rect 164250 6246 164302 6298
rect 164354 6246 164406 6298
rect 164458 6246 218624 6298
rect 1344 6212 218624 6246
rect 9550 6074 9602 6086
rect 9550 6010 9602 6022
rect 10670 6074 10722 6086
rect 10670 6010 10722 6022
rect 14422 6074 14474 6086
rect 14422 6010 14474 6022
rect 47070 6074 47122 6086
rect 47070 6010 47122 6022
rect 48638 6074 48690 6086
rect 48638 6010 48690 6022
rect 56590 6074 56642 6086
rect 56590 6010 56642 6022
rect 57374 6074 57426 6086
rect 57374 6010 57426 6022
rect 57710 6074 57762 6086
rect 57710 6010 57762 6022
rect 58382 6074 58434 6086
rect 58382 6010 58434 6022
rect 66894 6074 66946 6086
rect 66894 6010 66946 6022
rect 67902 6074 67954 6086
rect 67902 6010 67954 6022
rect 68350 6074 68402 6086
rect 68350 6010 68402 6022
rect 68798 6074 68850 6086
rect 70590 6074 70642 6086
rect 68798 6010 68850 6022
rect 70030 6018 70082 6030
rect 69918 5962 69970 5974
rect 12742 5906 12794 5918
rect 8810 5854 8822 5906
rect 8874 5854 8886 5906
rect 15866 5854 15878 5906
rect 15930 5854 15942 5906
rect 16886 5902 16938 5914
rect 12742 5842 12794 5854
rect 16886 5838 16938 5850
rect 17502 5850 17554 5862
rect 8138 5742 8150 5794
rect 8202 5742 8214 5794
rect 11946 5742 11958 5794
rect 12010 5742 12022 5794
rect 17502 5786 17554 5798
rect 18062 5850 18114 5862
rect 20010 5854 20022 5906
rect 20074 5854 20086 5906
rect 22250 5854 22262 5906
rect 22314 5854 22326 5906
rect 24714 5854 24726 5906
rect 24778 5854 24790 5906
rect 18062 5786 18114 5798
rect 25454 5850 25506 5862
rect 28186 5854 28198 5906
rect 28250 5854 28262 5906
rect 30426 5854 30438 5906
rect 30490 5854 30502 5906
rect 32666 5854 32678 5906
rect 32730 5854 32742 5906
rect 18890 5742 18902 5794
rect 18954 5742 18966 5794
rect 21130 5742 21142 5794
rect 21194 5742 21206 5794
rect 23370 5742 23382 5794
rect 23434 5742 23446 5794
rect 25454 5786 25506 5798
rect 33406 5850 33458 5862
rect 26842 5742 26854 5794
rect 26906 5742 26918 5794
rect 29082 5742 29094 5794
rect 29146 5742 29158 5794
rect 31434 5742 31446 5794
rect 31498 5742 31510 5794
rect 33406 5786 33458 5798
rect 33854 5850 33906 5862
rect 37034 5854 37046 5906
rect 37098 5854 37110 5906
rect 33854 5786 33906 5798
rect 37550 5850 37602 5862
rect 35802 5742 35814 5794
rect 35866 5742 35878 5794
rect 37550 5786 37602 5798
rect 42366 5850 42418 5862
rect 42366 5786 42418 5798
rect 43262 5850 43314 5862
rect 43262 5786 43314 5798
rect 43822 5850 43874 5862
rect 43822 5786 43874 5798
rect 44270 5850 44322 5862
rect 46554 5854 46566 5906
rect 46618 5854 46630 5906
rect 44270 5786 44322 5798
rect 48190 5850 48242 5862
rect 51034 5854 51046 5906
rect 51098 5854 51110 5906
rect 45210 5742 45222 5794
rect 45274 5742 45286 5794
rect 48190 5786 48242 5798
rect 51550 5850 51602 5862
rect 49802 5742 49814 5794
rect 49866 5742 49878 5794
rect 51550 5786 51602 5798
rect 52222 5850 52274 5862
rect 54506 5854 54518 5906
rect 54570 5854 54582 5906
rect 56198 5902 56250 5914
rect 69358 5906 69410 5918
rect 56198 5838 56250 5850
rect 58830 5850 58882 5862
rect 52222 5786 52274 5798
rect 58830 5786 58882 5798
rect 67454 5850 67506 5862
rect 71934 6074 71986 6086
rect 70590 6010 70642 6022
rect 71374 6018 71426 6030
rect 70030 5954 70082 5966
rect 71934 6010 71986 6022
rect 74286 6074 74338 6086
rect 77534 6074 77586 6086
rect 74286 6010 74338 6022
rect 74398 6018 74450 6030
rect 71374 5954 71426 5966
rect 75562 5966 75574 6018
rect 75626 5966 75638 6018
rect 77534 6010 77586 6022
rect 78094 6074 78146 6086
rect 78094 6010 78146 6022
rect 111470 6074 111522 6086
rect 81498 5966 81510 6018
rect 81562 5966 81574 6018
rect 83962 5966 83974 6018
rect 84026 5966 84038 6018
rect 99306 5966 99318 6018
rect 99370 5966 99382 6018
rect 111470 6010 111522 6022
rect 122446 6074 122498 6086
rect 117898 5966 117910 6018
rect 117962 5966 117974 6018
rect 122446 6010 122498 6022
rect 126702 6074 126754 6086
rect 126702 6010 126754 6022
rect 127038 6074 127090 6086
rect 127038 6010 127090 6022
rect 128270 6074 128322 6086
rect 128270 6010 128322 6022
rect 131070 6074 131122 6086
rect 74398 5954 74450 5966
rect 119758 5962 119810 5974
rect 129210 5966 129222 6018
rect 129274 5966 129286 6018
rect 131070 6010 131122 6022
rect 135102 6074 135154 6086
rect 135102 6010 135154 6022
rect 135998 6074 136050 6086
rect 135998 6010 136050 6022
rect 143726 6074 143778 6086
rect 145226 6078 145238 6130
rect 145290 6078 145302 6130
rect 69918 5898 69970 5910
rect 70702 5906 70754 5918
rect 69358 5842 69410 5854
rect 70702 5842 70754 5854
rect 72046 5906 72098 5918
rect 73390 5906 73442 5918
rect 72046 5842 72098 5854
rect 72606 5850 72658 5862
rect 67454 5786 67506 5798
rect 76906 5854 76918 5906
rect 76970 5854 76982 5906
rect 73390 5842 73442 5854
rect 78542 5850 78594 5862
rect 72606 5786 72658 5798
rect 78542 5786 78594 5798
rect 79774 5850 79826 5862
rect 82730 5854 82742 5906
rect 82794 5854 82806 5906
rect 85306 5854 85318 5906
rect 85370 5854 85382 5906
rect 79774 5786 79826 5798
rect 85822 5850 85874 5862
rect 85822 5786 85874 5798
rect 87950 5850 88002 5862
rect 100650 5854 100662 5906
rect 100714 5854 100726 5906
rect 87950 5786 88002 5798
rect 101278 5850 101330 5862
rect 101278 5786 101330 5798
rect 101726 5850 101778 5862
rect 101726 5786 101778 5798
rect 110910 5850 110962 5862
rect 119242 5854 119254 5906
rect 119306 5854 119318 5906
rect 119758 5898 119810 5910
rect 135550 5962 135602 5974
rect 137610 5966 137622 6018
rect 137674 5966 137686 6018
rect 143726 6010 143778 6022
rect 148766 6074 148818 6086
rect 152842 6078 152854 6130
rect 152906 6078 152918 6130
rect 130554 5854 130566 5906
rect 130618 5854 130630 5906
rect 110910 5786 110962 5798
rect 131630 5850 131682 5862
rect 131630 5786 131682 5798
rect 132078 5850 132130 5862
rect 132078 5786 132130 5798
rect 132526 5850 132578 5862
rect 134250 5854 134262 5906
rect 134314 5854 134326 5906
rect 135550 5898 135602 5910
rect 143390 5962 143442 5974
rect 146010 5966 146022 6018
rect 146074 5966 146086 6018
rect 148766 6010 148818 6022
rect 154702 6074 154754 6086
rect 149930 5966 149942 6018
rect 149994 5966 150006 6018
rect 154702 6010 154754 6022
rect 155262 6074 155314 6086
rect 155262 6010 155314 6022
rect 160638 6074 160690 6086
rect 167526 6074 167578 6086
rect 162250 6022 162262 6074
rect 162314 6022 162326 6074
rect 159450 5966 159462 6018
rect 159514 5966 159526 6018
rect 160638 6010 160690 6022
rect 167526 6010 167578 6022
rect 175142 6074 175194 6086
rect 175142 6010 175194 6022
rect 175478 6074 175530 6086
rect 182870 6074 182922 6086
rect 177482 6022 177494 6074
rect 177546 6022 177558 6074
rect 175478 6010 175530 6022
rect 182870 6010 182922 6022
rect 190878 6074 190930 6086
rect 192446 6074 192498 6086
rect 187338 5966 187350 6018
rect 187402 5966 187414 6018
rect 189242 5966 189254 6018
rect 189306 5966 189318 6018
rect 190878 6010 190930 6022
rect 190990 6018 191042 6030
rect 192446 6010 192498 6022
rect 192894 6074 192946 6086
rect 192894 6010 192946 6022
rect 193342 6074 193394 6086
rect 193342 6010 193394 6022
rect 193790 6074 193842 6086
rect 193790 6010 193842 6022
rect 195134 6074 195186 6086
rect 195134 6010 195186 6022
rect 199390 6074 199442 6086
rect 199390 6010 199442 6022
rect 200510 6074 200562 6086
rect 207566 6074 207618 6086
rect 202346 6022 202358 6074
rect 202410 6022 202422 6074
rect 200510 6010 200562 6022
rect 207566 6010 207618 6022
rect 212382 6074 212434 6086
rect 212382 6010 212434 6022
rect 213278 6074 213330 6086
rect 213278 6010 213330 6022
rect 138730 5854 138742 5906
rect 138794 5854 138806 5906
rect 139402 5854 139414 5906
rect 139466 5854 139478 5906
rect 140858 5854 140870 5906
rect 140922 5854 140934 5906
rect 141418 5854 141430 5906
rect 141482 5854 141494 5906
rect 142650 5854 142662 5906
rect 142714 5854 142726 5906
rect 143390 5898 143442 5910
rect 164838 5906 164890 5918
rect 167850 5910 167862 5962
rect 167914 5910 167926 5962
rect 145674 5854 145686 5906
rect 145738 5854 145750 5906
rect 146906 5854 146918 5906
rect 146970 5854 146982 5906
rect 147466 5854 147478 5906
rect 147530 5854 147542 5906
rect 132526 5786 132578 5798
rect 149214 5850 149266 5862
rect 150938 5854 150950 5906
rect 151002 5854 151014 5906
rect 69246 5738 69298 5750
rect 54170 5686 54182 5738
rect 54234 5686 54246 5738
rect 69246 5674 69298 5686
rect 71262 5738 71314 5750
rect 71262 5674 71314 5686
rect 73278 5738 73330 5750
rect 133130 5742 133142 5794
rect 133194 5742 133206 5794
rect 140074 5742 140086 5794
rect 140138 5742 140150 5794
rect 141306 5742 141318 5794
rect 141370 5742 141382 5794
rect 149214 5786 149266 5798
rect 151790 5850 151842 5862
rect 152842 5854 152854 5906
rect 152906 5854 152918 5906
rect 154298 5854 154310 5906
rect 154362 5854 154374 5906
rect 156090 5854 156102 5906
rect 156154 5854 156166 5906
rect 157546 5854 157558 5906
rect 157610 5854 157622 5906
rect 158106 5854 158118 5906
rect 158170 5854 158182 5906
rect 163818 5854 163830 5906
rect 163882 5854 163894 5906
rect 165386 5854 165398 5906
rect 165450 5854 165462 5906
rect 168746 5854 168758 5906
rect 168810 5854 168822 5906
rect 173002 5854 173014 5906
rect 173066 5854 173078 5906
rect 174570 5865 174582 5917
rect 174634 5865 174646 5917
rect 180182 5906 180234 5918
rect 183194 5910 183206 5962
rect 183258 5910 183270 5962
rect 190990 5954 191042 5966
rect 214174 5962 214226 5974
rect 178602 5854 178614 5906
rect 178666 5854 178678 5906
rect 181178 5854 181190 5906
rect 181242 5854 181254 5906
rect 164838 5842 164890 5854
rect 180182 5842 180234 5854
rect 183710 5850 183762 5862
rect 184650 5854 184662 5906
rect 184714 5854 184726 5906
rect 188010 5854 188022 5906
rect 188074 5854 188086 5906
rect 189578 5854 189590 5906
rect 189642 5854 189654 5906
rect 149706 5742 149718 5794
rect 149770 5742 149782 5794
rect 151790 5786 151842 5798
rect 166282 5742 166294 5794
rect 166346 5742 166358 5794
rect 169642 5742 169654 5794
rect 169706 5742 169718 5794
rect 181402 5742 181414 5794
rect 181466 5742 181478 5794
rect 183710 5786 183762 5798
rect 191438 5850 191490 5862
rect 184762 5742 184774 5794
rect 184826 5742 184838 5794
rect 186778 5742 186790 5794
rect 186842 5742 186854 5794
rect 191438 5786 191490 5798
rect 194238 5850 194290 5862
rect 194238 5786 194290 5798
rect 194686 5850 194738 5862
rect 194686 5786 194738 5798
rect 195582 5850 195634 5862
rect 197754 5854 197766 5906
rect 197818 5854 197830 5906
rect 195582 5786 195634 5798
rect 198494 5850 198546 5862
rect 196522 5742 196534 5794
rect 196586 5742 196598 5794
rect 198494 5786 198546 5798
rect 198942 5850 198994 5862
rect 198942 5786 198994 5798
rect 200846 5850 200898 5862
rect 203914 5854 203926 5906
rect 203978 5854 203990 5906
rect 204754 5854 204766 5906
rect 204818 5854 204830 5906
rect 205482 5854 205494 5906
rect 205546 5854 205558 5906
rect 210970 5854 210982 5906
rect 211034 5854 211046 5906
rect 211810 5854 211822 5906
rect 211874 5854 211886 5906
rect 214174 5898 214226 5910
rect 200846 5786 200898 5798
rect 212830 5850 212882 5862
rect 205818 5742 205830 5794
rect 205882 5742 205894 5794
rect 212830 5786 212882 5798
rect 213726 5850 213778 5862
rect 213726 5786 213778 5798
rect 214622 5850 214674 5862
rect 214622 5786 214674 5798
rect 215070 5850 215122 5862
rect 215070 5786 215122 5798
rect 208742 5738 208794 5750
rect 147802 5686 147814 5738
rect 147866 5686 147878 5738
rect 156986 5686 156998 5738
rect 157050 5686 157062 5738
rect 172666 5686 172678 5738
rect 172730 5686 172742 5738
rect 189802 5686 189814 5738
rect 189866 5686 189878 5738
rect 73278 5674 73330 5686
rect 208742 5674 208794 5686
rect 1344 5514 218624 5548
rect 1344 5462 28378 5514
rect 28430 5462 28482 5514
rect 28534 5462 28586 5514
rect 28638 5462 82706 5514
rect 82758 5462 82810 5514
rect 82862 5462 82914 5514
rect 82966 5462 137034 5514
rect 137086 5462 137138 5514
rect 137190 5462 137242 5514
rect 137294 5462 191362 5514
rect 191414 5462 191466 5514
rect 191518 5462 191570 5514
rect 191622 5462 218624 5514
rect 1344 5428 218624 5462
rect 204766 5290 204818 5302
rect 186890 5238 186902 5290
rect 186954 5238 186966 5290
rect 72538 5182 72550 5234
rect 72602 5182 72614 5234
rect 74622 5178 74674 5190
rect 8698 5070 8710 5122
rect 8762 5070 8774 5122
rect 11610 5070 11622 5122
rect 11674 5070 11686 5122
rect 15754 5070 15766 5122
rect 15818 5070 15830 5122
rect 20458 5070 20470 5122
rect 20522 5070 20534 5122
rect 24378 5070 24390 5122
rect 24442 5070 24454 5122
rect 28298 5070 28310 5122
rect 28362 5070 28374 5122
rect 31770 5070 31782 5122
rect 31834 5070 31846 5122
rect 35018 5070 35030 5122
rect 35082 5070 35094 5122
rect 38490 5070 38502 5122
rect 38554 5070 38566 5122
rect 43082 5070 43094 5122
rect 43146 5070 43158 5122
rect 46890 5070 46902 5122
rect 46954 5070 46966 5122
rect 51818 5070 51830 5122
rect 51882 5070 51894 5122
rect 55738 5070 55750 5122
rect 55802 5070 55814 5122
rect 58650 5070 58662 5122
rect 58714 5070 58726 5122
rect 63466 5070 63478 5122
rect 63530 5070 63542 5122
rect 66826 5070 66838 5122
rect 66890 5070 66902 5122
rect 70410 5070 70422 5122
rect 70474 5070 70486 5122
rect 73882 5070 73894 5122
rect 73946 5070 73958 5122
rect 74622 5114 74674 5126
rect 75182 5178 75234 5190
rect 91198 5178 91250 5190
rect 81386 5126 81398 5178
rect 81450 5175 81462 5178
rect 81450 5129 81559 5175
rect 81450 5126 81462 5129
rect 75182 5114 75234 5126
rect 79258 5070 79270 5122
rect 79322 5070 79334 5122
rect 8250 4958 8262 5010
rect 8314 4958 8326 5010
rect 9550 4954 9602 4966
rect 9550 4890 9602 4902
rect 10558 4954 10610 4966
rect 11162 4958 11174 5010
rect 11226 4958 11238 5010
rect 10558 4890 10610 4902
rect 13358 4954 13410 4966
rect 14410 4958 14422 5010
rect 14474 4958 14486 5010
rect 13358 4890 13410 4902
rect 16382 4954 16434 4966
rect 19898 4958 19910 5010
rect 19962 4958 19974 5010
rect 16382 4890 16434 4902
rect 21310 4954 21362 4966
rect 21310 4890 21362 4902
rect 21758 4954 21810 4966
rect 21758 4890 21810 4902
rect 22318 4954 22370 4966
rect 23034 4958 23046 5010
rect 23098 4958 23110 5010
rect 22318 4890 22370 4902
rect 25230 4954 25282 4966
rect 26954 4958 26966 5010
rect 27018 4958 27030 5010
rect 25230 4890 25282 4902
rect 29150 4954 29202 4966
rect 30874 4958 30886 5010
rect 30938 4958 30950 5010
rect 33898 4958 33910 5010
rect 33962 4958 33974 5010
rect 29150 4890 29202 4902
rect 35646 4954 35698 4966
rect 37258 4958 37270 5010
rect 37322 4958 37334 5010
rect 35646 4890 35698 4902
rect 39230 4954 39282 4966
rect 41738 4958 41750 5010
rect 41802 4958 41814 5010
rect 39230 4890 39282 4902
rect 43710 4954 43762 4966
rect 46554 4958 46566 5010
rect 46618 4958 46630 5010
rect 43710 4890 43762 4902
rect 48750 4954 48802 4966
rect 48750 4890 48802 4902
rect 49646 4954 49698 4966
rect 50474 4958 50486 5010
rect 50538 4958 50550 5010
rect 49646 4890 49698 4902
rect 52670 4954 52722 4966
rect 54730 4958 54742 5010
rect 54794 4958 54806 5010
rect 52670 4890 52722 4902
rect 56590 4954 56642 4966
rect 56590 4890 56642 4902
rect 57374 4954 57426 4966
rect 58314 4958 58326 5010
rect 58378 4958 58390 5010
rect 57374 4890 57426 4902
rect 60510 4954 60562 4966
rect 62234 4958 62246 5010
rect 62298 4958 62310 5010
rect 60510 4890 60562 4902
rect 64430 4954 64482 4966
rect 66042 4958 66054 5010
rect 66106 4958 66118 5010
rect 64430 4890 64482 4902
rect 68574 4954 68626 4966
rect 69178 4958 69190 5010
rect 69242 4958 69254 5010
rect 68574 4890 68626 4902
rect 71598 4954 71650 4966
rect 79034 4958 79046 5010
rect 79098 4958 79110 5010
rect 81513 5007 81559 5129
rect 83178 5070 83190 5122
rect 83242 5070 83254 5122
rect 87098 5070 87110 5122
rect 87162 5070 87174 5122
rect 90570 5070 90582 5122
rect 90634 5070 90646 5122
rect 91198 5114 91250 5126
rect 94782 5178 94834 5190
rect 93930 5070 93942 5122
rect 93994 5070 94006 5122
rect 94782 5114 94834 5126
rect 98030 5178 98082 5190
rect 102442 5182 102454 5234
rect 102506 5182 102518 5234
rect 97402 5070 97414 5122
rect 97466 5070 97478 5122
rect 98030 5114 98082 5126
rect 103630 5178 103682 5190
rect 105354 5182 105366 5234
rect 105418 5182 105430 5234
rect 102778 5070 102790 5122
rect 102842 5070 102854 5122
rect 103630 5114 103682 5126
rect 114158 5178 114210 5190
rect 106698 5070 106710 5122
rect 106762 5070 106774 5122
rect 110282 5070 110294 5122
rect 110346 5070 110358 5122
rect 113418 5070 113430 5122
rect 113482 5070 113494 5122
rect 114158 5114 114210 5126
rect 117630 5178 117682 5190
rect 120810 5182 120822 5234
rect 120874 5182 120886 5234
rect 117002 5070 117014 5122
rect 117066 5070 117078 5122
rect 117630 5114 117682 5126
rect 133870 5178 133922 5190
rect 122154 5070 122166 5122
rect 122218 5070 122230 5122
rect 123946 5070 123958 5122
rect 124010 5070 124022 5122
rect 128762 5070 128774 5122
rect 128826 5070 128838 5122
rect 132570 5070 132582 5122
rect 132634 5070 132646 5122
rect 133870 5114 133922 5126
rect 134318 5178 134370 5190
rect 134318 5114 134370 5126
rect 137566 5178 137618 5190
rect 139290 5182 139302 5234
rect 139354 5182 139366 5234
rect 144554 5182 144566 5234
rect 144618 5182 144630 5234
rect 136602 5070 136614 5122
rect 136666 5070 136678 5122
rect 137566 5114 137618 5126
rect 146750 5178 146802 5190
rect 151274 5182 151286 5234
rect 151338 5182 151350 5234
rect 162698 5182 162710 5234
rect 162762 5182 162774 5234
rect 204766 5226 204818 5238
rect 177214 5178 177266 5190
rect 140634 5070 140646 5122
rect 140698 5070 140710 5122
rect 145898 5070 145910 5122
rect 145962 5070 145974 5122
rect 146750 5114 146802 5126
rect 171894 5122 171946 5134
rect 148542 5066 148594 5078
rect 152618 5070 152630 5122
rect 152682 5070 152694 5122
rect 156090 5070 156102 5122
rect 156154 5070 156166 5122
rect 158554 5070 158566 5122
rect 158618 5070 158630 5122
rect 164042 5070 164054 5122
rect 164106 5070 164118 5122
rect 166394 5070 166406 5122
rect 166458 5070 166470 5122
rect 174234 5070 174246 5122
rect 174298 5070 174310 5122
rect 177214 5114 177266 5126
rect 211094 5122 211146 5134
rect 178154 5070 178166 5122
rect 178218 5070 178230 5122
rect 182634 5070 182646 5122
rect 182698 5070 182710 5122
rect 186218 5070 186230 5122
rect 186282 5070 186294 5122
rect 171894 5058 171946 5070
rect 188974 5066 189026 5078
rect 197978 5070 197990 5122
rect 198042 5070 198054 5122
rect 201674 5070 201686 5122
rect 201738 5070 201750 5122
rect 81610 5007 81622 5010
rect 71598 4890 71650 4902
rect 80110 4954 80162 4966
rect 81513 4961 81622 5007
rect 81610 4958 81622 4961
rect 81674 4958 81686 5010
rect 81834 4958 81846 5010
rect 81898 4958 81910 5010
rect 80110 4890 80162 4902
rect 83918 4954 83970 4966
rect 83918 4890 83970 4902
rect 84478 4954 84530 4966
rect 84478 4890 84530 4902
rect 84926 4954 84978 4966
rect 85754 4958 85766 5010
rect 85818 4958 85830 5010
rect 84926 4890 84978 4902
rect 87950 4954 88002 4966
rect 89226 4958 89238 5010
rect 89290 4958 89302 5010
rect 92810 4958 92822 5010
rect 92874 4958 92886 5010
rect 96058 4958 96070 5010
rect 96122 4958 96134 5010
rect 87950 4890 88002 4902
rect 107550 4954 107602 4966
rect 108938 4958 108950 5010
rect 109002 4958 109014 5010
rect 107550 4890 107602 4902
rect 111470 4954 111522 4966
rect 112186 4958 112198 5010
rect 112250 4958 112262 5010
rect 115658 4958 115670 5010
rect 115722 4958 115734 5010
rect 123498 4958 123510 5010
rect 123562 4958 123574 5010
rect 111470 4890 111522 4902
rect 125470 4954 125522 4966
rect 127418 4958 127430 5010
rect 127482 4958 127494 5010
rect 125470 4890 125522 4902
rect 129390 4954 129442 4966
rect 131450 4958 131462 5010
rect 131514 4958 131526 5010
rect 129390 4890 129442 4902
rect 133422 4954 133474 4966
rect 135258 4958 135270 5010
rect 135322 4958 135334 5010
rect 148542 5002 148594 5014
rect 133422 4890 133474 4902
rect 137118 4954 137170 4966
rect 137118 4890 137170 4902
rect 138126 4954 138178 4966
rect 138126 4890 138178 4902
rect 141150 4954 141202 4966
rect 141150 4890 141202 4902
rect 141598 4954 141650 4966
rect 141598 4890 141650 4902
rect 142158 4954 142210 4966
rect 142158 4890 142210 4902
rect 142830 4954 142882 4966
rect 142830 4890 142882 4902
rect 143278 4954 143330 4966
rect 143278 4890 143330 4902
rect 143614 4954 143666 4966
rect 143614 4890 143666 4902
rect 147086 4954 147138 4966
rect 147086 4890 147138 4902
rect 147646 4954 147698 4966
rect 147646 4890 147698 4902
rect 148094 4954 148146 4966
rect 148094 4890 148146 4902
rect 148878 4954 148930 4966
rect 148878 4890 148930 4902
rect 149438 4954 149490 4966
rect 149438 4890 149490 4902
rect 149774 4954 149826 4966
rect 149774 4890 149826 4902
rect 153134 4954 153186 4966
rect 153134 4890 153186 4902
rect 153582 4954 153634 4966
rect 153582 4890 153634 4902
rect 154478 4954 154530 4966
rect 154478 4890 154530 4902
rect 154926 4954 154978 4966
rect 154926 4890 154978 4902
rect 155374 4954 155426 4966
rect 156202 4958 156214 5010
rect 156266 4958 156278 5010
rect 158666 4958 158678 5010
rect 158730 4958 158742 5010
rect 155374 4890 155426 4902
rect 160750 4954 160802 4966
rect 160750 4890 160802 4902
rect 161086 4954 161138 4966
rect 161086 4890 161138 4902
rect 161534 4954 161586 4966
rect 161534 4890 161586 4902
rect 164558 4954 164610 4966
rect 164558 4890 164610 4902
rect 165118 4954 165170 4966
rect 165118 4890 165170 4902
rect 165454 4954 165506 4966
rect 166506 4958 166518 5010
rect 166570 4958 166582 5010
rect 165454 4890 165506 4902
rect 168646 4954 168698 4966
rect 168646 4890 168698 4902
rect 168982 4954 169034 4966
rect 168982 4890 169034 4902
rect 169486 4954 169538 4966
rect 170426 4958 170438 5010
rect 170490 4958 170502 5010
rect 169486 4890 169538 4902
rect 172678 4954 172730 4966
rect 172678 4890 172730 4902
rect 173014 4954 173066 4966
rect 174346 4958 174358 5010
rect 174410 4958 174422 5010
rect 173014 4890 173066 4902
rect 176374 4954 176426 4966
rect 176374 4890 176426 4902
rect 176710 4954 176762 4966
rect 178266 4958 178278 5010
rect 178330 4958 178342 5010
rect 176710 4890 176762 4902
rect 180294 4954 180346 4966
rect 180294 4890 180346 4902
rect 180630 4954 180682 4966
rect 180630 4890 180682 4902
rect 181134 4954 181186 4966
rect 182186 4958 182198 5010
rect 182250 4958 182262 5010
rect 181134 4890 181186 4902
rect 184214 4954 184266 4966
rect 184214 4890 184266 4902
rect 184550 4954 184602 4966
rect 184550 4890 184602 4902
rect 185166 4954 185218 4966
rect 186106 4958 186118 5010
rect 186170 4958 186182 5010
rect 188974 5002 189026 5014
rect 204654 5066 204706 5078
rect 205594 5070 205606 5122
rect 205658 5070 205670 5122
rect 185166 4890 185218 4902
rect 188022 4954 188074 4966
rect 188022 4890 188074 4902
rect 188358 4954 188410 4966
rect 188358 4890 188410 4902
rect 188862 4954 188914 4966
rect 188862 4890 188914 4902
rect 189758 4954 189810 4966
rect 189758 4890 189810 4902
rect 190206 4954 190258 4966
rect 190206 4890 190258 4902
rect 190654 4954 190706 4966
rect 190654 4890 190706 4902
rect 191102 4954 191154 4966
rect 191102 4890 191154 4902
rect 191550 4954 191602 4966
rect 191550 4890 191602 4902
rect 191998 4954 192050 4966
rect 191998 4890 192050 4902
rect 192446 4954 192498 4966
rect 192446 4890 192498 4902
rect 192894 4954 192946 4966
rect 192894 4890 192946 4902
rect 193678 4954 193730 4966
rect 193678 4890 193730 4902
rect 194126 4954 194178 4966
rect 194126 4890 194178 4902
rect 194574 4954 194626 4966
rect 194574 4890 194626 4902
rect 195022 4954 195074 4966
rect 195022 4890 195074 4902
rect 195470 4954 195522 4966
rect 195470 4890 195522 4902
rect 195918 4954 195970 4966
rect 195918 4890 195970 4902
rect 196366 4954 196418 4966
rect 196366 4890 196418 4902
rect 196814 4954 196866 4966
rect 197866 4958 197878 5010
rect 197930 4958 197942 5010
rect 196814 4890 196866 4902
rect 199838 4954 199890 4966
rect 199838 4890 199890 4902
rect 200286 4954 200338 4966
rect 200286 4890 200338 4902
rect 200734 4954 200786 4966
rect 201786 4958 201798 5010
rect 201850 4958 201862 5010
rect 204654 5002 204706 5014
rect 207790 5066 207842 5078
rect 200734 4890 200786 4902
rect 203758 4954 203810 4966
rect 205706 4958 205718 5010
rect 205770 4958 205782 5010
rect 207790 5002 207842 5014
rect 208574 5066 208626 5078
rect 211094 5058 211146 5070
rect 208574 5002 208626 5014
rect 203758 4890 203810 4902
rect 207902 4954 207954 4966
rect 207902 4890 207954 4902
rect 208462 4954 208514 4966
rect 209626 4958 209638 5010
rect 209690 4958 209702 5010
rect 208462 4890 208514 4902
rect 211598 4954 211650 4966
rect 211598 4890 211650 4902
rect 212046 4954 212098 4966
rect 212046 4890 212098 4902
rect 212494 4954 212546 4966
rect 212494 4890 212546 4902
rect 213278 4954 213330 4966
rect 213278 4890 213330 4902
rect 213726 4954 213778 4966
rect 213726 4890 213778 4902
rect 214174 4954 214226 4966
rect 214174 4890 214226 4902
rect 214622 4954 214674 4966
rect 214622 4890 214674 4902
rect 215070 4954 215122 4966
rect 215070 4890 215122 4902
rect 215518 4954 215570 4966
rect 215518 4890 215570 4902
rect 1344 4730 218624 4764
rect 1344 4678 55542 4730
rect 55594 4678 55646 4730
rect 55698 4678 55750 4730
rect 55802 4678 109870 4730
rect 109922 4678 109974 4730
rect 110026 4678 110078 4730
rect 110130 4678 164198 4730
rect 164250 4678 164302 4730
rect 164354 4678 164406 4730
rect 164458 4678 218624 4730
rect 1344 4644 218624 4678
rect 37706 4454 37718 4506
rect 37770 4503 37782 4506
rect 37770 4457 68119 4503
rect 37770 4454 37782 4457
rect 36138 4342 36150 4394
rect 36202 4391 36214 4394
rect 67946 4391 67958 4394
rect 36202 4345 67958 4391
rect 36202 4342 36214 4345
rect 67946 4342 67958 4345
rect 68010 4342 68022 4394
rect 68073 4391 68119 4457
rect 68562 4454 68574 4506
rect 68626 4503 68638 4506
rect 70410 4503 70422 4506
rect 68626 4457 70422 4503
rect 68626 4454 68638 4457
rect 70410 4454 70422 4457
rect 70474 4454 70486 4506
rect 71586 4454 71598 4506
rect 71650 4503 71662 4506
rect 72090 4503 72102 4506
rect 71650 4457 72102 4503
rect 71650 4454 71662 4457
rect 72090 4454 72102 4457
rect 72154 4503 72166 4506
rect 75674 4503 75686 4506
rect 72154 4457 75686 4503
rect 72154 4454 72166 4457
rect 75674 4454 75686 4457
rect 75738 4454 75750 4506
rect 75898 4454 75910 4506
rect 75962 4503 75974 4506
rect 79594 4503 79606 4506
rect 75962 4457 79606 4503
rect 75962 4454 75974 4457
rect 79594 4454 79606 4457
rect 79658 4454 79670 4506
rect 96058 4503 96070 4506
rect 79721 4457 96070 4503
rect 70634 4391 70646 4394
rect 68073 4345 70646 4391
rect 70634 4342 70646 4345
rect 70698 4342 70710 4394
rect 70858 4342 70870 4394
rect 70922 4391 70934 4394
rect 79721 4391 79767 4457
rect 96058 4454 96070 4457
rect 96122 4454 96134 4506
rect 96282 4454 96294 4506
rect 96346 4503 96358 4506
rect 99754 4503 99766 4506
rect 96346 4457 99766 4503
rect 96346 4454 96358 4457
rect 99754 4454 99766 4457
rect 99818 4454 99830 4506
rect 100090 4454 100102 4506
rect 100154 4503 100166 4506
rect 101994 4503 102006 4506
rect 100154 4457 102006 4503
rect 100154 4454 100166 4457
rect 101994 4454 102006 4457
rect 102058 4454 102070 4506
rect 102330 4454 102342 4506
rect 102394 4503 102406 4506
rect 115658 4503 115670 4506
rect 102394 4457 115670 4503
rect 102394 4454 102406 4457
rect 115658 4454 115670 4457
rect 115722 4454 115734 4506
rect 115994 4454 116006 4506
rect 116058 4503 116070 4506
rect 117786 4503 117798 4506
rect 116058 4457 117798 4503
rect 116058 4454 116070 4457
rect 117786 4454 117798 4457
rect 117850 4454 117862 4506
rect 118010 4454 118022 4506
rect 118074 4503 118086 4506
rect 123498 4503 123510 4506
rect 118074 4457 123510 4503
rect 118074 4454 118086 4457
rect 123498 4454 123510 4457
rect 123562 4454 123574 4506
rect 123946 4454 123958 4506
rect 124010 4503 124022 4506
rect 125458 4503 125470 4506
rect 124010 4457 125470 4503
rect 124010 4454 124022 4457
rect 125458 4454 125470 4457
rect 125522 4454 125534 4506
rect 128426 4454 128438 4506
rect 128490 4503 128502 4506
rect 133578 4503 133590 4506
rect 128490 4457 133590 4503
rect 128490 4454 128502 4457
rect 133578 4454 133590 4457
rect 133642 4454 133654 4506
rect 138282 4454 138294 4506
rect 138346 4503 138358 4506
rect 141978 4503 141990 4506
rect 138346 4457 141990 4503
rect 138346 4454 138358 4457
rect 141978 4454 141990 4457
rect 142042 4454 142054 4506
rect 142426 4454 142438 4506
rect 142490 4503 142502 4506
rect 145450 4503 145462 4506
rect 142490 4457 145462 4503
rect 142490 4454 142502 4457
rect 145450 4454 145462 4457
rect 145514 4454 145526 4506
rect 145674 4454 145686 4506
rect 145738 4503 145750 4506
rect 149482 4503 149494 4506
rect 145738 4457 149494 4503
rect 145738 4454 145750 4457
rect 149482 4454 149494 4457
rect 149546 4454 149558 4506
rect 180282 4503 180294 4506
rect 150281 4457 180294 4503
rect 70922 4345 79767 4391
rect 70922 4342 70934 4345
rect 79818 4342 79830 4394
rect 79882 4391 79894 4394
rect 80042 4391 80054 4394
rect 79882 4345 80054 4391
rect 79882 4342 79894 4345
rect 80042 4342 80054 4345
rect 80106 4342 80118 4394
rect 80266 4342 80278 4394
rect 80330 4391 80342 4394
rect 81386 4391 81398 4394
rect 80330 4345 81398 4391
rect 80330 4342 80342 4345
rect 81386 4342 81398 4345
rect 81450 4342 81462 4394
rect 82282 4342 82294 4394
rect 82346 4391 82358 4394
rect 115882 4391 115894 4394
rect 82346 4345 115894 4391
rect 82346 4342 82358 4345
rect 115882 4342 115894 4345
rect 115946 4342 115958 4394
rect 116106 4342 116118 4394
rect 116170 4391 116182 4394
rect 120026 4391 120038 4394
rect 116170 4345 120038 4391
rect 116170 4342 116182 4345
rect 120026 4342 120038 4345
rect 120090 4342 120102 4394
rect 120362 4342 120374 4394
rect 120426 4391 120438 4394
rect 120426 4345 121767 4391
rect 120426 4342 120438 4345
rect 36698 4230 36710 4282
rect 36762 4279 36774 4282
rect 104682 4279 104694 4282
rect 36762 4233 104694 4279
rect 36762 4230 36774 4233
rect 104682 4230 104694 4233
rect 104746 4230 104758 4282
rect 104906 4230 104918 4282
rect 104970 4279 104982 4282
rect 109050 4279 109062 4282
rect 104970 4233 109062 4279
rect 104970 4230 104982 4233
rect 109050 4230 109062 4233
rect 109114 4230 109126 4282
rect 109386 4230 109398 4282
rect 109450 4279 109462 4282
rect 113978 4279 113990 4282
rect 109450 4233 113990 4279
rect 109450 4230 109462 4233
rect 113978 4230 113990 4233
rect 114042 4230 114054 4282
rect 114314 4230 114326 4282
rect 114378 4279 114390 4282
rect 116330 4279 116342 4282
rect 114378 4233 116342 4279
rect 114378 4230 114390 4233
rect 116330 4230 116342 4233
rect 116394 4230 116406 4282
rect 117002 4230 117014 4282
rect 117066 4279 117078 4282
rect 119914 4279 119926 4282
rect 117066 4233 119926 4279
rect 117066 4230 117078 4233
rect 119914 4230 119926 4233
rect 119978 4230 119990 4282
rect 120250 4230 120262 4282
rect 120314 4279 120326 4282
rect 120314 4233 121655 4279
rect 120314 4230 120326 4233
rect 121609 4170 121655 4233
rect 37370 4118 37382 4170
rect 37434 4167 37446 4170
rect 120362 4167 120374 4170
rect 37434 4121 120374 4167
rect 37434 4118 37446 4121
rect 120362 4118 120374 4121
rect 120426 4118 120438 4170
rect 120545 4121 120983 4167
rect 57082 4006 57094 4058
rect 57146 4055 57158 4058
rect 58314 4055 58326 4058
rect 57146 4009 58326 4055
rect 57146 4006 57158 4009
rect 58314 4006 58326 4009
rect 58378 4006 58390 4058
rect 58650 4006 58662 4058
rect 58714 4055 58726 4058
rect 59434 4055 59446 4058
rect 58714 4009 59446 4055
rect 58714 4006 58726 4009
rect 59434 4006 59446 4009
rect 59498 4006 59510 4058
rect 65482 4055 65494 4058
rect 59561 4009 65494 4055
rect 49578 3894 49590 3946
rect 49642 3943 49654 3946
rect 59561 3943 59607 4009
rect 65482 4006 65494 4009
rect 65546 4006 65558 4058
rect 67233 4009 75511 4055
rect 49642 3897 59607 3943
rect 49642 3894 49654 3897
rect 65370 3894 65382 3946
rect 65434 3943 65446 3946
rect 67233 3943 67279 4009
rect 65434 3897 67279 3943
rect 65434 3894 65446 3897
rect 67946 3894 67958 3946
rect 68010 3943 68022 3946
rect 75338 3943 75350 3946
rect 68010 3897 75350 3943
rect 68010 3894 68022 3897
rect 75338 3894 75350 3897
rect 75402 3894 75414 3946
rect 75465 3943 75511 4009
rect 75562 4006 75574 4058
rect 75626 4055 75638 4058
rect 81834 4055 81846 4058
rect 75626 4009 81846 4055
rect 75626 4006 75638 4009
rect 81834 4006 81846 4009
rect 81898 4006 81910 4058
rect 82058 4006 82070 4058
rect 82122 4055 82134 4058
rect 85642 4055 85654 4058
rect 82122 4009 85654 4055
rect 82122 4006 82134 4009
rect 85642 4006 85654 4009
rect 85706 4006 85718 4058
rect 85866 4006 85878 4058
rect 85930 4055 85942 4058
rect 89226 4055 89238 4058
rect 85930 4009 89238 4055
rect 85930 4006 85942 4009
rect 89226 4006 89238 4009
rect 89290 4006 89302 4058
rect 89450 4006 89462 4058
rect 89514 4055 89526 4058
rect 91242 4055 91254 4058
rect 89514 4009 91254 4055
rect 89514 4006 89526 4009
rect 91242 4006 91254 4009
rect 91306 4006 91318 4058
rect 98186 4055 98198 4058
rect 91537 4009 98198 4055
rect 77354 3943 77366 3946
rect 75465 3897 77366 3943
rect 77354 3894 77366 3897
rect 77418 3894 77430 3946
rect 77578 3894 77590 3946
rect 77642 3943 77654 3946
rect 78026 3943 78038 3946
rect 77642 3897 78038 3943
rect 77642 3894 77654 3897
rect 78026 3894 78038 3897
rect 78090 3894 78102 3946
rect 78250 3894 78262 3946
rect 78314 3943 78326 3946
rect 80826 3943 80838 3946
rect 78314 3897 80838 3943
rect 78314 3894 78326 3897
rect 80826 3894 80838 3897
rect 80890 3894 80902 3946
rect 81386 3894 81398 3946
rect 81450 3943 81462 3946
rect 83738 3943 83750 3946
rect 81450 3897 83750 3943
rect 81450 3894 81462 3897
rect 83738 3894 83750 3897
rect 83802 3894 83814 3946
rect 84074 3894 84086 3946
rect 84138 3943 84150 3946
rect 91537 3943 91583 4009
rect 98186 4006 98198 4009
rect 98250 4006 98262 4058
rect 98410 4006 98422 4058
rect 98474 4055 98486 4058
rect 99306 4055 99318 4058
rect 98474 4009 99318 4055
rect 98474 4006 98486 4009
rect 99306 4006 99318 4009
rect 99370 4006 99382 4058
rect 99530 4006 99542 4058
rect 99594 4055 99606 4058
rect 99594 4009 102503 4055
rect 99594 4006 99606 4009
rect 84138 3897 91583 3943
rect 84138 3894 84150 3897
rect 91690 3894 91702 3946
rect 91754 3943 91766 3946
rect 102457 3943 102503 4009
rect 102554 4006 102566 4058
rect 102618 4055 102630 4058
rect 102618 4009 103399 4055
rect 102618 4006 102630 4009
rect 102890 3943 102902 3946
rect 91754 3897 102335 3943
rect 102457 3897 102902 3943
rect 91754 3894 91766 3897
rect 55066 3782 55078 3834
rect 55130 3831 55142 3834
rect 56634 3831 56646 3834
rect 55130 3785 56646 3831
rect 55130 3782 55142 3785
rect 56634 3782 56646 3785
rect 56698 3782 56710 3834
rect 66490 3831 66502 3834
rect 56761 3785 66502 3831
rect 52490 3670 52502 3722
rect 52554 3719 52566 3722
rect 56761 3719 56807 3785
rect 66490 3782 66502 3785
rect 66554 3782 66566 3834
rect 67050 3782 67062 3834
rect 67114 3831 67126 3834
rect 78698 3831 78710 3834
rect 67114 3785 78710 3831
rect 67114 3782 67126 3785
rect 78698 3782 78710 3785
rect 78762 3782 78774 3834
rect 79818 3782 79830 3834
rect 79882 3831 79894 3834
rect 81722 3831 81734 3834
rect 79882 3785 81734 3831
rect 79882 3782 79894 3785
rect 81722 3782 81734 3785
rect 81786 3782 81798 3834
rect 82282 3782 82294 3834
rect 82346 3831 82358 3834
rect 101994 3831 102006 3834
rect 82346 3785 102006 3831
rect 82346 3782 82358 3785
rect 101994 3782 102006 3785
rect 102058 3782 102070 3834
rect 102289 3831 102335 3897
rect 102890 3894 102902 3897
rect 102954 3894 102966 3946
rect 103353 3943 103399 4009
rect 103450 4006 103462 4058
rect 103514 4055 103526 4058
rect 104122 4055 104134 4058
rect 103514 4009 104134 4055
rect 103514 4006 103526 4009
rect 104122 4006 104134 4009
rect 104186 4006 104198 4058
rect 105802 4006 105814 4058
rect 105866 4055 105878 4058
rect 120138 4055 120150 4058
rect 105866 4009 120150 4055
rect 105866 4006 105878 4009
rect 120138 4006 120150 4009
rect 120202 4006 120214 4058
rect 120545 4055 120591 4121
rect 120265 4009 120591 4055
rect 114762 3943 114774 3946
rect 103353 3897 114774 3943
rect 114762 3894 114774 3897
rect 114826 3894 114838 3946
rect 115322 3894 115334 3946
rect 115386 3894 115398 3946
rect 120265 3943 120311 4009
rect 120937 3943 120983 4121
rect 121594 4118 121606 4170
rect 121658 4118 121670 4170
rect 121721 4167 121767 4345
rect 121818 4342 121830 4394
rect 121882 4391 121894 4394
rect 122602 4391 122614 4394
rect 121882 4345 122614 4391
rect 121882 4342 121894 4345
rect 122602 4342 122614 4345
rect 122666 4342 122678 4394
rect 124282 4342 124294 4394
rect 124346 4391 124358 4394
rect 133242 4391 133254 4394
rect 124346 4345 133254 4391
rect 124346 4342 124358 4345
rect 133242 4342 133254 4345
rect 133306 4342 133318 4394
rect 140298 4342 140310 4394
rect 140362 4391 140374 4394
rect 143266 4391 143278 4394
rect 140362 4345 143278 4391
rect 140362 4342 140374 4345
rect 143266 4342 143278 4345
rect 143330 4342 143342 4394
rect 143546 4342 143558 4394
rect 143610 4391 143622 4394
rect 150281 4391 150327 4457
rect 180282 4454 180294 4457
rect 180346 4454 180358 4506
rect 176362 4391 176374 4394
rect 143610 4345 150327 4391
rect 150393 4345 176374 4391
rect 143610 4342 143622 4345
rect 121930 4230 121942 4282
rect 121994 4279 122006 4282
rect 122826 4279 122838 4282
rect 121994 4233 122838 4279
rect 121994 4230 122006 4233
rect 122826 4230 122838 4233
rect 122890 4230 122902 4282
rect 124170 4230 124182 4282
rect 124234 4279 124246 4282
rect 150393 4279 150439 4345
rect 176362 4342 176374 4345
rect 176426 4342 176438 4394
rect 124234 4233 150439 4279
rect 124234 4230 124246 4233
rect 156090 4230 156102 4282
rect 156154 4279 156166 4282
rect 184202 4279 184214 4282
rect 156154 4233 184214 4279
rect 156154 4230 156166 4233
rect 184202 4230 184214 4233
rect 184266 4230 184278 4282
rect 127418 4167 127430 4170
rect 121721 4121 127430 4167
rect 127418 4118 127430 4121
rect 127482 4118 127494 4170
rect 127866 4118 127878 4170
rect 127930 4167 127942 4170
rect 131786 4167 131798 4170
rect 127930 4121 131798 4167
rect 127930 4118 127942 4121
rect 131786 4118 131798 4121
rect 131850 4118 131862 4170
rect 132010 4118 132022 4170
rect 132074 4167 132086 4170
rect 136154 4167 136166 4170
rect 132074 4121 136166 4167
rect 132074 4118 132086 4121
rect 136154 4118 136166 4121
rect 136218 4118 136230 4170
rect 137722 4118 137734 4170
rect 137786 4167 137798 4170
rect 139402 4167 139414 4170
rect 137786 4121 139414 4167
rect 137786 4118 137798 4121
rect 139402 4118 139414 4121
rect 139466 4118 139478 4170
rect 140634 4118 140646 4170
rect 140698 4167 140710 4170
rect 141194 4167 141206 4170
rect 140698 4121 141206 4167
rect 140698 4118 140710 4121
rect 141194 4118 141206 4121
rect 141258 4118 141270 4170
rect 143322 4118 143334 4170
rect 143386 4167 143398 4170
rect 148250 4167 148262 4170
rect 143386 4121 148262 4167
rect 143386 4118 143398 4121
rect 148250 4118 148262 4121
rect 148314 4118 148326 4170
rect 153402 4118 153414 4170
rect 153466 4167 153478 4170
rect 187002 4167 187014 4170
rect 153466 4121 187014 4167
rect 153466 4118 153478 4121
rect 187002 4118 187014 4121
rect 187066 4118 187078 4170
rect 121146 4006 121158 4058
rect 121210 4055 121222 4058
rect 134138 4055 134150 4058
rect 121210 4009 134150 4055
rect 121210 4006 121222 4009
rect 134138 4006 134150 4009
rect 134202 4006 134214 4058
rect 135818 4006 135830 4058
rect 135882 4055 135894 4058
rect 138170 4055 138182 4058
rect 135882 4009 138182 4055
rect 135882 4006 135894 4009
rect 138170 4006 138182 4009
rect 138234 4055 138246 4058
rect 143994 4055 144006 4058
rect 138234 4009 144006 4055
rect 138234 4006 138246 4009
rect 143994 4006 144006 4009
rect 144058 4006 144070 4058
rect 145450 4006 145462 4058
rect 145514 4055 145526 4058
rect 148138 4055 148150 4058
rect 145514 4009 148150 4055
rect 145514 4006 145526 4009
rect 148138 4006 148150 4009
rect 148202 4055 148214 4058
rect 150042 4055 150054 4058
rect 148202 4009 150054 4055
rect 148202 4006 148214 4009
rect 150042 4006 150054 4009
rect 150106 4006 150118 4058
rect 152618 4006 152630 4058
rect 152682 4055 152694 4058
rect 159114 4055 159126 4058
rect 152682 4009 159126 4055
rect 152682 4006 152694 4009
rect 159114 4006 159126 4009
rect 159178 4055 159190 4058
rect 161018 4055 161030 4058
rect 159178 4009 161030 4055
rect 159178 4006 159190 4009
rect 161018 4006 161030 4009
rect 161082 4006 161094 4058
rect 166394 4006 166406 4058
rect 166458 4055 166470 4058
rect 190138 4055 190150 4058
rect 166458 4009 190150 4055
rect 166458 4006 166470 4009
rect 190138 4006 190150 4009
rect 190202 4006 190214 4058
rect 191258 4006 191270 4058
rect 191322 4055 191334 4058
rect 193050 4055 193062 4058
rect 191322 4009 193062 4055
rect 191322 4006 191334 4009
rect 193050 4006 193062 4009
rect 193114 4006 193126 4058
rect 134250 3943 134262 3946
rect 115449 3897 120311 3943
rect 120489 3897 120759 3943
rect 120937 3897 134262 3943
rect 102289 3785 114263 3831
rect 52554 3673 56807 3719
rect 52554 3670 52566 3673
rect 59658 3670 59670 3722
rect 59722 3719 59734 3722
rect 66714 3719 66726 3722
rect 59722 3673 66726 3719
rect 59722 3670 59734 3673
rect 66714 3670 66726 3673
rect 66778 3670 66790 3722
rect 67162 3670 67174 3722
rect 67226 3719 67238 3722
rect 77130 3719 77142 3722
rect 67226 3673 77142 3719
rect 67226 3670 67238 3673
rect 77130 3670 77142 3673
rect 77194 3670 77206 3722
rect 77354 3670 77366 3722
rect 77418 3719 77430 3722
rect 78586 3719 78598 3722
rect 77418 3673 78598 3719
rect 77418 3670 77430 3673
rect 78586 3670 78598 3673
rect 78650 3670 78662 3722
rect 78810 3670 78822 3722
rect 78874 3719 78886 3722
rect 83066 3719 83078 3722
rect 78874 3673 83078 3719
rect 78874 3670 78886 3673
rect 83066 3670 83078 3673
rect 83130 3670 83142 3722
rect 83402 3670 83414 3722
rect 83466 3719 83478 3722
rect 99418 3719 99430 3722
rect 83466 3673 99430 3719
rect 83466 3670 83478 3673
rect 99418 3670 99430 3673
rect 99482 3670 99494 3722
rect 102666 3719 102678 3722
rect 99713 3673 102678 3719
rect 43418 3558 43430 3610
rect 43482 3607 43494 3610
rect 63914 3607 63926 3610
rect 43482 3561 63926 3607
rect 43482 3558 43494 3561
rect 63914 3558 63926 3561
rect 63978 3558 63990 3610
rect 68394 3558 68406 3610
rect 68458 3607 68470 3610
rect 68458 3561 79095 3607
rect 68458 3558 68470 3561
rect 79049 3498 79095 3561
rect 79258 3558 79270 3610
rect 79322 3607 79334 3610
rect 79322 3561 80103 3607
rect 79322 3558 79334 3561
rect 31882 3446 31894 3498
rect 31946 3495 31958 3498
rect 77354 3495 77366 3498
rect 31946 3449 77366 3495
rect 31946 3446 31958 3449
rect 77354 3446 77366 3449
rect 77418 3446 77430 3498
rect 78489 3449 78983 3495
rect 33002 3334 33014 3386
rect 33066 3383 33078 3386
rect 78489 3383 78535 3449
rect 78810 3383 78822 3386
rect 33066 3337 78535 3383
rect 78601 3337 78822 3383
rect 33066 3334 33078 3337
rect 21578 3222 21590 3274
rect 21642 3271 21654 3274
rect 56186 3271 56198 3274
rect 21642 3225 56198 3271
rect 21642 3222 21654 3225
rect 56186 3222 56198 3225
rect 56250 3222 56262 3274
rect 68954 3271 68966 3274
rect 66057 3225 68966 3271
rect 27514 3110 27526 3162
rect 27578 3159 27590 3162
rect 57866 3159 57878 3162
rect 27578 3113 57878 3159
rect 27578 3110 27590 3113
rect 57866 3110 57878 3113
rect 57930 3110 57942 3162
rect 58090 3110 58102 3162
rect 58154 3159 58166 3162
rect 66057 3159 66103 3225
rect 68954 3222 68966 3225
rect 69018 3222 69030 3274
rect 69402 3222 69414 3274
rect 69466 3271 69478 3274
rect 78601 3271 78647 3337
rect 78810 3334 78822 3337
rect 78874 3334 78886 3386
rect 78937 3383 78983 3449
rect 79034 3446 79046 3498
rect 79098 3446 79110 3498
rect 80057 3495 80103 3561
rect 80378 3558 80390 3610
rect 80442 3607 80454 3610
rect 85418 3607 85430 3610
rect 80442 3561 85430 3607
rect 80442 3558 80454 3561
rect 85418 3558 85430 3561
rect 85482 3558 85494 3610
rect 86202 3558 86214 3610
rect 86266 3607 86278 3610
rect 89226 3607 89238 3610
rect 86266 3561 89238 3607
rect 86266 3558 86278 3561
rect 89226 3558 89238 3561
rect 89290 3558 89302 3610
rect 89562 3558 89574 3610
rect 89626 3607 89638 3610
rect 98410 3607 98422 3610
rect 89626 3561 98422 3607
rect 89626 3558 89638 3561
rect 98410 3558 98422 3561
rect 98474 3558 98486 3610
rect 98634 3558 98646 3610
rect 98698 3607 98710 3610
rect 99713 3607 99759 3673
rect 102666 3670 102678 3673
rect 102730 3670 102742 3722
rect 104122 3670 104134 3722
rect 104186 3719 104198 3722
rect 110618 3719 110630 3722
rect 104186 3673 110630 3719
rect 104186 3670 104198 3673
rect 110618 3670 110630 3673
rect 110682 3670 110694 3722
rect 112746 3670 112758 3722
rect 112810 3670 112822 3722
rect 113194 3670 113206 3722
rect 113258 3719 113270 3722
rect 113642 3719 113654 3722
rect 113258 3673 113654 3719
rect 113258 3670 113270 3673
rect 113642 3670 113654 3673
rect 113706 3670 113718 3722
rect 113866 3670 113878 3722
rect 113930 3719 113942 3722
rect 114090 3719 114102 3722
rect 113930 3673 114102 3719
rect 113930 3670 113942 3673
rect 114090 3670 114102 3673
rect 114154 3670 114166 3722
rect 114217 3719 114263 3785
rect 114538 3782 114550 3834
rect 114602 3831 114614 3834
rect 115337 3831 115383 3894
rect 115449 3834 115495 3897
rect 114602 3785 115383 3831
rect 114602 3782 114614 3785
rect 115434 3782 115446 3834
rect 115498 3782 115510 3834
rect 115770 3782 115782 3834
rect 115834 3831 115846 3834
rect 115834 3785 118743 3831
rect 115834 3782 115846 3785
rect 114217 3673 114711 3719
rect 98698 3561 99759 3607
rect 98698 3558 98710 3561
rect 100986 3558 100998 3610
rect 101050 3607 101062 3610
rect 102330 3607 102342 3610
rect 101050 3561 102342 3607
rect 101050 3558 101062 3561
rect 102330 3558 102342 3561
rect 102394 3558 102406 3610
rect 104010 3558 104022 3610
rect 104074 3607 104086 3610
rect 112634 3607 112646 3610
rect 104074 3561 112646 3607
rect 104074 3558 104086 3561
rect 112634 3558 112646 3561
rect 112698 3558 112710 3610
rect 112761 3607 112807 3670
rect 113978 3607 113990 3610
rect 112761 3561 113990 3607
rect 113978 3558 113990 3561
rect 114042 3558 114054 3610
rect 114202 3558 114214 3610
rect 114266 3607 114278 3610
rect 114665 3607 114711 3673
rect 115098 3670 115110 3722
rect 115162 3719 115174 3722
rect 118570 3719 118582 3722
rect 115162 3673 118582 3719
rect 115162 3670 115174 3673
rect 118570 3670 118582 3673
rect 118634 3670 118646 3722
rect 118697 3719 118743 3785
rect 118794 3782 118806 3834
rect 118858 3831 118870 3834
rect 120489 3831 120535 3897
rect 118858 3785 120535 3831
rect 120713 3831 120759 3897
rect 134250 3894 134262 3897
rect 134314 3894 134326 3946
rect 139178 3894 139190 3946
rect 139242 3943 139254 3946
rect 140410 3943 140422 3946
rect 139242 3897 140422 3943
rect 139242 3894 139254 3897
rect 140410 3894 140422 3897
rect 140474 3943 140486 3946
rect 141530 3943 141542 3946
rect 140474 3897 141542 3943
rect 140474 3894 140486 3897
rect 141530 3894 141542 3897
rect 141594 3894 141606 3946
rect 145338 3894 145350 3946
rect 145402 3943 145414 3946
rect 149146 3943 149158 3946
rect 145402 3897 149158 3943
rect 145402 3894 145414 3897
rect 149146 3894 149158 3897
rect 149210 3894 149222 3946
rect 174234 3894 174246 3946
rect 174298 3943 174310 3946
rect 194170 3943 194182 3946
rect 174298 3897 194182 3943
rect 174298 3894 174310 3897
rect 194170 3894 194182 3897
rect 194234 3894 194246 3946
rect 131226 3831 131238 3834
rect 120713 3785 131238 3831
rect 118858 3782 118870 3785
rect 131226 3782 131238 3785
rect 131290 3782 131302 3834
rect 134362 3782 134374 3834
rect 134426 3831 134438 3834
rect 147914 3831 147926 3834
rect 134426 3785 147926 3831
rect 134426 3782 134438 3785
rect 147914 3782 147926 3785
rect 147978 3782 147990 3834
rect 158778 3782 158790 3834
rect 158842 3831 158854 3834
rect 159450 3831 159462 3834
rect 158842 3785 159462 3831
rect 158842 3782 158854 3785
rect 159450 3782 159462 3785
rect 159514 3782 159526 3834
rect 171882 3782 171894 3834
rect 171946 3831 171958 3834
rect 191482 3831 191494 3834
rect 171946 3785 191494 3831
rect 171946 3782 171958 3785
rect 191482 3782 191494 3785
rect 191546 3782 191558 3834
rect 118697 3673 120535 3719
rect 114266 3561 114599 3607
rect 114665 3561 120423 3607
rect 114266 3558 114278 3561
rect 84410 3495 84422 3498
rect 79161 3449 79991 3495
rect 80057 3449 84422 3495
rect 79161 3383 79207 3449
rect 79706 3383 79718 3386
rect 78937 3337 79207 3383
rect 79329 3337 79718 3383
rect 69466 3225 78647 3271
rect 69466 3222 69478 3225
rect 78698 3222 78710 3274
rect 78762 3271 78774 3274
rect 78762 3225 79095 3271
rect 78762 3222 78774 3225
rect 58154 3113 66103 3159
rect 58154 3110 58166 3113
rect 66602 3110 66614 3162
rect 66666 3159 66678 3162
rect 78922 3159 78934 3162
rect 66666 3113 78934 3159
rect 66666 3110 66678 3113
rect 78922 3110 78934 3113
rect 78986 3110 78998 3162
rect 79049 3159 79095 3225
rect 79329 3159 79375 3337
rect 79706 3334 79718 3337
rect 79770 3334 79782 3386
rect 79945 3383 79991 3449
rect 84410 3446 84422 3449
rect 84474 3446 84486 3498
rect 84634 3446 84646 3498
rect 84698 3495 84710 3498
rect 92810 3495 92822 3498
rect 84698 3449 92822 3495
rect 84698 3446 84710 3449
rect 92810 3446 92822 3449
rect 92874 3446 92886 3498
rect 93146 3446 93158 3498
rect 93210 3495 93222 3498
rect 103450 3495 103462 3498
rect 93210 3449 103462 3495
rect 93210 3446 93222 3449
rect 103450 3446 103462 3449
rect 103514 3446 103526 3498
rect 104682 3446 104694 3498
rect 104746 3495 104758 3498
rect 104746 3449 111799 3495
rect 104746 3446 104758 3449
rect 91690 3383 91702 3386
rect 79945 3337 91702 3383
rect 91690 3334 91702 3337
rect 91754 3334 91766 3386
rect 91914 3334 91926 3386
rect 91978 3383 91990 3386
rect 94378 3383 94390 3386
rect 91978 3337 94390 3383
rect 91978 3334 91990 3337
rect 94378 3334 94390 3337
rect 94442 3334 94454 3386
rect 96842 3334 96854 3386
rect 96906 3383 96918 3386
rect 101098 3383 101110 3386
rect 96906 3337 101110 3383
rect 96906 3334 96918 3337
rect 101098 3334 101110 3337
rect 101162 3334 101174 3386
rect 102330 3334 102342 3386
rect 102394 3383 102406 3386
rect 111626 3383 111638 3386
rect 102394 3337 111638 3383
rect 102394 3334 102406 3337
rect 111626 3334 111638 3337
rect 111690 3334 111702 3386
rect 111753 3383 111799 3449
rect 111850 3446 111862 3498
rect 111914 3495 111926 3498
rect 113530 3495 113542 3498
rect 111914 3449 113542 3495
rect 111914 3446 111926 3449
rect 113530 3446 113542 3449
rect 113594 3446 113606 3498
rect 114426 3495 114438 3498
rect 113881 3449 114438 3495
rect 113881 3383 113927 3449
rect 114426 3446 114438 3449
rect 114490 3446 114502 3498
rect 114553 3495 114599 3561
rect 120377 3498 120423 3561
rect 114874 3495 114886 3498
rect 114553 3449 114886 3495
rect 114874 3446 114886 3449
rect 114938 3446 114950 3498
rect 115210 3446 115222 3498
rect 115274 3495 115286 3498
rect 116890 3495 116902 3498
rect 115274 3449 116902 3495
rect 115274 3446 115286 3449
rect 116890 3446 116902 3449
rect 116954 3446 116966 3498
rect 117114 3446 117126 3498
rect 117178 3495 117190 3498
rect 119690 3495 119702 3498
rect 117178 3449 119702 3495
rect 117178 3446 117190 3449
rect 119690 3446 119702 3449
rect 119754 3446 119766 3498
rect 120362 3446 120374 3498
rect 120426 3446 120438 3498
rect 120489 3495 120535 3673
rect 120586 3670 120598 3722
rect 120650 3719 120662 3722
rect 132346 3719 132358 3722
rect 120650 3673 132358 3719
rect 120650 3670 120662 3673
rect 132346 3670 132358 3673
rect 132410 3670 132422 3722
rect 134026 3670 134038 3722
rect 134090 3719 134102 3722
rect 134810 3719 134822 3722
rect 134090 3673 134822 3719
rect 134090 3670 134102 3673
rect 134810 3670 134822 3673
rect 134874 3670 134886 3722
rect 135034 3670 135046 3722
rect 135098 3719 135110 3722
rect 143546 3719 143558 3722
rect 135098 3673 143558 3719
rect 135098 3670 135110 3673
rect 143546 3670 143558 3673
rect 143610 3670 143622 3722
rect 143994 3670 144006 3722
rect 144058 3719 144070 3722
rect 146122 3719 146134 3722
rect 144058 3673 146134 3719
rect 144058 3670 144070 3673
rect 146122 3670 146134 3673
rect 146186 3670 146198 3722
rect 153066 3670 153078 3722
rect 153130 3719 153142 3722
rect 153290 3719 153302 3722
rect 153130 3673 153302 3719
rect 153130 3670 153142 3673
rect 153290 3670 153302 3673
rect 153354 3670 153366 3722
rect 121146 3558 121158 3610
rect 121210 3607 121222 3610
rect 131450 3607 131462 3610
rect 121210 3561 131462 3607
rect 121210 3558 121222 3561
rect 131450 3558 131462 3561
rect 131514 3558 131526 3610
rect 132010 3558 132022 3610
rect 132074 3607 132086 3610
rect 132074 3561 139462 3607
rect 132074 3558 132086 3561
rect 121482 3495 121494 3498
rect 120489 3449 121494 3495
rect 121482 3446 121494 3449
rect 121546 3446 121558 3498
rect 122154 3446 122166 3498
rect 122218 3495 122230 3498
rect 127866 3495 127878 3498
rect 122218 3449 127878 3495
rect 122218 3446 122230 3449
rect 127866 3446 127878 3449
rect 127930 3446 127942 3498
rect 130890 3446 130902 3498
rect 130954 3495 130966 3498
rect 133466 3495 133478 3498
rect 130954 3449 133478 3495
rect 130954 3446 130966 3449
rect 133466 3446 133478 3449
rect 133530 3446 133542 3498
rect 111753 3337 113927 3383
rect 113978 3334 113990 3386
rect 114042 3383 114054 3386
rect 115770 3383 115782 3386
rect 114042 3337 115782 3383
rect 114042 3334 114054 3337
rect 115770 3334 115782 3337
rect 115834 3334 115846 3386
rect 116218 3334 116230 3386
rect 116282 3383 116294 3386
rect 116282 3337 117623 3383
rect 116282 3334 116294 3337
rect 85194 3271 85206 3274
rect 79049 3113 79375 3159
rect 79441 3225 85206 3271
rect 38490 2998 38502 3050
rect 38554 3047 38566 3050
rect 65258 3047 65270 3050
rect 38554 3001 65270 3047
rect 38554 2998 38566 3001
rect 65258 2998 65270 3001
rect 65322 2998 65334 3050
rect 65482 2998 65494 3050
rect 65546 3047 65558 3050
rect 78474 3047 78486 3050
rect 65546 3001 78486 3047
rect 65546 2998 65558 3001
rect 78474 2998 78486 3001
rect 78538 2998 78550 3050
rect 78698 2998 78710 3050
rect 78762 3047 78774 3050
rect 79034 3047 79046 3050
rect 78762 3001 79046 3047
rect 78762 2998 78774 3001
rect 79034 2998 79046 3001
rect 79098 2998 79110 3050
rect 51930 2886 51942 2938
rect 51994 2935 52006 2938
rect 79441 2935 79487 3225
rect 85194 3222 85206 3225
rect 85258 3222 85270 3274
rect 85418 3222 85430 3274
rect 85482 3271 85494 3274
rect 93146 3271 93158 3274
rect 85482 3225 93158 3271
rect 85482 3222 85494 3225
rect 93146 3222 93158 3225
rect 93210 3222 93222 3274
rect 94154 3222 94166 3274
rect 94218 3271 94230 3274
rect 95722 3271 95734 3274
rect 94218 3225 95734 3271
rect 94218 3222 94230 3225
rect 95722 3222 95734 3225
rect 95786 3222 95798 3274
rect 96058 3222 96070 3274
rect 96122 3271 96134 3274
rect 117338 3271 117350 3274
rect 96122 3225 100823 3271
rect 96122 3222 96134 3225
rect 79594 3110 79606 3162
rect 79658 3159 79670 3162
rect 81498 3159 81510 3162
rect 79658 3113 81510 3159
rect 79658 3110 79670 3113
rect 81498 3110 81510 3113
rect 81562 3159 81574 3162
rect 81946 3159 81958 3162
rect 81562 3113 81958 3159
rect 81562 3110 81574 3113
rect 81946 3110 81958 3113
rect 82010 3110 82022 3162
rect 82394 3110 82406 3162
rect 82458 3159 82470 3162
rect 82954 3159 82966 3162
rect 82458 3113 82966 3159
rect 82458 3110 82470 3113
rect 82954 3110 82966 3113
rect 83018 3110 83030 3162
rect 83178 3110 83190 3162
rect 83242 3159 83254 3162
rect 90906 3159 90918 3162
rect 83242 3113 90918 3159
rect 83242 3110 83254 3113
rect 90906 3110 90918 3113
rect 90970 3110 90982 3162
rect 91466 3110 91478 3162
rect 91530 3159 91542 3162
rect 100650 3159 100662 3162
rect 91530 3113 100662 3159
rect 91530 3110 91542 3113
rect 100650 3110 100662 3113
rect 100714 3110 100726 3162
rect 100777 3159 100823 3225
rect 101225 3225 117350 3271
rect 101225 3159 101271 3225
rect 117338 3222 117350 3225
rect 117402 3222 117414 3274
rect 117577 3271 117623 3337
rect 117674 3334 117686 3386
rect 117738 3383 117750 3386
rect 132794 3383 132806 3386
rect 117738 3337 132806 3383
rect 117738 3334 117750 3337
rect 132794 3334 132806 3337
rect 132858 3334 132870 3386
rect 139416 3383 139462 3561
rect 141082 3558 141094 3610
rect 141146 3607 141158 3610
rect 151050 3607 151062 3610
rect 141146 3561 151062 3607
rect 141146 3558 141158 3561
rect 151050 3558 151062 3561
rect 151114 3558 151126 3610
rect 152394 3558 152406 3610
rect 152458 3607 152470 3610
rect 156314 3607 156326 3610
rect 152458 3561 156326 3607
rect 152458 3558 152470 3561
rect 156314 3558 156326 3561
rect 156378 3558 156390 3610
rect 140970 3446 140982 3498
rect 141034 3495 141046 3498
rect 141034 3449 144502 3495
rect 141034 3446 141046 3449
rect 140186 3383 140198 3386
rect 132921 3337 133415 3383
rect 139416 3337 140198 3383
rect 132921 3271 132967 3337
rect 117577 3225 132967 3271
rect 133369 3271 133415 3337
rect 140186 3334 140198 3337
rect 140250 3383 140262 3386
rect 143098 3383 143110 3386
rect 140250 3337 143110 3383
rect 140250 3334 140262 3337
rect 143098 3334 143110 3337
rect 143162 3334 143174 3386
rect 144456 3383 144502 3449
rect 147802 3446 147814 3498
rect 147866 3495 147878 3498
rect 154858 3495 154870 3498
rect 147866 3449 154870 3495
rect 147866 3446 147878 3449
rect 154858 3446 154870 3449
rect 154922 3446 154934 3498
rect 156426 3446 156438 3498
rect 156490 3495 156502 3498
rect 189466 3495 189478 3498
rect 156490 3449 189478 3495
rect 156490 3446 156502 3449
rect 189466 3446 189478 3449
rect 189530 3446 189542 3498
rect 152506 3383 152518 3386
rect 144456 3337 152518 3383
rect 152506 3334 152518 3337
rect 152570 3334 152582 3386
rect 152842 3334 152854 3386
rect 152906 3383 152918 3386
rect 187562 3383 187574 3386
rect 152906 3337 187574 3383
rect 152906 3334 152918 3337
rect 187562 3334 187574 3337
rect 187626 3334 187638 3386
rect 150378 3271 150390 3274
rect 133369 3225 150390 3271
rect 150378 3222 150390 3225
rect 150442 3222 150454 3274
rect 178938 3222 178950 3274
rect 179002 3271 179014 3274
rect 191594 3271 191606 3274
rect 179002 3225 191606 3271
rect 179002 3222 179014 3225
rect 191594 3222 191606 3225
rect 191658 3222 191670 3274
rect 100777 3113 101271 3159
rect 101770 3110 101782 3162
rect 101834 3159 101846 3162
rect 107818 3159 107830 3162
rect 101834 3113 107830 3159
rect 101834 3110 101846 3113
rect 107818 3110 107830 3113
rect 107882 3110 107894 3162
rect 108490 3110 108502 3162
rect 108554 3159 108566 3162
rect 117562 3159 117574 3162
rect 108554 3113 117574 3159
rect 108554 3110 108566 3113
rect 117562 3110 117574 3113
rect 117626 3110 117638 3162
rect 117786 3110 117798 3162
rect 117850 3159 117862 3162
rect 119130 3159 119142 3162
rect 117850 3113 119142 3159
rect 117850 3110 117862 3113
rect 119130 3110 119142 3113
rect 119194 3159 119206 3162
rect 119578 3159 119590 3162
rect 119194 3113 119590 3159
rect 119194 3110 119206 3113
rect 119578 3110 119590 3113
rect 119642 3110 119654 3162
rect 120026 3110 120038 3162
rect 120090 3159 120102 3162
rect 138618 3159 138630 3162
rect 120090 3113 138630 3159
rect 120090 3110 120102 3113
rect 138618 3110 138630 3113
rect 138682 3110 138694 3162
rect 151498 3159 151510 3162
rect 138745 3113 151510 3159
rect 79706 2998 79718 3050
rect 79770 3047 79782 3050
rect 80154 3047 80166 3050
rect 79770 3001 80166 3047
rect 79770 2998 79782 3001
rect 80154 2998 80166 3001
rect 80218 2998 80230 3050
rect 80938 2998 80950 3050
rect 81002 3047 81014 3050
rect 82618 3047 82630 3050
rect 81002 3001 82630 3047
rect 81002 2998 81014 3001
rect 82618 2998 82630 3001
rect 82682 2998 82694 3050
rect 82842 2998 82854 3050
rect 82906 3047 82918 3050
rect 82906 3001 84471 3047
rect 82906 2998 82918 3001
rect 51994 2889 79487 2935
rect 51994 2886 52006 2889
rect 79594 2886 79606 2938
rect 79658 2935 79670 2938
rect 82282 2935 82294 2938
rect 79658 2889 82294 2935
rect 79658 2886 79670 2889
rect 82282 2886 82294 2889
rect 82346 2886 82358 2938
rect 82506 2886 82518 2938
rect 82570 2935 82582 2938
rect 84298 2935 84310 2938
rect 82570 2889 84310 2935
rect 82570 2886 82582 2889
rect 84298 2886 84310 2889
rect 84362 2886 84374 2938
rect 84425 2935 84471 3001
rect 84522 2998 84534 3050
rect 84586 3047 84598 3050
rect 85082 3047 85094 3050
rect 84586 3001 85094 3047
rect 84586 2998 84598 3001
rect 85082 2998 85094 3001
rect 85146 2998 85158 3050
rect 85306 2998 85318 3050
rect 85370 3047 85382 3050
rect 91914 3047 91926 3050
rect 85370 3001 91926 3047
rect 85370 2998 85382 3001
rect 91914 2998 91926 3001
rect 91978 2998 91990 3050
rect 92138 2998 92150 3050
rect 92202 3047 92214 3050
rect 99866 3047 99878 3050
rect 92202 3001 99878 3047
rect 92202 2998 92214 3001
rect 99866 2998 99878 3001
rect 99930 2998 99942 3050
rect 100202 2998 100214 3050
rect 100266 3047 100278 3050
rect 102442 3047 102454 3050
rect 100266 3001 102454 3047
rect 100266 2998 100278 3001
rect 102442 2998 102454 3001
rect 102506 2998 102518 3050
rect 102890 2998 102902 3050
rect 102954 3047 102966 3050
rect 104010 3047 104022 3050
rect 102954 3001 104022 3047
rect 102954 2998 102966 3001
rect 104010 2998 104022 3001
rect 104074 2998 104086 3050
rect 104234 2998 104246 3050
rect 104298 3047 104310 3050
rect 116442 3047 116454 3050
rect 104298 3001 116454 3047
rect 104298 2998 104310 3001
rect 116442 2998 116454 3001
rect 116506 2998 116518 3050
rect 117338 2998 117350 3050
rect 117402 3047 117414 3050
rect 117402 3001 132742 3047
rect 117402 2998 117414 3001
rect 90682 2935 90694 2938
rect 84425 2889 90694 2935
rect 90682 2886 90694 2889
rect 90746 2886 90758 2938
rect 90906 2886 90918 2938
rect 90970 2935 90982 2938
rect 95946 2935 95958 2938
rect 90970 2889 95958 2935
rect 90970 2886 90982 2889
rect 95946 2886 95958 2889
rect 96010 2886 96022 2938
rect 96170 2886 96182 2938
rect 96234 2935 96246 2938
rect 99306 2935 99318 2938
rect 96234 2889 99318 2935
rect 96234 2886 96246 2889
rect 99306 2886 99318 2889
rect 99370 2886 99382 2938
rect 99657 2889 100823 2935
rect 27514 2774 27526 2826
rect 27578 2823 27590 2826
rect 58650 2823 58662 2826
rect 27578 2777 58662 2823
rect 27578 2774 27590 2777
rect 58650 2774 58662 2777
rect 58714 2774 58726 2826
rect 61674 2774 61686 2826
rect 61738 2823 61750 2826
rect 99082 2823 99094 2826
rect 61738 2777 99094 2823
rect 61738 2774 61750 2777
rect 99082 2774 99094 2777
rect 99146 2774 99158 2826
rect 23258 2662 23270 2714
rect 23322 2711 23334 2714
rect 67386 2711 67398 2714
rect 23322 2665 67398 2711
rect 23322 2662 23334 2665
rect 67386 2662 67398 2665
rect 67450 2662 67462 2714
rect 79034 2711 79046 2714
rect 67513 2665 79046 2711
rect 22026 2550 22038 2602
rect 22090 2599 22102 2602
rect 58090 2599 58102 2602
rect 22090 2553 58102 2599
rect 22090 2550 22102 2553
rect 58090 2550 58102 2553
rect 58154 2550 58166 2602
rect 58874 2550 58886 2602
rect 58938 2599 58950 2602
rect 66266 2599 66278 2602
rect 58938 2553 66278 2599
rect 58938 2550 58950 2553
rect 66266 2550 66278 2553
rect 66330 2550 66342 2602
rect 66602 2550 66614 2602
rect 66666 2599 66678 2602
rect 67513 2599 67559 2665
rect 79034 2662 79046 2665
rect 79098 2662 79110 2714
rect 79482 2662 79494 2714
rect 79546 2711 79558 2714
rect 99657 2711 99703 2889
rect 100314 2774 100326 2826
rect 100378 2823 100390 2826
rect 100650 2823 100662 2826
rect 100378 2777 100662 2823
rect 100378 2774 100390 2777
rect 100650 2774 100662 2777
rect 100714 2774 100726 2826
rect 79546 2665 99703 2711
rect 79546 2662 79558 2665
rect 99754 2662 99766 2714
rect 99818 2711 99830 2714
rect 100777 2711 100823 2889
rect 101098 2886 101110 2938
rect 101162 2935 101174 2938
rect 132458 2935 132470 2938
rect 101162 2889 132470 2935
rect 101162 2886 101174 2889
rect 132458 2886 132470 2889
rect 132522 2886 132534 2938
rect 101882 2774 101894 2826
rect 101946 2823 101958 2826
rect 110842 2823 110854 2826
rect 101946 2777 110854 2823
rect 101946 2774 101958 2777
rect 110842 2774 110854 2777
rect 110906 2774 110918 2826
rect 115882 2823 115894 2826
rect 110969 2777 115894 2823
rect 110730 2711 110742 2714
rect 99818 2665 100375 2711
rect 100777 2665 110742 2711
rect 99818 2662 99830 2665
rect 66666 2553 67559 2599
rect 66666 2550 66678 2553
rect 68170 2550 68182 2602
rect 68234 2599 68246 2602
rect 79594 2599 79606 2602
rect 68234 2553 79606 2599
rect 68234 2550 68246 2553
rect 79594 2550 79606 2553
rect 79658 2550 79670 2602
rect 80154 2550 80166 2602
rect 80218 2599 80230 2602
rect 100202 2599 100214 2602
rect 80218 2553 100214 2599
rect 80218 2550 80230 2553
rect 100202 2550 100214 2553
rect 100266 2550 100278 2602
rect 100329 2599 100375 2665
rect 110730 2662 110742 2665
rect 110794 2662 110806 2714
rect 104906 2599 104918 2602
rect 100329 2553 104918 2599
rect 104906 2550 104918 2553
rect 104970 2550 104982 2602
rect 105130 2550 105142 2602
rect 105194 2599 105206 2602
rect 110969 2599 111015 2777
rect 115882 2774 115894 2777
rect 115946 2774 115958 2826
rect 116890 2774 116902 2826
rect 116954 2823 116966 2826
rect 117786 2823 117798 2826
rect 116954 2777 117798 2823
rect 116954 2774 116966 2777
rect 117786 2774 117798 2777
rect 117850 2774 117862 2826
rect 118458 2774 118470 2826
rect 118522 2823 118534 2826
rect 132696 2823 132742 3001
rect 133466 2998 133478 3050
rect 133530 3047 133542 3050
rect 138745 3047 138791 3113
rect 151498 3110 151510 3113
rect 151562 3110 151574 3162
rect 161018 3110 161030 3162
rect 161082 3159 161094 3162
rect 207722 3159 207734 3162
rect 161082 3113 207734 3159
rect 161082 3110 161094 3113
rect 207722 3110 207734 3113
rect 207786 3110 207798 3162
rect 133530 3001 138791 3047
rect 133530 2998 133542 3001
rect 150714 2998 150726 3050
rect 150778 3047 150790 3050
rect 150778 3001 153239 3047
rect 150778 2998 150790 3001
rect 132794 2886 132806 2938
rect 132858 2935 132870 2938
rect 153066 2935 153078 2938
rect 132858 2889 153078 2935
rect 132858 2886 132870 2889
rect 153066 2886 153078 2889
rect 153130 2886 153142 2938
rect 153193 2935 153239 3001
rect 154970 2998 154982 3050
rect 155034 3047 155046 3050
rect 189914 3047 189926 3050
rect 155034 3001 189926 3047
rect 155034 2998 155046 3001
rect 189914 2998 189926 3001
rect 189978 3047 189990 3050
rect 192266 3047 192278 3050
rect 189978 3001 192278 3047
rect 189978 2998 189990 3001
rect 192266 2998 192278 3001
rect 192330 2998 192342 3050
rect 186106 2935 186118 2938
rect 153193 2889 186118 2935
rect 186106 2886 186118 2889
rect 186170 2886 186182 2938
rect 154410 2823 154422 2826
rect 118522 2777 126919 2823
rect 132696 2777 154422 2823
rect 118522 2774 118534 2777
rect 111178 2662 111190 2714
rect 111242 2711 111254 2714
rect 117450 2711 117462 2714
rect 111242 2665 117462 2711
rect 111242 2662 111254 2665
rect 117450 2662 117462 2665
rect 117514 2662 117526 2714
rect 117674 2662 117686 2714
rect 117738 2711 117750 2714
rect 126746 2711 126758 2714
rect 117738 2665 126758 2711
rect 117738 2662 117750 2665
rect 126746 2662 126758 2665
rect 126810 2662 126822 2714
rect 105194 2553 111015 2599
rect 105194 2550 105206 2553
rect 111066 2550 111078 2602
rect 111130 2599 111142 2602
rect 126873 2599 126919 2777
rect 154410 2774 154422 2777
rect 154474 2774 154486 2826
rect 162698 2823 162710 2826
rect 161256 2777 162710 2823
rect 127306 2662 127318 2714
rect 127370 2711 127382 2714
rect 161256 2711 161302 2777
rect 162698 2774 162710 2777
rect 162762 2774 162774 2826
rect 185994 2774 186006 2826
rect 186058 2823 186070 2826
rect 186442 2823 186454 2826
rect 186058 2777 186454 2823
rect 186058 2774 186070 2777
rect 186442 2774 186454 2777
rect 186506 2774 186518 2826
rect 127370 2665 161302 2711
rect 127370 2662 127382 2665
rect 186554 2662 186566 2714
rect 186618 2711 186630 2714
rect 201562 2711 201574 2714
rect 186618 2665 201574 2711
rect 186618 2662 186630 2665
rect 201562 2662 201574 2665
rect 201626 2662 201638 2714
rect 174346 2599 174358 2602
rect 111130 2553 126807 2599
rect 126873 2553 174358 2599
rect 111130 2550 111142 2553
rect 21466 2438 21478 2490
rect 21530 2487 21542 2490
rect 65370 2487 65382 2490
rect 21530 2441 65382 2487
rect 21530 2438 21542 2441
rect 65370 2438 65382 2441
rect 65434 2438 65446 2490
rect 65930 2438 65942 2490
rect 65994 2487 66006 2490
rect 126761 2487 126807 2553
rect 174346 2550 174358 2553
rect 174410 2550 174422 2602
rect 175018 2550 175030 2602
rect 175082 2599 175094 2602
rect 196410 2599 196422 2602
rect 175082 2553 196422 2599
rect 175082 2550 175094 2553
rect 196410 2550 196422 2553
rect 196474 2550 196486 2602
rect 65994 2441 126695 2487
rect 126761 2441 134423 2487
rect 65994 2438 66006 2441
rect 37930 2326 37942 2378
rect 37994 2375 38006 2378
rect 62010 2375 62022 2378
rect 37994 2329 62022 2375
rect 37994 2326 38006 2329
rect 62010 2326 62022 2329
rect 62074 2326 62086 2378
rect 70298 2375 70310 2378
rect 62473 2329 70310 2375
rect 51370 2214 51382 2266
rect 51434 2263 51446 2266
rect 61898 2263 61910 2266
rect 51434 2217 61910 2263
rect 51434 2214 51446 2217
rect 61898 2214 61910 2217
rect 61962 2214 61974 2266
rect 62122 2214 62134 2266
rect 62186 2263 62198 2266
rect 62473 2263 62519 2329
rect 70298 2326 70310 2329
rect 70362 2326 70374 2378
rect 70522 2326 70534 2378
rect 70586 2375 70598 2378
rect 73434 2375 73446 2378
rect 70586 2329 73446 2375
rect 70586 2326 70598 2329
rect 73434 2326 73446 2329
rect 73498 2326 73510 2378
rect 76234 2375 76246 2378
rect 73896 2329 76246 2375
rect 62186 2217 62519 2263
rect 62186 2214 62198 2217
rect 62906 2214 62918 2266
rect 62970 2263 62982 2266
rect 73896 2263 73942 2329
rect 76234 2326 76246 2329
rect 76298 2326 76310 2378
rect 76458 2326 76470 2378
rect 76522 2375 76534 2378
rect 77802 2375 77814 2378
rect 76522 2329 77814 2375
rect 76522 2326 76534 2329
rect 77802 2326 77814 2329
rect 77866 2326 77878 2378
rect 78922 2326 78934 2378
rect 78986 2375 78998 2378
rect 81946 2375 81958 2378
rect 78986 2329 81958 2375
rect 78986 2326 78998 2329
rect 81946 2326 81958 2329
rect 82010 2326 82022 2378
rect 82170 2326 82182 2378
rect 82234 2375 82246 2378
rect 94154 2375 94166 2378
rect 82234 2329 94166 2375
rect 82234 2326 82246 2329
rect 94154 2326 94166 2329
rect 94218 2326 94230 2378
rect 100426 2375 100438 2378
rect 94281 2329 100438 2375
rect 62970 2217 73942 2263
rect 62970 2214 62982 2217
rect 73994 2214 74006 2266
rect 74058 2263 74070 2266
rect 75114 2263 75126 2266
rect 74058 2217 75126 2263
rect 74058 2214 74070 2217
rect 75114 2214 75126 2217
rect 75178 2214 75190 2266
rect 75241 2217 75735 2263
rect 49466 2102 49478 2154
rect 49530 2151 49542 2154
rect 59658 2151 59670 2154
rect 49530 2105 59670 2151
rect 49530 2102 49542 2105
rect 59658 2102 59670 2105
rect 59722 2102 59734 2154
rect 59882 2102 59894 2154
rect 59946 2151 59958 2154
rect 75241 2151 75287 2217
rect 59946 2105 75287 2151
rect 75689 2151 75735 2217
rect 75898 2214 75910 2266
rect 75962 2263 75974 2266
rect 83850 2263 83862 2266
rect 75962 2217 83862 2263
rect 75962 2214 75974 2217
rect 83850 2214 83862 2217
rect 83914 2214 83926 2266
rect 84186 2214 84198 2266
rect 84250 2263 84262 2266
rect 93930 2263 93942 2266
rect 84250 2217 93942 2263
rect 84250 2214 84262 2217
rect 93930 2214 93942 2217
rect 93994 2214 94006 2266
rect 94281 2263 94327 2329
rect 100426 2326 100438 2329
rect 100490 2326 100502 2378
rect 101546 2326 101558 2378
rect 101610 2375 101622 2378
rect 126410 2375 126422 2378
rect 101610 2329 126422 2375
rect 101610 2326 101622 2329
rect 126410 2326 126422 2329
rect 126474 2326 126486 2378
rect 94057 2217 94327 2263
rect 75689 2105 76071 2151
rect 59946 2102 59958 2105
rect 34906 1990 34918 2042
rect 34970 2039 34982 2042
rect 68170 2039 68182 2042
rect 34970 1993 68182 2039
rect 34970 1990 34982 1993
rect 68170 1990 68182 1993
rect 68234 1990 68246 2042
rect 68618 1990 68630 2042
rect 68682 2039 68694 2042
rect 75898 2039 75910 2042
rect 68682 1993 75910 2039
rect 68682 1990 68694 1993
rect 75898 1990 75910 1993
rect 75962 1990 75974 2042
rect 76025 2039 76071 2105
rect 76346 2102 76358 2154
rect 76410 2151 76422 2154
rect 83738 2151 83750 2154
rect 76410 2105 83750 2151
rect 76410 2102 76422 2105
rect 83738 2102 83750 2105
rect 83802 2102 83814 2154
rect 83962 2102 83974 2154
rect 84026 2151 84038 2154
rect 94057 2151 94103 2217
rect 95722 2214 95734 2266
rect 95786 2263 95798 2266
rect 125850 2263 125862 2266
rect 95786 2217 125862 2263
rect 95786 2214 95798 2217
rect 125850 2214 125862 2217
rect 125914 2214 125926 2266
rect 126649 2263 126695 2441
rect 126746 2326 126758 2378
rect 126810 2375 126822 2378
rect 134250 2375 134262 2378
rect 126810 2329 134262 2375
rect 126810 2326 126822 2329
rect 134250 2326 134262 2329
rect 134314 2326 134326 2378
rect 130890 2263 130902 2266
rect 126649 2217 130902 2263
rect 130890 2214 130902 2217
rect 130954 2214 130966 2266
rect 134377 2263 134423 2441
rect 138618 2438 138630 2490
rect 138682 2487 138694 2490
rect 152282 2487 152294 2490
rect 138682 2441 152294 2487
rect 138682 2438 138694 2441
rect 152282 2438 152294 2441
rect 152346 2438 152358 2490
rect 152618 2438 152630 2490
rect 152682 2487 152694 2490
rect 154186 2487 154198 2490
rect 152682 2441 154198 2487
rect 152682 2438 152694 2441
rect 154186 2438 154198 2441
rect 154250 2438 154262 2490
rect 154522 2438 154534 2490
rect 154586 2487 154598 2490
rect 204586 2487 204598 2490
rect 154586 2441 204598 2487
rect 154586 2438 154598 2441
rect 204586 2438 204598 2441
rect 204650 2438 204662 2490
rect 151274 2326 151286 2378
rect 151338 2375 151350 2378
rect 183082 2375 183094 2378
rect 151338 2329 183094 2375
rect 151338 2326 151350 2329
rect 183082 2326 183094 2329
rect 183146 2326 183158 2378
rect 185882 2326 185894 2378
rect 185946 2375 185958 2378
rect 190586 2375 190598 2378
rect 185946 2329 190598 2375
rect 185946 2326 185958 2329
rect 190586 2326 190598 2329
rect 190650 2326 190662 2378
rect 153850 2263 153862 2266
rect 134377 2217 153862 2263
rect 153850 2214 153862 2217
rect 153914 2214 153926 2266
rect 155642 2214 155654 2266
rect 155706 2263 155718 2266
rect 189354 2263 189366 2266
rect 155706 2217 189366 2263
rect 155706 2214 155718 2217
rect 189354 2214 189366 2217
rect 189418 2214 189430 2266
rect 95834 2151 95846 2154
rect 84026 2105 94103 2151
rect 94169 2105 95846 2151
rect 84026 2102 84038 2105
rect 88890 2039 88902 2042
rect 76025 1993 88902 2039
rect 88890 1990 88902 1993
rect 88954 1990 88966 2042
rect 89114 1990 89126 2042
rect 89178 2039 89190 2042
rect 89898 2039 89910 2042
rect 89178 1993 89910 2039
rect 89178 1990 89190 1993
rect 89898 1990 89910 1993
rect 89962 1990 89974 2042
rect 90682 1990 90694 2042
rect 90746 2039 90758 2042
rect 94169 2039 94215 2105
rect 95834 2102 95846 2105
rect 95898 2102 95910 2154
rect 96282 2102 96294 2154
rect 96346 2151 96358 2154
rect 101770 2151 101782 2154
rect 96346 2105 101782 2151
rect 96346 2102 96358 2105
rect 101770 2102 101782 2105
rect 101834 2102 101846 2154
rect 102554 2102 102566 2154
rect 102618 2151 102630 2154
rect 115434 2151 115446 2154
rect 102618 2105 115446 2151
rect 102618 2102 102630 2105
rect 115434 2102 115446 2105
rect 115498 2102 115510 2154
rect 115994 2102 116006 2154
rect 116058 2151 116070 2154
rect 117002 2151 117014 2154
rect 116058 2105 117014 2151
rect 116058 2102 116070 2105
rect 117002 2102 117014 2105
rect 117066 2102 117078 2154
rect 117226 2102 117238 2154
rect 117290 2151 117302 2154
rect 119354 2151 119366 2154
rect 117290 2105 119366 2151
rect 117290 2102 117302 2105
rect 119354 2102 119366 2105
rect 119418 2102 119430 2154
rect 119578 2102 119590 2154
rect 119642 2151 119654 2154
rect 126298 2151 126310 2154
rect 119642 2105 126310 2151
rect 119642 2102 119654 2105
rect 126298 2102 126310 2105
rect 126362 2102 126374 2154
rect 127642 2102 127654 2154
rect 127706 2151 127718 2154
rect 150266 2151 150278 2154
rect 127706 2105 150278 2151
rect 127706 2102 127718 2105
rect 150266 2102 150278 2105
rect 150330 2102 150342 2154
rect 154410 2102 154422 2154
rect 154474 2151 154486 2154
rect 188682 2151 188694 2154
rect 154474 2105 188694 2151
rect 154474 2102 154486 2105
rect 188682 2102 188694 2105
rect 188746 2102 188758 2154
rect 90746 1993 94215 2039
rect 90746 1990 90758 1993
rect 94490 1990 94502 2042
rect 94554 2039 94566 2042
rect 179050 2039 179062 2042
rect 94554 1993 102055 2039
rect 94554 1990 94566 1993
rect 61114 1878 61126 1930
rect 61178 1927 61190 1930
rect 62794 1927 62806 1930
rect 61178 1881 62806 1927
rect 61178 1878 61190 1881
rect 62794 1878 62806 1881
rect 62858 1878 62870 1930
rect 64698 1878 64710 1930
rect 64762 1927 64774 1930
rect 101098 1927 101110 1930
rect 64762 1881 101110 1927
rect 64762 1878 64774 1881
rect 101098 1878 101110 1881
rect 101162 1878 101174 1930
rect 102009 1927 102055 1993
rect 102233 1993 179062 2039
rect 102233 1927 102279 1993
rect 179050 1990 179062 1993
rect 179114 1990 179126 2042
rect 102009 1881 102279 1927
rect 102330 1878 102342 1930
rect 102394 1927 102406 1930
rect 151050 1927 151062 1930
rect 102394 1881 151062 1927
rect 102394 1878 102406 1881
rect 151050 1878 151062 1881
rect 151114 1878 151126 1930
rect 63578 1766 63590 1818
rect 63642 1815 63654 1818
rect 100650 1815 100662 1818
rect 63642 1769 100662 1815
rect 63642 1766 63654 1769
rect 100650 1766 100662 1769
rect 100714 1766 100726 1818
rect 100986 1766 100998 1818
rect 101050 1815 101062 1818
rect 102442 1815 102454 1818
rect 101050 1769 102454 1815
rect 101050 1766 101062 1769
rect 102442 1766 102454 1769
rect 102506 1766 102518 1818
rect 136378 1815 136390 1818
rect 102793 1769 136390 1815
rect 58090 1654 58102 1706
rect 58154 1703 58166 1706
rect 65146 1703 65158 1706
rect 58154 1657 65158 1703
rect 58154 1654 58166 1657
rect 65146 1654 65158 1657
rect 65210 1654 65222 1706
rect 65370 1654 65382 1706
rect 65434 1703 65446 1706
rect 100538 1703 100550 1706
rect 65434 1657 100550 1703
rect 65434 1654 65446 1657
rect 100538 1654 100550 1657
rect 100602 1654 100614 1706
rect 102793 1703 102839 1769
rect 136378 1766 136390 1769
rect 136442 1766 136454 1818
rect 155978 1766 155990 1818
rect 156042 1815 156054 1818
rect 156426 1815 156438 1818
rect 156042 1769 156438 1815
rect 156042 1766 156054 1769
rect 156426 1766 156438 1769
rect 156490 1766 156502 1818
rect 100665 1657 102839 1703
rect 32330 1542 32342 1594
rect 32394 1591 32406 1594
rect 75450 1591 75462 1594
rect 32394 1545 75462 1591
rect 32394 1542 32406 1545
rect 75450 1542 75462 1545
rect 75514 1542 75526 1594
rect 76794 1542 76806 1594
rect 76858 1591 76870 1594
rect 78250 1591 78262 1594
rect 76858 1545 78262 1591
rect 76858 1542 76870 1545
rect 78250 1542 78262 1545
rect 78314 1542 78326 1594
rect 78474 1542 78486 1594
rect 78538 1591 78550 1594
rect 82842 1591 82854 1594
rect 78538 1545 82854 1591
rect 78538 1542 78550 1545
rect 82842 1542 82854 1545
rect 82906 1542 82918 1594
rect 84746 1591 84758 1594
rect 83529 1545 84758 1591
rect 36362 1430 36374 1482
rect 36426 1479 36438 1482
rect 74778 1479 74790 1482
rect 36426 1433 74790 1479
rect 36426 1430 36438 1433
rect 74778 1430 74790 1433
rect 74842 1430 74854 1482
rect 75562 1430 75574 1482
rect 75626 1479 75638 1482
rect 83402 1479 83414 1482
rect 75626 1433 83414 1479
rect 75626 1430 75638 1433
rect 83402 1430 83414 1433
rect 83466 1430 83478 1482
rect 45994 1318 46006 1370
rect 46058 1367 46070 1370
rect 82058 1367 82070 1370
rect 46058 1321 82070 1367
rect 46058 1318 46070 1321
rect 82058 1318 82070 1321
rect 82122 1318 82134 1370
rect 82394 1318 82406 1370
rect 82458 1367 82470 1370
rect 82730 1367 82742 1370
rect 82458 1321 82742 1367
rect 82458 1318 82470 1321
rect 82730 1318 82742 1321
rect 82794 1367 82806 1370
rect 83529 1367 83575 1545
rect 84746 1542 84758 1545
rect 84810 1542 84822 1594
rect 85082 1542 85094 1594
rect 85146 1591 85158 1594
rect 88442 1591 88454 1594
rect 85146 1545 88454 1591
rect 85146 1542 85158 1545
rect 88442 1542 88454 1545
rect 88506 1542 88518 1594
rect 88778 1542 88790 1594
rect 88842 1591 88854 1594
rect 92138 1591 92150 1594
rect 88842 1545 92150 1591
rect 88842 1542 88854 1545
rect 92138 1542 92150 1545
rect 92202 1542 92214 1594
rect 92362 1542 92374 1594
rect 92426 1591 92438 1594
rect 97626 1591 97638 1594
rect 92426 1545 97638 1591
rect 92426 1542 92438 1545
rect 97626 1542 97638 1545
rect 97690 1542 97702 1594
rect 98298 1542 98310 1594
rect 98362 1591 98374 1594
rect 100314 1591 100326 1594
rect 98362 1545 100326 1591
rect 98362 1542 98374 1545
rect 100314 1542 100326 1545
rect 100378 1542 100390 1594
rect 83962 1430 83974 1482
rect 84026 1479 84038 1482
rect 100665 1479 100711 1657
rect 102890 1654 102902 1706
rect 102954 1703 102966 1706
rect 102954 1657 107431 1703
rect 102954 1654 102966 1657
rect 100762 1542 100774 1594
rect 100826 1591 100838 1594
rect 101770 1591 101782 1594
rect 100826 1545 101782 1591
rect 100826 1542 100838 1545
rect 101770 1542 101782 1545
rect 101834 1542 101846 1594
rect 101994 1542 102006 1594
rect 102058 1591 102070 1594
rect 105242 1591 105254 1594
rect 102058 1545 105254 1591
rect 102058 1542 102070 1545
rect 105242 1542 105254 1545
rect 105306 1542 105318 1594
rect 105914 1542 105926 1594
rect 105978 1591 105990 1594
rect 106922 1591 106934 1594
rect 105978 1545 106934 1591
rect 105978 1542 105990 1545
rect 106922 1542 106934 1545
rect 106986 1542 106998 1594
rect 107385 1591 107431 1657
rect 107482 1654 107494 1706
rect 107546 1703 107558 1706
rect 108154 1703 108166 1706
rect 107546 1657 108166 1703
rect 107546 1654 107558 1657
rect 108154 1654 108166 1657
rect 108218 1654 108230 1706
rect 150266 1703 150278 1706
rect 108281 1657 150278 1703
rect 108281 1591 108327 1657
rect 150266 1654 150278 1657
rect 150330 1654 150342 1706
rect 107385 1545 108327 1591
rect 108378 1542 108390 1594
rect 108442 1591 108454 1594
rect 109946 1591 109958 1594
rect 108442 1545 109958 1591
rect 108442 1542 108454 1545
rect 109946 1542 109958 1545
rect 110010 1542 110022 1594
rect 112634 1591 112646 1594
rect 110073 1545 112646 1591
rect 106698 1479 106710 1482
rect 84026 1433 100711 1479
rect 100777 1433 106710 1479
rect 84026 1430 84038 1433
rect 82794 1321 83575 1367
rect 82794 1318 82806 1321
rect 84410 1318 84422 1370
rect 84474 1367 84486 1370
rect 90570 1367 90582 1370
rect 84474 1321 90582 1367
rect 84474 1318 84486 1321
rect 90570 1318 90582 1321
rect 90634 1318 90646 1370
rect 91242 1318 91254 1370
rect 91306 1367 91318 1370
rect 94602 1367 94614 1370
rect 91306 1321 94614 1367
rect 91306 1318 91318 1321
rect 94602 1318 94614 1321
rect 94666 1318 94678 1370
rect 97402 1318 97414 1370
rect 97466 1367 97478 1370
rect 100777 1367 100823 1433
rect 106698 1430 106710 1433
rect 106762 1430 106774 1482
rect 109722 1430 109734 1482
rect 109786 1479 109798 1482
rect 110073 1479 110119 1545
rect 112634 1542 112646 1545
rect 112698 1542 112710 1594
rect 112858 1542 112870 1594
rect 112922 1591 112934 1594
rect 112922 1545 117511 1591
rect 112922 1542 112934 1545
rect 117338 1479 117350 1482
rect 109786 1433 110119 1479
rect 111305 1433 117350 1479
rect 109786 1430 109798 1433
rect 97466 1321 100823 1367
rect 97466 1318 97478 1321
rect 100874 1318 100886 1370
rect 100938 1367 100950 1370
rect 111305 1367 111351 1433
rect 117338 1430 117350 1433
rect 117402 1430 117414 1482
rect 117465 1479 117511 1545
rect 118010 1542 118022 1594
rect 118074 1591 118086 1594
rect 120250 1591 120262 1594
rect 118074 1545 120262 1591
rect 118074 1542 118086 1545
rect 120250 1542 120262 1545
rect 120314 1542 120326 1594
rect 120474 1542 120486 1594
rect 120538 1591 120550 1594
rect 123386 1591 123398 1594
rect 120538 1545 123398 1591
rect 120538 1542 120550 1545
rect 123386 1542 123398 1545
rect 123450 1542 123462 1594
rect 123610 1542 123622 1594
rect 123674 1591 123686 1594
rect 132458 1591 132470 1594
rect 123674 1545 132470 1591
rect 123674 1542 123686 1545
rect 132458 1542 132470 1545
rect 132522 1542 132534 1594
rect 144778 1542 144790 1594
rect 144842 1591 144854 1594
rect 147466 1591 147478 1594
rect 144842 1545 147478 1591
rect 144842 1542 144854 1545
rect 147466 1542 147478 1545
rect 147530 1542 147542 1594
rect 118122 1479 118134 1482
rect 117465 1433 118134 1479
rect 118122 1430 118134 1433
rect 118186 1430 118198 1482
rect 119802 1430 119814 1482
rect 119866 1479 119878 1482
rect 136490 1479 136502 1482
rect 119866 1433 136502 1479
rect 119866 1430 119878 1433
rect 136490 1430 136502 1433
rect 136554 1430 136566 1482
rect 100938 1321 111351 1367
rect 100938 1318 100950 1321
rect 111402 1318 111414 1370
rect 111466 1367 111478 1370
rect 116666 1367 116678 1370
rect 111466 1321 116678 1367
rect 111466 1318 111478 1321
rect 116666 1318 116678 1321
rect 116730 1318 116742 1370
rect 117002 1318 117014 1370
rect 117066 1367 117078 1370
rect 119466 1367 119478 1370
rect 117066 1321 119478 1367
rect 117066 1318 117078 1321
rect 119466 1318 119478 1321
rect 119530 1318 119542 1370
rect 119690 1318 119702 1370
rect 119754 1367 119766 1370
rect 120474 1367 120486 1370
rect 119754 1321 120486 1367
rect 119754 1318 119766 1321
rect 120474 1318 120486 1321
rect 120538 1318 120550 1370
rect 120698 1318 120710 1370
rect 120762 1367 120774 1370
rect 121594 1367 121606 1370
rect 120762 1321 121606 1367
rect 120762 1318 120774 1321
rect 121594 1318 121606 1321
rect 121658 1318 121670 1370
rect 122938 1318 122950 1370
rect 123002 1367 123014 1370
rect 135034 1367 135046 1370
rect 123002 1321 135046 1367
rect 123002 1318 123014 1321
rect 135034 1318 135046 1321
rect 135098 1318 135110 1370
rect 44762 1206 44774 1258
rect 44826 1255 44838 1258
rect 69962 1255 69974 1258
rect 44826 1209 69974 1255
rect 44826 1206 44838 1209
rect 69962 1206 69974 1209
rect 70026 1206 70038 1258
rect 70522 1206 70534 1258
rect 70586 1255 70598 1258
rect 70586 1209 132742 1255
rect 70586 1206 70598 1209
rect 10154 1094 10166 1146
rect 10218 1143 10230 1146
rect 71978 1143 71990 1146
rect 10218 1097 71990 1143
rect 10218 1094 10230 1097
rect 71978 1094 71990 1097
rect 72042 1094 72054 1146
rect 75114 1094 75126 1146
rect 75178 1143 75190 1146
rect 81722 1143 81734 1146
rect 75178 1097 81734 1143
rect 75178 1094 75190 1097
rect 81722 1094 81734 1097
rect 81786 1094 81798 1146
rect 81946 1094 81958 1146
rect 82010 1143 82022 1146
rect 84074 1143 84086 1146
rect 82010 1097 84086 1143
rect 82010 1094 82022 1097
rect 84074 1094 84086 1097
rect 84138 1094 84150 1146
rect 85418 1094 85430 1146
rect 85482 1143 85494 1146
rect 86762 1143 86774 1146
rect 85482 1097 86774 1143
rect 85482 1094 85494 1097
rect 86762 1094 86774 1097
rect 86826 1094 86838 1146
rect 87210 1094 87222 1146
rect 87274 1143 87286 1146
rect 87434 1143 87446 1146
rect 87274 1097 87446 1143
rect 87274 1094 87286 1097
rect 87434 1094 87446 1097
rect 87498 1094 87510 1146
rect 87882 1094 87894 1146
rect 87946 1143 87958 1146
rect 89674 1143 89686 1146
rect 87946 1097 89686 1143
rect 87946 1094 87958 1097
rect 89674 1094 89686 1097
rect 89738 1094 89750 1146
rect 89898 1094 89910 1146
rect 89962 1143 89974 1146
rect 97962 1143 97974 1146
rect 89962 1097 97974 1143
rect 89962 1094 89974 1097
rect 97962 1094 97974 1097
rect 98026 1094 98038 1146
rect 100762 1094 100774 1146
rect 100826 1143 100838 1146
rect 101434 1143 101446 1146
rect 100826 1097 101446 1143
rect 100826 1094 100838 1097
rect 101434 1094 101446 1097
rect 101498 1094 101510 1146
rect 101770 1094 101782 1146
rect 101834 1143 101846 1146
rect 110282 1143 110294 1146
rect 101834 1097 110294 1143
rect 101834 1094 101846 1097
rect 110282 1094 110294 1097
rect 110346 1094 110358 1146
rect 111066 1094 111078 1146
rect 111130 1143 111142 1146
rect 111850 1143 111862 1146
rect 111130 1097 111862 1143
rect 111130 1094 111142 1097
rect 111850 1094 111862 1097
rect 111914 1094 111926 1146
rect 112074 1094 112086 1146
rect 112138 1143 112150 1146
rect 114650 1143 114662 1146
rect 112138 1097 114662 1143
rect 112138 1094 112150 1097
rect 114650 1094 114662 1097
rect 114714 1094 114726 1146
rect 117898 1143 117910 1146
rect 114777 1097 117910 1143
rect 42522 982 42534 1034
rect 42586 1031 42598 1034
rect 74890 1031 74902 1034
rect 42586 985 74902 1031
rect 42586 982 42598 985
rect 74890 982 74902 985
rect 74954 982 74966 1034
rect 75226 982 75238 1034
rect 75290 1031 75302 1034
rect 77242 1031 77254 1034
rect 75290 985 77254 1031
rect 75290 982 75302 985
rect 77242 982 77254 985
rect 77306 982 77318 1034
rect 81274 1031 81286 1034
rect 77817 985 81286 1031
rect 5562 870 5574 922
rect 5626 870 5638 922
rect 13514 870 13526 922
rect 13578 919 13590 922
rect 37258 919 37270 922
rect 13578 873 37270 919
rect 13578 870 13590 873
rect 37258 870 37270 873
rect 37322 870 37334 922
rect 43418 870 43430 922
rect 43482 870 43494 922
rect 63690 870 63702 922
rect 63754 870 63766 922
rect 63914 870 63926 922
rect 63978 919 63990 922
rect 68954 919 68966 922
rect 63978 873 68966 919
rect 63978 870 63990 873
rect 68954 870 68966 873
rect 69018 870 69030 922
rect 71418 870 71430 922
rect 71482 919 71494 922
rect 77817 919 77863 985
rect 81274 982 81286 985
rect 81338 982 81350 1034
rect 81498 982 81510 1034
rect 81562 1031 81574 1034
rect 82730 1031 82742 1034
rect 81562 985 82742 1031
rect 81562 982 81574 985
rect 82730 982 82742 985
rect 82794 982 82806 1034
rect 83514 982 83526 1034
rect 83578 1031 83590 1034
rect 84858 1031 84870 1034
rect 83578 985 84870 1031
rect 83578 982 83590 985
rect 84858 982 84870 985
rect 84922 982 84934 1034
rect 86986 982 86998 1034
rect 87050 1031 87062 1034
rect 92138 1031 92150 1034
rect 87050 985 92150 1031
rect 87050 982 87062 985
rect 92138 982 92150 985
rect 92202 1031 92214 1034
rect 96618 1031 96630 1034
rect 92202 985 96630 1031
rect 92202 982 92214 985
rect 96618 982 96630 985
rect 96682 982 96694 1034
rect 96842 982 96854 1034
rect 96906 1031 96918 1034
rect 96906 985 98695 1031
rect 96906 982 96918 985
rect 71482 873 77863 919
rect 71482 870 71494 873
rect 77914 870 77926 922
rect 77978 919 77990 922
rect 88218 919 88230 922
rect 77978 873 88230 919
rect 77978 870 77990 873
rect 88218 870 88230 873
rect 88282 870 88294 922
rect 88442 870 88454 922
rect 88506 919 88518 922
rect 90346 919 90358 922
rect 88506 873 90358 919
rect 88506 870 88518 873
rect 90346 870 90358 873
rect 90410 919 90422 922
rect 98522 919 98534 922
rect 90410 873 98534 919
rect 90410 870 90422 873
rect 98522 870 98534 873
rect 98586 870 98598 922
rect 98649 919 98695 985
rect 99418 982 99430 1034
rect 99482 1031 99494 1034
rect 106138 1031 106150 1034
rect 99482 985 106150 1031
rect 99482 982 99494 985
rect 106138 982 106150 985
rect 106202 982 106214 1034
rect 106362 982 106374 1034
rect 106426 1031 106438 1034
rect 106426 985 110679 1031
rect 106426 982 106438 985
rect 99866 919 99878 922
rect 98649 873 99878 919
rect 99866 870 99878 873
rect 99930 870 99942 922
rect 100986 870 100998 922
rect 101050 919 101062 922
rect 109722 919 109734 922
rect 101050 873 109734 919
rect 101050 870 101062 873
rect 109722 870 109734 873
rect 109786 870 109798 922
rect 110633 919 110679 985
rect 110730 982 110742 1034
rect 110794 1031 110806 1034
rect 111626 1031 111638 1034
rect 110794 985 111638 1031
rect 110794 982 110806 985
rect 111626 982 111638 985
rect 111690 982 111702 1034
rect 112634 982 112646 1034
rect 112698 1031 112710 1034
rect 114777 1031 114823 1097
rect 117898 1094 117910 1097
rect 117962 1094 117974 1146
rect 118458 1094 118470 1146
rect 118522 1143 118534 1146
rect 121258 1143 121270 1146
rect 118522 1097 121270 1143
rect 118522 1094 118534 1097
rect 121258 1094 121270 1097
rect 121322 1094 121334 1146
rect 121706 1094 121718 1146
rect 121770 1143 121782 1146
rect 125290 1143 125302 1146
rect 121770 1097 125302 1143
rect 121770 1094 121782 1097
rect 125290 1094 125302 1097
rect 125354 1094 125366 1146
rect 125514 1094 125526 1146
rect 125578 1143 125590 1146
rect 126298 1143 126310 1146
rect 125578 1097 126310 1143
rect 125578 1094 125590 1097
rect 126298 1094 126310 1097
rect 126362 1094 126374 1146
rect 132696 1143 132742 1209
rect 202570 1143 202582 1146
rect 132696 1097 202582 1143
rect 202570 1094 202582 1097
rect 202634 1094 202646 1146
rect 112698 985 114823 1031
rect 112698 982 112710 985
rect 114874 982 114886 1034
rect 114938 1031 114950 1034
rect 116442 1031 116454 1034
rect 114938 985 116454 1031
rect 114938 982 114950 985
rect 116442 982 116454 985
rect 116506 982 116518 1034
rect 116778 982 116790 1034
rect 116842 1031 116854 1034
rect 129994 1031 130006 1034
rect 116842 985 130006 1031
rect 116842 982 116854 985
rect 129994 982 130006 985
rect 130058 982 130070 1034
rect 133914 982 133926 1034
rect 133978 1031 133990 1034
rect 193386 1031 193398 1034
rect 133978 985 193398 1031
rect 133978 982 133990 985
rect 193386 982 193398 985
rect 193450 982 193462 1034
rect 116106 919 116118 922
rect 110633 873 116118 919
rect 116106 870 116118 873
rect 116170 870 116182 922
rect 118234 870 118246 922
rect 118298 919 118310 922
rect 218362 919 218374 922
rect 118298 873 218374 919
rect 118298 870 118310 873
rect 218362 870 218374 873
rect 218426 870 218438 922
rect 5577 807 5623 870
rect 28970 807 28982 810
rect 5577 761 28982 807
rect 28970 758 28982 761
rect 29034 758 29046 810
rect 16202 646 16214 698
rect 16266 695 16278 698
rect 43433 695 43479 870
rect 16266 649 43479 695
rect 16266 646 16278 649
rect 7242 534 7254 586
rect 7306 583 7318 586
rect 33898 583 33910 586
rect 7306 537 33910 583
rect 7306 534 7318 537
rect 33898 534 33910 537
rect 33962 534 33974 586
rect 63705 583 63751 870
rect 69962 758 69974 810
rect 70026 807 70038 810
rect 76122 807 76134 810
rect 70026 761 76134 807
rect 70026 758 70038 761
rect 76122 758 76134 761
rect 76186 758 76198 810
rect 76682 758 76694 810
rect 76746 807 76758 810
rect 77130 807 77142 810
rect 76746 761 77142 807
rect 76746 758 76758 761
rect 77130 758 77142 761
rect 77194 758 77206 810
rect 77354 758 77366 810
rect 77418 807 77430 810
rect 81498 807 81510 810
rect 77418 761 81510 807
rect 77418 758 77430 761
rect 81498 758 81510 761
rect 81562 758 81574 810
rect 82058 807 82070 810
rect 81625 761 82070 807
rect 70410 646 70422 698
rect 70474 695 70486 698
rect 77914 695 77926 698
rect 70474 649 77926 695
rect 70474 646 70486 649
rect 77914 646 77926 649
rect 77978 646 77990 698
rect 78362 646 78374 698
rect 78426 695 78438 698
rect 81625 695 81671 761
rect 82058 758 82070 761
rect 82122 758 82134 810
rect 82730 758 82742 810
rect 82794 807 82806 810
rect 82794 761 83351 807
rect 82794 758 82806 761
rect 83305 695 83351 761
rect 83850 758 83862 810
rect 83914 807 83926 810
rect 83914 761 85479 807
rect 83914 758 83926 761
rect 85306 695 85318 698
rect 78426 649 81671 695
rect 81737 649 83183 695
rect 83305 649 85318 695
rect 78426 646 78438 649
rect 81737 583 81783 649
rect 63705 537 81783 583
rect 82058 534 82070 586
rect 82122 583 82134 586
rect 83137 583 83183 649
rect 85306 646 85318 649
rect 85370 646 85382 698
rect 85433 695 85479 761
rect 85754 758 85766 810
rect 85818 807 85830 810
rect 196186 807 196198 810
rect 85818 761 196198 807
rect 85818 758 85830 761
rect 196186 758 196198 761
rect 196250 758 196262 810
rect 215674 807 215686 810
rect 203256 761 215686 807
rect 203256 695 203302 761
rect 215674 758 215686 761
rect 215738 758 215750 810
rect 85433 649 203302 695
rect 195402 583 195414 586
rect 82122 537 83071 583
rect 83137 537 195414 583
rect 82122 534 82134 537
rect 8922 422 8934 474
rect 8986 471 8998 474
rect 42522 471 42534 474
rect 8986 425 42534 471
rect 8986 422 8998 425
rect 42522 422 42534 425
rect 42586 422 42598 474
rect 49914 422 49926 474
rect 49978 471 49990 474
rect 68730 471 68742 474
rect 49978 425 68742 471
rect 49978 422 49990 425
rect 68730 422 68742 425
rect 68794 422 68806 474
rect 69290 422 69302 474
rect 69354 471 69366 474
rect 81386 471 81398 474
rect 69354 425 81398 471
rect 69354 422 69366 425
rect 81386 422 81398 425
rect 81450 422 81462 474
rect 83025 471 83071 537
rect 195402 534 195414 537
rect 195466 534 195478 586
rect 216122 471 216134 474
rect 81513 425 82959 471
rect 83025 425 216134 471
rect 24266 310 24278 362
rect 24330 359 24342 362
rect 73546 359 73558 362
rect 24330 313 73558 359
rect 24330 310 24342 313
rect 73546 310 73558 313
rect 73610 310 73622 362
rect 74890 310 74902 362
rect 74954 359 74966 362
rect 81513 359 81559 425
rect 74954 313 81559 359
rect 82913 359 82959 425
rect 216122 422 216134 425
rect 216186 422 216198 474
rect 207050 359 207062 362
rect 82913 313 207062 359
rect 74954 310 74966 313
rect 207050 310 207062 313
rect 207114 310 207126 362
rect 21298 198 21310 250
rect 21362 247 21374 250
rect 66826 247 66838 250
rect 21362 201 66838 247
rect 21362 198 21374 201
rect 66826 198 66838 201
rect 66890 198 66902 250
rect 68842 198 68854 250
rect 68906 247 68918 250
rect 77354 247 77366 250
rect 68906 201 77366 247
rect 68906 198 68918 201
rect 77354 198 77366 201
rect 77418 198 77430 250
rect 77802 198 77814 250
rect 77866 247 77878 250
rect 83850 247 83862 250
rect 77866 201 83862 247
rect 77866 198 77878 201
rect 83850 198 83862 201
rect 83914 198 83926 250
rect 84074 198 84086 250
rect 84138 247 84150 250
rect 215002 247 215014 250
rect 84138 201 215014 247
rect 84138 198 84150 201
rect 215002 198 215014 201
rect 215066 198 215078 250
rect 17602 86 17614 138
rect 17666 135 17678 138
rect 54730 135 54742 138
rect 17666 89 54742 135
rect 17666 86 17678 89
rect 54730 86 54742 89
rect 54794 86 54806 138
rect 56522 86 56534 138
rect 56586 135 56598 138
rect 208282 135 208294 138
rect 56586 89 208294 135
rect 56586 86 56598 89
rect 208282 86 208294 89
rect 208346 86 208358 138
<< via1 >>
rect 11622 14870 11674 14922
rect 63254 14870 63306 14922
rect 68406 14758 68458 14810
rect 73334 14870 73386 14922
rect 79494 14870 79546 14922
rect 80726 14870 80778 14922
rect 103238 14870 103290 14922
rect 9494 14646 9546 14698
rect 63142 14646 63194 14698
rect 64038 14646 64090 14698
rect 73334 14646 73386 14698
rect 73558 14646 73610 14698
rect 78710 14646 78762 14698
rect 10054 14534 10106 14586
rect 79270 14646 79322 14698
rect 79942 14646 79994 14698
rect 80166 14646 80218 14698
rect 80726 14646 80778 14698
rect 80950 14646 81002 14698
rect 82854 14646 82906 14698
rect 83078 14646 83130 14698
rect 84422 14646 84474 14698
rect 84982 14646 85034 14698
rect 90806 14646 90858 14698
rect 91030 14646 91082 14698
rect 102678 14646 102730 14698
rect 104022 14758 104074 14810
rect 104806 14870 104858 14922
rect 115670 14646 115722 14698
rect 51046 14422 51098 14474
rect 74902 14422 74954 14474
rect 75574 14422 75626 14474
rect 79494 14534 79546 14586
rect 81510 14534 81562 14586
rect 79382 14422 79434 14474
rect 103910 14534 103962 14586
rect 104694 14534 104746 14586
rect 113430 14534 113482 14586
rect 8486 14310 8538 14362
rect 53062 14198 53114 14250
rect 73558 14198 73610 14250
rect 1878 14086 1930 14138
rect 57542 14086 57594 14138
rect 61686 14086 61738 14138
rect 64150 14086 64202 14138
rect 65942 14086 65994 14138
rect 80726 14198 80778 14250
rect 80950 14310 81002 14362
rect 83078 14310 83130 14362
rect 84534 14310 84586 14362
rect 91590 14310 91642 14362
rect 98310 14422 98362 14474
rect 102006 14310 102058 14362
rect 74006 14086 74058 14138
rect 75574 14086 75626 14138
rect 76918 14086 76970 14138
rect 77366 14086 77418 14138
rect 77590 14086 77642 14138
rect 78038 14086 78090 14138
rect 78374 14086 78426 14138
rect 78822 14086 78874 14138
rect 79046 14086 79098 14138
rect 45446 13974 45498 14026
rect 64038 13974 64090 14026
rect 64486 13974 64538 14026
rect 70422 13974 70474 14026
rect 71654 13974 71706 14026
rect 74678 13974 74730 14026
rect 75014 13974 75066 14026
rect 80502 14086 80554 14138
rect 81734 14086 81786 14138
rect 82182 14086 82234 14138
rect 88230 14198 88282 14250
rect 88678 14198 88730 14250
rect 100998 14198 101050 14250
rect 102566 14422 102618 14474
rect 102454 14310 102506 14362
rect 102678 14198 102730 14250
rect 104246 14310 104298 14362
rect 114886 14422 114938 14474
rect 114998 14310 115050 14362
rect 115894 14758 115946 14810
rect 120262 14758 120314 14810
rect 121046 14870 121098 14922
rect 127430 14870 127482 14922
rect 131126 14870 131178 14922
rect 148598 14870 148650 14922
rect 121494 14758 121546 14810
rect 122502 14758 122554 14810
rect 151510 14758 151562 14810
rect 116342 14646 116394 14698
rect 148374 14646 148426 14698
rect 116566 14534 116618 14586
rect 116678 14422 116730 14474
rect 117126 14422 117178 14474
rect 138966 14534 139018 14586
rect 167526 14534 167578 14586
rect 118806 14310 118858 14362
rect 120710 14310 120762 14362
rect 121606 14310 121658 14362
rect 136278 14310 136330 14362
rect 149830 14422 149882 14474
rect 141094 14310 141146 14362
rect 147926 14310 147978 14362
rect 114214 14198 114266 14250
rect 116342 14198 116394 14250
rect 43654 13862 43706 13914
rect 75126 13862 75178 13914
rect 80838 13974 80890 14026
rect 81062 13974 81114 14026
rect 83750 14086 83802 14138
rect 84310 14086 84362 14138
rect 91030 14086 91082 14138
rect 83526 13974 83578 14026
rect 87222 13974 87274 14026
rect 88230 13974 88282 14026
rect 90022 13974 90074 14026
rect 92710 14086 92762 14138
rect 92934 14086 92986 14138
rect 97526 14086 97578 14138
rect 98086 14086 98138 14138
rect 99206 14086 99258 14138
rect 99430 14086 99482 14138
rect 116678 14086 116730 14138
rect 117350 14086 117402 14138
rect 118694 14198 118746 14250
rect 148710 14198 148762 14250
rect 149270 14198 149322 14250
rect 119254 14086 119306 14138
rect 149382 14086 149434 14138
rect 91590 13974 91642 14026
rect 102566 13974 102618 14026
rect 103910 13974 103962 14026
rect 111190 13974 111242 14026
rect 111974 13974 112026 14026
rect 112982 13974 113034 14026
rect 113430 13974 113482 14026
rect 114214 13974 114266 14026
rect 114998 13974 115050 14026
rect 120038 13974 120090 14026
rect 47574 13750 47626 13802
rect 75462 13750 75514 13802
rect 6806 13638 6858 13690
rect 55750 13638 55802 13690
rect 58214 13638 58266 13690
rect 75686 13750 75738 13802
rect 79606 13750 79658 13802
rect 82518 13750 82570 13802
rect 75798 13638 75850 13690
rect 82070 13638 82122 13690
rect 54406 13526 54458 13578
rect 82406 13638 82458 13690
rect 82742 13750 82794 13802
rect 82966 13750 83018 13802
rect 84310 13750 84362 13802
rect 84534 13750 84586 13802
rect 117126 13862 117178 13914
rect 117350 13862 117402 13914
rect 119926 13862 119978 13914
rect 134150 13974 134202 14026
rect 138518 13974 138570 14026
rect 176374 14086 176426 14138
rect 196422 14086 196474 14138
rect 197206 13974 197258 14026
rect 82854 13526 82906 13578
rect 90134 13526 90186 13578
rect 90358 13526 90410 13578
rect 100550 13638 100602 13690
rect 100998 13750 101050 13802
rect 101334 13750 101386 13802
rect 101782 13750 101834 13802
rect 102118 13750 102170 13802
rect 102454 13638 102506 13690
rect 104582 13750 104634 13802
rect 119366 13750 119418 13802
rect 119590 13750 119642 13802
rect 121046 13862 121098 13914
rect 122502 13862 122554 13914
rect 122950 13862 123002 13914
rect 125974 13862 126026 13914
rect 126198 13862 126250 13914
rect 134262 13862 134314 13914
rect 134710 13862 134762 13914
rect 142886 13862 142938 13914
rect 143222 13862 143274 13914
rect 212774 13862 212826 13914
rect 120262 13750 120314 13802
rect 91030 13526 91082 13578
rect 103462 13638 103514 13690
rect 118470 13638 118522 13690
rect 118694 13638 118746 13690
rect 116230 13526 116282 13578
rect 116454 13526 116506 13578
rect 138518 13526 138570 13578
rect 53846 13414 53898 13466
rect 75798 13414 75850 13466
rect 76022 13414 76074 13466
rect 49814 13302 49866 13354
rect 55974 13190 56026 13242
rect 86 13078 138 13130
rect 67510 13078 67562 13130
rect 41078 12966 41130 13018
rect 67846 12966 67898 13018
rect 68406 13190 68458 13242
rect 79046 13190 79098 13242
rect 79606 13190 79658 13242
rect 80838 13190 80890 13242
rect 81174 13190 81226 13242
rect 81734 13190 81786 13242
rect 68070 13078 68122 13130
rect 80726 13078 80778 13130
rect 73782 12966 73834 13018
rect 43206 12854 43258 12906
rect 68070 12854 68122 12906
rect 69974 12854 70026 12906
rect 74454 12966 74506 13018
rect 75126 12966 75178 13018
rect 78710 12966 78762 13018
rect 78934 12966 78986 13018
rect 82182 13078 82234 13130
rect 83190 13414 83242 13466
rect 90246 13414 90298 13466
rect 90806 13414 90858 13466
rect 103350 13414 103402 13466
rect 104134 13414 104186 13466
rect 139078 13526 139130 13578
rect 139526 13526 139578 13578
rect 143222 13526 143274 13578
rect 138742 13414 138794 13466
rect 140646 13414 140698 13466
rect 149158 13750 149210 13802
rect 153190 13750 153242 13802
rect 159238 13750 159290 13802
rect 178278 13750 178330 13802
rect 149382 13638 149434 13690
rect 210422 13638 210474 13690
rect 148374 13414 148426 13466
rect 161254 13526 161306 13578
rect 182534 13526 182586 13578
rect 184550 13414 184602 13466
rect 82742 13302 82794 13354
rect 84198 13302 84250 13354
rect 84422 13302 84474 13354
rect 103238 13190 103290 13242
rect 82742 13078 82794 13130
rect 101110 13078 101162 13130
rect 102566 13078 102618 13130
rect 114662 13190 114714 13242
rect 115222 13302 115274 13354
rect 149158 13302 149210 13354
rect 149382 13302 149434 13354
rect 211654 13302 211706 13354
rect 138966 13190 139018 13242
rect 144454 13190 144506 13242
rect 149494 13190 149546 13242
rect 151062 13190 151114 13242
rect 155318 13190 155370 13242
rect 165062 13190 165114 13242
rect 173686 13190 173738 13242
rect 103462 13078 103514 13130
rect 120598 13078 120650 13130
rect 120822 13078 120874 13130
rect 126198 13078 126250 13130
rect 126758 13078 126810 13130
rect 142662 13078 142714 13130
rect 149270 13078 149322 13130
rect 185894 13078 185946 13130
rect 74006 12854 74058 12906
rect 77366 12854 77418 12906
rect 77814 12854 77866 12906
rect 81958 12854 82010 12906
rect 99430 12966 99482 13018
rect 88454 12854 88506 12906
rect 88678 12854 88730 12906
rect 89462 12854 89514 12906
rect 89798 12854 89850 12906
rect 102790 12966 102842 13018
rect 103014 12966 103066 13018
rect 103798 12966 103850 13018
rect 104022 12966 104074 13018
rect 117238 12966 117290 13018
rect 117462 12966 117514 13018
rect 122278 12966 122330 13018
rect 122502 12966 122554 13018
rect 138182 12966 138234 13018
rect 138406 12966 138458 13018
rect 142326 12966 142378 13018
rect 148598 12966 148650 13018
rect 186566 12966 186618 13018
rect 99654 12854 99706 12906
rect 102342 12854 102394 12906
rect 102566 12854 102618 12906
rect 102902 12854 102954 12906
rect 5350 12742 5402 12794
rect 56982 12742 57034 12794
rect 58550 12742 58602 12794
rect 82406 12742 82458 12794
rect 104806 12854 104858 12906
rect 109174 12854 109226 12906
rect 109846 12854 109898 12906
rect 110854 12854 110906 12906
rect 114438 12854 114490 12906
rect 114662 12854 114714 12906
rect 121606 12854 121658 12906
rect 125862 12854 125914 12906
rect 126758 12854 126810 12906
rect 127430 12854 127482 12906
rect 149046 12854 149098 12906
rect 149270 12854 149322 12906
rect 188470 12854 188522 12906
rect 103126 12742 103178 12794
rect 114550 12742 114602 12794
rect 29430 12630 29482 12682
rect 71766 12630 71818 12682
rect 71990 12630 72042 12682
rect 76806 12630 76858 12682
rect 56422 12518 56474 12570
rect 78710 12630 78762 12682
rect 80614 12630 80666 12682
rect 80838 12630 80890 12682
rect 81398 12630 81450 12682
rect 84534 12630 84586 12682
rect 84870 12630 84922 12682
rect 102678 12630 102730 12682
rect 51942 12406 51994 12458
rect 54182 12294 54234 12346
rect 75238 12294 75290 12346
rect 77926 12406 77978 12458
rect 79942 12406 79994 12458
rect 80614 12406 80666 12458
rect 81062 12406 81114 12458
rect 82294 12518 82346 12570
rect 83078 12518 83130 12570
rect 87894 12518 87946 12570
rect 103574 12630 103626 12682
rect 4678 12182 4730 12234
rect 64486 12182 64538 12234
rect 67734 12182 67786 12234
rect 69638 12182 69690 12234
rect 69862 12182 69914 12234
rect 78262 12294 78314 12346
rect 76694 12182 76746 12234
rect 78374 12182 78426 12234
rect 78598 12294 78650 12346
rect 80278 12294 80330 12346
rect 81734 12406 81786 12458
rect 89798 12406 89850 12458
rect 102902 12518 102954 12570
rect 114998 12630 115050 12682
rect 115558 12742 115610 12794
rect 142662 12742 142714 12794
rect 142886 12742 142938 12794
rect 188582 12742 188634 12794
rect 138406 12630 138458 12682
rect 139078 12630 139130 12682
rect 189814 12630 189866 12682
rect 104134 12518 104186 12570
rect 114886 12518 114938 12570
rect 116566 12518 116618 12570
rect 119590 12518 119642 12570
rect 119926 12518 119978 12570
rect 120822 12518 120874 12570
rect 20694 12070 20746 12122
rect 63702 12070 63754 12122
rect 65158 12070 65210 12122
rect 80726 12182 80778 12234
rect 81958 12182 82010 12234
rect 116790 12406 116842 12458
rect 118470 12406 118522 12458
rect 118694 12406 118746 12458
rect 121046 12406 121098 12458
rect 145126 12406 145178 12458
rect 90246 12294 90298 12346
rect 103350 12294 103402 12346
rect 103686 12294 103738 12346
rect 148710 12518 148762 12570
rect 149270 12518 149322 12570
rect 152854 12518 152906 12570
rect 196310 12518 196362 12570
rect 145350 12406 145402 12458
rect 150390 12406 150442 12458
rect 162822 12406 162874 12458
rect 209302 12406 209354 12458
rect 43542 11958 43594 12010
rect 58326 11958 58378 12010
rect 61238 11958 61290 12010
rect 68294 11958 68346 12010
rect 69526 11958 69578 12010
rect 55190 11846 55242 11898
rect 67846 11846 67898 11898
rect 33798 11734 33850 11786
rect 57094 11734 57146 11786
rect 56982 11622 57034 11674
rect 65718 11734 65770 11786
rect 73222 11846 73274 11898
rect 68070 11734 68122 11786
rect 74118 11846 74170 11898
rect 74678 11846 74730 11898
rect 77590 11846 77642 11898
rect 77814 11958 77866 12010
rect 79606 11958 79658 12010
rect 80838 12070 80890 12122
rect 80614 11958 80666 12010
rect 82070 12070 82122 12122
rect 81062 11958 81114 12010
rect 81958 11958 82010 12010
rect 90134 12182 90186 12234
rect 98198 12182 98250 12234
rect 98534 12182 98586 12234
rect 103238 12182 103290 12234
rect 103462 12182 103514 12234
rect 115222 12182 115274 12234
rect 116678 12182 116730 12234
rect 117014 12182 117066 12234
rect 117238 12182 117290 12234
rect 144454 12182 144506 12234
rect 193062 12294 193114 12346
rect 148598 12182 148650 12234
rect 158790 12182 158842 12234
rect 175926 12182 175978 12234
rect 82742 12070 82794 12122
rect 83302 12070 83354 12122
rect 83750 12070 83802 12122
rect 91366 12070 91418 12122
rect 73558 11734 73610 11786
rect 80278 11846 80330 11898
rect 81286 11846 81338 11898
rect 81846 11846 81898 11898
rect 82518 11958 82570 12010
rect 102902 12070 102954 12122
rect 103126 12070 103178 12122
rect 114550 12070 114602 12122
rect 114774 12070 114826 12122
rect 115670 12070 115722 12122
rect 115894 12070 115946 12122
rect 122502 12070 122554 12122
rect 122726 12070 122778 12122
rect 131126 12070 131178 12122
rect 136278 12070 136330 12122
rect 82406 11846 82458 11898
rect 117462 11958 117514 12010
rect 91702 11846 91754 11898
rect 97750 11846 97802 11898
rect 98310 11846 98362 11898
rect 99206 11846 99258 11898
rect 51046 11510 51098 11562
rect 68182 11622 68234 11674
rect 79606 11622 79658 11674
rect 80502 11734 80554 11786
rect 92934 11734 92986 11786
rect 93158 11734 93210 11786
rect 64038 11510 64090 11562
rect 80166 11510 80218 11562
rect 80390 11622 80442 11674
rect 81398 11622 81450 11674
rect 81734 11622 81786 11674
rect 100438 11734 100490 11786
rect 100998 11846 101050 11898
rect 102566 11846 102618 11898
rect 103014 11846 103066 11898
rect 102230 11734 102282 11786
rect 102454 11734 102506 11786
rect 103686 11734 103738 11786
rect 104022 11846 104074 11898
rect 108726 11846 108778 11898
rect 108950 11846 109002 11898
rect 110966 11846 111018 11898
rect 111190 11846 111242 11898
rect 138854 11958 138906 12010
rect 139190 12070 139242 12122
rect 144230 12070 144282 12122
rect 159574 12070 159626 12122
rect 139750 11958 139802 12010
rect 141094 11958 141146 12010
rect 162374 11958 162426 12010
rect 170998 12070 171050 12122
rect 192054 12070 192106 12122
rect 213670 11958 213722 12010
rect 118246 11846 118298 11898
rect 118470 11846 118522 11898
rect 104582 11734 104634 11786
rect 105814 11734 105866 11786
rect 114998 11734 115050 11786
rect 115222 11734 115274 11786
rect 119254 11734 119306 11786
rect 120374 11734 120426 11786
rect 120598 11734 120650 11786
rect 125862 11734 125914 11786
rect 126086 11846 126138 11898
rect 148150 11846 148202 11898
rect 148934 11846 148986 11898
rect 151510 11846 151562 11898
rect 154870 11846 154922 11898
rect 170662 11846 170714 11898
rect 192390 11846 192442 11898
rect 141094 11734 141146 11786
rect 164614 11734 164666 11786
rect 191718 11734 191770 11786
rect 82070 11510 82122 11562
rect 50598 11398 50650 11450
rect 66950 11398 67002 11450
rect 67622 11398 67674 11450
rect 69078 11398 69130 11450
rect 69414 11398 69466 11450
rect 71878 11398 71930 11450
rect 72102 11398 72154 11450
rect 82854 11398 82906 11450
rect 83414 11398 83466 11450
rect 83974 11510 84026 11562
rect 90582 11510 90634 11562
rect 90806 11510 90858 11562
rect 91926 11510 91978 11562
rect 92934 11510 92986 11562
rect 94726 11510 94778 11562
rect 94950 11510 95002 11562
rect 98086 11510 98138 11562
rect 100998 11622 101050 11674
rect 101558 11622 101610 11674
rect 109286 11622 109338 11674
rect 109734 11622 109786 11674
rect 127766 11622 127818 11674
rect 134038 11622 134090 11674
rect 138294 11622 138346 11674
rect 138518 11622 138570 11674
rect 151286 11622 151338 11674
rect 99654 11510 99706 11562
rect 112086 11510 112138 11562
rect 98310 11398 98362 11450
rect 103350 11398 103402 11450
rect 103574 11398 103626 11450
rect 108054 11398 108106 11450
rect 49030 11286 49082 11338
rect 61798 11286 61850 11338
rect 62358 11286 62410 11338
rect 113654 11398 113706 11450
rect 109286 11286 109338 11338
rect 113878 11398 113930 11450
rect 117238 11398 117290 11450
rect 117462 11398 117514 11450
rect 114102 11286 114154 11338
rect 116454 11286 116506 11338
rect 16326 11174 16378 11226
rect 79158 11174 79210 11226
rect 79494 11174 79546 11226
rect 80614 11174 80666 11226
rect 80838 11174 80890 11226
rect 82518 11174 82570 11226
rect 82742 11174 82794 11226
rect 86438 11174 86490 11226
rect 86662 11174 86714 11226
rect 88790 11174 88842 11226
rect 89014 11174 89066 11226
rect 119030 11510 119082 11562
rect 119590 11510 119642 11562
rect 126310 11510 126362 11562
rect 126534 11510 126586 11562
rect 117798 11398 117850 11450
rect 124406 11398 124458 11450
rect 129222 11398 129274 11450
rect 135382 11398 135434 11450
rect 135718 11510 135770 11562
rect 147478 11510 147530 11562
rect 138630 11398 138682 11450
rect 150054 11398 150106 11450
rect 153526 11398 153578 11450
rect 117686 11286 117738 11338
rect 117910 11286 117962 11338
rect 121046 11286 121098 11338
rect 121830 11286 121882 11338
rect 136614 11286 136666 11338
rect 118358 11174 118410 11226
rect 118582 11174 118634 11226
rect 124966 11174 125018 11226
rect 127766 11174 127818 11226
rect 151174 11286 151226 11338
rect 138070 11174 138122 11226
rect 138966 11174 139018 11226
rect 139526 11174 139578 11226
rect 53398 11062 53450 11114
rect 130006 11062 130058 11114
rect 130454 11062 130506 11114
rect 132918 11062 132970 11114
rect 133590 11062 133642 11114
rect 135158 11062 135210 11114
rect 135382 11062 135434 11114
rect 140870 11062 140922 11114
rect 143334 11174 143386 11226
rect 146022 11174 146074 11226
rect 150390 11062 150442 11114
rect 166630 11062 166682 11114
rect 206390 11062 206442 11114
rect 6470 10950 6522 11002
rect 83638 10950 83690 11002
rect 84310 10950 84362 11002
rect 85094 10950 85146 11002
rect 85318 10950 85370 11002
rect 89574 10950 89626 11002
rect 90022 10950 90074 11002
rect 98758 10950 98810 11002
rect 98982 10950 99034 11002
rect 103014 10950 103066 11002
rect 103350 10950 103402 11002
rect 135718 10950 135770 11002
rect 135942 10950 135994 11002
rect 150278 10950 150330 11002
rect 151062 10950 151114 11002
rect 190038 10950 190090 11002
rect 21814 10838 21866 10890
rect 125526 10838 125578 10890
rect 125750 10838 125802 10890
rect 138518 10838 138570 10890
rect 138966 10838 139018 10890
rect 41302 10726 41354 10778
rect 60790 10726 60842 10778
rect 61014 10726 61066 10778
rect 65270 10726 65322 10778
rect 65494 10726 65546 10778
rect 69302 10726 69354 10778
rect 71318 10726 71370 10778
rect 73446 10726 73498 10778
rect 73782 10726 73834 10778
rect 125638 10726 125690 10778
rect 125862 10726 125914 10778
rect 134822 10726 134874 10778
rect 136390 10726 136442 10778
rect 143558 10726 143610 10778
rect 151398 10838 151450 10890
rect 194518 10838 194570 10890
rect 187798 10726 187850 10778
rect 54294 10614 54346 10666
rect 109734 10614 109786 10666
rect 109958 10614 110010 10666
rect 114214 10614 114266 10666
rect 114438 10614 114490 10666
rect 117350 10614 117402 10666
rect 117686 10614 117738 10666
rect 120486 10614 120538 10666
rect 121606 10614 121658 10666
rect 129110 10614 129162 10666
rect 130902 10614 130954 10666
rect 50038 10502 50090 10554
rect 133926 10502 133978 10554
rect 21590 10390 21642 10442
rect 83750 10390 83802 10442
rect 83974 10390 84026 10442
rect 89350 10390 89402 10442
rect 89574 10390 89626 10442
rect 134262 10390 134314 10442
rect 181078 10614 181130 10666
rect 186566 10614 186618 10666
rect 200902 10614 200954 10666
rect 137734 10502 137786 10554
rect 194966 10502 195018 10554
rect 136838 10390 136890 10442
rect 143334 10390 143386 10442
rect 143558 10390 143610 10442
rect 211430 10390 211482 10442
rect 28378 10166 28430 10218
rect 28482 10166 28534 10218
rect 28586 10166 28638 10218
rect 82706 10166 82758 10218
rect 82810 10166 82862 10218
rect 82914 10166 82966 10218
rect 137034 10166 137086 10218
rect 137138 10166 137190 10218
rect 137242 10166 137294 10218
rect 191362 10166 191414 10218
rect 191466 10166 191518 10218
rect 191570 10166 191622 10218
rect 9830 9942 9882 9994
rect 10726 9942 10778 9994
rect 11622 9942 11674 9994
rect 45558 9942 45610 9994
rect 54518 9942 54570 9994
rect 76582 9942 76634 9994
rect 77590 9942 77642 9994
rect 78374 9998 78426 10050
rect 42590 9830 42642 9882
rect 43486 9830 43538 9882
rect 47966 9830 48018 9882
rect 48862 9830 48914 9882
rect 50542 9830 50594 9882
rect 52782 9830 52834 9882
rect 70926 9830 70978 9882
rect 55190 9774 55242 9826
rect 55414 9774 55466 9826
rect 8318 9718 8370 9770
rect 11062 9718 11114 9770
rect 53566 9718 53618 9770
rect 56590 9718 56642 9770
rect 8878 9606 8930 9658
rect 10166 9606 10218 9658
rect 11958 9606 12010 9658
rect 12574 9606 12626 9658
rect 22542 9606 22594 9658
rect 25230 9606 25282 9658
rect 43934 9606 43986 9658
rect 45222 9606 45274 9658
rect 46062 9606 46114 9658
rect 46510 9606 46562 9658
rect 47070 9606 47122 9658
rect 57038 9606 57090 9658
rect 57374 9606 57426 9658
rect 58046 9606 58098 9658
rect 76246 9606 76298 9658
rect 79270 9942 79322 9994
rect 80950 9942 81002 9994
rect 81846 9942 81898 9994
rect 86774 9942 86826 9994
rect 104022 9942 104074 9994
rect 109958 9942 110010 9994
rect 111862 9942 111914 9994
rect 115782 9942 115834 9994
rect 121382 9942 121434 9994
rect 129222 9942 129274 9994
rect 131574 9942 131626 9994
rect 132582 9942 132634 9994
rect 135494 9942 135546 9994
rect 137398 9942 137450 9994
rect 139302 9942 139354 9994
rect 143222 9942 143274 9994
rect 144118 9942 144170 9994
rect 147142 9942 147194 9994
rect 151062 9942 151114 9994
rect 154982 9942 155034 9994
rect 165622 9942 165674 9994
rect 172454 9942 172506 9994
rect 176934 9942 176986 9994
rect 180070 9942 180122 9994
rect 182534 9942 182586 9994
rect 183990 9942 184042 9994
rect 187910 9942 187962 9994
rect 191830 9942 191882 9994
rect 109062 9830 109114 9882
rect 114718 9830 114770 9882
rect 137790 9830 137842 9882
rect 78934 9718 78986 9770
rect 80110 9718 80162 9770
rect 80614 9718 80666 9770
rect 82406 9718 82458 9770
rect 83134 9718 83186 9770
rect 132022 9774 132074 9826
rect 133478 9774 133530 9826
rect 134934 9774 134986 9826
rect 141710 9830 141762 9882
rect 139750 9774 139802 9826
rect 144510 9830 144562 9882
rect 147534 9830 147586 9882
rect 147982 9830 148034 9882
rect 148430 9830 148482 9882
rect 149774 9830 149826 9882
rect 151454 9830 151506 9882
rect 153022 9830 153074 9882
rect 155374 9830 155426 9882
rect 161422 9830 161474 9882
rect 156326 9774 156378 9826
rect 157782 9774 157834 9826
rect 159350 9774 159402 9826
rect 160806 9774 160858 9826
rect 164334 9830 164386 9882
rect 162374 9774 162426 9826
rect 168702 9830 168754 9882
rect 166630 9774 166682 9826
rect 173294 9830 173346 9882
rect 191382 9886 191434 9938
rect 193734 9942 193786 9994
rect 195078 9942 195130 9994
rect 195974 9942 196026 9994
rect 196422 9942 196474 9994
rect 198102 9942 198154 9994
rect 199446 9942 199498 9994
rect 202022 9942 202074 9994
rect 204822 9942 204874 9994
rect 206166 9942 206218 9994
rect 211878 9942 211930 9994
rect 171222 9774 171274 9826
rect 188750 9830 188802 9882
rect 174806 9774 174858 9826
rect 179622 9774 179674 9826
rect 181134 9774 181186 9826
rect 182758 9774 182810 9826
rect 185054 9774 185106 9826
rect 185894 9774 185946 9826
rect 198494 9830 198546 9882
rect 189814 9774 189866 9826
rect 200398 9830 200450 9882
rect 200734 9830 200786 9882
rect 202414 9830 202466 9882
rect 208182 9886 208234 9938
rect 213782 9942 213834 9994
rect 203310 9830 203362 9882
rect 208070 9774 208122 9826
rect 210982 9774 211034 9826
rect 102958 9718 103010 9770
rect 103686 9718 103738 9770
rect 108726 9718 108778 9770
rect 111526 9718 111578 9770
rect 115446 9718 115498 9770
rect 120542 9718 120594 9770
rect 121046 9718 121098 9770
rect 130006 9718 130058 9770
rect 131238 9718 131290 9770
rect 137062 9718 137114 9770
rect 142886 9718 142938 9770
rect 144958 9718 145010 9770
rect 146806 9718 146858 9770
rect 150726 9718 150778 9770
rect 154646 9718 154698 9770
rect 165286 9718 165338 9770
rect 172790 9718 172842 9770
rect 174190 9718 174242 9770
rect 177270 9718 177322 9770
rect 180406 9718 180458 9770
rect 192166 9718 192218 9770
rect 194742 9718 194794 9770
rect 204486 9718 204538 9770
rect 217310 9718 217362 9770
rect 77254 9606 77306 9658
rect 78262 9606 78314 9658
rect 78430 9606 78482 9658
rect 81510 9606 81562 9658
rect 82742 9606 82794 9658
rect 83918 9606 83970 9658
rect 85934 9606 85986 9658
rect 86438 9606 86490 9658
rect 96014 9606 96066 9658
rect 98926 9606 98978 9658
rect 99710 9606 99762 9658
rect 100046 9606 100098 9658
rect 106878 9606 106930 9658
rect 107830 9606 107882 9658
rect 108166 9606 108218 9658
rect 109622 9606 109674 9658
rect 110798 9606 110850 9658
rect 128382 9606 128434 9658
rect 128886 9606 128938 9658
rect 130342 9606 130394 9658
rect 135942 9662 135994 9714
rect 134094 9606 134146 9658
rect 140758 9662 140810 9714
rect 138966 9606 139018 9658
rect 143782 9606 143834 9658
rect 140982 9550 141034 9602
rect 145518 9606 145570 9658
rect 145966 9606 146018 9658
rect 148878 9606 148930 9658
rect 149438 9606 149490 9658
rect 152238 9606 152290 9658
rect 152686 9606 152738 9658
rect 153582 9606 153634 9658
rect 158566 9606 158618 9658
rect 156326 9550 156378 9602
rect 163718 9662 163770 9714
rect 166742 9662 166794 9714
rect 158902 9606 158954 9658
rect 171670 9662 171722 9714
rect 175142 9662 175194 9714
rect 178278 9662 178330 9714
rect 169150 9606 169202 9658
rect 160582 9550 160634 9602
rect 163606 9550 163658 9602
rect 182086 9662 182138 9714
rect 181022 9606 181074 9658
rect 170326 9550 170378 9602
rect 178166 9550 178218 9602
rect 184326 9606 184378 9658
rect 186006 9662 186058 9714
rect 184942 9606 184994 9658
rect 189926 9662 189978 9714
rect 188246 9606 188298 9658
rect 187350 9550 187402 9602
rect 192782 9606 192834 9658
rect 194070 9606 194122 9658
rect 195638 9606 195690 9658
rect 196758 9606 196810 9658
rect 197766 9606 197818 9658
rect 199110 9606 199162 9658
rect 199950 9606 200002 9658
rect 201686 9606 201738 9658
rect 202862 9606 202914 9658
rect 203870 9606 203922 9658
rect 210758 9662 210810 9714
rect 205830 9606 205882 9658
rect 211542 9606 211594 9658
rect 209526 9550 209578 9602
rect 212270 9606 212322 9658
rect 213446 9606 213498 9658
rect 214174 9606 214226 9658
rect 214622 9606 214674 9658
rect 215070 9606 215122 9658
rect 215518 9606 215570 9658
rect 215966 9606 216018 9658
rect 216414 9606 216466 9658
rect 55542 9382 55594 9434
rect 55646 9382 55698 9434
rect 55750 9382 55802 9434
rect 109870 9382 109922 9434
rect 109974 9382 110026 9434
rect 110078 9382 110130 9434
rect 164198 9382 164250 9434
rect 164302 9382 164354 9434
rect 164406 9382 164458 9434
rect 9718 9158 9770 9210
rect 10614 9158 10666 9210
rect 15598 9158 15650 9210
rect 17782 9158 17834 9210
rect 18118 9158 18170 9210
rect 18510 9158 18562 9210
rect 19910 9158 19962 9210
rect 20246 9158 20298 9210
rect 20638 9158 20690 9210
rect 22262 9158 22314 9210
rect 25958 9158 26010 9210
rect 41974 9158 42026 9210
rect 42310 9158 42362 9210
rect 43206 9158 43258 9210
rect 44046 9158 44098 9210
rect 44550 9158 44602 9210
rect 44886 9158 44938 9210
rect 45390 9158 45442 9210
rect 47350 9158 47402 9210
rect 47686 9158 47738 9210
rect 48582 9158 48634 9210
rect 49926 9158 49978 9210
rect 50262 9158 50314 9210
rect 50822 9158 50874 9210
rect 51158 9158 51210 9210
rect 51550 9158 51602 9210
rect 52166 9158 52218 9210
rect 52502 9158 52554 9210
rect 57766 9158 57818 9210
rect 61238 9158 61290 9210
rect 61574 9158 61626 9210
rect 61966 9158 62018 9210
rect 70198 9158 70250 9210
rect 74118 9158 74170 9210
rect 74454 9158 74506 9210
rect 76750 9158 76802 9210
rect 78654 9158 78706 9210
rect 79606 9158 79658 9210
rect 80502 9158 80554 9210
rect 82518 9158 82570 9210
rect 8990 9046 9042 9098
rect 10054 9046 10106 9098
rect 10950 9046 11002 9098
rect 21926 9046 21978 9098
rect 25622 9046 25674 9098
rect 42870 9046 42922 9098
rect 45894 9046 45946 9098
rect 46846 9046 46898 9098
rect 48246 9046 48298 9098
rect 14086 8990 14138 9042
rect 15094 8990 15146 9042
rect 23382 8990 23434 9042
rect 16046 8934 16098 8986
rect 26350 8934 26402 8986
rect 23046 8878 23098 8930
rect 36990 8934 37042 8986
rect 38110 8934 38162 8986
rect 41470 8934 41522 8986
rect 54854 8990 54906 9042
rect 56422 9001 56474 9053
rect 57430 9046 57482 9098
rect 58382 9046 58434 9098
rect 86046 9102 86098 9154
rect 86494 9158 86546 9210
rect 87726 9158 87778 9210
rect 90694 9158 90746 9210
rect 92206 9158 92258 9210
rect 92822 9158 92874 9210
rect 93158 9158 93210 9210
rect 97750 9214 97802 9266
rect 94894 9158 94946 9210
rect 99766 9158 99818 9210
rect 99094 9102 99146 9154
rect 104302 9158 104354 9210
rect 105142 9158 105194 9210
rect 108334 9158 108386 9210
rect 118414 9158 118466 9210
rect 118526 9102 118578 9154
rect 129614 9158 129666 9210
rect 130846 9158 130898 9210
rect 131406 9158 131458 9210
rect 141318 9158 141370 9210
rect 141710 9158 141762 9210
rect 146974 9158 147026 9210
rect 159182 9158 159234 9210
rect 153078 9102 153130 9154
rect 159630 9158 159682 9210
rect 161310 9158 161362 9210
rect 166462 9158 166514 9210
rect 58830 9046 58882 9098
rect 62806 9046 62858 9098
rect 69862 9046 69914 9098
rect 71262 9046 71314 9098
rect 79270 9046 79322 9098
rect 80166 9046 80218 9098
rect 81286 9046 81338 9098
rect 82182 9046 82234 9098
rect 90358 9046 90410 9098
rect 49310 8934 49362 8986
rect 59390 8934 59442 8986
rect 63534 8934 63586 8986
rect 65326 8934 65378 8986
rect 68686 8934 68738 8986
rect 70590 8934 70642 8986
rect 72046 8934 72098 8986
rect 73278 8934 73330 8986
rect 74846 8934 74898 8986
rect 77758 8934 77810 8986
rect 83078 8990 83130 9042
rect 78206 8934 78258 8986
rect 83806 8934 83858 8986
rect 84254 8934 84306 8986
rect 84702 8934 84754 8986
rect 87054 8934 87106 8986
rect 88398 8990 88450 9042
rect 95958 9046 96010 9098
rect 140982 9046 141034 9098
rect 89070 8934 89122 8986
rect 89742 8934 89794 8986
rect 91310 8990 91362 9042
rect 91758 8934 91810 8986
rect 98982 8990 99034 9042
rect 100830 8990 100882 9042
rect 95342 8934 95394 8986
rect 101278 8934 101330 8986
rect 109230 8934 109282 8986
rect 118974 8934 119026 8986
rect 131798 8990 131850 9042
rect 133254 8990 133306 9042
rect 134262 8990 134314 9042
rect 135270 8990 135322 9042
rect 124798 8934 124850 8986
rect 137622 8990 137674 9042
rect 138294 8990 138346 9042
rect 138854 8990 138906 9042
rect 140310 8990 140362 9042
rect 142326 8990 142378 9042
rect 143782 8990 143834 9042
rect 145126 8990 145178 9042
rect 146470 8990 146522 9042
rect 135774 8934 135826 8986
rect 13078 8822 13130 8874
rect 46230 8822 46282 8874
rect 53286 8822 53338 8874
rect 58270 8822 58322 8874
rect 63142 8822 63194 8874
rect 81622 8822 81674 8874
rect 83414 8822 83466 8874
rect 85934 8822 85986 8874
rect 88286 8822 88338 8874
rect 91198 8822 91250 8874
rect 96294 8822 96346 8874
rect 100102 8822 100154 8874
rect 100718 8822 100770 8874
rect 133142 8878 133194 8930
rect 135382 8878 135434 8930
rect 148150 8990 148202 9042
rect 149494 8990 149546 9042
rect 150502 8990 150554 9042
rect 151846 8990 151898 9042
rect 152966 8990 153018 9042
rect 155206 8990 155258 9042
rect 156326 8990 156378 9042
rect 157222 8990 157274 9042
rect 158678 8990 158730 9042
rect 160862 8990 160914 9042
rect 161758 9046 161810 9098
rect 167918 9102 167970 9154
rect 172566 9158 172618 9210
rect 175478 9158 175530 9210
rect 181862 9214 181914 9266
rect 176598 9158 176650 9210
rect 190598 9158 190650 9210
rect 170830 9046 170882 9098
rect 164390 8990 164442 9042
rect 166070 8990 166122 9042
rect 147422 8934 147474 8986
rect 168870 8990 168922 9042
rect 170102 8990 170154 9042
rect 182758 9102 182810 9154
rect 185110 9102 185162 9154
rect 186678 9102 186730 9154
rect 188694 9102 188746 9154
rect 190934 9158 190986 9210
rect 191438 9158 191490 9210
rect 194518 9158 194570 9210
rect 192838 9102 192890 9154
rect 195414 9158 195466 9210
rect 196310 9158 196362 9210
rect 197206 9158 197258 9210
rect 198046 9158 198098 9210
rect 198494 9158 198546 9210
rect 199390 9158 199442 9210
rect 200398 9158 200450 9210
rect 200846 9158 200898 9210
rect 201294 9158 201346 9210
rect 202190 9158 202242 9210
rect 203254 9158 203306 9210
rect 212774 9158 212826 9210
rect 207510 9102 207562 9154
rect 209862 9102 209914 9154
rect 211094 9102 211146 9154
rect 213110 9158 213162 9210
rect 214846 9158 214898 9210
rect 216750 9158 216802 9210
rect 170942 9046 170994 9098
rect 173350 8990 173402 9042
rect 175814 9046 175866 9098
rect 176934 9046 176986 9098
rect 140422 8878 140474 8930
rect 143894 8878 143946 8930
rect 166910 8934 166962 8986
rect 175030 8986 175082 9038
rect 179622 8990 179674 9042
rect 194854 9046 194906 9098
rect 195750 9046 195802 9098
rect 196646 9046 196698 9098
rect 197542 9046 197594 9098
rect 202918 9046 202970 9098
rect 216302 9046 216354 9098
rect 181302 8986 181354 9038
rect 182982 8990 183034 9042
rect 184550 8990 184602 9042
rect 186566 8990 186618 9042
rect 188582 8990 188634 9042
rect 193062 8990 193114 9042
rect 154422 8878 154474 8930
rect 183710 8934 183762 8986
rect 198942 8934 198994 8986
rect 105478 8822 105530 8874
rect 137398 8822 137450 8874
rect 145574 8822 145626 8874
rect 148598 8822 148650 8874
rect 150950 8822 151002 8874
rect 155430 8822 155482 8874
rect 157782 8822 157834 8874
rect 160750 8822 160802 8874
rect 162822 8822 162874 8874
rect 186118 8878 186170 8930
rect 187910 8878 187962 8930
rect 192726 8878 192778 8930
rect 204038 8990 204090 9042
rect 206502 8990 206554 9042
rect 209526 8990 209578 9042
rect 211430 8990 211482 9042
rect 201742 8934 201794 8986
rect 213502 8934 213554 8986
rect 204150 8878 204202 8930
rect 211990 8878 212042 8930
rect 213950 8934 214002 8986
rect 214398 8934 214450 8986
rect 215294 8934 215346 8986
rect 167806 8822 167858 8874
rect 169206 8822 169258 8874
rect 179286 8822 179338 8874
rect 189142 8822 189194 8874
rect 206726 8822 206778 8874
rect 28378 8598 28430 8650
rect 28482 8598 28534 8650
rect 28586 8598 28638 8650
rect 82706 8598 82758 8650
rect 82810 8598 82862 8650
rect 82914 8598 82966 8650
rect 137034 8598 137086 8650
rect 137138 8598 137190 8650
rect 137242 8598 137294 8650
rect 191362 8598 191414 8650
rect 191466 8598 191518 8650
rect 191570 8598 191622 8650
rect 16326 8374 16378 8426
rect 21814 8374 21866 8426
rect 56422 8374 56474 8426
rect 70198 8374 70250 8426
rect 71766 8374 71818 8426
rect 87726 8374 87778 8426
rect 90414 8374 90466 8426
rect 98310 8374 98362 8426
rect 118918 8374 118970 8426
rect 139526 8374 139578 8426
rect 145686 8374 145738 8426
rect 149270 8374 149322 8426
rect 153974 8374 154026 8426
rect 158902 8374 158954 8426
rect 171334 8374 171386 8426
rect 179062 8374 179114 8426
rect 181526 8374 181578 8426
rect 183542 8374 183594 8426
rect 185558 8374 185610 8426
rect 186566 8374 186618 8426
rect 10278 8262 10330 8314
rect 11622 8206 11674 8258
rect 12854 8210 12906 8262
rect 13582 8262 13634 8314
rect 16662 8206 16714 8258
rect 18342 8206 18394 8258
rect 23382 8206 23434 8258
rect 25062 8206 25114 8258
rect 26966 8262 27018 8314
rect 29878 8262 29930 8314
rect 31894 8262 31946 8314
rect 34358 8262 34410 8314
rect 35254 8262 35306 8314
rect 36710 8262 36762 8314
rect 37830 8262 37882 8314
rect 39062 8262 39114 8314
rect 39958 8262 40010 8314
rect 41078 8262 41130 8314
rect 41974 8262 42026 8314
rect 42870 8262 42922 8314
rect 43766 8262 43818 8314
rect 44662 8262 44714 8314
rect 45894 8262 45946 8314
rect 46790 8262 46842 8314
rect 47686 8262 47738 8314
rect 48582 8262 48634 8314
rect 50038 8262 50090 8314
rect 51606 8206 51658 8258
rect 52614 8206 52666 8258
rect 54406 8262 54458 8314
rect 56758 8206 56810 8258
rect 58438 8206 58490 8258
rect 59334 8262 59386 8314
rect 62358 8262 62410 8314
rect 63254 8206 63306 8258
rect 64934 8210 64986 8262
rect 66558 8262 66610 8314
rect 67398 8262 67450 8314
rect 73782 8262 73834 8314
rect 26630 8150 26682 8202
rect 29542 8150 29594 8202
rect 31558 8150 31610 8202
rect 34918 8150 34970 8202
rect 45558 8150 45610 8202
rect 48246 8150 48298 8202
rect 58998 8150 59050 8202
rect 65718 8150 65770 8202
rect 66054 8150 66106 8202
rect 68462 8206 68514 8258
rect 70758 8206 70810 8258
rect 74790 8206 74842 8258
rect 76470 8206 76522 8258
rect 77982 8262 78034 8314
rect 93942 8318 93994 8370
rect 101670 8318 101722 8370
rect 199670 8374 199722 8426
rect 83302 8206 83354 8258
rect 84422 8206 84474 8258
rect 71430 8150 71482 8202
rect 88510 8206 88562 8258
rect 89910 8262 89962 8314
rect 13918 8038 13970 8090
rect 18734 8038 18786 8090
rect 19182 8038 19234 8090
rect 25454 8038 25506 8090
rect 25902 8038 25954 8090
rect 27470 8038 27522 8090
rect 30382 8038 30434 8090
rect 32398 8038 32450 8090
rect 34022 8038 34074 8090
rect 35758 8038 35810 8090
rect 36374 8038 36426 8090
rect 37494 8038 37546 8090
rect 38726 8038 38778 8090
rect 39622 8038 39674 8090
rect 40742 8038 40794 8090
rect 41638 8038 41690 8090
rect 42534 8038 42586 8090
rect 43430 8038 43482 8090
rect 44326 8038 44378 8090
rect 46454 8038 46506 8090
rect 47350 8038 47402 8090
rect 53566 8038 53618 8090
rect 54070 8038 54122 8090
rect 59838 8038 59890 8090
rect 59950 8094 60002 8146
rect 60510 8038 60562 8090
rect 67062 8038 67114 8090
rect 67902 8038 67954 8090
rect 70646 8094 70698 8146
rect 68350 8038 68402 8090
rect 72382 8038 72434 8090
rect 78318 8038 78370 8090
rect 78878 8038 78930 8090
rect 79326 8038 79378 8090
rect 79438 8094 79490 8146
rect 86550 8150 86602 8202
rect 80054 8038 80106 8090
rect 80390 8038 80442 8090
rect 81958 8038 82010 8090
rect 85262 8038 85314 8090
rect 85710 8038 85762 8090
rect 85822 8094 85874 8146
rect 86886 8038 86938 8090
rect 87838 8094 87890 8146
rect 88398 8038 88450 8090
rect 89070 8038 89122 8090
rect 89574 8038 89626 8090
rect 90526 8094 90578 8146
rect 91198 8150 91250 8202
rect 94838 8206 94890 8258
rect 98646 8206 98698 8258
rect 100326 8210 100378 8262
rect 107886 8262 107938 8314
rect 91646 8150 91698 8202
rect 102566 8206 102618 8258
rect 110462 8206 110514 8258
rect 117014 8225 117066 8277
rect 117910 8206 117962 8258
rect 125078 8225 125130 8277
rect 125974 8206 126026 8258
rect 130510 8206 130562 8258
rect 132078 8262 132130 8314
rect 133590 8262 133642 8314
rect 133982 8262 134034 8314
rect 147086 8262 147138 8314
rect 116174 8150 116226 8202
rect 95398 8094 95450 8146
rect 91086 8038 91138 8090
rect 103014 8094 103066 8146
rect 96238 8038 96290 8090
rect 103630 8038 103682 8090
rect 104078 8038 104130 8090
rect 104526 8038 104578 8090
rect 107550 8038 107602 8090
rect 110350 8038 110402 8090
rect 110910 8038 110962 8090
rect 121662 8038 121714 8090
rect 123230 8038 123282 8090
rect 123342 8094 123394 8146
rect 130958 8150 131010 8202
rect 133254 8150 133306 8202
rect 134598 8195 134650 8247
rect 135494 8206 135546 8258
rect 139190 8206 139242 8258
rect 143334 8206 143386 8258
rect 144230 8195 144282 8247
rect 145126 8206 145178 8258
rect 146582 8206 146634 8258
rect 147534 8262 147586 8314
rect 151118 8262 151170 8314
rect 148710 8206 148762 8258
rect 190486 8262 190538 8314
rect 150670 8150 150722 8202
rect 151902 8206 151954 8258
rect 154310 8206 154362 8258
rect 155990 8206 156042 8258
rect 159238 8206 159290 8258
rect 160918 8206 160970 8258
rect 161478 8206 161530 8258
rect 163886 8206 163938 8258
rect 164726 8206 164778 8258
rect 166966 8206 167018 8258
rect 170774 8206 170826 8258
rect 175926 8206 175978 8258
rect 177606 8206 177658 8258
rect 179174 8206 179226 8258
rect 181190 8206 181242 8258
rect 182870 8206 182922 8258
rect 186118 8206 186170 8258
rect 123790 8038 123842 8090
rect 127542 8038 127594 8090
rect 129054 8038 129106 8090
rect 130398 8038 130450 8090
rect 138966 8094 139018 8146
rect 131630 8038 131682 8090
rect 137286 8038 137338 8090
rect 141878 8038 141930 8090
rect 150054 8094 150106 8146
rect 187518 8150 187570 8202
rect 187630 8206 187682 8258
rect 188470 8206 188522 8258
rect 200398 8262 200450 8314
rect 192278 8195 192330 8247
rect 193622 8206 193674 8258
rect 196422 8206 196474 8258
rect 197542 8206 197594 8258
rect 201406 8262 201458 8314
rect 204318 8262 204370 8314
rect 209862 8318 209914 8370
rect 205942 8262 205994 8314
rect 211262 8262 211314 8314
rect 206950 8206 207002 8258
rect 208630 8206 208682 8258
rect 209190 8206 209242 8258
rect 215070 8262 215122 8314
rect 215518 8262 215570 8314
rect 147982 8038 148034 8090
rect 151790 8038 151842 8090
rect 162374 8094 162426 8146
rect 156606 8038 156658 8090
rect 166070 8094 166122 8146
rect 167414 8094 167466 8146
rect 169318 8094 169370 8146
rect 163774 8038 163826 8090
rect 171670 8038 171722 8090
rect 172566 8038 172618 8090
rect 172902 8038 172954 8090
rect 179398 8094 179450 8146
rect 180966 8094 181018 8146
rect 182982 8094 183034 8146
rect 185894 8094 185946 8146
rect 202190 8150 202242 8202
rect 188694 8094 188746 8146
rect 214510 8150 214562 8202
rect 173406 8038 173458 8090
rect 175030 8038 175082 8090
rect 186902 8038 186954 8090
rect 190822 8038 190874 8090
rect 189366 7982 189418 8034
rect 191326 8038 191378 8090
rect 194630 8038 194682 8090
rect 200846 8038 200898 8090
rect 201742 8038 201794 8090
rect 202638 8038 202690 8090
rect 203086 8038 203138 8090
rect 203646 8038 203698 8090
rect 212270 8038 212322 8090
rect 212718 8038 212770 8090
rect 213166 8038 213218 8090
rect 213614 8038 213666 8090
rect 214062 8038 214114 8090
rect 215854 8038 215906 8090
rect 216302 8038 216354 8090
rect 55542 7814 55594 7866
rect 55646 7814 55698 7866
rect 55750 7814 55802 7866
rect 109870 7814 109922 7866
rect 109974 7814 110026 7866
rect 110078 7814 110130 7866
rect 164198 7814 164250 7866
rect 164302 7814 164354 7866
rect 164406 7814 164458 7866
rect 6470 7590 6522 7642
rect 9550 7590 9602 7642
rect 21590 7590 21642 7642
rect 26854 7590 26906 7642
rect 40798 7590 40850 7642
rect 42198 7590 42250 7642
rect 43094 7590 43146 7642
rect 46230 7590 46282 7642
rect 50710 7646 50762 7698
rect 49814 7590 49866 7642
rect 59502 7590 59554 7642
rect 51942 7534 51994 7586
rect 58662 7534 58714 7586
rect 63422 7590 63474 7642
rect 62918 7534 62970 7586
rect 63870 7590 63922 7642
rect 79438 7590 79490 7642
rect 66726 7534 66778 7586
rect 74678 7534 74730 7586
rect 78374 7534 78426 7586
rect 118806 7646 118858 7698
rect 88510 7590 88562 7642
rect 95622 7590 95674 7642
rect 115950 7590 116002 7642
rect 84870 7534 84922 7586
rect 87222 7534 87274 7586
rect 90358 7534 90410 7586
rect 104134 7534 104186 7586
rect 107158 7534 107210 7586
rect 115446 7534 115498 7586
rect 120878 7590 120930 7642
rect 117798 7534 117850 7586
rect 119926 7534 119978 7586
rect 126702 7590 126754 7642
rect 126814 7534 126866 7586
rect 127262 7590 127314 7642
rect 135214 7590 135266 7642
rect 133590 7534 133642 7586
rect 135998 7590 136050 7642
rect 142830 7590 142882 7642
rect 139974 7534 140026 7586
rect 143726 7590 143778 7642
rect 145294 7590 145346 7642
rect 150446 7590 150498 7642
rect 151006 7590 151058 7642
rect 151342 7590 151394 7642
rect 151790 7590 151842 7642
rect 157166 7590 157218 7642
rect 7926 7422 7978 7474
rect 8934 7422 8986 7474
rect 12742 7422 12794 7474
rect 15878 7422 15930 7474
rect 10334 7366 10386 7418
rect 16886 7418 16938 7470
rect 17614 7366 17666 7418
rect 11398 7310 11450 7362
rect 18062 7366 18114 7418
rect 18622 7366 18674 7418
rect 23046 7422 23098 7474
rect 19182 7366 19234 7418
rect 24054 7418 24106 7470
rect 24558 7366 24610 7418
rect 28198 7422 28250 7474
rect 41862 7478 41914 7530
rect 42758 7478 42810 7530
rect 43654 7478 43706 7530
rect 49478 7478 49530 7530
rect 80166 7478 80218 7530
rect 152966 7534 153018 7586
rect 156102 7534 156154 7586
rect 166966 7590 167018 7642
rect 169430 7590 169482 7642
rect 174918 7590 174970 7642
rect 177718 7590 177770 7642
rect 184774 7646 184826 7698
rect 25566 7366 25618 7418
rect 29654 7418 29706 7470
rect 30158 7366 30210 7418
rect 30606 7366 30658 7418
rect 37830 7422 37882 7474
rect 34526 7366 34578 7418
rect 38726 7403 38778 7455
rect 39230 7366 39282 7418
rect 39790 7366 39842 7418
rect 40126 7366 40178 7418
rect 47686 7422 47738 7474
rect 44606 7366 44658 7418
rect 48582 7403 48634 7455
rect 52166 7422 52218 7474
rect 54966 7422 55018 7474
rect 56646 7422 56698 7474
rect 58998 7422 59050 7474
rect 52670 7366 52722 7418
rect 63030 7422 63082 7474
rect 66390 7422 66442 7474
rect 60174 7366 60226 7418
rect 14870 7254 14922 7306
rect 36822 7254 36874 7306
rect 43990 7254 44042 7306
rect 57430 7310 57482 7362
rect 67230 7366 67282 7418
rect 68126 7366 68178 7418
rect 70870 7422 70922 7474
rect 72550 7422 72602 7474
rect 74566 7422 74618 7474
rect 68574 7366 68626 7418
rect 75182 7366 75234 7418
rect 75630 7366 75682 7418
rect 78038 7422 78090 7474
rect 76078 7366 76130 7418
rect 78878 7366 78930 7418
rect 79550 7422 79602 7474
rect 81286 7422 81338 7474
rect 81846 7422 81898 7474
rect 84982 7422 85034 7474
rect 87446 7422 87498 7474
rect 85374 7366 85426 7418
rect 81174 7310 81226 7362
rect 90582 7422 90634 7474
rect 87950 7366 88002 7418
rect 85990 7310 86042 7362
rect 91086 7366 91138 7418
rect 89126 7310 89178 7362
rect 91534 7366 91586 7418
rect 92430 7366 92482 7418
rect 92822 7418 92874 7470
rect 93830 7422 93882 7474
rect 97694 7366 97746 7418
rect 98086 7418 98138 7470
rect 99094 7422 99146 7474
rect 104246 7422 104298 7474
rect 100662 7366 100714 7418
rect 107270 7422 107322 7474
rect 104974 7366 105026 7418
rect 107830 7403 107882 7455
rect 108726 7422 108778 7474
rect 115558 7422 115610 7474
rect 118134 7422 118186 7474
rect 120262 7422 120314 7474
rect 121942 7433 121994 7485
rect 122838 7422 122890 7474
rect 102790 7310 102842 7362
rect 121326 7366 121378 7418
rect 105702 7310 105754 7362
rect 113990 7310 114042 7362
rect 117014 7310 117066 7362
rect 129390 7422 129442 7474
rect 130230 7422 130282 7474
rect 133366 7422 133418 7474
rect 136110 7422 136162 7474
rect 136950 7422 137002 7474
rect 138294 7422 138346 7474
rect 140310 7422 140362 7474
rect 140982 7422 141034 7474
rect 142438 7422 142490 7474
rect 143614 7422 143666 7474
rect 128270 7366 128322 7418
rect 147926 7422 147978 7474
rect 144734 7366 144786 7418
rect 149606 7418 149658 7470
rect 149998 7478 150050 7530
rect 167302 7478 167354 7530
rect 153414 7422 153466 7474
rect 155542 7422 155594 7474
rect 156718 7366 156770 7418
rect 159462 7422 159514 7474
rect 162598 7422 162650 7474
rect 164278 7422 164330 7474
rect 164838 7422 164890 7474
rect 157614 7366 157666 7418
rect 170662 7422 170714 7474
rect 172230 7422 172282 7474
rect 167806 7366 167858 7418
rect 175254 7478 175306 7530
rect 175758 7478 175810 7530
rect 180798 7534 180850 7586
rect 183710 7590 183762 7642
rect 190598 7590 190650 7642
rect 183822 7534 183874 7586
rect 189926 7534 189978 7586
rect 190934 7590 190986 7642
rect 191774 7534 191826 7586
rect 192446 7590 192498 7642
rect 192894 7590 192946 7642
rect 193790 7590 193842 7642
rect 193902 7534 193954 7586
rect 195022 7534 195074 7586
rect 195134 7590 195186 7642
rect 195582 7590 195634 7642
rect 196030 7590 196082 7642
rect 196926 7590 196978 7642
rect 197374 7590 197426 7642
rect 198270 7590 198322 7642
rect 198718 7590 198770 7642
rect 203086 7590 203138 7642
rect 210870 7590 210922 7642
rect 209638 7534 209690 7586
rect 211710 7590 211762 7642
rect 212158 7590 212210 7642
rect 212606 7590 212658 7642
rect 213054 7590 213106 7642
rect 215294 7590 215346 7642
rect 174358 7422 174410 7474
rect 178502 7422 178554 7474
rect 199614 7478 199666 7530
rect 180182 7418 180234 7470
rect 182982 7422 183034 7474
rect 184662 7422 184714 7474
rect 185782 7422 185834 7474
rect 186678 7422 186730 7474
rect 188022 7422 188074 7474
rect 189702 7422 189754 7474
rect 158454 7310 158506 7362
rect 166182 7310 166234 7362
rect 194350 7366 194402 7418
rect 173126 7310 173178 7362
rect 53398 7254 53450 7306
rect 62470 7254 62522 7306
rect 66278 7254 66330 7306
rect 70534 7254 70586 7306
rect 74230 7254 74282 7306
rect 77926 7254 77978 7306
rect 80502 7254 80554 7306
rect 84422 7254 84474 7306
rect 110966 7254 111018 7306
rect 123846 7254 123898 7306
rect 132470 7254 132522 7306
rect 133814 7254 133866 7306
rect 137398 7254 137450 7306
rect 139862 7254 139914 7306
rect 141878 7254 141930 7306
rect 147590 7254 147642 7306
rect 153750 7254 153802 7306
rect 155318 7254 155370 7306
rect 161030 7254 161082 7306
rect 181638 7310 181690 7362
rect 186566 7310 186618 7362
rect 196478 7366 196530 7418
rect 197822 7366 197874 7418
rect 200566 7422 200618 7474
rect 199166 7366 199218 7418
rect 202638 7366 202690 7418
rect 201574 7310 201626 7362
rect 206054 7422 206106 7474
rect 210534 7478 210586 7530
rect 213950 7478 214002 7530
rect 203534 7366 203586 7418
rect 207734 7418 207786 7470
rect 209862 7422 209914 7474
rect 211262 7366 211314 7418
rect 180686 7254 180738 7306
rect 189590 7254 189642 7306
rect 191662 7254 191714 7306
rect 208406 7310 208458 7362
rect 213502 7366 213554 7418
rect 214398 7366 214450 7418
rect 214846 7366 214898 7418
rect 204486 7254 204538 7306
rect 28378 7030 28430 7082
rect 28482 7030 28534 7082
rect 28586 7030 28638 7082
rect 82706 7030 82758 7082
rect 82810 7030 82862 7082
rect 82914 7030 82966 7082
rect 137034 7030 137086 7082
rect 137138 7030 137190 7082
rect 137242 7030 137294 7082
rect 191362 7030 191414 7082
rect 191466 7030 191518 7082
rect 191570 7030 191622 7082
rect 10838 6806 10890 6858
rect 16214 6806 16266 6858
rect 32678 6806 32730 6858
rect 41414 6806 41466 6858
rect 48358 6806 48410 6858
rect 58046 6806 58098 6858
rect 63814 6806 63866 6858
rect 69358 6806 69410 6858
rect 72214 6806 72266 6858
rect 105478 6806 105530 6858
rect 105702 6806 105754 6858
rect 127990 6806 128042 6858
rect 137846 6806 137898 6858
rect 141766 6806 141818 6858
rect 145798 6806 145850 6858
rect 152182 6806 152234 6858
rect 157334 6806 157386 6858
rect 174134 6806 174186 6858
rect 182646 6806 182698 6858
rect 187126 6806 187178 6858
rect 200566 6806 200618 6858
rect 210702 6806 210754 6858
rect 43934 6694 43986 6746
rect 11510 6638 11562 6690
rect 12854 6638 12906 6690
rect 16662 6638 16714 6690
rect 18230 6638 18282 6690
rect 20694 6638 20746 6690
rect 24390 6638 24442 6690
rect 27750 6638 27802 6690
rect 13582 6582 13634 6634
rect 28702 6582 28754 6634
rect 8766 6470 8818 6522
rect 19350 6526 19402 6578
rect 14030 6470 14082 6522
rect 23046 6526 23098 6578
rect 21534 6470 21586 6522
rect 26406 6526 26458 6578
rect 33462 6638 33514 6690
rect 34694 6638 34746 6690
rect 41862 6638 41914 6690
rect 47406 6694 47458 6746
rect 49870 6694 49922 6746
rect 30606 6582 30658 6634
rect 43318 6627 43370 6679
rect 49030 6638 49082 6690
rect 50542 6638 50594 6690
rect 50990 6694 51042 6746
rect 51774 6694 51826 6746
rect 54294 6694 54346 6746
rect 55190 6638 55242 6690
rect 56758 6627 56810 6679
rect 25006 6470 25058 6522
rect 28366 6470 28418 6522
rect 35086 6470 35138 6522
rect 35534 6470 35586 6522
rect 39006 6470 39058 6522
rect 48358 6526 48410 6578
rect 44382 6470 44434 6522
rect 50430 6470 50482 6522
rect 52110 6470 52162 6522
rect 52558 6470 52610 6522
rect 57374 6470 57426 6522
rect 57486 6526 57538 6578
rect 58158 6526 58210 6578
rect 58606 6582 58658 6634
rect 64150 6638 64202 6690
rect 65830 6642 65882 6694
rect 66558 6694 66610 6746
rect 67902 6694 67954 6746
rect 70030 6694 70082 6746
rect 59390 6582 59442 6634
rect 70142 6638 70194 6690
rect 72550 6638 72602 6690
rect 74230 6638 74282 6690
rect 75070 6638 75122 6690
rect 59950 6470 60002 6522
rect 61742 6470 61794 6522
rect 67006 6470 67058 6522
rect 67454 6470 67506 6522
rect 68350 6470 68402 6522
rect 68462 6526 68514 6578
rect 69470 6526 69522 6578
rect 75182 6582 75234 6634
rect 75854 6638 75906 6690
rect 76302 6694 76354 6746
rect 77198 6638 77250 6690
rect 78318 6694 78370 6746
rect 81510 6694 81562 6746
rect 78822 6638 78874 6690
rect 79830 6638 79882 6690
rect 82910 6638 82962 6690
rect 83470 6694 83522 6746
rect 84030 6694 84082 6746
rect 98758 6750 98810 6802
rect 86662 6638 86714 6690
rect 87670 6638 87722 6690
rect 90750 6638 90802 6690
rect 91758 6694 91810 6746
rect 113262 6694 113314 6746
rect 97414 6638 97466 6690
rect 100326 6638 100378 6690
rect 102118 6638 102170 6690
rect 103126 6638 103178 6690
rect 110518 6638 110570 6690
rect 112758 6638 112810 6690
rect 121046 6750 121098 6802
rect 124854 6750 124906 6802
rect 129334 6750 129386 6802
rect 132806 6750 132858 6802
rect 134822 6750 134874 6802
rect 115950 6694 116002 6746
rect 142774 6750 142826 6802
rect 148710 6750 148762 6802
rect 170214 6750 170266 6802
rect 177158 6750 177210 6802
rect 138798 6694 138850 6746
rect 185110 6750 185162 6802
rect 188470 6750 188522 6802
rect 75742 6470 75794 6522
rect 77310 6470 77362 6522
rect 77982 6470 78034 6522
rect 83022 6470 83074 6522
rect 84478 6470 84530 6522
rect 85150 6526 85202 6578
rect 90862 6582 90914 6634
rect 122614 6638 122666 6690
rect 126422 6638 126474 6690
rect 128550 6638 128602 6690
rect 130902 6638 130954 6690
rect 118414 6582 118466 6634
rect 85262 6470 85314 6522
rect 85822 6470 85874 6522
rect 97302 6526 97354 6578
rect 86158 6470 86210 6522
rect 89462 6470 89514 6522
rect 91422 6470 91474 6522
rect 97918 6470 97970 6522
rect 95958 6414 96010 6466
rect 100214 6526 100266 6578
rect 98366 6470 98418 6522
rect 101054 6470 101106 6522
rect 110406 6526 110458 6578
rect 112310 6526 112362 6578
rect 134374 6638 134426 6690
rect 135830 6638 135882 6690
rect 136950 6638 137002 6690
rect 137174 6638 137226 6690
rect 131406 6582 131458 6634
rect 101614 6470 101666 6522
rect 104918 6470 104970 6522
rect 107662 6470 107714 6522
rect 113710 6470 113762 6522
rect 109286 6414 109338 6466
rect 111302 6414 111354 6466
rect 122502 6526 122554 6578
rect 118750 6470 118802 6522
rect 123118 6470 123170 6522
rect 126310 6526 126362 6578
rect 128438 6526 128490 6578
rect 130790 6526 130842 6578
rect 142326 6638 142378 6690
rect 144342 6638 144394 6690
rect 146358 6638 146410 6690
rect 150278 6638 150330 6690
rect 139694 6582 139746 6634
rect 123566 6470 123618 6522
rect 133814 6526 133866 6578
rect 135382 6526 135434 6578
rect 151734 6638 151786 6690
rect 153078 6638 153130 6690
rect 150782 6582 150834 6634
rect 131854 6470 131906 6522
rect 140982 6526 141034 6578
rect 142998 6526 143050 6578
rect 145350 6526 145402 6578
rect 139246 6470 139298 6522
rect 146750 6470 146802 6522
rect 147198 6470 147250 6522
rect 149270 6526 149322 6578
rect 155990 6638 156042 6690
rect 156774 6638 156826 6690
rect 158230 6638 158282 6690
rect 159350 6638 159402 6690
rect 161142 6638 161194 6690
rect 153694 6582 153746 6634
rect 167638 6638 167690 6690
rect 169206 6657 169258 6709
rect 180462 6694 180514 6746
rect 171222 6638 171274 6690
rect 174470 6638 174522 6690
rect 176150 6638 176202 6690
rect 177942 6638 177994 6690
rect 163326 6582 163378 6634
rect 147646 6470 147698 6522
rect 155430 6526 155482 6578
rect 159014 6526 159066 6578
rect 162486 6526 162538 6578
rect 178838 6582 178890 6634
rect 182982 6638 183034 6690
rect 184494 6638 184546 6690
rect 185670 6638 185722 6690
rect 189478 6638 189530 6690
rect 190654 6638 190706 6690
rect 193118 6694 193170 6746
rect 195694 6694 195746 6746
rect 196814 6694 196866 6746
rect 179678 6582 179730 6634
rect 151118 6470 151170 6522
rect 163662 6470 163714 6522
rect 154534 6414 154586 6466
rect 164558 6470 164610 6522
rect 165006 6470 165058 6522
rect 166854 6470 166906 6522
rect 186342 6526 186394 6578
rect 179174 6470 179226 6522
rect 188694 6526 188746 6578
rect 187462 6470 187514 6522
rect 190542 6470 190594 6522
rect 191214 6470 191266 6522
rect 191326 6526 191378 6578
rect 191774 6582 191826 6634
rect 192222 6470 192274 6522
rect 192670 6470 192722 6522
rect 193566 6470 193618 6522
rect 194238 6470 194290 6522
rect 194350 6526 194402 6578
rect 196366 6582 196418 6634
rect 200902 6638 200954 6690
rect 202582 6638 202634 6690
rect 205270 6694 205322 6746
rect 197262 6582 197314 6634
rect 206502 6638 206554 6690
rect 207958 6638 208010 6690
rect 209862 6638 209914 6690
rect 203086 6582 203138 6634
rect 194798 6470 194850 6522
rect 195246 6470 195298 6522
rect 197710 6470 197762 6522
rect 198158 6470 198210 6522
rect 203198 6526 203250 6578
rect 209750 6526 209802 6578
rect 210814 6526 210866 6578
rect 203646 6470 203698 6522
rect 211374 6526 211426 6578
rect 214510 6582 214562 6634
rect 211486 6470 211538 6522
rect 212270 6470 212322 6522
rect 212718 6470 212770 6522
rect 213166 6470 213218 6522
rect 213614 6470 213666 6522
rect 214062 6470 214114 6522
rect 214958 6470 215010 6522
rect 215406 6470 215458 6522
rect 55542 6246 55594 6298
rect 55646 6246 55698 6298
rect 55750 6246 55802 6298
rect 109870 6246 109922 6298
rect 109974 6246 110026 6298
rect 110078 6246 110130 6298
rect 164198 6246 164250 6298
rect 164302 6246 164354 6298
rect 164406 6246 164458 6298
rect 9550 6022 9602 6074
rect 10670 6022 10722 6074
rect 14422 6022 14474 6074
rect 47070 6022 47122 6074
rect 48638 6022 48690 6074
rect 56590 6022 56642 6074
rect 57374 6022 57426 6074
rect 57710 6022 57762 6074
rect 58382 6022 58434 6074
rect 66894 6022 66946 6074
rect 67902 6022 67954 6074
rect 68350 6022 68402 6074
rect 68798 6022 68850 6074
rect 8822 5854 8874 5906
rect 12742 5854 12794 5906
rect 15878 5854 15930 5906
rect 16886 5850 16938 5902
rect 17502 5798 17554 5850
rect 8150 5742 8202 5794
rect 11958 5742 12010 5794
rect 20022 5854 20074 5906
rect 22262 5854 22314 5906
rect 24726 5854 24778 5906
rect 18062 5798 18114 5850
rect 28198 5854 28250 5906
rect 30438 5854 30490 5906
rect 32678 5854 32730 5906
rect 25454 5798 25506 5850
rect 18902 5742 18954 5794
rect 21142 5742 21194 5794
rect 23382 5742 23434 5794
rect 33406 5798 33458 5850
rect 26854 5742 26906 5794
rect 29094 5742 29146 5794
rect 31446 5742 31498 5794
rect 37046 5854 37098 5906
rect 33854 5798 33906 5850
rect 37550 5798 37602 5850
rect 35814 5742 35866 5794
rect 42366 5798 42418 5850
rect 43262 5798 43314 5850
rect 43822 5798 43874 5850
rect 46566 5854 46618 5906
rect 44270 5798 44322 5850
rect 51046 5854 51098 5906
rect 48190 5798 48242 5850
rect 45222 5742 45274 5794
rect 51550 5798 51602 5850
rect 49814 5742 49866 5794
rect 54518 5854 54570 5906
rect 52222 5798 52274 5850
rect 56198 5850 56250 5902
rect 58830 5798 58882 5850
rect 67454 5798 67506 5850
rect 69358 5854 69410 5906
rect 69918 5910 69970 5962
rect 70030 5966 70082 6018
rect 70590 6022 70642 6074
rect 71374 5966 71426 6018
rect 71934 6022 71986 6074
rect 74286 6022 74338 6074
rect 77534 6022 77586 6074
rect 74398 5966 74450 6018
rect 75574 5966 75626 6018
rect 78094 6022 78146 6074
rect 111470 6022 111522 6074
rect 81510 5966 81562 6018
rect 83974 5966 84026 6018
rect 99318 5966 99370 6018
rect 122446 6022 122498 6074
rect 117910 5966 117962 6018
rect 126702 6022 126754 6074
rect 127038 6022 127090 6074
rect 128270 6022 128322 6074
rect 131070 6022 131122 6074
rect 129222 5966 129274 6018
rect 135102 6022 135154 6074
rect 135998 6022 136050 6074
rect 145238 6078 145290 6130
rect 143726 6022 143778 6074
rect 70702 5854 70754 5906
rect 72046 5854 72098 5906
rect 119758 5910 119810 5962
rect 72606 5798 72658 5850
rect 73390 5854 73442 5906
rect 76918 5854 76970 5906
rect 78542 5798 78594 5850
rect 82742 5854 82794 5906
rect 85318 5854 85370 5906
rect 79774 5798 79826 5850
rect 85822 5798 85874 5850
rect 100662 5854 100714 5906
rect 87950 5798 88002 5850
rect 101278 5798 101330 5850
rect 101726 5798 101778 5850
rect 119254 5854 119306 5906
rect 137622 5966 137674 6018
rect 152854 6078 152906 6130
rect 148766 6022 148818 6074
rect 135550 5910 135602 5962
rect 130566 5854 130618 5906
rect 110910 5798 110962 5850
rect 131630 5798 131682 5850
rect 132078 5798 132130 5850
rect 134262 5854 134314 5906
rect 146022 5966 146074 6018
rect 154702 6022 154754 6074
rect 149942 5966 149994 6018
rect 155262 6022 155314 6074
rect 160638 6022 160690 6074
rect 162262 6022 162314 6074
rect 167526 6022 167578 6074
rect 159462 5966 159514 6018
rect 175142 6022 175194 6074
rect 175478 6022 175530 6074
rect 177494 6022 177546 6074
rect 182870 6022 182922 6074
rect 190878 6022 190930 6074
rect 187350 5966 187402 6018
rect 189254 5966 189306 6018
rect 190990 5966 191042 6018
rect 192446 6022 192498 6074
rect 192894 6022 192946 6074
rect 193342 6022 193394 6074
rect 193790 6022 193842 6074
rect 195134 6022 195186 6074
rect 199390 6022 199442 6074
rect 200510 6022 200562 6074
rect 202358 6022 202410 6074
rect 207566 6022 207618 6074
rect 212382 6022 212434 6074
rect 213278 6022 213330 6074
rect 143390 5910 143442 5962
rect 138742 5854 138794 5906
rect 139414 5854 139466 5906
rect 140870 5854 140922 5906
rect 141430 5854 141482 5906
rect 142662 5854 142714 5906
rect 167862 5910 167914 5962
rect 145686 5854 145738 5906
rect 146918 5854 146970 5906
rect 147478 5854 147530 5906
rect 132526 5798 132578 5850
rect 150950 5854 151002 5906
rect 149214 5798 149266 5850
rect 54182 5686 54234 5738
rect 69246 5686 69298 5738
rect 71262 5686 71314 5738
rect 133142 5742 133194 5794
rect 140086 5742 140138 5794
rect 141318 5742 141370 5794
rect 152854 5854 152906 5906
rect 154310 5854 154362 5906
rect 156102 5854 156154 5906
rect 157558 5854 157610 5906
rect 158118 5854 158170 5906
rect 163830 5854 163882 5906
rect 164838 5854 164890 5906
rect 165398 5854 165450 5906
rect 168758 5854 168810 5906
rect 173014 5854 173066 5906
rect 174582 5865 174634 5917
rect 183206 5910 183258 5962
rect 214174 5910 214226 5962
rect 178614 5854 178666 5906
rect 180182 5854 180234 5906
rect 181190 5854 181242 5906
rect 151790 5798 151842 5850
rect 184662 5854 184714 5906
rect 188022 5854 188074 5906
rect 189590 5854 189642 5906
rect 149718 5742 149770 5794
rect 183710 5798 183762 5850
rect 166294 5742 166346 5794
rect 169654 5742 169706 5794
rect 181414 5742 181466 5794
rect 191438 5798 191490 5850
rect 184774 5742 184826 5794
rect 186790 5742 186842 5794
rect 194238 5798 194290 5850
rect 194686 5798 194738 5850
rect 197766 5854 197818 5906
rect 195582 5798 195634 5850
rect 198494 5798 198546 5850
rect 196534 5742 196586 5794
rect 198942 5798 198994 5850
rect 203926 5854 203978 5906
rect 204766 5854 204818 5906
rect 205494 5854 205546 5906
rect 210982 5854 211034 5906
rect 211822 5854 211874 5906
rect 200846 5798 200898 5850
rect 212830 5798 212882 5850
rect 205830 5742 205882 5794
rect 213726 5798 213778 5850
rect 214622 5798 214674 5850
rect 215070 5798 215122 5850
rect 73278 5686 73330 5738
rect 147814 5686 147866 5738
rect 156998 5686 157050 5738
rect 172678 5686 172730 5738
rect 189814 5686 189866 5738
rect 208742 5686 208794 5738
rect 28378 5462 28430 5514
rect 28482 5462 28534 5514
rect 28586 5462 28638 5514
rect 82706 5462 82758 5514
rect 82810 5462 82862 5514
rect 82914 5462 82966 5514
rect 137034 5462 137086 5514
rect 137138 5462 137190 5514
rect 137242 5462 137294 5514
rect 191362 5462 191414 5514
rect 191466 5462 191518 5514
rect 191570 5462 191622 5514
rect 186902 5238 186954 5290
rect 204766 5238 204818 5290
rect 72550 5182 72602 5234
rect 74622 5126 74674 5178
rect 8710 5070 8762 5122
rect 11622 5070 11674 5122
rect 15766 5070 15818 5122
rect 20470 5070 20522 5122
rect 24390 5070 24442 5122
rect 28310 5070 28362 5122
rect 31782 5070 31834 5122
rect 35030 5070 35082 5122
rect 38502 5070 38554 5122
rect 43094 5070 43146 5122
rect 46902 5070 46954 5122
rect 51830 5070 51882 5122
rect 55750 5070 55802 5122
rect 58662 5070 58714 5122
rect 63478 5070 63530 5122
rect 66838 5070 66890 5122
rect 70422 5070 70474 5122
rect 73894 5070 73946 5122
rect 75182 5126 75234 5178
rect 81398 5126 81450 5178
rect 79270 5070 79322 5122
rect 8262 4958 8314 5010
rect 9550 4902 9602 4954
rect 11174 4958 11226 5010
rect 10558 4902 10610 4954
rect 14422 4958 14474 5010
rect 13358 4902 13410 4954
rect 19910 4958 19962 5010
rect 16382 4902 16434 4954
rect 21310 4902 21362 4954
rect 21758 4902 21810 4954
rect 23046 4958 23098 5010
rect 22318 4902 22370 4954
rect 26966 4958 27018 5010
rect 25230 4902 25282 4954
rect 30886 4958 30938 5010
rect 33910 4958 33962 5010
rect 29150 4902 29202 4954
rect 37270 4958 37322 5010
rect 35646 4902 35698 4954
rect 41750 4958 41802 5010
rect 39230 4902 39282 4954
rect 46566 4958 46618 5010
rect 43710 4902 43762 4954
rect 48750 4902 48802 4954
rect 50486 4958 50538 5010
rect 49646 4902 49698 4954
rect 54742 4958 54794 5010
rect 52670 4902 52722 4954
rect 56590 4902 56642 4954
rect 58326 4958 58378 5010
rect 57374 4902 57426 4954
rect 62246 4958 62298 5010
rect 60510 4902 60562 4954
rect 66054 4958 66106 5010
rect 64430 4902 64482 4954
rect 69190 4958 69242 5010
rect 68574 4902 68626 4954
rect 79046 4958 79098 5010
rect 91198 5126 91250 5178
rect 83190 5070 83242 5122
rect 87110 5070 87162 5122
rect 90582 5070 90634 5122
rect 94782 5126 94834 5178
rect 93942 5070 93994 5122
rect 102454 5182 102506 5234
rect 98030 5126 98082 5178
rect 97414 5070 97466 5122
rect 105366 5182 105418 5234
rect 103630 5126 103682 5178
rect 102790 5070 102842 5122
rect 114158 5126 114210 5178
rect 106710 5070 106762 5122
rect 110294 5070 110346 5122
rect 113430 5070 113482 5122
rect 120822 5182 120874 5234
rect 117630 5126 117682 5178
rect 117014 5070 117066 5122
rect 133870 5126 133922 5178
rect 122166 5070 122218 5122
rect 123958 5070 124010 5122
rect 128774 5070 128826 5122
rect 132582 5070 132634 5122
rect 134318 5126 134370 5178
rect 139302 5182 139354 5234
rect 144566 5182 144618 5234
rect 137566 5126 137618 5178
rect 136614 5070 136666 5122
rect 151286 5182 151338 5234
rect 162710 5182 162762 5234
rect 146750 5126 146802 5178
rect 140646 5070 140698 5122
rect 145910 5070 145962 5122
rect 177214 5126 177266 5178
rect 152630 5070 152682 5122
rect 156102 5070 156154 5122
rect 158566 5070 158618 5122
rect 164054 5070 164106 5122
rect 166406 5070 166458 5122
rect 171894 5070 171946 5122
rect 174246 5070 174298 5122
rect 178166 5070 178218 5122
rect 182646 5070 182698 5122
rect 186230 5070 186282 5122
rect 148542 5014 148594 5066
rect 197990 5070 198042 5122
rect 201686 5070 201738 5122
rect 71598 4902 71650 4954
rect 81622 4958 81674 5010
rect 81846 4958 81898 5010
rect 80110 4902 80162 4954
rect 83918 4902 83970 4954
rect 84478 4902 84530 4954
rect 85766 4958 85818 5010
rect 84926 4902 84978 4954
rect 89238 4958 89290 5010
rect 92822 4958 92874 5010
rect 96070 4958 96122 5010
rect 87950 4902 88002 4954
rect 108950 4958 109002 5010
rect 107550 4902 107602 4954
rect 112198 4958 112250 5010
rect 115670 4958 115722 5010
rect 123510 4958 123562 5010
rect 111470 4902 111522 4954
rect 127430 4958 127482 5010
rect 125470 4902 125522 4954
rect 131462 4958 131514 5010
rect 129390 4902 129442 4954
rect 135270 4958 135322 5010
rect 188974 5014 189026 5066
rect 133422 4902 133474 4954
rect 137118 4902 137170 4954
rect 138126 4902 138178 4954
rect 141150 4902 141202 4954
rect 141598 4902 141650 4954
rect 142158 4902 142210 4954
rect 142830 4902 142882 4954
rect 143278 4902 143330 4954
rect 143614 4902 143666 4954
rect 147086 4902 147138 4954
rect 147646 4902 147698 4954
rect 148094 4902 148146 4954
rect 148878 4902 148930 4954
rect 149438 4902 149490 4954
rect 149774 4902 149826 4954
rect 153134 4902 153186 4954
rect 153582 4902 153634 4954
rect 154478 4902 154530 4954
rect 154926 4902 154978 4954
rect 156214 4958 156266 5010
rect 158678 4958 158730 5010
rect 155374 4902 155426 4954
rect 160750 4902 160802 4954
rect 161086 4902 161138 4954
rect 161534 4902 161586 4954
rect 164558 4902 164610 4954
rect 165118 4902 165170 4954
rect 166518 4958 166570 5010
rect 165454 4902 165506 4954
rect 168646 4902 168698 4954
rect 168982 4902 169034 4954
rect 170438 4958 170490 5010
rect 169486 4902 169538 4954
rect 172678 4902 172730 4954
rect 174358 4958 174410 5010
rect 173014 4902 173066 4954
rect 176374 4902 176426 4954
rect 178278 4958 178330 5010
rect 176710 4902 176762 4954
rect 180294 4902 180346 4954
rect 180630 4902 180682 4954
rect 182198 4958 182250 5010
rect 181134 4902 181186 4954
rect 184214 4902 184266 4954
rect 184550 4902 184602 4954
rect 186118 4958 186170 5010
rect 205606 5070 205658 5122
rect 204654 5014 204706 5066
rect 185166 4902 185218 4954
rect 188022 4902 188074 4954
rect 188358 4902 188410 4954
rect 188862 4902 188914 4954
rect 189758 4902 189810 4954
rect 190206 4902 190258 4954
rect 190654 4902 190706 4954
rect 191102 4902 191154 4954
rect 191550 4902 191602 4954
rect 191998 4902 192050 4954
rect 192446 4902 192498 4954
rect 192894 4902 192946 4954
rect 193678 4902 193730 4954
rect 194126 4902 194178 4954
rect 194574 4902 194626 4954
rect 195022 4902 195074 4954
rect 195470 4902 195522 4954
rect 195918 4902 195970 4954
rect 196366 4902 196418 4954
rect 197878 4958 197930 5010
rect 196814 4902 196866 4954
rect 199838 4902 199890 4954
rect 200286 4902 200338 4954
rect 201798 4958 201850 5010
rect 207790 5014 207842 5066
rect 200734 4902 200786 4954
rect 205718 4958 205770 5010
rect 208574 5014 208626 5066
rect 211094 5070 211146 5122
rect 203758 4902 203810 4954
rect 207902 4902 207954 4954
rect 209638 4958 209690 5010
rect 208462 4902 208514 4954
rect 211598 4902 211650 4954
rect 212046 4902 212098 4954
rect 212494 4902 212546 4954
rect 213278 4902 213330 4954
rect 213726 4902 213778 4954
rect 214174 4902 214226 4954
rect 214622 4902 214674 4954
rect 215070 4902 215122 4954
rect 215518 4902 215570 4954
rect 55542 4678 55594 4730
rect 55646 4678 55698 4730
rect 55750 4678 55802 4730
rect 109870 4678 109922 4730
rect 109974 4678 110026 4730
rect 110078 4678 110130 4730
rect 164198 4678 164250 4730
rect 164302 4678 164354 4730
rect 164406 4678 164458 4730
rect 37718 4454 37770 4506
rect 36150 4342 36202 4394
rect 67958 4342 68010 4394
rect 68574 4454 68626 4506
rect 70422 4454 70474 4506
rect 71598 4454 71650 4506
rect 72102 4454 72154 4506
rect 75686 4454 75738 4506
rect 75910 4454 75962 4506
rect 79606 4454 79658 4506
rect 70646 4342 70698 4394
rect 70870 4342 70922 4394
rect 96070 4454 96122 4506
rect 96294 4454 96346 4506
rect 99766 4454 99818 4506
rect 100102 4454 100154 4506
rect 102006 4454 102058 4506
rect 102342 4454 102394 4506
rect 115670 4454 115722 4506
rect 116006 4454 116058 4506
rect 117798 4454 117850 4506
rect 118022 4454 118074 4506
rect 123510 4454 123562 4506
rect 123958 4454 124010 4506
rect 125470 4454 125522 4506
rect 128438 4454 128490 4506
rect 133590 4454 133642 4506
rect 138294 4454 138346 4506
rect 141990 4454 142042 4506
rect 142438 4454 142490 4506
rect 145462 4454 145514 4506
rect 145686 4454 145738 4506
rect 149494 4454 149546 4506
rect 79830 4342 79882 4394
rect 80054 4342 80106 4394
rect 80278 4342 80330 4394
rect 81398 4342 81450 4394
rect 82294 4342 82346 4394
rect 115894 4342 115946 4394
rect 116118 4342 116170 4394
rect 120038 4342 120090 4394
rect 120374 4342 120426 4394
rect 36710 4230 36762 4282
rect 104694 4230 104746 4282
rect 104918 4230 104970 4282
rect 109062 4230 109114 4282
rect 109398 4230 109450 4282
rect 113990 4230 114042 4282
rect 114326 4230 114378 4282
rect 116342 4230 116394 4282
rect 117014 4230 117066 4282
rect 119926 4230 119978 4282
rect 120262 4230 120314 4282
rect 37382 4118 37434 4170
rect 120374 4118 120426 4170
rect 57094 4006 57146 4058
rect 58326 4006 58378 4058
rect 58662 4006 58714 4058
rect 59446 4006 59498 4058
rect 49590 3894 49642 3946
rect 65494 4006 65546 4058
rect 65382 3894 65434 3946
rect 67958 3894 68010 3946
rect 75350 3894 75402 3946
rect 75574 4006 75626 4058
rect 81846 4006 81898 4058
rect 82070 4006 82122 4058
rect 85654 4006 85706 4058
rect 85878 4006 85930 4058
rect 89238 4006 89290 4058
rect 89462 4006 89514 4058
rect 91254 4006 91306 4058
rect 77366 3894 77418 3946
rect 77590 3894 77642 3946
rect 78038 3894 78090 3946
rect 78262 3894 78314 3946
rect 80838 3894 80890 3946
rect 81398 3894 81450 3946
rect 83750 3894 83802 3946
rect 84086 3894 84138 3946
rect 98198 4006 98250 4058
rect 98422 4006 98474 4058
rect 99318 4006 99370 4058
rect 99542 4006 99594 4058
rect 91702 3894 91754 3946
rect 102566 4006 102618 4058
rect 55078 3782 55130 3834
rect 56646 3782 56698 3834
rect 52502 3670 52554 3722
rect 66502 3782 66554 3834
rect 67062 3782 67114 3834
rect 78710 3782 78762 3834
rect 79830 3782 79882 3834
rect 81734 3782 81786 3834
rect 82294 3782 82346 3834
rect 102006 3782 102058 3834
rect 102902 3894 102954 3946
rect 103462 4006 103514 4058
rect 104134 4006 104186 4058
rect 105814 4006 105866 4058
rect 120150 4006 120202 4058
rect 114774 3894 114826 3946
rect 115334 3894 115386 3946
rect 121606 4118 121658 4170
rect 121830 4342 121882 4394
rect 122614 4342 122666 4394
rect 124294 4342 124346 4394
rect 133254 4342 133306 4394
rect 140310 4342 140362 4394
rect 143278 4342 143330 4394
rect 143558 4342 143610 4394
rect 180294 4454 180346 4506
rect 121942 4230 121994 4282
rect 122838 4230 122890 4282
rect 124182 4230 124234 4282
rect 176374 4342 176426 4394
rect 156102 4230 156154 4282
rect 184214 4230 184266 4282
rect 127430 4118 127482 4170
rect 127878 4118 127930 4170
rect 131798 4118 131850 4170
rect 132022 4118 132074 4170
rect 136166 4118 136218 4170
rect 137734 4118 137786 4170
rect 139414 4118 139466 4170
rect 140646 4118 140698 4170
rect 141206 4118 141258 4170
rect 143334 4118 143386 4170
rect 148262 4118 148314 4170
rect 153414 4118 153466 4170
rect 187014 4118 187066 4170
rect 121158 4006 121210 4058
rect 134150 4006 134202 4058
rect 135830 4006 135882 4058
rect 138182 4006 138234 4058
rect 144006 4006 144058 4058
rect 145462 4006 145514 4058
rect 148150 4006 148202 4058
rect 150054 4006 150106 4058
rect 152630 4006 152682 4058
rect 159126 4006 159178 4058
rect 161030 4006 161082 4058
rect 166406 4006 166458 4058
rect 190150 4006 190202 4058
rect 191270 4006 191322 4058
rect 193062 4006 193114 4058
rect 59670 3670 59722 3722
rect 66726 3670 66778 3722
rect 67174 3670 67226 3722
rect 77142 3670 77194 3722
rect 77366 3670 77418 3722
rect 78598 3670 78650 3722
rect 78822 3670 78874 3722
rect 83078 3670 83130 3722
rect 83414 3670 83466 3722
rect 99430 3670 99482 3722
rect 43430 3558 43482 3610
rect 63926 3558 63978 3610
rect 68406 3558 68458 3610
rect 79270 3558 79322 3610
rect 31894 3446 31946 3498
rect 77366 3446 77418 3498
rect 33014 3334 33066 3386
rect 21590 3222 21642 3274
rect 56198 3222 56250 3274
rect 27526 3110 27578 3162
rect 57878 3110 57930 3162
rect 58102 3110 58154 3162
rect 68966 3222 69018 3274
rect 69414 3222 69466 3274
rect 78822 3334 78874 3386
rect 79046 3446 79098 3498
rect 80390 3558 80442 3610
rect 85430 3558 85482 3610
rect 86214 3558 86266 3610
rect 89238 3558 89290 3610
rect 89574 3558 89626 3610
rect 98422 3558 98474 3610
rect 98646 3558 98698 3610
rect 102678 3670 102730 3722
rect 104134 3670 104186 3722
rect 110630 3670 110682 3722
rect 112758 3670 112810 3722
rect 113206 3670 113258 3722
rect 113654 3670 113706 3722
rect 113878 3670 113930 3722
rect 114102 3670 114154 3722
rect 114550 3782 114602 3834
rect 115446 3782 115498 3834
rect 115782 3782 115834 3834
rect 100998 3558 101050 3610
rect 102342 3558 102394 3610
rect 104022 3558 104074 3610
rect 112646 3558 112698 3610
rect 113990 3558 114042 3610
rect 114214 3558 114266 3610
rect 115110 3670 115162 3722
rect 118582 3670 118634 3722
rect 118806 3782 118858 3834
rect 134262 3894 134314 3946
rect 139190 3894 139242 3946
rect 140422 3894 140474 3946
rect 141542 3894 141594 3946
rect 145350 3894 145402 3946
rect 149158 3894 149210 3946
rect 174246 3894 174298 3946
rect 194182 3894 194234 3946
rect 131238 3782 131290 3834
rect 134374 3782 134426 3834
rect 147926 3782 147978 3834
rect 158790 3782 158842 3834
rect 159462 3782 159514 3834
rect 171894 3782 171946 3834
rect 191494 3782 191546 3834
rect 78710 3222 78762 3274
rect 66614 3110 66666 3162
rect 78934 3110 78986 3162
rect 79718 3334 79770 3386
rect 84422 3446 84474 3498
rect 84646 3446 84698 3498
rect 92822 3446 92874 3498
rect 93158 3446 93210 3498
rect 103462 3446 103514 3498
rect 104694 3446 104746 3498
rect 91702 3334 91754 3386
rect 91926 3334 91978 3386
rect 94390 3334 94442 3386
rect 96854 3334 96906 3386
rect 101110 3334 101162 3386
rect 102342 3334 102394 3386
rect 111638 3334 111690 3386
rect 111862 3446 111914 3498
rect 113542 3446 113594 3498
rect 114438 3446 114490 3498
rect 114886 3446 114938 3498
rect 115222 3446 115274 3498
rect 116902 3446 116954 3498
rect 117126 3446 117178 3498
rect 119702 3446 119754 3498
rect 120374 3446 120426 3498
rect 120598 3670 120650 3722
rect 132358 3670 132410 3722
rect 134038 3670 134090 3722
rect 134822 3670 134874 3722
rect 135046 3670 135098 3722
rect 143558 3670 143610 3722
rect 144006 3670 144058 3722
rect 146134 3670 146186 3722
rect 153078 3670 153130 3722
rect 153302 3670 153354 3722
rect 121158 3558 121210 3610
rect 131462 3558 131514 3610
rect 132022 3558 132074 3610
rect 121494 3446 121546 3498
rect 122166 3446 122218 3498
rect 127878 3446 127930 3498
rect 130902 3446 130954 3498
rect 133478 3446 133530 3498
rect 113990 3334 114042 3386
rect 115782 3334 115834 3386
rect 116230 3334 116282 3386
rect 38502 2998 38554 3050
rect 65270 2998 65322 3050
rect 65494 2998 65546 3050
rect 78486 2998 78538 3050
rect 78710 2998 78762 3050
rect 79046 2998 79098 3050
rect 51942 2886 51994 2938
rect 85206 3222 85258 3274
rect 85430 3222 85482 3274
rect 93158 3222 93210 3274
rect 94166 3222 94218 3274
rect 95734 3222 95786 3274
rect 96070 3222 96122 3274
rect 79606 3110 79658 3162
rect 81510 3110 81562 3162
rect 81958 3110 82010 3162
rect 82406 3110 82458 3162
rect 82966 3110 83018 3162
rect 83190 3110 83242 3162
rect 90918 3110 90970 3162
rect 91478 3110 91530 3162
rect 100662 3110 100714 3162
rect 117350 3222 117402 3274
rect 117686 3334 117738 3386
rect 132806 3334 132858 3386
rect 141094 3558 141146 3610
rect 151062 3558 151114 3610
rect 152406 3558 152458 3610
rect 156326 3558 156378 3610
rect 140982 3446 141034 3498
rect 140198 3334 140250 3386
rect 143110 3334 143162 3386
rect 147814 3446 147866 3498
rect 154870 3446 154922 3498
rect 156438 3446 156490 3498
rect 189478 3446 189530 3498
rect 152518 3334 152570 3386
rect 152854 3334 152906 3386
rect 187574 3334 187626 3386
rect 150390 3222 150442 3274
rect 178950 3222 179002 3274
rect 191606 3222 191658 3274
rect 101782 3110 101834 3162
rect 107830 3110 107882 3162
rect 108502 3110 108554 3162
rect 117574 3110 117626 3162
rect 117798 3110 117850 3162
rect 119142 3110 119194 3162
rect 119590 3110 119642 3162
rect 120038 3110 120090 3162
rect 138630 3110 138682 3162
rect 79718 2998 79770 3050
rect 80166 2998 80218 3050
rect 80950 2998 81002 3050
rect 82630 2998 82682 3050
rect 82854 2998 82906 3050
rect 79606 2886 79658 2938
rect 82294 2886 82346 2938
rect 82518 2886 82570 2938
rect 84310 2886 84362 2938
rect 84534 2998 84586 3050
rect 85094 2998 85146 3050
rect 85318 2998 85370 3050
rect 91926 2998 91978 3050
rect 92150 2998 92202 3050
rect 99878 2998 99930 3050
rect 100214 2998 100266 3050
rect 102454 2998 102506 3050
rect 102902 2998 102954 3050
rect 104022 2998 104074 3050
rect 104246 2998 104298 3050
rect 116454 2998 116506 3050
rect 117350 2998 117402 3050
rect 90694 2886 90746 2938
rect 90918 2886 90970 2938
rect 95958 2886 96010 2938
rect 96182 2886 96234 2938
rect 99318 2886 99370 2938
rect 27526 2774 27578 2826
rect 58662 2774 58714 2826
rect 61686 2774 61738 2826
rect 99094 2774 99146 2826
rect 23270 2662 23322 2714
rect 67398 2662 67450 2714
rect 22038 2550 22090 2602
rect 58102 2550 58154 2602
rect 58886 2550 58938 2602
rect 66278 2550 66330 2602
rect 66614 2550 66666 2602
rect 79046 2662 79098 2714
rect 79494 2662 79546 2714
rect 100326 2774 100378 2826
rect 100662 2774 100714 2826
rect 99766 2662 99818 2714
rect 101110 2886 101162 2938
rect 132470 2886 132522 2938
rect 101894 2774 101946 2826
rect 110854 2774 110906 2826
rect 68182 2550 68234 2602
rect 79606 2550 79658 2602
rect 80166 2550 80218 2602
rect 100214 2550 100266 2602
rect 110742 2662 110794 2714
rect 104918 2550 104970 2602
rect 105142 2550 105194 2602
rect 115894 2774 115946 2826
rect 116902 2774 116954 2826
rect 117798 2774 117850 2826
rect 118470 2774 118522 2826
rect 133478 2998 133530 3050
rect 151510 3110 151562 3162
rect 161030 3110 161082 3162
rect 207734 3110 207786 3162
rect 150726 2998 150778 3050
rect 132806 2886 132858 2938
rect 153078 2886 153130 2938
rect 154982 2998 155034 3050
rect 189926 2998 189978 3050
rect 192278 2998 192330 3050
rect 186118 2886 186170 2938
rect 111190 2662 111242 2714
rect 117462 2662 117514 2714
rect 117686 2662 117738 2714
rect 126758 2662 126810 2714
rect 111078 2550 111130 2602
rect 154422 2774 154474 2826
rect 127318 2662 127370 2714
rect 162710 2774 162762 2826
rect 186006 2774 186058 2826
rect 186454 2774 186506 2826
rect 186566 2662 186618 2714
rect 201574 2662 201626 2714
rect 21478 2438 21530 2490
rect 65382 2438 65434 2490
rect 65942 2438 65994 2490
rect 174358 2550 174410 2602
rect 175030 2550 175082 2602
rect 196422 2550 196474 2602
rect 37942 2326 37994 2378
rect 62022 2326 62074 2378
rect 51382 2214 51434 2266
rect 61910 2214 61962 2266
rect 62134 2214 62186 2266
rect 70310 2326 70362 2378
rect 70534 2326 70586 2378
rect 73446 2326 73498 2378
rect 62918 2214 62970 2266
rect 76246 2326 76298 2378
rect 76470 2326 76522 2378
rect 77814 2326 77866 2378
rect 78934 2326 78986 2378
rect 81958 2326 82010 2378
rect 82182 2326 82234 2378
rect 94166 2326 94218 2378
rect 74006 2214 74058 2266
rect 75126 2214 75178 2266
rect 49478 2102 49530 2154
rect 59670 2102 59722 2154
rect 59894 2102 59946 2154
rect 75910 2214 75962 2266
rect 83862 2214 83914 2266
rect 84198 2214 84250 2266
rect 93942 2214 93994 2266
rect 100438 2326 100490 2378
rect 101558 2326 101610 2378
rect 126422 2326 126474 2378
rect 34918 1990 34970 2042
rect 68182 1990 68234 2042
rect 68630 1990 68682 2042
rect 75910 1990 75962 2042
rect 76358 2102 76410 2154
rect 83750 2102 83802 2154
rect 83974 2102 84026 2154
rect 95734 2214 95786 2266
rect 125862 2214 125914 2266
rect 126758 2326 126810 2378
rect 134262 2326 134314 2378
rect 130902 2214 130954 2266
rect 138630 2438 138682 2490
rect 152294 2438 152346 2490
rect 152630 2438 152682 2490
rect 154198 2438 154250 2490
rect 154534 2438 154586 2490
rect 204598 2438 204650 2490
rect 151286 2326 151338 2378
rect 183094 2326 183146 2378
rect 185894 2326 185946 2378
rect 190598 2326 190650 2378
rect 153862 2214 153914 2266
rect 155654 2214 155706 2266
rect 189366 2214 189418 2266
rect 88902 1990 88954 2042
rect 89126 1990 89178 2042
rect 89910 1990 89962 2042
rect 90694 1990 90746 2042
rect 95846 2102 95898 2154
rect 96294 2102 96346 2154
rect 101782 2102 101834 2154
rect 102566 2102 102618 2154
rect 115446 2102 115498 2154
rect 116006 2102 116058 2154
rect 117014 2102 117066 2154
rect 117238 2102 117290 2154
rect 119366 2102 119418 2154
rect 119590 2102 119642 2154
rect 126310 2102 126362 2154
rect 127654 2102 127706 2154
rect 150278 2102 150330 2154
rect 154422 2102 154474 2154
rect 188694 2102 188746 2154
rect 94502 1990 94554 2042
rect 61126 1878 61178 1930
rect 62806 1878 62858 1930
rect 64710 1878 64762 1930
rect 101110 1878 101162 1930
rect 179062 1990 179114 2042
rect 102342 1878 102394 1930
rect 151062 1878 151114 1930
rect 63590 1766 63642 1818
rect 100662 1766 100714 1818
rect 100998 1766 101050 1818
rect 102454 1766 102506 1818
rect 58102 1654 58154 1706
rect 65158 1654 65210 1706
rect 65382 1654 65434 1706
rect 100550 1654 100602 1706
rect 136390 1766 136442 1818
rect 155990 1766 156042 1818
rect 156438 1766 156490 1818
rect 32342 1542 32394 1594
rect 75462 1542 75514 1594
rect 76806 1542 76858 1594
rect 78262 1542 78314 1594
rect 78486 1542 78538 1594
rect 82854 1542 82906 1594
rect 36374 1430 36426 1482
rect 74790 1430 74842 1482
rect 75574 1430 75626 1482
rect 83414 1430 83466 1482
rect 46006 1318 46058 1370
rect 82070 1318 82122 1370
rect 82406 1318 82458 1370
rect 82742 1318 82794 1370
rect 84758 1542 84810 1594
rect 85094 1542 85146 1594
rect 88454 1542 88506 1594
rect 88790 1542 88842 1594
rect 92150 1542 92202 1594
rect 92374 1542 92426 1594
rect 97638 1542 97690 1594
rect 98310 1542 98362 1594
rect 100326 1542 100378 1594
rect 83974 1430 84026 1482
rect 102902 1654 102954 1706
rect 100774 1542 100826 1594
rect 101782 1542 101834 1594
rect 102006 1542 102058 1594
rect 105254 1542 105306 1594
rect 105926 1542 105978 1594
rect 106934 1542 106986 1594
rect 107494 1654 107546 1706
rect 108166 1654 108218 1706
rect 150278 1654 150330 1706
rect 108390 1542 108442 1594
rect 109958 1542 110010 1594
rect 84422 1318 84474 1370
rect 90582 1318 90634 1370
rect 91254 1318 91306 1370
rect 94614 1318 94666 1370
rect 97414 1318 97466 1370
rect 106710 1430 106762 1482
rect 109734 1430 109786 1482
rect 112646 1542 112698 1594
rect 112870 1542 112922 1594
rect 100886 1318 100938 1370
rect 117350 1430 117402 1482
rect 118022 1542 118074 1594
rect 120262 1542 120314 1594
rect 120486 1542 120538 1594
rect 123398 1542 123450 1594
rect 123622 1542 123674 1594
rect 132470 1542 132522 1594
rect 144790 1542 144842 1594
rect 147478 1542 147530 1594
rect 118134 1430 118186 1482
rect 119814 1430 119866 1482
rect 136502 1430 136554 1482
rect 111414 1318 111466 1370
rect 116678 1318 116730 1370
rect 117014 1318 117066 1370
rect 119478 1318 119530 1370
rect 119702 1318 119754 1370
rect 120486 1318 120538 1370
rect 120710 1318 120762 1370
rect 121606 1318 121658 1370
rect 122950 1318 123002 1370
rect 135046 1318 135098 1370
rect 44774 1206 44826 1258
rect 69974 1206 70026 1258
rect 70534 1206 70586 1258
rect 10166 1094 10218 1146
rect 71990 1094 72042 1146
rect 75126 1094 75178 1146
rect 81734 1094 81786 1146
rect 81958 1094 82010 1146
rect 84086 1094 84138 1146
rect 85430 1094 85482 1146
rect 86774 1094 86826 1146
rect 87222 1094 87274 1146
rect 87446 1094 87498 1146
rect 87894 1094 87946 1146
rect 89686 1094 89738 1146
rect 89910 1094 89962 1146
rect 97974 1094 98026 1146
rect 100774 1094 100826 1146
rect 101446 1094 101498 1146
rect 101782 1094 101834 1146
rect 110294 1094 110346 1146
rect 111078 1094 111130 1146
rect 111862 1094 111914 1146
rect 112086 1094 112138 1146
rect 114662 1094 114714 1146
rect 42534 982 42586 1034
rect 74902 982 74954 1034
rect 75238 982 75290 1034
rect 77254 982 77306 1034
rect 5574 870 5626 922
rect 13526 870 13578 922
rect 37270 870 37322 922
rect 43430 870 43482 922
rect 63702 870 63754 922
rect 63926 870 63978 922
rect 68966 870 69018 922
rect 71430 870 71482 922
rect 81286 982 81338 1034
rect 81510 982 81562 1034
rect 82742 982 82794 1034
rect 83526 982 83578 1034
rect 84870 982 84922 1034
rect 86998 982 87050 1034
rect 92150 982 92202 1034
rect 96630 982 96682 1034
rect 96854 982 96906 1034
rect 77926 870 77978 922
rect 88230 870 88282 922
rect 88454 870 88506 922
rect 90358 870 90410 922
rect 98534 870 98586 922
rect 99430 982 99482 1034
rect 106150 982 106202 1034
rect 106374 982 106426 1034
rect 99878 870 99930 922
rect 100998 870 101050 922
rect 109734 870 109786 922
rect 110742 982 110794 1034
rect 111638 982 111690 1034
rect 112646 982 112698 1034
rect 117910 1094 117962 1146
rect 118470 1094 118522 1146
rect 121270 1094 121322 1146
rect 121718 1094 121770 1146
rect 125302 1094 125354 1146
rect 125526 1094 125578 1146
rect 126310 1094 126362 1146
rect 202582 1094 202634 1146
rect 114886 982 114938 1034
rect 116454 982 116506 1034
rect 116790 982 116842 1034
rect 130006 982 130058 1034
rect 133926 982 133978 1034
rect 193398 982 193450 1034
rect 116118 870 116170 922
rect 118246 870 118298 922
rect 218374 870 218426 922
rect 28982 758 29034 810
rect 16214 646 16266 698
rect 7254 534 7306 586
rect 33910 534 33962 586
rect 69974 758 70026 810
rect 76134 758 76186 810
rect 76694 758 76746 810
rect 77142 758 77194 810
rect 77366 758 77418 810
rect 81510 758 81562 810
rect 70422 646 70474 698
rect 77926 646 77978 698
rect 78374 646 78426 698
rect 82070 758 82122 810
rect 82742 758 82794 810
rect 83862 758 83914 810
rect 82070 534 82122 586
rect 85318 646 85370 698
rect 85766 758 85818 810
rect 196198 758 196250 810
rect 215686 758 215738 810
rect 8934 422 8986 474
rect 42534 422 42586 474
rect 49926 422 49978 474
rect 68742 422 68794 474
rect 69302 422 69354 474
rect 81398 422 81450 474
rect 195414 534 195466 586
rect 24278 310 24330 362
rect 73558 310 73610 362
rect 74902 310 74954 362
rect 216134 422 216186 474
rect 207062 310 207114 362
rect 21310 198 21362 250
rect 66838 198 66890 250
rect 68854 198 68906 250
rect 77366 198 77418 250
rect 77814 198 77866 250
rect 83862 198 83914 250
rect 84086 198 84138 250
rect 215014 198 215066 250
rect 17614 86 17666 138
rect 54742 86 54794 138
rect 56534 86 56586 138
rect 208294 86 208346 138
<< metal2 >>
rect 280 14200 392 15000
rect 952 14200 1064 15000
rect 1736 14200 1848 15000
rect 2408 14200 2520 15000
rect 3192 14200 3304 15000
rect 3864 14200 3976 15000
rect 4648 14200 4760 15000
rect 5320 14200 5432 15000
rect 6104 14200 6216 15000
rect 6776 14200 6888 15000
rect 7560 14200 7672 15000
rect 8232 14200 8344 15000
rect 8484 14362 8540 14374
rect 8484 14310 8486 14362
rect 8538 14310 8540 14362
rect 308 13356 364 14200
rect 308 13290 364 13300
rect 980 13244 1036 14200
rect 1764 14140 1820 14200
rect 1876 14140 1932 14150
rect 1764 14138 1932 14140
rect 1764 14086 1878 14138
rect 1930 14086 1932 14138
rect 1764 14084 1932 14086
rect 1876 14074 1932 14084
rect 980 13178 1036 13188
rect 84 13130 140 13142
rect 84 13078 86 13130
rect 138 13078 140 13130
rect 84 7980 140 13078
rect 2436 12348 2492 14200
rect 3220 13020 3276 14200
rect 3892 13132 3948 14200
rect 3892 13066 3948 13076
rect 3220 12954 3276 12964
rect 2436 12282 2492 12292
rect 4676 12234 4732 14200
rect 5348 12794 5404 14200
rect 6132 12908 6188 14200
rect 6804 13690 6860 14200
rect 7588 14140 7644 14200
rect 7700 14140 7756 14150
rect 7588 14084 7700 14140
rect 8260 14140 8316 14200
rect 8484 14140 8540 14310
rect 9016 14200 9128 15000
rect 9492 14698 9548 14710
rect 9492 14646 9494 14698
rect 9546 14646 9548 14698
rect 9492 14364 9548 14646
rect 9268 14308 9548 14364
rect 8260 14084 8540 14140
rect 9044 14140 9100 14200
rect 9268 14140 9324 14308
rect 9688 14200 9800 15000
rect 10052 14586 10108 14598
rect 10052 14534 10054 14586
rect 10106 14534 10108 14586
rect 10052 14364 10108 14534
rect 9940 14308 10108 14364
rect 9044 14084 9324 14140
rect 9716 14140 9772 14200
rect 9940 14140 9996 14308
rect 10472 14200 10584 15000
rect 11144 14200 11256 15000
rect 11620 14922 11676 14934
rect 11620 14870 11622 14922
rect 11674 14870 11676 14922
rect 11620 14364 11676 14870
rect 11396 14308 11676 14364
rect 9716 14084 9996 14140
rect 7700 14074 7756 14084
rect 6804 13638 6806 13690
rect 6858 13638 6860 13690
rect 6804 13626 6860 13638
rect 10500 13580 10556 14200
rect 11172 14140 11228 14200
rect 11396 14140 11452 14308
rect 11928 14200 12040 15000
rect 12600 14200 12712 15000
rect 13384 14200 13496 15000
rect 14056 14200 14168 15000
rect 14840 14200 14952 15000
rect 15512 14200 15624 15000
rect 16296 14200 16408 15000
rect 16660 14476 16716 14486
rect 16660 14364 16716 14420
rect 16548 14308 16716 14364
rect 11172 14084 11452 14140
rect 10500 13514 10556 13524
rect 10612 13356 10668 13366
rect 6132 12842 6188 12852
rect 9828 13020 9884 13030
rect 5348 12742 5350 12794
rect 5402 12742 5404 12794
rect 5348 12730 5404 12742
rect 4676 12182 4678 12234
rect 4730 12182 4732 12234
rect 4676 12170 4732 12182
rect 6692 12460 6748 12470
rect 84 7914 140 7924
rect 6468 11002 6524 11014
rect 6468 10950 6470 11002
rect 6522 10950 6524 11002
rect 6468 7642 6524 10950
rect 6692 9772 6748 12404
rect 9716 12348 9772 12358
rect 6692 9706 6748 9716
rect 8316 9772 8372 9782
rect 8316 9678 8372 9716
rect 8876 9660 8932 9670
rect 8876 9566 8932 9604
rect 9716 9210 9772 12292
rect 9828 9994 9884 12964
rect 9828 9942 9830 9994
rect 9882 9942 9884 9994
rect 9828 9930 9884 9942
rect 10164 9660 10220 9670
rect 10164 9566 10220 9604
rect 9716 9158 9718 9210
rect 9770 9158 9772 9210
rect 9716 9146 9772 9158
rect 10612 9210 10668 13300
rect 10724 13244 10780 13254
rect 10724 9994 10780 13188
rect 11620 13132 11676 13142
rect 10724 9942 10726 9994
rect 10778 9942 10780 9994
rect 10724 9930 10780 9942
rect 10836 11004 10892 11014
rect 10612 9158 10614 9210
rect 10666 9158 10668 9210
rect 10612 9146 10668 9158
rect 8988 9100 9044 9110
rect 8988 9006 9044 9044
rect 10052 9100 10108 9110
rect 10052 9006 10108 9044
rect 9716 8428 9772 8438
rect 6468 7590 6470 7642
rect 6522 7590 6524 7642
rect 6468 7578 6524 7590
rect 8932 7644 8988 7654
rect 7924 7474 7980 7486
rect 7924 7422 7926 7474
rect 7978 7422 7980 7474
rect 7924 7308 7980 7422
rect 8932 7474 8988 7588
rect 9548 7644 9604 7654
rect 9548 7550 9604 7588
rect 8932 7422 8934 7474
rect 8986 7422 8988 7474
rect 8932 7410 8988 7422
rect 7924 7242 7980 7252
rect 8764 7308 8820 7318
rect 8764 6522 8820 7252
rect 9716 6524 9772 8372
rect 10276 8316 10332 8326
rect 10276 8222 10332 8260
rect 10332 7420 10388 7430
rect 8764 6470 8766 6522
rect 8818 6470 8820 6522
rect 4452 6412 4508 6422
rect 3780 4844 3836 4854
rect 756 924 812 934
rect 196 868 476 924
rect 196 800 252 868
rect 168 0 280 800
rect 420 588 476 868
rect 756 800 812 868
rect 1316 924 1372 934
rect 1316 800 1372 868
rect 1988 924 2044 934
rect 1988 800 2044 868
rect 2548 924 2604 934
rect 2548 800 2604 868
rect 3220 924 3276 934
rect 3220 800 3276 868
rect 3780 800 3836 4788
rect 4452 800 4508 6356
rect 8764 6300 8820 6470
rect 9548 6468 9772 6524
rect 10276 7364 10332 7420
rect 10276 7288 10388 7364
rect 8764 6244 8988 6300
rect 8820 6076 8876 6086
rect 8820 5906 8876 6020
rect 8820 5854 8822 5906
rect 8874 5854 8876 5906
rect 8820 5842 8876 5854
rect 8148 5794 8204 5806
rect 8148 5742 8150 5794
rect 8202 5742 8204 5794
rect 5012 4732 5068 4742
rect 5012 800 5068 4676
rect 8148 1484 8204 5742
rect 8708 5122 8764 5134
rect 8708 5070 8710 5122
rect 8762 5070 8764 5122
rect 8260 5010 8316 5022
rect 8260 4958 8262 5010
rect 8314 4958 8316 5010
rect 8260 1596 8316 4958
rect 8708 4956 8764 5070
rect 8708 4890 8764 4900
rect 8260 1530 8316 1540
rect 8708 3388 8764 3398
rect 8148 1418 8204 1428
rect 8036 1372 8092 1382
rect 5572 922 5628 934
rect 5572 870 5574 922
rect 5626 870 5628 922
rect 5572 800 5628 870
rect 6244 868 6524 924
rect 6244 800 6300 868
rect 420 532 588 588
rect 532 252 588 532
rect 532 186 588 196
rect 728 0 840 800
rect 1288 0 1400 800
rect 1960 0 2072 800
rect 2520 0 2632 800
rect 3192 0 3304 800
rect 3752 0 3864 800
rect 4424 0 4536 800
rect 4984 0 5096 800
rect 5544 0 5656 800
rect 6216 0 6328 800
rect 6468 700 6524 868
rect 6804 868 7084 924
rect 6804 800 6860 868
rect 6468 644 6636 700
rect 6580 588 6636 644
rect 6580 522 6636 532
rect 6776 0 6888 800
rect 7028 700 7084 868
rect 7476 868 7756 924
rect 7476 800 7532 868
rect 7028 644 7308 700
rect 7252 586 7308 644
rect 7252 534 7254 586
rect 7306 534 7308 586
rect 7252 522 7308 534
rect 7448 0 7560 800
rect 7700 588 7756 868
rect 8036 800 8092 1316
rect 8708 800 8764 3332
rect 7700 532 7868 588
rect 7812 364 7868 532
rect 7812 298 7868 308
rect 8008 0 8120 800
rect 8680 0 8792 800
rect 8932 474 8988 6244
rect 9548 6076 9604 6468
rect 9548 5944 9604 6020
rect 9548 4956 9604 4966
rect 9548 4862 9604 4900
rect 10276 2604 10332 7288
rect 10836 6858 10892 10948
rect 11620 9994 11676 13076
rect 11956 12684 12012 14200
rect 12628 13804 12684 14200
rect 12628 13738 12684 13748
rect 11956 12618 12012 12628
rect 13412 12460 13468 14200
rect 14084 13916 14140 14200
rect 14868 14028 14924 14200
rect 14868 13962 14924 13972
rect 14084 13850 14140 13860
rect 15540 13132 15596 14200
rect 16324 14140 16380 14200
rect 16548 14140 16604 14308
rect 16968 14200 17080 15000
rect 17752 14200 17864 15000
rect 18424 14200 18536 15000
rect 19208 14200 19320 15000
rect 19880 14200 19992 15000
rect 20664 14200 20776 15000
rect 21336 14200 21448 15000
rect 22120 14200 22232 15000
rect 22792 14200 22904 15000
rect 23380 14812 23436 14822
rect 23380 14588 23436 14756
rect 23044 14532 23436 14588
rect 16324 14084 16604 14140
rect 16996 14140 17052 14200
rect 17108 14140 17164 14150
rect 16996 14084 17108 14140
rect 17108 14074 17164 14084
rect 17780 14028 17836 14200
rect 17780 13962 17836 13972
rect 18452 13244 18508 14200
rect 19236 13356 19292 14200
rect 19236 13290 19292 13300
rect 18452 13178 18508 13188
rect 15540 13066 15596 13076
rect 13412 12394 13468 12404
rect 18116 11788 18172 11798
rect 16324 11226 16380 11238
rect 16324 11174 16326 11226
rect 16378 11174 16380 11226
rect 14420 11116 14476 11126
rect 11620 9942 11622 9994
rect 11674 9942 11676 9994
rect 11620 9930 11676 9942
rect 13076 10892 13132 10902
rect 11060 9772 11116 9782
rect 11060 9678 11116 9716
rect 11956 9658 12012 9670
rect 11956 9606 11958 9658
rect 12010 9606 12012 9658
rect 11956 9436 12012 9606
rect 11956 9370 12012 9380
rect 12572 9658 12628 9670
rect 12572 9606 12574 9658
rect 12626 9606 12628 9658
rect 12572 9436 12628 9606
rect 12572 9370 12628 9380
rect 10948 9098 11004 9110
rect 10948 9046 10950 9098
rect 11002 9046 11004 9098
rect 10948 7420 11004 9046
rect 13076 8874 13132 10836
rect 13748 9884 13804 9894
rect 13076 8822 13078 8874
rect 13130 8822 13132 8874
rect 13076 8810 13132 8822
rect 13636 8876 13692 8886
rect 13636 8427 13692 8820
rect 13580 8371 13692 8427
rect 12852 8316 12908 8326
rect 11620 8258 11676 8270
rect 11620 8206 11622 8258
rect 11674 8206 11676 8258
rect 11620 8092 11676 8206
rect 12852 8210 12854 8260
rect 12906 8210 12908 8260
rect 13580 8316 13636 8371
rect 13580 8222 13636 8260
rect 12852 8198 12908 8210
rect 11620 8026 11676 8036
rect 12740 7532 12796 7542
rect 12740 7474 12796 7476
rect 12740 7422 12742 7474
rect 12794 7422 12796 7474
rect 12740 7410 12796 7422
rect 13748 7532 13804 9828
rect 14084 9042 14140 9054
rect 14084 8990 14086 9042
rect 14138 8990 14140 9042
rect 14084 8988 14140 8990
rect 14084 8922 14140 8932
rect 13916 8092 13972 8102
rect 13916 7998 13972 8036
rect 10948 7354 11004 7364
rect 11396 7362 11452 7374
rect 10836 6806 10838 6858
rect 10890 6806 10892 6858
rect 10836 6794 10892 6806
rect 11396 7310 11398 7362
rect 11450 7310 11452 7362
rect 10668 6076 10724 6086
rect 10668 5982 10724 6020
rect 11172 5010 11228 5022
rect 10556 4956 10612 4966
rect 10556 4862 10612 4900
rect 11172 4958 11174 5010
rect 11226 4958 11228 5010
rect 11172 3388 11228 4958
rect 11172 3322 11228 3332
rect 10276 2538 10332 2548
rect 9940 1596 9996 1606
rect 9268 1260 9324 1270
rect 9268 800 9324 1204
rect 9940 800 9996 1540
rect 11060 1596 11116 1606
rect 10500 1484 10556 1494
rect 10164 1148 10220 1158
rect 10164 1054 10220 1092
rect 10500 800 10556 1428
rect 11060 800 11116 1540
rect 11396 1260 11452 7310
rect 13748 7308 13804 7476
rect 13580 7252 13804 7308
rect 11508 6690 11564 6702
rect 11508 6638 11510 6690
rect 11562 6638 11564 6690
rect 11508 4620 11564 6638
rect 12852 6690 12908 6702
rect 12852 6638 12854 6690
rect 12906 6638 12908 6690
rect 12852 6524 12908 6638
rect 13580 6634 13636 7252
rect 13580 6582 13582 6634
rect 13634 6582 13636 6634
rect 13580 6570 13636 6582
rect 12852 6458 12908 6468
rect 14028 6524 14084 6534
rect 14084 6468 14140 6524
rect 14028 6392 14140 6468
rect 12740 6076 12796 6086
rect 12740 5906 12796 6020
rect 12740 5854 12742 5906
rect 12794 5854 12796 5906
rect 12740 5842 12796 5854
rect 11956 5794 12012 5806
rect 11956 5742 11958 5794
rect 12010 5742 12012 5794
rect 11620 5122 11676 5134
rect 11620 5070 11622 5122
rect 11674 5070 11676 5122
rect 11620 4956 11676 5070
rect 11620 4890 11676 4900
rect 11508 4554 11564 4564
rect 11396 1194 11452 1204
rect 11732 1484 11788 1494
rect 11732 800 11788 1428
rect 11956 1372 12012 5742
rect 14084 5292 14140 6392
rect 14420 6074 14476 11060
rect 14868 10668 14924 10678
rect 14868 7306 14924 10612
rect 16212 10108 16268 10118
rect 15596 9772 15652 9782
rect 15092 9212 15148 9222
rect 15092 9042 15148 9156
rect 15596 9212 15652 9716
rect 15596 9080 15652 9156
rect 15092 8990 15094 9042
rect 15146 8990 15148 9042
rect 15092 8978 15148 8990
rect 16044 8988 16100 8998
rect 16044 8427 16100 8932
rect 16044 8371 16156 8427
rect 15876 7474 15932 7486
rect 15876 7422 15878 7474
rect 15930 7422 15932 7474
rect 15876 7420 15932 7422
rect 15876 7354 15932 7364
rect 14868 7254 14870 7306
rect 14922 7254 14924 7306
rect 14868 7242 14924 7254
rect 16100 6188 16156 8371
rect 16212 6858 16268 10052
rect 16324 8426 16380 11174
rect 17780 9212 17836 9222
rect 17780 9118 17836 9156
rect 18116 9210 18172 11732
rect 19908 11788 19964 14200
rect 20692 12122 20748 14200
rect 21364 14140 21420 14200
rect 21476 14140 21532 14150
rect 21364 14084 21476 14140
rect 21476 14074 21532 14084
rect 20692 12070 20694 12122
rect 20746 12070 20748 12122
rect 20692 12058 20748 12070
rect 19908 11722 19964 11732
rect 20244 11788 20300 11798
rect 19908 9324 19964 9334
rect 18116 9158 18118 9210
rect 18170 9158 18172 9210
rect 18116 9146 18172 9158
rect 18508 9212 18564 9222
rect 18508 9118 18564 9156
rect 19908 9210 19964 9268
rect 19908 9158 19910 9210
rect 19962 9158 19964 9210
rect 19908 9146 19964 9158
rect 20244 9210 20300 11732
rect 22148 11788 22204 14200
rect 22820 14140 22876 14200
rect 23044 14140 23100 14532
rect 23576 14200 23688 15000
rect 24248 14200 24360 15000
rect 25032 14200 25144 15000
rect 25704 14200 25816 15000
rect 25956 14308 26348 14364
rect 22820 14084 23100 14140
rect 23604 13244 23660 14200
rect 23604 13178 23660 13188
rect 22148 11722 22204 11732
rect 22260 11900 22316 11910
rect 21812 10890 21868 10902
rect 21812 10838 21814 10890
rect 21866 10838 21868 10890
rect 21588 10442 21644 10454
rect 21588 10390 21590 10442
rect 21642 10390 21644 10442
rect 20244 9158 20246 9210
rect 20298 9158 20300 9210
rect 20244 9146 20300 9158
rect 20636 9324 20692 9334
rect 20636 9210 20692 9268
rect 20636 9158 20638 9210
rect 20690 9158 20692 9210
rect 20636 9146 20692 9158
rect 16324 8374 16326 8426
rect 16378 8374 16380 8426
rect 16324 8362 16380 8374
rect 16660 8258 16716 8270
rect 16660 8206 16662 8258
rect 16714 8206 16716 8258
rect 16660 8092 16716 8206
rect 18340 8258 18396 8270
rect 18340 8206 18342 8258
rect 18394 8206 18396 8258
rect 18340 8092 18396 8206
rect 18732 8092 18788 8102
rect 19180 8092 19236 8102
rect 18340 8090 18844 8092
rect 18340 8038 18734 8090
rect 18786 8038 18844 8090
rect 18340 8036 18844 8038
rect 16660 8026 16716 8036
rect 18732 8026 18844 8036
rect 16884 7470 16940 7482
rect 16884 7418 16886 7470
rect 16938 7418 16940 7470
rect 16884 7308 16940 7418
rect 16884 7242 16940 7252
rect 17612 7418 17668 7430
rect 17612 7366 17614 7418
rect 17666 7366 17668 7418
rect 17612 7308 17668 7366
rect 18060 7420 18116 7430
rect 18620 7420 18676 7430
rect 18060 7326 18116 7364
rect 18452 7364 18620 7420
rect 17612 7242 17668 7252
rect 16212 6806 16214 6858
rect 16266 6806 16268 6858
rect 16212 6794 16268 6806
rect 16660 6690 16716 6702
rect 16660 6638 16662 6690
rect 16714 6638 16716 6690
rect 16660 6636 16716 6638
rect 18228 6690 18284 6702
rect 18228 6638 18230 6690
rect 18282 6638 18284 6690
rect 18228 6636 18284 6638
rect 18452 6636 18508 7364
rect 18620 7326 18676 7364
rect 18228 6580 18508 6636
rect 16660 6570 16716 6580
rect 16100 6132 16268 6188
rect 14420 6022 14422 6074
rect 14474 6022 14476 6074
rect 14420 6010 14476 6022
rect 15876 5906 15932 5918
rect 15876 5854 15878 5906
rect 15930 5854 15932 5906
rect 15876 5740 15932 5854
rect 15876 5674 15932 5684
rect 14084 5226 14140 5236
rect 15764 5122 15820 5134
rect 15764 5070 15766 5122
rect 15818 5070 15820 5122
rect 14420 5010 14476 5022
rect 13356 4956 13412 4966
rect 13300 4954 13412 4956
rect 13300 4902 13358 4954
rect 13410 4902 13412 4954
rect 13300 4890 13412 4902
rect 14420 4958 14422 5010
rect 14474 4958 14476 5010
rect 13300 4620 13356 4890
rect 11956 1306 12012 1316
rect 12964 4508 13020 4518
rect 12292 1148 12348 1158
rect 12292 800 12348 1092
rect 12964 800 13020 4452
rect 13300 4060 13356 4564
rect 13300 3994 13356 4004
rect 14196 3052 14252 3062
rect 13524 922 13580 934
rect 13524 870 13526 922
rect 13578 870 13580 922
rect 13524 800 13580 870
rect 14196 800 14252 2996
rect 14420 1596 14476 4958
rect 15764 4956 15820 5070
rect 15764 4890 15820 4900
rect 14420 1530 14476 1540
rect 14756 2716 14812 2726
rect 14756 800 14812 2660
rect 15428 2604 15484 2614
rect 15428 800 15484 2548
rect 15988 924 16044 934
rect 15988 800 16044 868
rect 8932 422 8934 474
rect 8986 422 8988 474
rect 8932 410 8988 422
rect 9240 0 9352 800
rect 9912 0 10024 800
rect 10472 0 10584 800
rect 11032 0 11144 800
rect 11704 0 11816 800
rect 12264 0 12376 800
rect 12936 0 13048 800
rect 13496 0 13608 800
rect 14168 0 14280 800
rect 14728 0 14840 800
rect 15400 0 15512 800
rect 15960 0 16072 800
rect 16212 698 16268 6132
rect 16884 5902 16940 5914
rect 16884 5852 16886 5902
rect 16938 5852 16940 5902
rect 16884 5786 16940 5796
rect 17500 5852 17556 5862
rect 17500 5758 17556 5796
rect 18060 5850 18116 5862
rect 18060 5798 18062 5850
rect 18114 5798 18116 5850
rect 18060 5740 18116 5798
rect 18060 5674 18116 5684
rect 18788 5628 18844 8026
rect 19180 7998 19236 8036
rect 21476 7756 21532 7766
rect 19180 7420 19236 7430
rect 19180 7418 19292 7420
rect 19180 7366 19182 7418
rect 19234 7366 19292 7418
rect 19180 7354 19292 7366
rect 19236 6636 19292 7354
rect 20020 6748 20076 6758
rect 21476 6748 21532 7700
rect 21588 7642 21644 10390
rect 21812 8426 21868 10838
rect 22260 9210 22316 11844
rect 24276 11900 24332 14200
rect 25060 13916 25116 14200
rect 25060 13850 25116 13860
rect 25732 13468 25788 14200
rect 25732 13402 25788 13412
rect 24276 11834 24332 11844
rect 25732 10444 25788 10454
rect 22260 9158 22262 9210
rect 22314 9158 22316 9210
rect 22260 9146 22316 9158
rect 22372 9996 22428 10006
rect 21924 9098 21980 9110
rect 21924 9046 21926 9098
rect 21978 9046 21980 9098
rect 21924 8764 21980 9046
rect 21924 8698 21980 8708
rect 22372 8427 22428 9940
rect 22540 9660 22596 9670
rect 22484 9658 22596 9660
rect 22484 9606 22542 9658
rect 22594 9606 22596 9658
rect 22484 9594 22596 9606
rect 25228 9658 25284 9670
rect 25228 9606 25230 9658
rect 25282 9606 25284 9658
rect 22484 8764 22540 9594
rect 23380 9548 23436 9558
rect 23380 9042 23436 9492
rect 25228 9548 25284 9606
rect 25228 9482 25284 9492
rect 23380 8990 23382 9042
rect 23434 8990 23436 9042
rect 23380 8978 23436 8990
rect 25620 9098 25676 9110
rect 25620 9046 25622 9098
rect 25674 9046 25676 9098
rect 25620 8988 25676 9046
rect 22484 8698 22540 8708
rect 23044 8930 23100 8942
rect 23044 8878 23046 8930
rect 23098 8878 23100 8930
rect 25620 8922 25676 8932
rect 23044 8427 23100 8878
rect 21812 8374 21814 8426
rect 21866 8374 21868 8426
rect 21812 8362 21868 8374
rect 22260 8371 22428 8427
rect 22932 8371 23100 8427
rect 21588 7590 21590 7642
rect 21642 7590 21644 7642
rect 21588 7578 21644 7590
rect 18788 5562 18844 5572
rect 18900 5794 18956 5806
rect 18900 5742 18902 5794
rect 18954 5742 18956 5794
rect 16380 4956 16436 4966
rect 16380 4862 16436 4900
rect 16548 2492 16604 2502
rect 16548 800 16604 2436
rect 17780 1596 17836 1606
rect 17220 868 17500 924
rect 17220 800 17276 868
rect 16212 646 16214 698
rect 16266 646 16268 698
rect 16212 634 16268 646
rect 16520 0 16632 800
rect 17192 0 17304 800
rect 17444 252 17500 868
rect 17780 800 17836 1540
rect 18452 1036 18508 1046
rect 18452 800 18508 980
rect 18900 924 18956 5742
rect 19236 5180 19292 6580
rect 19236 5114 19292 5124
rect 19348 6578 19404 6590
rect 19348 6526 19350 6578
rect 19402 6526 19404 6578
rect 19348 1484 19404 6526
rect 20020 5906 20076 6692
rect 20692 6690 20748 6702
rect 20692 6638 20694 6690
rect 20746 6638 20748 6690
rect 20692 6524 20748 6638
rect 20692 6458 20748 6468
rect 21364 6692 21476 6748
rect 20020 5854 20022 5906
rect 20074 5854 20076 5906
rect 20020 5842 20076 5854
rect 21140 5794 21196 5806
rect 21140 5742 21142 5794
rect 21194 5742 21196 5794
rect 20468 5180 20524 5190
rect 20468 5122 20524 5124
rect 20468 5070 20470 5122
rect 20522 5070 20524 5122
rect 20468 5058 20524 5070
rect 21140 5068 21196 5742
rect 19348 1418 19404 1428
rect 19908 5010 19964 5022
rect 19908 4958 19910 5010
rect 19962 4958 19964 5010
rect 21140 5002 21196 5012
rect 21364 4966 21420 6692
rect 21476 6682 21532 6692
rect 21700 6860 21756 6870
rect 21532 6524 21588 6534
rect 21588 6468 21644 6524
rect 21532 6392 21644 6468
rect 19684 924 19740 934
rect 18900 858 18956 868
rect 19012 868 19292 924
rect 19012 800 19068 868
rect 17444 196 17612 252
rect 17556 150 17612 196
rect 17556 138 17668 150
rect 17556 86 17614 138
rect 17666 86 17668 138
rect 17556 84 17668 86
rect 17612 74 17668 84
rect 17752 0 17864 800
rect 18424 0 18536 800
rect 18984 0 19096 800
rect 19236 140 19292 868
rect 19684 800 19740 868
rect 19236 74 19292 84
rect 19656 0 19768 800
rect 19908 252 19964 4958
rect 21308 4954 21420 4966
rect 21308 4902 21310 4954
rect 21362 4902 21420 4954
rect 21308 4900 21420 4902
rect 21308 4890 21364 4900
rect 21588 3274 21644 6392
rect 21700 5180 21756 6804
rect 21700 4966 21756 5124
rect 22260 5906 22316 8371
rect 22260 5854 22262 5906
rect 22314 5854 22316 5906
rect 22260 4966 22316 5854
rect 21700 4954 21812 4966
rect 21700 4902 21758 4954
rect 21810 4902 21812 4954
rect 21700 4900 21812 4902
rect 22260 4954 22372 4966
rect 22260 4902 22318 4954
rect 22370 4902 22372 4954
rect 22260 4900 22372 4902
rect 21756 4890 21812 4900
rect 22316 4890 22372 4900
rect 21588 3222 21590 3274
rect 21642 3222 21644 3274
rect 21588 3210 21644 3222
rect 22036 2602 22092 2614
rect 22036 2550 22038 2602
rect 22090 2550 22092 2602
rect 21476 2490 21532 2502
rect 21476 2438 21478 2490
rect 21530 2438 21532 2490
rect 20244 868 20524 924
rect 20244 800 20300 868
rect 19908 186 19964 196
rect 20216 0 20328 800
rect 20468 364 20524 868
rect 20916 868 21196 924
rect 20916 800 20972 868
rect 20468 308 20748 364
rect 20692 252 20748 308
rect 20692 186 20748 196
rect 20888 0 21000 800
rect 21140 364 21196 868
rect 21476 800 21532 2438
rect 22036 800 22092 2550
rect 22708 1596 22764 1606
rect 22708 800 22764 1540
rect 21140 308 21308 364
rect 21252 262 21308 308
rect 21252 250 21364 262
rect 21252 198 21310 250
rect 21362 198 21364 250
rect 21252 196 21364 198
rect 21308 186 21364 196
rect 21448 0 21560 800
rect 22008 0 22120 800
rect 22680 0 22792 800
rect 22932 700 22988 8371
rect 23380 8258 23436 8270
rect 23380 8206 23382 8258
rect 23434 8206 23436 8258
rect 23380 7980 23436 8206
rect 25060 8258 25116 8270
rect 25060 8206 25062 8258
rect 25114 8206 25116 8258
rect 25060 8092 25116 8206
rect 25060 8026 25116 8036
rect 25452 8092 25508 8102
rect 25452 7998 25508 8036
rect 23380 7914 23436 7924
rect 23044 7474 23100 7486
rect 23044 7422 23046 7474
rect 23098 7422 23100 7474
rect 23044 7196 23100 7422
rect 24052 7470 24108 7482
rect 24052 7418 24054 7470
rect 24106 7420 24108 7470
rect 24556 7420 24612 7430
rect 24106 7418 24668 7420
rect 24052 7366 24558 7418
rect 24610 7366 24668 7418
rect 24052 7364 24668 7366
rect 24556 7354 24668 7364
rect 23044 7130 23100 7140
rect 24388 6690 24444 6702
rect 24388 6638 24390 6690
rect 24442 6638 24444 6690
rect 23044 6578 23100 6590
rect 23044 6526 23046 6578
rect 23098 6526 23100 6578
rect 23044 5180 23100 6526
rect 24388 6300 24444 6638
rect 24612 6524 24668 7354
rect 25564 7418 25620 7430
rect 25564 7366 25566 7418
rect 25618 7366 25620 7418
rect 25564 7196 25620 7366
rect 25564 7130 25620 7140
rect 24612 6458 24668 6468
rect 25004 6522 25060 6534
rect 25004 6470 25006 6522
rect 25058 6470 25060 6522
rect 24388 6234 24444 6244
rect 25004 6300 25060 6470
rect 25004 6234 25060 6244
rect 24724 5964 24780 5974
rect 24724 5906 24780 5908
rect 24724 5854 24726 5906
rect 24778 5854 24780 5906
rect 24724 5842 24780 5854
rect 25452 5964 25508 5974
rect 25452 5850 25508 5908
rect 23044 5114 23100 5124
rect 23380 5794 23436 5806
rect 23380 5742 23382 5794
rect 23434 5742 23436 5794
rect 23380 5068 23436 5742
rect 25452 5798 25454 5850
rect 25506 5798 25508 5850
rect 25452 5404 25508 5798
rect 25452 5338 25508 5348
rect 23044 5010 23100 5022
rect 23044 4958 23046 5010
rect 23098 4958 23100 5010
rect 23380 5002 23436 5012
rect 24388 5122 24444 5134
rect 24388 5070 24390 5122
rect 24442 5070 24444 5122
rect 24388 5068 24444 5070
rect 24388 5002 24444 5012
rect 25228 5068 25284 5078
rect 23044 4844 23100 4958
rect 25228 4956 25284 5012
rect 25228 4954 25340 4956
rect 25228 4902 25230 4954
rect 25282 4902 25340 4954
rect 25228 4890 25340 4902
rect 23044 4778 23100 4788
rect 25284 3612 25340 4890
rect 25284 3546 25340 3556
rect 24500 3164 24556 3174
rect 23268 2714 23324 2726
rect 23268 2662 23270 2714
rect 23322 2662 23324 2714
rect 23268 800 23324 2662
rect 23940 868 24220 924
rect 23940 800 23996 868
rect 22932 634 22988 644
rect 23240 0 23352 800
rect 23912 0 24024 800
rect 24164 476 24220 868
rect 24500 800 24556 3108
rect 25172 1484 25228 1494
rect 25172 800 25228 1428
rect 25732 800 25788 10388
rect 25956 9210 26012 14308
rect 26292 14140 26348 14308
rect 26488 14200 26600 15000
rect 27160 14200 27272 15000
rect 27944 14200 28056 15000
rect 28616 14200 28728 15000
rect 29400 14200 29512 15000
rect 30072 14200 30184 15000
rect 30856 14200 30968 15000
rect 31528 14200 31640 15000
rect 32312 14200 32424 15000
rect 32984 14200 33096 15000
rect 33768 14200 33880 15000
rect 34440 14200 34552 15000
rect 35224 14200 35336 15000
rect 35896 14200 36008 15000
rect 36680 14200 36792 15000
rect 37352 14200 37464 15000
rect 38136 14200 38248 15000
rect 38808 14200 38920 15000
rect 39592 14200 39704 15000
rect 40264 14200 40376 15000
rect 41048 14200 41160 15000
rect 41720 14200 41832 15000
rect 42308 14924 42364 14934
rect 26516 14140 26572 14200
rect 26292 14084 26572 14140
rect 27188 12796 27244 14200
rect 27972 13020 28028 14200
rect 27972 12954 28028 12964
rect 27188 12730 27244 12740
rect 26964 11788 27020 11798
rect 25956 9158 25958 9210
rect 26010 9158 26012 9210
rect 25956 9146 26012 9158
rect 26740 10108 26796 10118
rect 26348 8988 26404 8998
rect 26348 8894 26404 8932
rect 26628 8204 26684 8214
rect 26628 8110 26684 8148
rect 25900 8090 25956 8102
rect 25900 8038 25902 8090
rect 25954 8038 25956 8090
rect 25900 7980 25956 8038
rect 25900 7914 25956 7924
rect 26740 7644 26796 10052
rect 26964 8314 27020 11732
rect 28644 11788 28700 14200
rect 29428 12682 29484 14200
rect 29428 12630 29430 12682
rect 29482 12630 29484 12682
rect 29428 12618 29484 12630
rect 30100 12572 30156 14200
rect 30100 12506 30156 12516
rect 28644 11722 28700 11732
rect 29876 11788 29932 11798
rect 28376 10220 28640 10230
rect 28432 10164 28480 10220
rect 28536 10164 28584 10220
rect 28376 10154 28640 10164
rect 28376 8652 28640 8662
rect 28432 8596 28480 8652
rect 28536 8596 28584 8652
rect 28376 8586 28640 8596
rect 26964 8262 26966 8314
rect 27018 8262 27020 8314
rect 26964 8250 27020 8262
rect 29876 8314 29932 11732
rect 30884 11788 30940 14200
rect 31556 12572 31612 14200
rect 32340 13692 32396 14200
rect 32340 13626 32396 13636
rect 31556 12506 31612 12516
rect 30884 11722 30940 11732
rect 33012 11340 33068 14200
rect 33796 11786 33852 14200
rect 34468 13020 34524 14200
rect 34468 12954 34524 12964
rect 33796 11734 33798 11786
rect 33850 11734 33852 11786
rect 33796 11722 33852 11734
rect 34356 11788 34412 11798
rect 29876 8262 29878 8314
rect 29930 8262 29932 8314
rect 29876 8250 29932 8262
rect 31892 11284 33068 11340
rect 31892 8314 31948 11284
rect 31892 8262 31894 8314
rect 31946 8262 31948 8314
rect 31892 8250 31948 8262
rect 32676 10220 32732 10230
rect 27468 8204 27524 8214
rect 27468 8092 27524 8148
rect 29540 8204 29596 8214
rect 29540 8110 29596 8148
rect 30324 8204 30380 8214
rect 30324 8102 30380 8148
rect 31556 8204 31612 8214
rect 31556 8110 31612 8148
rect 32340 8204 32396 8214
rect 32340 8102 32396 8148
rect 27468 8090 27580 8092
rect 27468 8038 27470 8090
rect 27522 8038 27580 8090
rect 27468 8026 27580 8038
rect 26852 7644 26908 7654
rect 26740 7642 26908 7644
rect 26740 7590 26854 7642
rect 26906 7590 26908 7642
rect 26740 7588 26908 7590
rect 26852 7578 26908 7588
rect 26404 6578 26460 6590
rect 26404 6526 26406 6578
rect 26458 6526 26460 6578
rect 26404 6412 26460 6526
rect 26404 6346 26460 6356
rect 26852 5794 26908 5806
rect 26852 5742 26854 5794
rect 26906 5742 26908 5794
rect 26404 1708 26460 1718
rect 26404 800 26460 1652
rect 26852 1148 26908 5742
rect 26964 5010 27020 5022
rect 26964 4958 26966 5010
rect 27018 4958 27020 5010
rect 26964 4732 27020 4958
rect 26964 4666 27020 4676
rect 27524 3162 27580 8026
rect 30324 8090 30436 8102
rect 30324 8038 30382 8090
rect 30434 8038 30436 8090
rect 30324 8026 30436 8038
rect 32340 8090 32452 8102
rect 32340 8038 32398 8090
rect 32450 8038 32452 8090
rect 32340 8026 32452 8038
rect 28196 7474 28252 7486
rect 28196 7422 28198 7474
rect 28250 7422 28252 7474
rect 28196 7196 28252 7422
rect 29652 7470 29708 7482
rect 29652 7418 29654 7470
rect 29706 7420 29708 7470
rect 30156 7420 30212 7430
rect 29706 7418 30212 7420
rect 29652 7366 30158 7418
rect 30210 7366 30212 7418
rect 29652 7364 30212 7366
rect 28196 7130 28252 7140
rect 30100 7354 30212 7364
rect 28376 7084 28640 7094
rect 28432 7028 28480 7084
rect 28536 7028 28584 7084
rect 28376 7018 28640 7028
rect 27748 6690 27804 6702
rect 27748 6638 27750 6690
rect 27802 6638 27804 6690
rect 27748 6188 27804 6638
rect 28700 6636 28756 6646
rect 28532 6580 28700 6636
rect 27748 6122 27804 6132
rect 28364 6522 28420 6534
rect 28364 6470 28366 6522
rect 28418 6470 28420 6522
rect 28364 6188 28420 6470
rect 28364 6122 28420 6132
rect 28196 5908 28252 5918
rect 28532 5908 28588 6580
rect 28700 6542 28756 6580
rect 30100 6076 30156 7354
rect 30100 6010 30156 6020
rect 28196 5906 28588 5908
rect 28196 5854 28198 5906
rect 28250 5854 28588 5906
rect 28196 5852 28588 5854
rect 28196 5842 28252 5852
rect 29092 5794 29148 5806
rect 29092 5742 29094 5794
rect 29146 5742 29148 5794
rect 28376 5516 28640 5526
rect 28432 5460 28480 5516
rect 28536 5460 28584 5516
rect 28376 5450 28640 5460
rect 29092 5180 29148 5742
rect 28308 5122 28364 5134
rect 28308 5070 28310 5122
rect 28362 5070 28364 5122
rect 28308 4956 28364 5070
rect 28308 4890 28364 4900
rect 28980 5124 29148 5180
rect 27524 3110 27526 3162
rect 27578 3110 27580 3162
rect 27524 3098 27580 3110
rect 28196 2940 28252 2950
rect 26852 1082 26908 1092
rect 26964 2828 27020 2838
rect 26964 800 27020 2772
rect 27524 2826 27580 2838
rect 27524 2774 27526 2826
rect 27578 2774 27580 2826
rect 27524 800 27580 2774
rect 28196 800 28252 2884
rect 28756 1596 28812 1606
rect 28756 800 28812 1540
rect 28980 810 29036 5124
rect 29148 4956 29204 4966
rect 29204 4900 29260 4956
rect 29148 4824 29260 4900
rect 29204 3948 29260 4824
rect 30324 4284 30380 8026
rect 30604 7418 30660 7430
rect 30604 7366 30606 7418
rect 30658 7366 30660 7418
rect 30604 7196 30660 7366
rect 30604 7130 30660 7140
rect 30604 6972 30660 6982
rect 30604 6636 30660 6916
rect 30436 6634 30660 6636
rect 30436 6582 30606 6634
rect 30658 6582 30660 6634
rect 30436 6580 30660 6582
rect 30436 5906 30492 6580
rect 30604 6570 30660 6580
rect 30436 5854 30438 5906
rect 30490 5854 30492 5906
rect 30436 5842 30492 5854
rect 31444 5794 31500 5806
rect 31444 5742 31446 5794
rect 31498 5742 31500 5794
rect 30884 5010 30940 5022
rect 30884 4958 30886 5010
rect 30938 4958 30940 5010
rect 30884 4620 30940 4958
rect 30884 4554 30940 4564
rect 30324 4218 30380 4228
rect 29204 3882 29260 3892
rect 31220 3500 31276 3510
rect 30660 3388 30716 3398
rect 29988 1596 30044 1606
rect 24164 420 24332 476
rect 24276 362 24332 420
rect 24276 310 24278 362
rect 24330 310 24332 362
rect 24276 298 24332 310
rect 24472 0 24584 800
rect 25144 0 25256 800
rect 25704 0 25816 800
rect 26376 0 26488 800
rect 26936 0 27048 800
rect 27496 0 27608 800
rect 28168 0 28280 800
rect 28728 0 28840 800
rect 28980 758 28982 810
rect 29034 758 29036 810
rect 29428 868 29708 924
rect 29428 800 29484 868
rect 28980 746 29036 758
rect 29400 0 29512 800
rect 29652 700 29708 868
rect 29988 800 30044 1540
rect 30660 800 30716 3332
rect 31220 800 31276 3444
rect 29652 634 29708 644
rect 29960 0 30072 800
rect 30632 0 30744 800
rect 31192 0 31304 800
rect 31444 588 31500 5742
rect 31780 5516 31836 5526
rect 31780 5122 31836 5460
rect 31780 5070 31782 5122
rect 31834 5070 31836 5122
rect 31780 5058 31836 5070
rect 31892 3498 31948 3510
rect 31892 3446 31894 3498
rect 31946 3446 31948 3498
rect 31892 800 31948 3446
rect 32340 1594 32396 8026
rect 32676 6858 32732 10164
rect 34356 8314 34412 11732
rect 35252 11788 35308 14200
rect 35252 11722 35308 11732
rect 35924 8427 35980 14200
rect 36708 12796 36764 14200
rect 36708 12730 36764 12740
rect 34356 8262 34358 8314
rect 34410 8262 34412 8314
rect 34356 8250 34412 8262
rect 35252 8371 35980 8427
rect 36708 11788 36764 11798
rect 35252 8314 35308 8371
rect 35252 8262 35254 8314
rect 35306 8262 35308 8314
rect 35252 8250 35308 8262
rect 36708 8314 36764 11732
rect 37380 11788 37436 14200
rect 37380 11722 37436 11732
rect 38164 11452 38220 14200
rect 38836 13580 38892 14200
rect 38836 13514 38892 13524
rect 37828 11396 38220 11452
rect 36708 8262 36710 8314
rect 36762 8262 36764 8314
rect 36708 8250 36764 8262
rect 36820 10108 36876 10118
rect 34916 8204 34972 8214
rect 34916 8110 34972 8148
rect 35756 8204 35812 8214
rect 34020 8090 34076 8102
rect 34020 8038 34022 8090
rect 34074 8038 34076 8090
rect 34020 7196 34076 8038
rect 35756 8092 35812 8148
rect 36372 8204 36428 8214
rect 35756 8090 35980 8092
rect 35756 8038 35758 8090
rect 35810 8038 35980 8090
rect 35756 8036 35980 8038
rect 35756 8026 35812 8036
rect 34020 7130 34076 7140
rect 34524 7418 34580 7430
rect 34524 7366 34526 7418
rect 34578 7366 34580 7418
rect 34524 7196 34580 7366
rect 34524 7130 34580 7140
rect 32676 6806 32678 6858
rect 32730 6806 32732 6858
rect 32676 6794 32732 6806
rect 33460 6690 33516 6702
rect 33460 6638 33462 6690
rect 33514 6638 33516 6690
rect 33460 6076 33516 6638
rect 34692 6690 34748 6702
rect 34692 6638 34694 6690
rect 34746 6638 34748 6690
rect 34692 6412 34748 6638
rect 34692 6346 34748 6356
rect 35084 6522 35140 6534
rect 35084 6470 35086 6522
rect 35138 6470 35140 6522
rect 35084 6412 35140 6470
rect 35084 6346 35140 6356
rect 35532 6522 35588 6534
rect 35532 6470 35534 6522
rect 35586 6470 35588 6522
rect 33460 6010 33516 6020
rect 35532 6076 35588 6470
rect 35532 6010 35588 6020
rect 32676 5906 32732 5918
rect 32676 5854 32678 5906
rect 32730 5854 32732 5906
rect 32676 5740 32732 5854
rect 33404 5852 33460 5862
rect 33404 5850 33516 5852
rect 33404 5798 33406 5850
rect 33458 5798 33516 5850
rect 33404 5786 33516 5798
rect 32676 5674 32732 5684
rect 33460 5740 33516 5786
rect 33460 4732 33516 5684
rect 33852 5850 33908 5862
rect 33852 5798 33854 5850
rect 33906 5798 33908 5850
rect 33852 5740 33908 5798
rect 33852 5674 33908 5684
rect 35812 5794 35868 5806
rect 35812 5742 35814 5794
rect 35866 5742 35868 5794
rect 35028 5122 35084 5134
rect 35028 5070 35030 5122
rect 35082 5070 35084 5122
rect 33460 4666 33516 4676
rect 33908 5010 33964 5022
rect 33908 4958 33910 5010
rect 33962 4958 33964 5010
rect 33012 3386 33068 3398
rect 33012 3334 33014 3386
rect 33066 3334 33068 3386
rect 32340 1542 32342 1594
rect 32394 1542 32396 1594
rect 32340 1530 32396 1542
rect 32452 3276 32508 3286
rect 32452 800 32508 3220
rect 33012 800 33068 3334
rect 33684 1260 33740 1270
rect 33684 800 33740 1204
rect 31444 522 31500 532
rect 31864 0 31976 800
rect 32424 0 32536 800
rect 32984 0 33096 800
rect 33656 0 33768 800
rect 33908 586 33964 4958
rect 35028 4956 35084 5070
rect 35028 4890 35084 4900
rect 35644 4956 35700 4966
rect 35644 4862 35700 4900
rect 34916 2042 34972 2054
rect 34916 1990 34918 2042
rect 34970 1990 34972 2042
rect 34244 1596 34300 1606
rect 34244 800 34300 1540
rect 34916 800 34972 1990
rect 35476 1596 35532 1606
rect 35476 800 35532 1540
rect 33908 534 33910 586
rect 33962 534 33964 586
rect 33908 522 33964 534
rect 34216 0 34328 800
rect 34888 0 35000 800
rect 35448 0 35560 800
rect 35812 364 35868 5742
rect 35924 4508 35980 8036
rect 35924 4442 35980 4452
rect 36372 8090 36428 8148
rect 36372 8038 36374 8090
rect 36426 8038 36428 8090
rect 36148 4394 36204 4406
rect 36148 4342 36150 4394
rect 36202 4342 36204 4394
rect 36148 800 36204 4342
rect 36372 1482 36428 8038
rect 36820 7306 36876 10052
rect 36988 8986 37044 8998
rect 36988 8934 36990 8986
rect 37042 8934 37044 8986
rect 36988 8427 37044 8934
rect 36932 8371 37044 8427
rect 36932 8204 36988 8371
rect 37828 8314 37884 11396
rect 39620 11228 39676 14200
rect 40292 11788 40348 14200
rect 41076 13018 41132 14200
rect 41076 12966 41078 13018
rect 41130 12966 41132 13018
rect 41076 12954 41132 12966
rect 39060 11172 39676 11228
rect 39956 11732 40348 11788
rect 38108 8986 38164 8998
rect 38108 8934 38110 8986
rect 38162 8934 38164 8986
rect 38108 8427 38164 8934
rect 37828 8262 37830 8314
rect 37882 8262 37884 8314
rect 37828 8250 37884 8262
rect 38052 8371 38164 8427
rect 36932 8138 36988 8148
rect 37492 8092 37548 8102
rect 38052 8092 38108 8371
rect 39060 8314 39116 11172
rect 39060 8262 39062 8314
rect 39114 8262 39116 8314
rect 39060 8250 39116 8262
rect 39956 8314 40012 11732
rect 41748 11340 41804 14200
rect 39956 8262 39958 8314
rect 40010 8262 40012 8314
rect 39956 8250 40012 8262
rect 41076 11284 41804 11340
rect 41076 8314 41132 11284
rect 41076 8262 41078 8314
rect 41130 8262 41132 8314
rect 41076 8250 41132 8262
rect 41300 10778 41356 10790
rect 41300 10726 41302 10778
rect 41354 10726 41356 10778
rect 37492 8090 38108 8092
rect 37492 8038 37494 8090
rect 37546 8038 38108 8090
rect 37492 8036 38108 8038
rect 38724 8092 38780 8102
rect 39620 8092 39676 8102
rect 38724 8090 38892 8092
rect 38724 8038 38726 8090
rect 38778 8038 38892 8090
rect 38724 8036 38892 8038
rect 37492 8026 37548 8036
rect 36820 7254 36822 7306
rect 36874 7254 36876 7306
rect 36820 7242 36876 7254
rect 37044 5906 37100 5918
rect 37044 5854 37046 5906
rect 37098 5854 37100 5906
rect 37044 5852 37100 5854
rect 37548 5852 37604 5862
rect 37044 5850 37660 5852
rect 37044 5798 37550 5850
rect 37602 5798 37660 5850
rect 37044 5796 37660 5798
rect 37548 5786 37660 5796
rect 37268 5010 37324 5022
rect 37268 4958 37270 5010
rect 37322 4958 37324 5010
rect 36372 1430 36374 1482
rect 36426 1430 36428 1482
rect 36372 1418 36428 1430
rect 36708 4282 36764 4294
rect 36708 4230 36710 4282
rect 36762 4230 36764 4282
rect 36708 800 36764 4230
rect 37268 922 37324 4958
rect 37268 870 37270 922
rect 37322 870 37324 922
rect 37268 858 37324 870
rect 37380 4170 37436 4182
rect 37380 4118 37382 4170
rect 37434 4118 37436 4170
rect 37380 800 37436 4118
rect 37604 2380 37660 5786
rect 37716 4506 37772 8036
rect 38724 8026 38780 8036
rect 37828 7474 37884 7486
rect 37828 7422 37830 7474
rect 37882 7422 37884 7474
rect 37828 6636 37884 7422
rect 38724 7455 38780 7467
rect 38724 7403 38726 7455
rect 38778 7403 38780 7455
rect 38724 7084 38780 7403
rect 38836 7420 38892 8036
rect 39620 8090 40012 8092
rect 39620 8038 39622 8090
rect 39674 8038 40012 8090
rect 39620 8036 40012 8038
rect 39620 8026 39676 8036
rect 39228 7420 39284 7430
rect 38836 7418 39452 7420
rect 38836 7366 39230 7418
rect 39282 7366 39452 7418
rect 38836 7364 39452 7366
rect 39228 7354 39284 7364
rect 38724 7018 38780 7028
rect 37828 6570 37884 6580
rect 39004 6636 39060 6646
rect 39004 6524 39060 6580
rect 39004 6522 39116 6524
rect 39004 6470 39006 6522
rect 39058 6470 39116 6522
rect 39004 6458 39116 6470
rect 38500 5628 38556 5638
rect 38500 5122 38556 5572
rect 38500 5070 38502 5122
rect 38554 5070 38556 5122
rect 38500 5058 38556 5070
rect 37716 4454 37718 4506
rect 37770 4454 37772 4506
rect 37716 4442 37772 4454
rect 38500 3050 38556 3062
rect 38500 2998 38502 3050
rect 38554 2998 38556 3050
rect 37604 2314 37660 2324
rect 37940 2378 37996 2390
rect 37940 2326 37942 2378
rect 37994 2326 37996 2378
rect 37940 800 37996 2326
rect 38500 800 38556 2998
rect 39060 1484 39116 6458
rect 39228 5628 39284 5638
rect 39228 4954 39284 5572
rect 39228 4902 39230 4954
rect 39282 4902 39284 4954
rect 39228 4890 39284 4902
rect 39060 1418 39116 1428
rect 39172 1036 39228 1046
rect 39172 800 39228 980
rect 39396 812 39452 7364
rect 39788 7418 39844 7430
rect 39788 7366 39790 7418
rect 39842 7366 39844 7418
rect 39788 7084 39844 7366
rect 39956 7420 40012 8036
rect 40740 8090 40796 8102
rect 40740 8038 40742 8090
rect 40794 8038 40796 8090
rect 40740 7980 40796 8038
rect 40740 7654 40796 7924
rect 40740 7642 40852 7654
rect 40740 7590 40798 7642
rect 40850 7590 40852 7642
rect 40740 7588 40852 7590
rect 40796 7578 40852 7588
rect 40124 7420 40180 7430
rect 39956 7418 40236 7420
rect 39956 7366 40126 7418
rect 40178 7366 40236 7418
rect 39956 7364 40236 7366
rect 40124 7354 40236 7364
rect 39788 7018 39844 7028
rect 40068 6188 40124 6198
rect 40068 5628 40124 6132
rect 40068 5562 40124 5572
rect 40180 4284 40236 7354
rect 41300 6860 41356 10726
rect 41972 10108 42028 10118
rect 41972 9210 42028 10052
rect 41972 9158 41974 9210
rect 42026 9158 42028 9210
rect 41972 9146 42028 9158
rect 42308 9210 42364 14868
rect 42504 14200 42616 15000
rect 42980 14700 43036 14710
rect 42532 10332 42588 14200
rect 42980 12012 43036 14644
rect 43176 14200 43288 15000
rect 43960 14200 44072 15000
rect 44632 14200 44744 15000
rect 45416 14200 45528 15000
rect 45668 14588 45724 14598
rect 43204 12906 43260 14200
rect 43204 12854 43206 12906
rect 43258 12854 43260 12906
rect 43204 12842 43260 12854
rect 43652 13914 43708 13926
rect 43652 13862 43654 13914
rect 43706 13862 43708 13914
rect 43652 12684 43708 13862
rect 43652 12618 43708 12628
rect 42980 11956 43148 12012
rect 42980 11788 43036 11798
rect 42308 9158 42310 9210
rect 42362 9158 42364 9210
rect 42308 9146 42364 9158
rect 42420 10276 42588 10332
rect 42644 11340 42700 11350
rect 41468 8988 41524 8998
rect 42420 8988 42476 10276
rect 42644 10108 42700 11284
rect 42644 9894 42700 10052
rect 42588 9882 42700 9894
rect 42588 9830 42590 9882
rect 42642 9830 42700 9882
rect 42588 9828 42700 9830
rect 42588 9818 42644 9828
rect 41468 8986 41580 8988
rect 41468 8934 41470 8986
rect 41522 8934 41580 8986
rect 41468 8922 41580 8934
rect 41524 8092 41580 8922
rect 41972 8932 42476 8988
rect 42532 9324 42588 9334
rect 41972 8314 42028 8932
rect 41972 8262 41974 8314
rect 42026 8262 42028 8314
rect 41972 8250 42028 8262
rect 41636 8092 41692 8102
rect 41524 8090 41692 8092
rect 41524 8038 41638 8090
rect 41690 8038 41692 8090
rect 41524 8036 41692 8038
rect 41412 6860 41468 6870
rect 41300 6858 41468 6860
rect 41300 6806 41414 6858
rect 41466 6806 41468 6858
rect 41300 6804 41468 6806
rect 41412 6794 41468 6804
rect 40180 4218 40236 4228
rect 41636 2268 41692 8036
rect 42532 8090 42588 9268
rect 42868 9100 42924 9110
rect 42868 9006 42924 9044
rect 42868 8316 42924 8326
rect 42980 8316 43036 11732
rect 42868 8314 43036 8316
rect 42868 8262 42870 8314
rect 42922 8262 43036 8314
rect 42868 8260 43036 8262
rect 42868 8250 42924 8260
rect 42532 8038 42534 8090
rect 42586 8038 42588 8090
rect 42196 7644 42252 7654
rect 42196 7550 42252 7588
rect 41860 7532 41916 7542
rect 41860 7530 42028 7532
rect 41860 7478 41862 7530
rect 41914 7478 42028 7530
rect 41860 7476 42028 7478
rect 41860 7466 41916 7476
rect 41860 6690 41916 6702
rect 41860 6638 41862 6690
rect 41914 6638 41916 6690
rect 41748 5010 41804 5022
rect 41748 4958 41750 5010
rect 41802 4958 41804 5010
rect 41748 3052 41804 4958
rect 41860 4732 41916 6638
rect 41972 5852 42028 7476
rect 41972 5786 42028 5796
rect 42364 5852 42420 5862
rect 42364 5758 42420 5796
rect 41860 4666 41916 4676
rect 41748 2986 41804 2996
rect 42196 4060 42252 4070
rect 41636 2202 41692 2212
rect 35812 298 35868 308
rect 36120 0 36232 800
rect 36680 0 36792 800
rect 37352 0 37464 800
rect 37912 0 38024 800
rect 38472 0 38584 800
rect 39144 0 39256 800
rect 39732 924 39788 934
rect 39732 800 39788 868
rect 40404 924 40460 934
rect 40404 800 40460 868
rect 40964 924 41020 934
rect 40964 800 41020 868
rect 41412 868 41692 924
rect 39396 746 39452 756
rect 39704 0 39816 800
rect 40376 0 40488 800
rect 40936 0 41048 800
rect 41412 588 41468 868
rect 41636 800 41692 868
rect 42196 800 42252 4004
rect 42532 1034 42588 8038
rect 43092 7642 43148 11956
rect 43540 12010 43596 12022
rect 43540 11958 43542 12010
rect 43594 11958 43596 12010
rect 43540 9894 43596 11958
rect 43988 11788 44044 14200
rect 44660 12012 44716 14200
rect 45444 14026 45500 14200
rect 45444 13974 45446 14026
rect 45498 13974 45500 14026
rect 45444 13962 45500 13974
rect 43988 11722 44044 11732
rect 44100 11956 44716 12012
rect 44884 12124 44940 12134
rect 45668 12124 45724 14532
rect 46088 14200 46200 15000
rect 46872 14200 46984 15000
rect 47544 14200 47656 15000
rect 48328 14200 48440 15000
rect 49000 14200 49112 15000
rect 49784 14200 49896 15000
rect 50456 14200 50568 15000
rect 51044 14474 51100 14486
rect 51044 14422 51046 14474
rect 51098 14422 51100 14474
rect 44100 11340 44156 11956
rect 43484 9882 43596 9894
rect 43484 9830 43486 9882
rect 43538 9830 43596 9882
rect 43484 9828 43596 9830
rect 43764 11284 44156 11340
rect 44660 11788 44716 11798
rect 43204 9660 43260 9670
rect 43204 9210 43260 9604
rect 43204 9158 43206 9210
rect 43258 9158 43260 9210
rect 43204 9146 43260 9158
rect 43484 9100 43540 9828
rect 43484 9034 43540 9044
rect 43092 7590 43094 7642
rect 43146 7590 43148 7642
rect 43092 7578 43148 7590
rect 43204 8316 43260 8326
rect 42756 7530 42812 7542
rect 42756 7478 42758 7530
rect 42810 7478 42812 7530
rect 42756 5852 42812 7478
rect 43204 6188 43260 8260
rect 43764 8314 43820 11284
rect 43932 9658 43988 9670
rect 43932 9606 43934 9658
rect 43986 9606 43988 9658
rect 43932 9324 43988 9606
rect 43932 9258 43988 9268
rect 44100 9324 44156 9334
rect 44100 9222 44156 9268
rect 44044 9210 44156 9222
rect 44044 9158 44046 9210
rect 44098 9158 44156 9210
rect 44044 9156 44156 9158
rect 44548 9324 44604 9334
rect 44548 9210 44604 9268
rect 44548 9158 44550 9210
rect 44602 9158 44604 9210
rect 44044 9146 44100 9156
rect 44548 9146 44604 9158
rect 43764 8262 43766 8314
rect 43818 8262 43820 8314
rect 43764 8250 43820 8262
rect 44660 8314 44716 11732
rect 44884 9210 44940 12068
rect 45556 12068 45724 12124
rect 45444 11452 45500 11462
rect 45220 9660 45276 9670
rect 45220 9566 45276 9604
rect 45444 9222 45500 11396
rect 45556 9994 45612 12068
rect 46116 11788 46172 14200
rect 46900 13244 46956 14200
rect 47572 13802 47628 14200
rect 47572 13750 47574 13802
rect 47626 13750 47628 13802
rect 47572 13738 47628 13750
rect 46116 11722 46172 11732
rect 46228 13188 46956 13244
rect 46228 11228 46284 13188
rect 45556 9942 45558 9994
rect 45610 9942 45612 9994
rect 45556 9930 45612 9942
rect 45780 11172 46284 11228
rect 46452 13020 46508 13030
rect 44884 9158 44886 9210
rect 44938 9158 44940 9210
rect 44884 9146 44940 9158
rect 45388 9210 45500 9222
rect 45388 9158 45390 9210
rect 45442 9158 45500 9210
rect 45388 9146 45500 9158
rect 44660 8262 44662 8314
rect 44714 8262 44716 8314
rect 44660 8250 44716 8262
rect 45444 8204 45500 9146
rect 45780 8316 45836 11172
rect 46452 10892 46508 12964
rect 47684 12348 47740 12358
rect 46228 10836 46508 10892
rect 46900 11900 46956 11910
rect 46060 9660 46116 9670
rect 46060 9566 46116 9604
rect 45892 9100 45948 9110
rect 45892 9098 46060 9100
rect 45892 9046 45894 9098
rect 45946 9046 46060 9098
rect 45892 9044 46060 9046
rect 45892 9034 45948 9044
rect 46004 8652 46060 9044
rect 46228 8874 46284 10836
rect 46508 9660 46564 9670
rect 46228 8822 46230 8874
rect 46282 8822 46284 8874
rect 46228 8810 46284 8822
rect 46452 9658 46564 9660
rect 46452 9606 46510 9658
rect 46562 9606 46564 9658
rect 46452 9594 46564 9606
rect 46676 9660 46732 9670
rect 46452 8652 46508 9594
rect 46004 8596 46508 8652
rect 45892 8316 45948 8326
rect 45780 8314 45948 8316
rect 45780 8262 45894 8314
rect 45946 8262 45948 8314
rect 45780 8260 45948 8262
rect 45892 8250 45948 8260
rect 45556 8204 45612 8214
rect 45444 8202 45612 8204
rect 45444 8150 45558 8202
rect 45610 8150 45612 8202
rect 45444 8148 45612 8150
rect 45556 8138 45612 8148
rect 43428 8090 43484 8102
rect 43428 8038 43430 8090
rect 43482 8038 43484 8090
rect 43428 6748 43484 8038
rect 44324 8090 44380 8102
rect 44324 8038 44326 8090
rect 44378 8038 44380 8090
rect 43316 6679 43372 6691
rect 43316 6636 43318 6679
rect 43370 6636 43372 6679
rect 43316 6570 43372 6580
rect 43204 6122 43260 6132
rect 42756 5786 42812 5796
rect 43260 5852 43316 5862
rect 43316 5796 43372 5852
rect 43260 5720 43372 5796
rect 43092 5122 43148 5134
rect 43092 5070 43094 5122
rect 43146 5070 43148 5122
rect 43092 4844 43148 5070
rect 43092 4778 43148 4788
rect 43316 2044 43372 5720
rect 43428 3610 43484 6692
rect 43652 7530 43708 7542
rect 43652 7478 43654 7530
rect 43706 7478 43708 7530
rect 43652 6524 43708 7478
rect 44324 7420 44380 8038
rect 44604 7420 44660 7430
rect 44324 7418 44660 7420
rect 44324 7366 44606 7418
rect 44658 7366 44660 7418
rect 44324 7364 44660 7366
rect 43988 7308 44044 7318
rect 43988 7306 44156 7308
rect 43988 7254 43990 7306
rect 44042 7254 44156 7306
rect 43988 7252 44156 7254
rect 43988 7242 44044 7252
rect 43932 6748 43988 6758
rect 43932 6654 43988 6692
rect 43652 6458 43708 6468
rect 43820 6636 43876 6646
rect 43820 5852 43876 6580
rect 43820 5850 43932 5852
rect 43820 5798 43822 5850
rect 43874 5798 43932 5850
rect 43820 5786 43932 5798
rect 43876 5180 43932 5786
rect 43876 5114 43932 5124
rect 43708 4954 43764 4966
rect 43708 4902 43710 4954
rect 43762 4902 43764 4954
rect 43708 4844 43764 4902
rect 43708 4778 43764 4788
rect 43428 3558 43430 3610
rect 43482 3558 43484 3610
rect 43428 3546 43484 3558
rect 43316 1978 43372 1988
rect 42532 982 42534 1034
rect 42586 982 42588 1034
rect 42532 970 42588 982
rect 43988 1372 44044 1382
rect 42644 868 42924 924
rect 41188 532 41468 588
rect 41188 476 41244 532
rect 41188 410 41244 420
rect 41608 0 41720 800
rect 42168 0 42280 800
rect 42644 588 42700 868
rect 42868 800 42924 868
rect 43428 922 43484 934
rect 43428 870 43430 922
rect 43482 870 43484 922
rect 43428 800 43484 870
rect 43988 800 44044 1316
rect 44100 924 44156 7252
rect 44604 7196 44660 7364
rect 44604 7130 44660 7140
rect 44380 6524 44436 6534
rect 44436 6468 44828 6524
rect 44380 6392 44436 6468
rect 44268 5852 44324 5862
rect 44268 5850 44380 5852
rect 44268 5798 44270 5850
rect 44322 5798 44380 5850
rect 44268 5786 44380 5798
rect 44324 4732 44380 5786
rect 44324 4666 44380 4676
rect 44772 1258 44828 6468
rect 45220 5794 45276 5806
rect 45220 5742 45222 5794
rect 45274 5742 45276 5794
rect 45108 4844 45164 4854
rect 45108 3052 45164 4788
rect 45108 2986 45164 2996
rect 45220 2716 45276 5742
rect 45220 2650 45276 2660
rect 45892 1484 45948 1494
rect 44772 1206 44774 1258
rect 44826 1206 44828 1258
rect 44772 1194 44828 1206
rect 45220 1372 45276 1382
rect 44660 1148 44716 1158
rect 44100 868 44268 924
rect 42532 532 42700 588
rect 42532 474 42588 532
rect 42532 422 42534 474
rect 42586 422 42588 474
rect 42532 410 42588 422
rect 42840 0 42952 800
rect 43400 0 43512 800
rect 43960 0 44072 800
rect 44212 364 44268 868
rect 44660 800 44716 1092
rect 45220 800 45276 1316
rect 45892 800 45948 1428
rect 46004 1370 46060 8596
rect 46452 8092 46508 8102
rect 46676 8092 46732 9604
rect 46900 9324 46956 11844
rect 47348 10332 47404 10342
rect 47068 9660 47124 9670
rect 47068 9566 47124 9604
rect 46900 9268 47068 9324
rect 46844 9100 46900 9110
rect 46844 9006 46900 9044
rect 47012 8764 47068 9268
rect 47348 9210 47404 10276
rect 47348 9158 47350 9210
rect 47402 9158 47404 9210
rect 47348 9146 47404 9158
rect 47684 9210 47740 12292
rect 48356 11900 48412 14200
rect 48580 12236 48636 12246
rect 48356 11834 48412 11844
rect 48468 12012 48524 12022
rect 47684 9158 47686 9210
rect 47738 9158 47740 9210
rect 47684 9146 47740 9158
rect 47796 11788 47852 11798
rect 46788 8708 47068 8764
rect 46788 8314 46844 8708
rect 46788 8262 46790 8314
rect 46842 8262 46844 8314
rect 46788 8250 46844 8262
rect 47684 8316 47740 8326
rect 47796 8316 47852 11732
rect 48020 11228 48076 11238
rect 48020 10332 48076 11172
rect 48020 9894 48076 10276
rect 47964 9882 48076 9894
rect 47964 9830 47966 9882
rect 48018 9830 48076 9882
rect 47964 9828 48076 9830
rect 47964 9818 48020 9828
rect 48244 9098 48300 9110
rect 48244 9046 48246 9098
rect 48298 9046 48300 9098
rect 48244 8988 48300 9046
rect 48244 8922 48300 8932
rect 47684 8314 47852 8316
rect 47684 8262 47686 8314
rect 47738 8262 47852 8314
rect 47684 8260 47852 8262
rect 48244 8652 48300 8662
rect 47684 8250 47740 8260
rect 48244 8202 48300 8596
rect 48468 8316 48524 11956
rect 48580 9210 48636 12180
rect 49028 11788 49084 14200
rect 49812 13354 49868 14200
rect 50484 13468 50540 14200
rect 49812 13302 49814 13354
rect 49866 13302 49868 13354
rect 49812 13290 49868 13302
rect 50372 13412 50540 13468
rect 50260 11900 50316 11910
rect 49028 11722 49084 11732
rect 49812 11788 49868 11798
rect 49028 11338 49084 11350
rect 49028 11286 49030 11338
rect 49082 11286 49084 11338
rect 48860 10332 48916 10342
rect 48860 9884 48916 10276
rect 48580 9158 48582 9210
rect 48634 9158 48636 9210
rect 48580 9146 48636 9158
rect 48804 9882 48916 9884
rect 48804 9830 48862 9882
rect 48914 9830 48916 9882
rect 48804 9818 48916 9830
rect 48804 8652 48860 9818
rect 48804 8586 48860 8596
rect 48580 8316 48636 8326
rect 48468 8314 48636 8316
rect 48468 8262 48582 8314
rect 48634 8262 48636 8314
rect 48468 8260 48636 8262
rect 48580 8250 48636 8260
rect 48244 8150 48246 8202
rect 48298 8150 48300 8202
rect 48244 8138 48300 8150
rect 46452 8090 46732 8092
rect 46452 8038 46454 8090
rect 46506 8038 46732 8090
rect 46452 8036 46732 8038
rect 46452 8026 46508 8036
rect 46228 7644 46284 7654
rect 46228 7550 46284 7588
rect 46564 5906 46620 5918
rect 46564 5854 46566 5906
rect 46618 5854 46620 5906
rect 46564 5852 46620 5854
rect 46564 5786 46620 5796
rect 46564 5010 46620 5022
rect 46564 4958 46566 5010
rect 46618 4958 46620 5010
rect 46564 2604 46620 4958
rect 46564 2538 46620 2548
rect 46004 1318 46006 1370
rect 46058 1318 46060 1370
rect 46004 1306 46060 1318
rect 46452 1596 46508 1606
rect 46452 800 46508 1540
rect 44212 298 44268 308
rect 44632 0 44744 800
rect 45192 0 45304 800
rect 45864 0 45976 800
rect 46424 0 46536 800
rect 46676 588 46732 8036
rect 47348 8092 47404 8102
rect 47348 7998 47404 8036
rect 47124 7644 47180 7654
rect 47124 6086 47180 7588
rect 47684 7474 47740 7486
rect 47684 7422 47686 7474
rect 47738 7422 47740 7474
rect 47404 6748 47460 6758
rect 47404 6654 47460 6692
rect 47068 6074 47180 6086
rect 47068 6022 47070 6074
rect 47122 6022 47180 6074
rect 47068 6020 47180 6022
rect 47068 5852 47124 6020
rect 47684 5852 47740 7422
rect 48580 7455 48636 7467
rect 48580 7403 48582 7455
rect 48634 7403 48636 7455
rect 48356 6860 48412 6870
rect 48356 6766 48412 6804
rect 48356 6578 48412 6590
rect 48356 6526 48358 6578
rect 48410 6526 48412 6578
rect 48188 5852 48244 5862
rect 47684 5850 48244 5852
rect 47684 5798 48190 5850
rect 48242 5798 48244 5850
rect 47684 5796 48244 5798
rect 47068 5786 47124 5796
rect 48132 5786 48244 5796
rect 46900 5122 46956 5134
rect 46900 5070 46902 5122
rect 46954 5070 46956 5122
rect 46900 4620 46956 5070
rect 46900 4554 46956 4564
rect 48132 3387 48188 5786
rect 48356 4844 48412 6526
rect 48580 6198 48636 7403
rect 49028 6748 49084 11286
rect 49308 8988 49364 8998
rect 49308 8894 49364 8932
rect 49812 7642 49868 11732
rect 50036 10554 50092 10566
rect 50036 10502 50038 10554
rect 50090 10502 50092 10554
rect 49924 9324 49980 9334
rect 49924 9210 49980 9268
rect 49924 9158 49926 9210
rect 49978 9158 49980 9210
rect 49924 9146 49980 9158
rect 50036 8314 50092 10502
rect 50260 9210 50316 11844
rect 50372 11788 50428 13412
rect 51044 13244 51100 14422
rect 51240 14200 51352 15000
rect 51912 14200 52024 15000
rect 52696 14200 52808 15000
rect 52948 14700 53004 14710
rect 52948 14588 53004 14644
rect 52948 14532 53228 14588
rect 53060 14250 53116 14262
rect 51044 13178 51100 13188
rect 51268 12012 51324 14200
rect 51940 12458 51996 14200
rect 51940 12406 51942 12458
rect 51994 12406 51996 12458
rect 51940 12394 51996 12406
rect 52724 12124 52780 14200
rect 53060 14198 53062 14250
rect 53114 14198 53116 14250
rect 53060 13244 53116 14198
rect 53172 14140 53228 14532
rect 53368 14200 53480 15000
rect 53620 14700 53676 14710
rect 53396 14140 53452 14200
rect 53172 14084 53452 14140
rect 53060 13178 53116 13188
rect 52724 12058 52780 12068
rect 51268 11946 51324 11956
rect 52500 12012 52556 12022
rect 50372 11722 50428 11732
rect 51156 11676 51212 11686
rect 51044 11562 51100 11574
rect 51044 11510 51046 11562
rect 51098 11510 51100 11562
rect 50596 11450 50652 11462
rect 50596 11398 50598 11450
rect 50650 11398 50652 11450
rect 50596 9894 50652 11398
rect 50540 9882 50652 9894
rect 50540 9830 50542 9882
rect 50594 9830 50652 9882
rect 50540 9828 50652 9830
rect 50820 10332 50876 10342
rect 50540 9324 50596 9828
rect 50540 9258 50596 9268
rect 50708 9548 50764 9558
rect 50260 9158 50262 9210
rect 50314 9158 50316 9210
rect 50260 9146 50316 9158
rect 50036 8262 50038 8314
rect 50090 8262 50092 8314
rect 50036 8250 50092 8262
rect 49812 7590 49814 7642
rect 49866 7590 49868 7642
rect 50708 7698 50764 9492
rect 50820 9210 50876 10276
rect 50820 9158 50822 9210
rect 50874 9158 50876 9210
rect 50820 9146 50876 9158
rect 50708 7646 50710 7698
rect 50762 7646 50764 7698
rect 50708 7634 50764 7646
rect 49812 7578 49868 7590
rect 49028 6690 49084 6692
rect 49028 6638 49030 6690
rect 49082 6638 49084 6690
rect 49028 6616 49084 6638
rect 49476 7530 49532 7542
rect 49476 7478 49478 7530
rect 49530 7478 49532 7530
rect 49476 6748 49532 7478
rect 51044 6758 51100 11510
rect 51156 9210 51212 11620
rect 51828 10444 51884 10454
rect 51604 10332 51660 10342
rect 51604 9222 51660 10276
rect 51156 9158 51158 9210
rect 51210 9158 51212 9210
rect 51156 9146 51212 9158
rect 51548 9210 51660 9222
rect 51548 9158 51550 9210
rect 51602 9158 51660 9210
rect 51548 9156 51660 9158
rect 51548 9146 51604 9156
rect 51604 8258 51660 8270
rect 51604 8206 51606 8258
rect 51658 8206 51660 8258
rect 51604 6860 51660 8206
rect 51828 8204 51884 10388
rect 52164 10108 52220 10118
rect 52164 9210 52220 10052
rect 52164 9158 52166 9210
rect 52218 9158 52220 9210
rect 52164 9146 52220 9158
rect 52500 9210 52556 11956
rect 53620 12012 53676 14644
rect 54152 14200 54264 15000
rect 54404 14924 54460 14934
rect 54404 14812 54460 14868
rect 54404 14756 54684 14812
rect 53844 13468 53900 13478
rect 53844 13374 53900 13412
rect 54180 12346 54236 14200
rect 54628 14140 54684 14756
rect 54824 14200 54936 15000
rect 55608 14200 55720 15000
rect 56392 14200 56504 15000
rect 57064 14200 57176 15000
rect 57848 14200 57960 15000
rect 58324 14364 58380 14374
rect 54852 14140 54908 14200
rect 54628 14084 54908 14140
rect 54404 13578 54460 13590
rect 54404 13526 54406 13578
rect 54458 13526 54460 13578
rect 54404 13356 54460 13526
rect 54404 13290 54460 13300
rect 54180 12294 54182 12346
rect 54234 12294 54236 12346
rect 54180 12282 54236 12294
rect 55636 12348 55692 14200
rect 55748 13690 55804 13702
rect 55748 13638 55750 13690
rect 55802 13638 55804 13690
rect 55748 13356 55804 13638
rect 55748 13290 55804 13300
rect 55972 13242 56028 13254
rect 55972 13190 55974 13242
rect 56026 13190 56028 13242
rect 55972 12908 56028 13190
rect 55972 12842 56028 12852
rect 56420 12570 56476 14200
rect 57092 13804 57148 14200
rect 57092 13738 57148 13748
rect 57540 14138 57596 14150
rect 57540 14086 57542 14138
rect 57594 14086 57596 14138
rect 56420 12518 56422 12570
rect 56474 12518 56476 12570
rect 56420 12506 56476 12518
rect 56980 12794 57036 12806
rect 56980 12742 56982 12794
rect 57034 12742 57036 12794
rect 55636 12282 55692 12292
rect 53620 11946 53676 11956
rect 54404 12012 54460 12022
rect 53396 11114 53452 11126
rect 53396 11062 53398 11114
rect 53450 11062 53452 11114
rect 53284 10556 53340 10566
rect 52780 10108 52836 10118
rect 52780 9882 52836 10052
rect 52780 9830 52782 9882
rect 52834 9830 52836 9882
rect 52780 9818 52836 9830
rect 52500 9158 52502 9210
rect 52554 9158 52556 9210
rect 52500 9146 52556 9158
rect 52500 8988 52556 8998
rect 52388 8932 52500 8988
rect 51828 8138 51884 8148
rect 52164 8540 52220 8550
rect 51940 7586 51996 7598
rect 51940 7534 51942 7586
rect 51994 7534 51996 7586
rect 51940 7532 51996 7534
rect 51940 7476 52108 7532
rect 51604 6794 51660 6804
rect 49868 6748 49924 6758
rect 50988 6748 51100 6758
rect 49476 6746 49924 6748
rect 49476 6694 49870 6746
rect 49922 6694 49924 6746
rect 49476 6692 49924 6694
rect 48580 6188 48692 6198
rect 48580 6132 48636 6188
rect 48636 6074 48692 6132
rect 48636 6022 48638 6074
rect 48690 6022 48692 6074
rect 48636 6010 48692 6022
rect 48356 4778 48412 4788
rect 48748 4954 48804 4966
rect 48748 4902 48750 4954
rect 48802 4902 48804 4954
rect 48748 4620 48804 4902
rect 48748 4554 48804 4564
rect 47124 3331 48188 3387
rect 47124 800 47180 3331
rect 49476 2154 49532 6692
rect 49868 6682 49924 6692
rect 50540 6746 51100 6748
rect 50540 6694 50990 6746
rect 51042 6694 51100 6746
rect 50540 6692 51100 6694
rect 51772 6748 51828 6758
rect 50540 6690 50596 6692
rect 50540 6638 50542 6690
rect 50594 6638 50596 6690
rect 50988 6682 51044 6692
rect 51772 6654 51828 6692
rect 50540 6626 50596 6638
rect 52052 6534 52108 7476
rect 52164 7474 52220 8484
rect 52164 7422 52166 7474
rect 52218 7422 52220 7474
rect 52164 6748 52220 7422
rect 52164 6682 52220 6692
rect 50428 6524 50484 6534
rect 50372 6522 50484 6524
rect 50372 6470 50430 6522
rect 50482 6470 50484 6522
rect 50372 6458 50484 6470
rect 52052 6522 52164 6534
rect 52052 6470 52110 6522
rect 52162 6470 52164 6522
rect 52052 6458 52164 6470
rect 50372 5852 50428 6458
rect 49812 5794 49868 5806
rect 49812 5742 49814 5794
rect 49866 5742 49868 5794
rect 50372 5786 50428 5796
rect 51044 5906 51100 5918
rect 51044 5854 51046 5906
rect 51098 5854 51100 5906
rect 51044 5852 51100 5854
rect 51044 5786 51100 5796
rect 51548 5852 51604 5862
rect 51548 5758 51604 5796
rect 49812 5068 49868 5742
rect 52052 5628 52108 6458
rect 52220 5852 52276 5862
rect 52220 5850 52332 5852
rect 52220 5798 52222 5850
rect 52274 5798 52332 5850
rect 52220 5786 52332 5798
rect 52052 5562 52108 5572
rect 51828 5122 51884 5134
rect 51828 5070 51830 5122
rect 51882 5070 51884 5122
rect 49812 5002 49868 5012
rect 50484 5010 50540 5022
rect 49644 4954 49700 4966
rect 49644 4902 49646 4954
rect 49698 4902 49700 4954
rect 49644 4844 49700 4902
rect 50484 4958 50486 5010
rect 50538 4958 50540 5010
rect 49700 4788 49756 4844
rect 49644 4778 49756 4788
rect 49588 3946 49644 3958
rect 49588 3894 49590 3946
rect 49642 3894 49644 3946
rect 49588 2940 49644 3894
rect 49700 3724 49756 4778
rect 49700 3658 49756 3668
rect 49588 2874 49644 2884
rect 50484 2492 50540 4958
rect 51828 5012 51884 5070
rect 51828 4956 52108 5012
rect 52052 4732 52108 4956
rect 52052 4666 52108 4676
rect 52276 4844 52332 5786
rect 52276 3387 52332 4788
rect 52388 3948 52444 8932
rect 52500 8922 52556 8932
rect 53284 8874 53340 10500
rect 53284 8822 53286 8874
rect 53338 8822 53340 8874
rect 53284 8810 53340 8822
rect 52612 8258 52668 8270
rect 52612 8206 52614 8258
rect 52666 8206 52668 8258
rect 52612 7430 52668 8206
rect 52612 7418 52724 7430
rect 52612 7366 52670 7418
rect 52722 7366 52724 7418
rect 52612 7364 52724 7366
rect 52668 7084 52724 7364
rect 53396 7306 53452 11062
rect 54292 10666 54348 10678
rect 54292 10614 54294 10666
rect 54346 10614 54348 10666
rect 54180 10332 54236 10342
rect 53564 9772 53620 9782
rect 53564 9678 53620 9716
rect 53564 8092 53620 8102
rect 54068 8092 54124 8102
rect 53564 8090 54124 8092
rect 53564 8038 53566 8090
rect 53618 8038 54070 8090
rect 54122 8038 54124 8090
rect 53564 8036 54124 8038
rect 53564 8026 53620 8036
rect 54068 7980 54124 8036
rect 54068 7914 54124 7924
rect 53396 7254 53398 7306
rect 53450 7254 53452 7306
rect 53396 7242 53452 7254
rect 52668 7018 52724 7028
rect 52556 6860 52612 6870
rect 52556 6524 52612 6804
rect 52556 6430 52612 6468
rect 53844 6636 53900 6646
rect 52668 4956 52724 4966
rect 52668 4954 52780 4956
rect 52668 4902 52670 4954
rect 52722 4902 52780 4954
rect 52668 4890 52780 4902
rect 52388 3882 52444 3892
rect 52724 4732 52780 4890
rect 52724 3948 52780 4676
rect 52724 3882 52780 3892
rect 52164 3331 52332 3387
rect 52500 3722 52556 3734
rect 52500 3670 52502 3722
rect 52554 3670 52556 3722
rect 51940 2938 51996 2950
rect 51940 2886 51942 2938
rect 51994 2886 51996 2938
rect 50484 2426 50540 2436
rect 50708 2604 50764 2614
rect 49476 2102 49478 2154
rect 49530 2102 49532 2154
rect 49476 2090 49532 2102
rect 48356 1932 48412 1942
rect 47684 1596 47740 1606
rect 47684 800 47740 1540
rect 48356 800 48412 1876
rect 49476 1484 49532 1494
rect 48916 1372 48972 1382
rect 48916 800 48972 1316
rect 49476 800 49532 1428
rect 50148 1148 50204 1158
rect 50148 800 50204 1092
rect 50708 800 50764 2548
rect 51380 2266 51436 2278
rect 51380 2214 51382 2266
rect 51434 2214 51436 2266
rect 51380 800 51436 2214
rect 51940 800 51996 2886
rect 52164 1596 52220 3331
rect 52500 3164 52556 3670
rect 52500 3098 52556 3108
rect 52164 1530 52220 1540
rect 53172 1708 53228 1718
rect 52388 868 52668 924
rect 46676 522 46732 532
rect 47096 0 47208 800
rect 47656 0 47768 800
rect 48328 0 48440 800
rect 48888 0 49000 800
rect 49448 0 49560 800
rect 49924 476 49980 486
rect 49924 382 49980 420
rect 50120 0 50232 800
rect 50680 0 50792 800
rect 51352 0 51464 800
rect 51912 0 52024 800
rect 52388 700 52444 868
rect 52612 800 52668 868
rect 53172 800 53228 1652
rect 53844 800 53900 6580
rect 54180 5738 54236 10276
rect 54292 6746 54348 10614
rect 54404 8314 54460 11956
rect 55188 11898 55244 11910
rect 55188 11846 55190 11898
rect 55242 11846 55244 11898
rect 54516 9996 54572 10006
rect 54516 9902 54572 9940
rect 55188 9826 55244 11846
rect 56980 11674 57036 12742
rect 57092 12124 57148 12134
rect 57092 11786 57148 12068
rect 57092 11734 57094 11786
rect 57146 11734 57148 11786
rect 57092 11722 57148 11734
rect 56980 11622 56982 11674
rect 57034 11622 57036 11674
rect 56980 11610 57036 11622
rect 56308 10444 56364 10454
rect 55188 9774 55190 9826
rect 55242 9774 55244 9826
rect 55188 9772 55244 9774
rect 55188 9696 55244 9716
rect 55412 9826 55468 9838
rect 55412 9774 55414 9826
rect 55466 9774 55468 9826
rect 55412 9772 55468 9774
rect 55412 9706 55468 9716
rect 55540 9436 55804 9446
rect 55596 9380 55644 9436
rect 55700 9380 55748 9436
rect 55540 9370 55804 9380
rect 54404 8262 54406 8314
rect 54458 8262 54460 8314
rect 54404 8250 54460 8262
rect 54852 9212 54908 9222
rect 54852 9042 54908 9156
rect 54852 8990 54854 9042
rect 54906 8990 54908 9042
rect 54852 7308 54908 8990
rect 56308 8428 56364 10388
rect 56588 9772 56644 9782
rect 56588 9678 56644 9716
rect 57036 9658 57092 9670
rect 57372 9660 57428 9670
rect 57036 9606 57038 9658
rect 57090 9606 57092 9658
rect 56420 9548 56476 9558
rect 56420 9053 56476 9492
rect 57036 9548 57092 9606
rect 57036 9482 57092 9492
rect 57316 9658 57428 9660
rect 57316 9606 57374 9658
rect 57426 9606 57428 9658
rect 57316 9594 57428 9606
rect 57316 9212 57372 9594
rect 57316 9146 57372 9156
rect 56420 9001 56422 9053
rect 56474 9001 56476 9053
rect 56420 8989 56476 9001
rect 57428 9098 57484 9110
rect 57428 9046 57430 9098
rect 57482 9046 57484 9098
rect 57428 8988 57484 9046
rect 57428 8922 57484 8932
rect 56420 8428 56476 8438
rect 56308 8426 56476 8428
rect 56308 8374 56422 8426
rect 56474 8374 56476 8426
rect 56308 8372 56476 8374
rect 56420 8362 56476 8372
rect 56756 8258 56812 8270
rect 56756 8206 56758 8258
rect 56810 8206 56812 8258
rect 56644 7980 56700 7990
rect 55540 7868 55804 7878
rect 55596 7812 55644 7868
rect 55700 7812 55748 7868
rect 55540 7802 55804 7812
rect 54292 6694 54294 6746
rect 54346 6694 54348 6746
rect 54292 6682 54348 6694
rect 54404 7252 54908 7308
rect 54964 7474 55020 7486
rect 54964 7422 54966 7474
rect 55018 7422 55020 7474
rect 54180 5686 54182 5738
rect 54234 5686 54236 5738
rect 54180 5674 54236 5686
rect 54404 800 54460 7252
rect 54964 6636 55020 7422
rect 56644 7474 56700 7924
rect 56644 7422 56646 7474
rect 56698 7422 56700 7474
rect 56644 7410 56700 7422
rect 56756 7308 56812 8206
rect 56084 7252 56812 7308
rect 54964 6570 55020 6580
rect 55188 6690 55244 6702
rect 55188 6638 55190 6690
rect 55242 6638 55244 6690
rect 54516 5906 54572 5918
rect 54516 5854 54518 5906
rect 54570 5854 54572 5906
rect 54516 4844 54572 5854
rect 54516 4778 54572 4788
rect 54740 5010 54796 5022
rect 54740 4958 54742 5010
rect 54794 4958 54796 5010
rect 54628 4732 54684 4742
rect 54628 1708 54684 4676
rect 54628 1642 54684 1652
rect 52164 644 52444 700
rect 52164 588 52220 644
rect 52164 522 52220 532
rect 52584 0 52696 800
rect 53144 0 53256 800
rect 53816 0 53928 800
rect 54376 0 54488 800
rect 54740 138 54796 4958
rect 55188 4732 55244 6638
rect 55540 6300 55804 6310
rect 55596 6244 55644 6300
rect 55700 6244 55748 6300
rect 55540 6234 55804 6244
rect 55748 5180 55804 5190
rect 55748 5122 55804 5124
rect 55748 5070 55750 5122
rect 55802 5070 55804 5122
rect 55748 5058 55804 5070
rect 55188 4284 55244 4676
rect 55540 4732 55804 4742
rect 55596 4676 55644 4732
rect 55700 4676 55748 4732
rect 55540 4666 55804 4676
rect 55188 4218 55244 4228
rect 55076 3836 55132 3846
rect 55076 3742 55132 3780
rect 55636 1820 55692 1830
rect 55076 1596 55132 1606
rect 54964 1540 55076 1596
rect 54964 800 55020 1540
rect 55076 1530 55132 1540
rect 55636 800 55692 1764
rect 56084 1708 56140 7252
rect 56756 6860 56812 7252
rect 56756 6794 56812 6804
rect 56868 7756 56924 7766
rect 56756 6679 56812 6691
rect 56588 6636 56644 6646
rect 56420 6524 56476 6534
rect 56196 5902 56252 5914
rect 56196 5850 56198 5902
rect 56250 5850 56252 5902
rect 56196 5628 56252 5850
rect 56196 5562 56252 5572
rect 56196 5180 56252 5190
rect 56196 4060 56252 5124
rect 56196 3994 56252 4004
rect 56196 3276 56252 3286
rect 56196 3182 56252 3220
rect 55972 1652 56140 1708
rect 56196 1932 56252 1942
rect 55972 1596 56028 1652
rect 55972 1530 56028 1540
rect 56196 800 56252 1876
rect 56420 1708 56476 6468
rect 56588 6074 56644 6580
rect 56756 6627 56758 6679
rect 56810 6627 56812 6679
rect 56756 6412 56812 6627
rect 56868 6636 56924 7700
rect 57540 7756 57596 14086
rect 57764 13244 57820 13254
rect 57540 7690 57596 7700
rect 57652 10780 57708 10790
rect 57428 7362 57484 7374
rect 57428 7310 57430 7362
rect 57482 7310 57484 7362
rect 57428 6860 57484 7310
rect 57092 6804 57484 6860
rect 56868 6570 56924 6580
rect 56980 6748 57036 6758
rect 56980 6412 57036 6692
rect 56756 6356 57036 6412
rect 56588 6022 56590 6074
rect 56642 6022 56644 6074
rect 56588 6010 56644 6022
rect 56980 5068 57036 6356
rect 57092 5404 57148 6804
rect 57484 6580 57540 6590
rect 57652 6580 57708 10724
rect 57764 9210 57820 13188
rect 57876 11788 57932 14200
rect 58324 14140 58380 14308
rect 58520 14200 58632 15000
rect 58772 14588 58828 14598
rect 58772 14476 58828 14532
rect 58772 14420 59164 14476
rect 58324 14074 58380 14084
rect 58212 13690 58268 13702
rect 58212 13638 58214 13690
rect 58266 13638 58268 13690
rect 58212 13132 58268 13638
rect 58212 13066 58268 13076
rect 58548 12794 58604 14200
rect 59108 14140 59164 14420
rect 59304 14200 59416 15000
rect 59976 14200 60088 15000
rect 60760 14200 60872 15000
rect 61432 14200 61544 15000
rect 62216 14200 62328 15000
rect 62888 14200 63000 15000
rect 63140 14924 63196 14934
rect 63140 14698 63196 14868
rect 63140 14646 63142 14698
rect 63194 14646 63196 14698
rect 63140 14634 63196 14646
rect 63252 14922 63308 14934
rect 63252 14870 63254 14922
rect 63306 14870 63308 14922
rect 59332 14140 59388 14200
rect 59108 14084 59388 14140
rect 60004 13020 60060 14200
rect 60004 12954 60060 12964
rect 60452 13468 60508 13478
rect 58548 12742 58550 12794
rect 58602 12742 58604 12794
rect 58548 12730 58604 12742
rect 59220 12684 59276 12694
rect 58324 12010 58380 12022
rect 58324 11958 58326 12010
rect 58378 11958 58380 12010
rect 57876 11722 57932 11732
rect 58100 11788 58156 11798
rect 58100 11340 58156 11732
rect 58100 11274 58156 11284
rect 58324 11340 58380 11958
rect 58324 11274 58380 11284
rect 58044 9660 58100 9670
rect 57764 9158 57766 9210
rect 57818 9158 57820 9210
rect 57764 9146 57820 9158
rect 57988 9658 58100 9660
rect 57988 9606 58046 9658
rect 58098 9606 58100 9658
rect 57988 9594 58100 9606
rect 57988 8988 58044 9594
rect 58380 9100 58436 9110
rect 58828 9100 58884 9110
rect 58380 9098 58828 9100
rect 58380 9046 58382 9098
rect 58434 9046 58828 9098
rect 58380 9044 58828 9046
rect 58380 9034 58436 9044
rect 58828 8968 58884 9044
rect 57988 8922 58044 8932
rect 58268 8876 58324 8886
rect 58268 8782 58324 8820
rect 58996 8428 59052 8438
rect 58436 8258 58492 8270
rect 58436 8206 58438 8258
rect 58490 8206 58492 8258
rect 58436 7868 58492 8206
rect 58996 8202 59052 8372
rect 59220 8316 59276 12628
rect 60452 11900 60508 13412
rect 60788 13020 60844 14200
rect 60788 12954 60844 12964
rect 61236 13692 61292 13702
rect 61236 12010 61292 13636
rect 61460 12236 61516 14200
rect 61460 12170 61516 12180
rect 61684 14138 61740 14150
rect 61684 14086 61686 14138
rect 61738 14086 61740 14138
rect 61236 11958 61238 12010
rect 61290 11958 61292 12010
rect 61236 11946 61292 11958
rect 60452 11834 60508 11844
rect 60788 10778 60844 10790
rect 60788 10726 60790 10778
rect 60842 10726 60844 10778
rect 60788 10668 60844 10726
rect 60788 10602 60844 10612
rect 61012 10778 61068 10790
rect 61012 10726 61014 10778
rect 61066 10726 61068 10778
rect 60788 10108 60844 10118
rect 60564 9772 60620 9782
rect 60452 9100 60508 9110
rect 59388 8988 59444 8998
rect 59388 8894 59444 8932
rect 60452 8540 60508 9044
rect 60564 8652 60620 9716
rect 60564 8586 60620 8596
rect 60788 8652 60844 10052
rect 61012 9212 61068 10726
rect 61012 9146 61068 9156
rect 61236 9212 61292 9222
rect 61236 9118 61292 9156
rect 61572 9212 61628 9222
rect 61684 9212 61740 14086
rect 61796 13692 61852 13702
rect 61796 11338 61852 13636
rect 62244 12908 62300 14200
rect 62916 14140 62972 14200
rect 63252 14140 63308 14870
rect 63672 14200 63784 15000
rect 64036 14698 64092 14710
rect 64036 14646 64038 14698
rect 64090 14646 64092 14698
rect 62916 14084 63308 14140
rect 63700 13468 63756 14200
rect 64036 14026 64092 14646
rect 64148 14364 64204 14374
rect 64148 14138 64204 14308
rect 64344 14200 64456 15000
rect 65128 14200 65240 15000
rect 65380 14588 65436 14598
rect 65380 14476 65436 14532
rect 65380 14420 65660 14476
rect 64148 14086 64150 14138
rect 64202 14086 64204 14138
rect 64148 14074 64204 14086
rect 64036 13974 64038 14026
rect 64090 13974 64092 14026
rect 64036 13962 64092 13974
rect 63700 13402 63756 13412
rect 64260 13580 64316 13590
rect 62244 12842 62300 12852
rect 63700 12124 63756 12134
rect 63700 12030 63756 12068
rect 63364 11900 63420 11910
rect 62356 11788 62412 11798
rect 62356 11564 62412 11732
rect 62356 11498 62412 11508
rect 61796 11286 61798 11338
rect 61850 11286 61852 11338
rect 61796 11274 61852 11286
rect 62356 11338 62412 11350
rect 62356 11286 62358 11338
rect 62410 11286 62412 11338
rect 61572 9210 61740 9212
rect 61572 9158 61574 9210
rect 61626 9158 61740 9210
rect 61572 9156 61740 9158
rect 61964 9212 62020 9222
rect 61572 9146 61628 9156
rect 61964 9118 62020 9156
rect 60788 8586 60844 8596
rect 60452 8474 60508 8484
rect 59444 8428 59500 8438
rect 59332 8316 59388 8326
rect 59220 8314 59388 8316
rect 59220 8262 59334 8314
rect 59386 8262 59388 8314
rect 59220 8260 59388 8262
rect 59332 8250 59388 8260
rect 58996 8150 58998 8202
rect 59050 8150 59052 8202
rect 58996 8138 59052 8150
rect 58436 7802 58492 7812
rect 58324 7756 58380 7766
rect 58044 7308 58100 7318
rect 58044 6858 58100 7252
rect 58324 7308 58380 7700
rect 58660 7756 58716 7766
rect 58660 7586 58716 7700
rect 58660 7534 58662 7586
rect 58714 7534 58716 7586
rect 58660 7522 58716 7534
rect 59332 7756 59388 7766
rect 58324 7242 58380 7252
rect 58996 7474 59052 7486
rect 58996 7422 58998 7474
rect 59050 7422 59052 7474
rect 58044 6806 58046 6858
rect 58098 6806 58100 6858
rect 58044 6794 58100 6806
rect 58604 6860 58660 6870
rect 58604 6634 58660 6804
rect 57484 6578 57708 6580
rect 57372 6524 57428 6534
rect 57204 6522 57428 6524
rect 57204 6470 57374 6522
rect 57426 6470 57428 6522
rect 57484 6526 57486 6578
rect 57538 6526 57708 6578
rect 57484 6524 57708 6526
rect 57484 6514 57540 6524
rect 57204 6468 57428 6470
rect 57204 5516 57260 6468
rect 57372 6458 57428 6468
rect 57372 6300 57428 6310
rect 57372 6074 57428 6244
rect 57372 6022 57374 6074
rect 57426 6022 57428 6074
rect 57372 6010 57428 6022
rect 57652 6086 57708 6524
rect 58156 6578 58212 6590
rect 58156 6526 58158 6578
rect 58210 6526 58212 6578
rect 58604 6582 58606 6634
rect 58658 6582 58660 6634
rect 58604 6570 58660 6582
rect 58156 6300 58212 6526
rect 58996 6524 59052 7422
rect 59332 6646 59388 7700
rect 59444 7654 59500 8372
rect 62356 8314 62412 11286
rect 62804 9098 62860 9110
rect 62804 9046 62806 9098
rect 62858 9046 62860 9098
rect 62804 8652 62860 9046
rect 63140 8876 63196 8886
rect 63364 8876 63420 11844
rect 63924 11564 63980 11574
rect 63532 8988 63588 8998
rect 63532 8986 63644 8988
rect 63532 8934 63534 8986
rect 63586 8934 63644 8986
rect 63532 8922 63644 8934
rect 63140 8874 63420 8876
rect 63140 8822 63142 8874
rect 63194 8822 63420 8874
rect 63140 8820 63420 8822
rect 63140 8810 63196 8820
rect 63588 8652 63644 8922
rect 62804 8596 63644 8652
rect 62356 8262 62358 8314
rect 62410 8262 62412 8314
rect 62356 8250 62412 8262
rect 63252 8258 63308 8270
rect 60508 8204 60564 8214
rect 59948 8146 60004 8158
rect 59836 8092 59892 8102
rect 59780 8090 59892 8092
rect 59780 8038 59838 8090
rect 59890 8038 59892 8090
rect 59780 8026 59892 8038
rect 59948 8094 59950 8146
rect 60002 8094 60004 8146
rect 59444 7642 59556 7654
rect 59444 7590 59502 7642
rect 59554 7590 59556 7642
rect 59444 7588 59556 7590
rect 59500 7578 59556 7588
rect 59780 7420 59836 8026
rect 59948 7644 60004 8094
rect 60508 8090 60564 8148
rect 63252 8206 63254 8258
rect 63306 8206 63308 8258
rect 63252 8204 63308 8206
rect 63252 8138 63308 8148
rect 60508 8038 60510 8090
rect 60562 8038 60564 8090
rect 59948 7588 60060 7644
rect 60004 7420 60060 7588
rect 60508 7532 60564 8038
rect 62916 7756 62972 7766
rect 62916 7586 62972 7700
rect 62916 7534 62918 7586
rect 62970 7534 62972 7586
rect 63420 7756 63476 7766
rect 63420 7642 63476 7700
rect 63420 7590 63422 7642
rect 63474 7590 63476 7642
rect 63420 7578 63476 7590
rect 60508 7476 60844 7532
rect 62916 7522 62972 7534
rect 60172 7420 60228 7430
rect 60004 7418 60228 7420
rect 60004 7366 60174 7418
rect 60226 7366 60228 7418
rect 60004 7364 60228 7366
rect 59780 7354 59836 7364
rect 60116 7354 60228 7364
rect 59332 6634 59444 6646
rect 59332 6582 59390 6634
rect 59442 6582 59444 6634
rect 59332 6580 59444 6582
rect 59388 6570 59444 6580
rect 58996 6458 59052 6468
rect 59948 6524 60004 6534
rect 59948 6430 60004 6468
rect 58380 6300 58436 6310
rect 60116 6300 60172 7354
rect 60676 6636 60732 6646
rect 58156 6244 58380 6300
rect 57652 6074 57764 6086
rect 57652 6022 57710 6074
rect 57762 6022 57764 6074
rect 57652 6020 57764 6022
rect 57708 6010 57764 6020
rect 58380 6074 58436 6244
rect 58380 6022 58382 6074
rect 58434 6022 58436 6074
rect 58380 6010 58436 6022
rect 60004 6244 60172 6300
rect 60228 6580 60676 6636
rect 58828 5852 58884 5862
rect 57204 5450 57260 5460
rect 58772 5850 58884 5852
rect 58772 5798 58830 5850
rect 58882 5798 58884 5850
rect 58772 5786 58884 5798
rect 57092 5338 57148 5348
rect 58660 5404 58716 5414
rect 58660 5122 58716 5348
rect 58660 5070 58662 5122
rect 58714 5070 58716 5122
rect 56980 5012 57148 5068
rect 58660 5058 58716 5070
rect 56588 4956 56644 4966
rect 57092 4956 57148 5012
rect 58324 5010 58380 5022
rect 57372 4956 57428 4966
rect 57092 4954 57428 4956
rect 57092 4902 57374 4954
rect 57426 4902 57428 4954
rect 57092 4900 57428 4902
rect 56588 4862 56644 4900
rect 57372 4890 57428 4900
rect 57988 4956 58044 4966
rect 57092 4060 57148 4070
rect 57092 3966 57148 4004
rect 57316 4060 57372 4070
rect 56644 3834 56700 3846
rect 56644 3782 56646 3834
rect 56698 3782 56700 3834
rect 56644 2492 56700 3782
rect 57316 3612 57372 4004
rect 57316 3546 57372 3556
rect 57876 3162 57932 3174
rect 57876 3110 57878 3162
rect 57930 3110 57932 3162
rect 56980 2716 57036 2726
rect 56980 2492 57036 2660
rect 56644 2436 57036 2492
rect 56420 1642 56476 1652
rect 56868 2268 56924 2278
rect 56868 800 56924 2212
rect 57876 2044 57932 3110
rect 57988 2156 58044 4900
rect 58324 4958 58326 5010
rect 58378 4958 58380 5010
rect 58324 4058 58380 4958
rect 58772 4284 58828 5786
rect 58772 4218 58828 4228
rect 58884 4172 58940 4182
rect 58324 4006 58326 4058
rect 58378 4006 58380 4058
rect 58324 3994 58380 4006
rect 58660 4058 58716 4070
rect 58660 4006 58662 4058
rect 58714 4006 58716 4058
rect 58100 3162 58156 3174
rect 58100 3110 58102 3162
rect 58154 3110 58156 3162
rect 58100 2602 58156 3110
rect 58660 2826 58716 4006
rect 58660 2774 58662 2826
rect 58714 2774 58716 2826
rect 58660 2762 58716 2774
rect 58100 2550 58102 2602
rect 58154 2550 58156 2602
rect 58100 2538 58156 2550
rect 58884 2602 58940 4116
rect 59444 4172 59500 4182
rect 59444 4058 59500 4116
rect 59444 4006 59446 4058
rect 59498 4006 59500 4058
rect 59444 3994 59500 4006
rect 58884 2550 58886 2602
rect 58938 2550 58940 2602
rect 58884 2538 58940 2550
rect 59668 3722 59724 3734
rect 59668 3670 59670 3722
rect 59722 3670 59724 3722
rect 59668 2604 59724 3670
rect 60004 3387 60060 6244
rect 60228 5012 60284 6580
rect 60676 6570 60732 6580
rect 59892 3331 60060 3387
rect 60116 4956 60284 5012
rect 60508 5404 60564 5414
rect 59892 2716 59948 3331
rect 60116 3052 60172 4956
rect 60508 4954 60564 5348
rect 60508 4902 60510 4954
rect 60562 4902 60564 4954
rect 60508 4890 60564 4902
rect 60676 5180 60732 5190
rect 60228 4732 60284 4742
rect 60228 3164 60284 4676
rect 60676 4060 60732 5124
rect 60676 3994 60732 4004
rect 60340 3836 60396 3846
rect 60340 3276 60396 3780
rect 60788 3387 60844 7476
rect 63028 7474 63084 7486
rect 63028 7422 63030 7474
rect 63082 7422 63084 7474
rect 63028 7420 63084 7422
rect 63028 7354 63084 7364
rect 60340 3210 60396 3220
rect 60676 3331 60844 3387
rect 60900 7308 60956 7318
rect 60228 3098 60284 3108
rect 60116 2986 60172 2996
rect 59892 2650 59948 2660
rect 59668 2538 59724 2548
rect 60116 2492 60172 2502
rect 57988 2090 58044 2100
rect 58660 2268 58716 2278
rect 57876 1978 57932 1988
rect 57428 1708 57484 1718
rect 57428 800 57484 1652
rect 58100 1706 58156 1718
rect 58100 1654 58102 1706
rect 58154 1654 58156 1706
rect 58100 800 58156 1654
rect 58660 800 58716 2212
rect 59668 2154 59724 2166
rect 59668 2102 59670 2154
rect 59722 2102 59724 2154
rect 59220 1260 59276 1270
rect 59220 800 59276 1204
rect 54740 86 54742 138
rect 54794 86 54796 138
rect 54740 74 54796 86
rect 54936 0 55048 800
rect 55608 0 55720 800
rect 56168 0 56280 800
rect 56532 476 56588 486
rect 56532 138 56588 420
rect 56532 86 56534 138
rect 56586 86 56588 138
rect 56532 74 56588 86
rect 56840 0 56952 800
rect 57400 0 57512 800
rect 58072 0 58184 800
rect 58632 0 58744 800
rect 59192 0 59304 800
rect 59668 364 59724 2102
rect 59892 2154 59948 2166
rect 59892 2102 59894 2154
rect 59946 2102 59948 2154
rect 59892 800 59948 2102
rect 60116 1932 60172 2436
rect 60116 1866 60172 1876
rect 60676 1820 60732 3331
rect 60900 3052 60956 7252
rect 62356 7308 62412 7318
rect 62244 6860 62300 6870
rect 62356 6860 62412 7252
rect 62300 6804 62412 6860
rect 62468 7306 62524 7318
rect 62468 7254 62470 7306
rect 62522 7254 62524 7306
rect 62244 6794 62300 6804
rect 61740 6522 61796 6534
rect 61740 6470 61742 6522
rect 61794 6470 61796 6522
rect 61740 6300 61796 6470
rect 61740 6234 61796 6244
rect 62468 6188 62524 7254
rect 62692 6748 62748 6758
rect 62692 6300 62748 6692
rect 62692 6234 62748 6244
rect 62468 6122 62524 6132
rect 63476 5122 63532 5134
rect 63476 5070 63478 5122
rect 63530 5070 63532 5122
rect 60900 2986 60956 2996
rect 62244 5010 62300 5022
rect 62244 4958 62246 5010
rect 62298 4958 62300 5010
rect 61684 2826 61740 2838
rect 61684 2774 61686 2826
rect 61738 2774 61740 2826
rect 60676 1754 60732 1764
rect 61124 1930 61180 1942
rect 61124 1878 61126 1930
rect 61178 1878 61180 1930
rect 60452 1708 60508 1718
rect 60452 800 60508 1652
rect 61124 800 61180 1878
rect 61684 800 61740 2774
rect 61908 2492 61964 2502
rect 61796 2380 61852 2390
rect 61796 2044 61852 2324
rect 61908 2266 61964 2436
rect 62020 2380 62076 2390
rect 62020 2286 62076 2324
rect 61908 2214 61910 2266
rect 61962 2214 61964 2266
rect 61908 2202 61964 2214
rect 62132 2266 62188 2278
rect 62132 2214 62134 2266
rect 62186 2214 62188 2266
rect 62132 2156 62188 2214
rect 62132 2090 62188 2100
rect 61796 1978 61852 1988
rect 62244 1596 62300 4958
rect 63476 4844 63532 5070
rect 63476 4778 63532 4788
rect 62804 4172 62860 4182
rect 62804 3388 62860 4116
rect 62804 3322 62860 3332
rect 63588 3387 63644 8596
rect 63924 7654 63980 11508
rect 63868 7642 63980 7654
rect 63868 7590 63870 7642
rect 63922 7590 63980 7642
rect 63868 7588 63980 7590
rect 64036 11562 64092 11574
rect 64036 11510 64038 11562
rect 64090 11510 64092 11562
rect 63868 7420 63924 7588
rect 63868 7354 63924 7364
rect 63812 6860 63868 6870
rect 64036 6860 64092 11510
rect 64260 8316 64316 13524
rect 64372 11788 64428 14200
rect 64484 14026 64540 14038
rect 64484 13974 64486 14026
rect 64538 13974 64540 14026
rect 64484 12234 64540 13974
rect 64484 12182 64486 12234
rect 64538 12182 64540 12234
rect 64484 12170 64540 12182
rect 65156 12122 65212 14200
rect 65604 14140 65660 14420
rect 65800 14200 65912 15000
rect 66584 14200 66696 15000
rect 67256 14200 67368 15000
rect 67900 14924 67956 14934
rect 67844 14868 67900 14924
rect 67844 14858 67956 14868
rect 67844 14364 67900 14858
rect 67508 14308 67900 14364
rect 65828 14140 65884 14200
rect 65604 14084 65884 14140
rect 65940 14138 65996 14150
rect 65940 14086 65942 14138
rect 65994 14086 65996 14138
rect 65940 13692 65996 14086
rect 65940 13626 65996 13636
rect 66500 13132 66556 13142
rect 66276 13076 66500 13132
rect 65716 12348 65772 12358
rect 65156 12070 65158 12122
rect 65210 12070 65212 12122
rect 65156 12058 65212 12070
rect 65268 12124 65324 12134
rect 64372 11722 64428 11732
rect 65268 10778 65324 12068
rect 65716 11786 65772 12292
rect 65716 11734 65718 11786
rect 65770 11734 65772 11786
rect 65716 11722 65772 11734
rect 66276 11228 66332 13076
rect 66500 13066 66556 13076
rect 66612 12012 66668 14200
rect 67284 14140 67340 14200
rect 67508 14140 67564 14308
rect 68040 14200 68152 15000
rect 68404 14810 68460 14822
rect 68404 14758 68406 14810
rect 68458 14758 68460 14810
rect 67284 14084 67564 14140
rect 66724 13692 66780 13702
rect 66724 12348 66780 13636
rect 68068 13580 68124 14200
rect 68068 13514 68124 13524
rect 68292 13244 68348 13254
rect 67508 13188 67788 13244
rect 67508 13130 67564 13188
rect 67508 13078 67510 13130
rect 67562 13078 67564 13130
rect 67508 13066 67564 13078
rect 66724 12282 66780 12292
rect 66948 12348 67004 12358
rect 66612 11946 66668 11956
rect 66948 11450 67004 12292
rect 67732 12234 67788 13188
rect 68068 13130 68124 13142
rect 68068 13078 68070 13130
rect 68122 13078 68124 13130
rect 67732 12182 67734 12234
rect 67786 12182 67788 12234
rect 67732 12170 67788 12182
rect 67844 13018 67900 13030
rect 67844 12966 67846 13018
rect 67898 12966 67900 13018
rect 67844 12236 67900 12966
rect 68068 12906 68124 13078
rect 68068 12854 68070 12906
rect 68122 12854 68124 12906
rect 68068 12842 68124 12854
rect 67844 12170 67900 12180
rect 66948 11398 66950 11450
rect 67002 11398 67004 11450
rect 66948 11386 67004 11398
rect 67396 12012 67452 12022
rect 66276 11162 66332 11172
rect 66500 11228 66556 11238
rect 65268 10726 65270 10778
rect 65322 10726 65324 10778
rect 65268 10714 65324 10726
rect 65492 10778 65548 10790
rect 65492 10726 65494 10778
rect 65546 10726 65548 10778
rect 64260 8250 64316 8260
rect 64932 8988 64988 8998
rect 64932 8262 64988 8932
rect 65324 8988 65380 8998
rect 65324 8894 65380 8932
rect 64932 8210 64934 8262
rect 64986 8210 64988 8262
rect 64932 8198 64988 8210
rect 63812 6858 64092 6860
rect 63812 6806 63814 6858
rect 63866 6806 64092 6858
rect 63812 6804 64092 6806
rect 63812 6794 63868 6804
rect 64148 6748 64204 6758
rect 64148 6690 64204 6692
rect 64148 6638 64150 6690
rect 64202 6638 64204 6690
rect 64148 6626 64204 6638
rect 63812 5180 63868 5190
rect 63700 3612 63756 3622
rect 63812 3612 63868 5124
rect 64428 4954 64484 4966
rect 64428 4902 64430 4954
rect 64482 4902 64484 4954
rect 64428 4844 64484 4902
rect 64428 4778 64484 4788
rect 65268 4732 65324 4742
rect 64820 4676 65268 4732
rect 64820 4620 64876 4676
rect 65268 4666 65324 4676
rect 64820 4554 64876 4564
rect 65492 4058 65548 10726
rect 66500 10332 66556 11172
rect 67060 10668 67116 10678
rect 67284 10668 67340 10678
rect 67116 10612 67228 10668
rect 67060 10602 67116 10612
rect 66500 10266 66556 10276
rect 67172 9996 67228 10612
rect 67172 9930 67228 9940
rect 66388 9324 66444 9334
rect 65604 8428 65660 8438
rect 65604 5852 65660 8372
rect 65716 8316 65772 8326
rect 65716 8202 65772 8260
rect 65716 8150 65718 8202
rect 65770 8150 65772 8202
rect 65716 8138 65772 8150
rect 66052 8204 66108 8214
rect 66052 8110 66108 8148
rect 66388 7476 66444 9268
rect 67284 8652 67340 10612
rect 66724 8596 67340 8652
rect 66556 8316 66612 8326
rect 66556 8222 66612 8260
rect 66724 7756 66780 8596
rect 66724 7690 66780 7700
rect 66836 8428 66892 8438
rect 66724 7586 66780 7598
rect 66724 7534 66726 7586
rect 66778 7534 66780 7586
rect 66388 7474 66556 7476
rect 66388 7422 66390 7474
rect 66442 7422 66556 7474
rect 66388 7420 66556 7422
rect 66388 7410 66444 7420
rect 66276 7306 66332 7318
rect 66276 7254 66278 7306
rect 66330 7254 66332 7306
rect 66276 6860 66332 7254
rect 66276 6794 66332 6804
rect 66500 6758 66556 7420
rect 66724 6860 66780 7534
rect 66724 6794 66780 6804
rect 65828 6748 65884 6758
rect 66500 6746 66612 6758
rect 66500 6694 66558 6746
rect 66610 6694 66612 6746
rect 66500 6692 66612 6694
rect 65828 6642 65830 6692
rect 65882 6642 65884 6692
rect 66556 6682 66612 6692
rect 65828 6630 65884 6642
rect 65604 5786 65660 5796
rect 66724 6188 66780 6198
rect 65492 4006 65494 4058
rect 65546 4006 65548 4058
rect 65492 3994 65548 4006
rect 66052 5010 66108 5022
rect 66052 4958 66054 5010
rect 66106 4958 66108 5010
rect 65380 3946 65436 3958
rect 65380 3894 65382 3946
rect 65434 3894 65436 3946
rect 63756 3556 63868 3612
rect 63924 3610 63980 3622
rect 63924 3558 63926 3610
rect 63978 3558 63980 3610
rect 63700 3546 63756 3556
rect 63588 3331 63756 3387
rect 62580 2940 62636 2950
rect 62468 2604 62524 2614
rect 62468 1932 62524 2548
rect 62580 2268 62636 2884
rect 62580 2202 62636 2212
rect 62916 2266 62972 2278
rect 62916 2214 62918 2266
rect 62970 2214 62972 2266
rect 62468 1866 62524 1876
rect 62804 1932 62860 1942
rect 62804 1838 62860 1876
rect 62244 1530 62300 1540
rect 62468 1596 62524 1606
rect 62244 1372 62300 1382
rect 62468 1372 62524 1540
rect 62300 1316 62524 1372
rect 62244 1306 62300 1316
rect 62580 1260 62636 1270
rect 62356 1204 62580 1260
rect 62356 800 62412 1204
rect 62580 1194 62636 1204
rect 62916 800 62972 2214
rect 63588 1818 63644 1830
rect 63588 1766 63590 1818
rect 63642 1766 63644 1818
rect 63588 800 63644 1766
rect 63700 922 63756 3331
rect 63700 870 63702 922
rect 63754 870 63756 922
rect 63700 858 63756 870
rect 63924 922 63980 3558
rect 65268 3050 65324 3062
rect 65268 2998 65270 3050
rect 65322 2998 65324 3050
rect 65156 2044 65212 2054
rect 64708 1930 64764 1942
rect 64708 1878 64710 1930
rect 64762 1878 64764 1930
rect 63924 870 63926 922
rect 63978 870 63980 922
rect 63924 858 63980 870
rect 64148 1036 64204 1046
rect 64148 800 64204 980
rect 64708 800 64764 1878
rect 65156 1706 65212 1988
rect 65268 1932 65324 2998
rect 65380 2490 65436 3894
rect 66052 3164 66108 4958
rect 66724 4844 66780 6132
rect 66836 6086 66892 8372
rect 67396 8314 67452 11956
rect 68292 12010 68348 13188
rect 68404 13242 68460 14758
rect 68712 14200 68824 15000
rect 69496 14200 69608 15000
rect 69860 14364 69916 14374
rect 68404 13190 68406 13242
rect 68458 13190 68460 13242
rect 68404 13178 68460 13190
rect 68740 12908 68796 14200
rect 68628 12852 68796 12908
rect 68628 12684 68684 12852
rect 68628 12618 68684 12628
rect 68292 11958 68294 12010
rect 68346 11958 68348 12010
rect 68292 11946 68348 11958
rect 69076 12124 69132 12134
rect 67844 11898 67900 11910
rect 67844 11846 67846 11898
rect 67898 11846 67900 11898
rect 67844 11788 67900 11846
rect 68068 11788 68124 11798
rect 67844 11786 68124 11788
rect 67844 11734 68070 11786
rect 68122 11734 68124 11786
rect 67844 11732 68124 11734
rect 68068 11722 68124 11732
rect 68180 11674 68236 11686
rect 68180 11622 68182 11674
rect 68234 11622 68236 11674
rect 67620 11450 67676 11462
rect 67620 11398 67622 11450
rect 67674 11398 67676 11450
rect 67620 10444 67676 11398
rect 68180 11228 68236 11622
rect 69076 11450 69132 12068
rect 69524 12010 69580 14200
rect 69860 14140 69916 14308
rect 70168 14200 70280 15000
rect 70420 14812 70476 14822
rect 70196 14140 70252 14200
rect 69860 14084 70252 14140
rect 70420 14026 70476 14756
rect 70952 14200 71064 15000
rect 71624 14200 71736 15000
rect 71876 14812 71932 14822
rect 70420 13974 70422 14026
rect 70474 13974 70476 14026
rect 70420 13962 70476 13974
rect 69972 12906 70028 12918
rect 69972 12854 69974 12906
rect 70026 12854 70028 12906
rect 69524 11958 69526 12010
rect 69578 11958 69580 12010
rect 69524 11946 69580 11958
rect 69636 12234 69692 12246
rect 69636 12182 69638 12234
rect 69690 12182 69692 12234
rect 69076 11398 69078 11450
rect 69130 11398 69132 11450
rect 69076 11386 69132 11398
rect 69412 11450 69468 11462
rect 69412 11398 69414 11450
rect 69466 11398 69468 11450
rect 68180 11162 68236 11172
rect 69188 11340 69244 11350
rect 67620 10378 67676 10388
rect 67844 10444 67900 10454
rect 67508 9324 67564 9334
rect 67508 9156 67564 9268
rect 67844 9156 67900 10388
rect 68964 10444 69020 10454
rect 68964 10220 69020 10388
rect 68964 10154 69020 10164
rect 69188 9884 69244 11284
rect 69300 10778 69356 10790
rect 69300 10726 69302 10778
rect 69354 10726 69356 10778
rect 69300 10220 69356 10726
rect 69300 10154 69356 10164
rect 69188 9818 69244 9828
rect 67508 9100 67900 9156
rect 69300 9660 69356 9670
rect 68684 8986 68740 8998
rect 68684 8934 68686 8986
rect 68738 8934 68740 8986
rect 67956 8428 68012 8438
rect 67396 8262 67398 8314
rect 67450 8262 67452 8314
rect 67396 8250 67452 8262
rect 67732 8372 67956 8428
rect 67060 8090 67116 8102
rect 67060 8038 67062 8090
rect 67114 8038 67116 8090
rect 67060 7756 67116 8038
rect 67060 7690 67116 7700
rect 67228 7420 67284 7430
rect 67172 7418 67284 7420
rect 67172 7366 67230 7418
rect 67282 7366 67284 7418
rect 67172 7354 67284 7366
rect 67172 6860 67228 7354
rect 67004 6524 67060 6534
rect 67004 6522 67116 6524
rect 67004 6470 67006 6522
rect 67058 6470 67116 6522
rect 67004 6458 67116 6470
rect 66836 6074 66948 6086
rect 66836 6022 66894 6074
rect 66946 6022 66948 6074
rect 66836 6010 66948 6022
rect 66836 5122 66892 6010
rect 66836 5070 66838 5122
rect 66890 5070 66892 5122
rect 66836 5058 66892 5070
rect 67060 4956 67116 6458
rect 67172 5516 67228 6804
rect 67452 6522 67508 6534
rect 67452 6470 67454 6522
rect 67506 6470 67508 6522
rect 67452 6188 67508 6470
rect 67452 6132 67676 6188
rect 67452 5852 67508 5862
rect 67452 5758 67508 5796
rect 67172 5460 67340 5516
rect 67060 4890 67116 4900
rect 66724 4788 66892 4844
rect 66612 4284 66668 4294
rect 66500 4060 66556 4070
rect 66500 3834 66556 4004
rect 66500 3782 66502 3834
rect 66554 3782 66556 3834
rect 66500 3770 66556 3782
rect 66052 3098 66108 3108
rect 66164 3388 66220 3398
rect 65380 2438 65382 2490
rect 65434 2438 65436 2490
rect 65380 2426 65436 2438
rect 65492 3050 65548 3062
rect 65492 2998 65494 3050
rect 65546 2998 65548 3050
rect 65492 2380 65548 2998
rect 65492 2314 65548 2324
rect 65940 2490 65996 2502
rect 65940 2438 65942 2490
rect 65994 2438 65996 2490
rect 65268 1866 65324 1876
rect 65156 1654 65158 1706
rect 65210 1654 65212 1706
rect 65156 1642 65212 1654
rect 65380 1706 65436 1718
rect 65380 1654 65382 1706
rect 65434 1654 65436 1706
rect 65380 800 65436 1654
rect 65940 800 65996 2438
rect 66164 812 66220 3332
rect 66612 3162 66668 4228
rect 66724 3836 66780 3846
rect 66724 3722 66780 3780
rect 66724 3670 66726 3722
rect 66778 3670 66780 3722
rect 66724 3658 66780 3670
rect 66612 3110 66614 3162
rect 66666 3110 66668 3162
rect 66612 3098 66668 3110
rect 66276 2602 66332 2614
rect 66276 2550 66278 2602
rect 66330 2550 66332 2602
rect 66276 1596 66332 2550
rect 66276 1530 66332 1540
rect 66612 2602 66668 2614
rect 66612 2550 66614 2602
rect 66666 2550 66668 2602
rect 59668 298 59724 308
rect 59864 0 59976 800
rect 60424 0 60536 800
rect 61096 0 61208 800
rect 61656 0 61768 800
rect 62328 0 62440 800
rect 62888 0 63000 800
rect 63560 0 63672 800
rect 64120 0 64232 800
rect 64680 0 64792 800
rect 65352 0 65464 800
rect 65912 0 66024 800
rect 66612 800 66668 2550
rect 66164 746 66220 756
rect 66584 0 66696 800
rect 66836 250 66892 4788
rect 67060 3836 67116 3846
rect 67060 3742 67116 3780
rect 67172 3722 67228 3734
rect 67172 3670 67174 3722
rect 67226 3670 67228 3722
rect 67172 800 67228 3670
rect 67284 3500 67340 5460
rect 67620 4844 67676 6132
rect 67732 6076 67788 8372
rect 67956 8362 68012 8372
rect 68684 8316 68740 8934
rect 68460 8260 69132 8316
rect 68460 8258 68516 8260
rect 68460 8206 68462 8258
rect 68514 8206 68516 8258
rect 68460 8194 68516 8206
rect 67900 8090 67956 8102
rect 67900 8038 67902 8090
rect 67954 8038 67956 8090
rect 67900 7756 67956 8038
rect 67900 7690 67956 7700
rect 68348 8090 68404 8102
rect 68348 8038 68350 8090
rect 68402 8038 68404 8090
rect 68348 7532 68404 8038
rect 68348 7466 68404 7476
rect 68964 7756 69020 7766
rect 68124 7420 68180 7430
rect 68068 7364 68124 7420
rect 68068 7288 68180 7364
rect 68572 7420 68628 7430
rect 68572 7418 68684 7420
rect 68572 7366 68574 7418
rect 68626 7366 68684 7418
rect 68572 7354 68684 7366
rect 67900 6860 67956 6870
rect 67900 6746 67956 6804
rect 67900 6694 67902 6746
rect 67954 6694 67956 6746
rect 67900 6682 67956 6694
rect 67900 6076 67956 6086
rect 67732 6074 67956 6076
rect 67732 6022 67902 6074
rect 67954 6022 67956 6074
rect 67732 6020 67956 6022
rect 67900 6010 67956 6020
rect 68068 5124 68124 7288
rect 68460 6578 68516 6590
rect 68348 6524 68404 6534
rect 68180 6522 68404 6524
rect 68180 6470 68350 6522
rect 68402 6470 68404 6522
rect 68180 6468 68404 6470
rect 68180 5292 68236 6468
rect 68348 6458 68404 6468
rect 68460 6526 68462 6578
rect 68514 6526 68516 6578
rect 68348 6300 68404 6310
rect 68348 6074 68404 6244
rect 68348 6022 68350 6074
rect 68402 6022 68404 6074
rect 68348 6010 68404 6022
rect 68460 5908 68516 6526
rect 68180 5226 68236 5236
rect 68404 5852 68516 5908
rect 68628 5852 68684 7354
rect 68796 6188 68852 6198
rect 68796 6074 68852 6132
rect 68796 6022 68798 6074
rect 68850 6022 68852 6074
rect 68796 6010 68852 6022
rect 68068 5068 68348 5124
rect 67620 4778 67676 4788
rect 67956 4394 68012 4406
rect 67956 4342 67958 4394
rect 68010 4342 68012 4394
rect 67284 3434 67340 3444
rect 67396 4060 67452 4070
rect 67396 2714 67452 4004
rect 67956 3946 68012 4342
rect 67956 3894 67958 3946
rect 68010 3894 68012 3946
rect 67956 3882 68012 3894
rect 67396 2662 67398 2714
rect 67450 2662 67452 2714
rect 67396 2650 67452 2662
rect 68180 2602 68236 2614
rect 68180 2550 68182 2602
rect 68234 2550 68236 2602
rect 67844 2268 67900 2278
rect 67844 800 67900 2212
rect 68180 2042 68236 2550
rect 68292 2156 68348 5068
rect 68404 4956 68460 5852
rect 68628 5796 68796 5852
rect 68404 4284 68460 4900
rect 68572 4954 68628 4966
rect 68572 4902 68574 4954
rect 68626 4902 68628 4954
rect 68572 4506 68628 4902
rect 68572 4454 68574 4506
rect 68626 4454 68628 4506
rect 68572 4442 68628 4454
rect 68404 4228 68572 4284
rect 68404 3612 68460 3622
rect 68404 3518 68460 3556
rect 68292 2090 68348 2100
rect 68404 2828 68460 2838
rect 68180 1990 68182 2042
rect 68234 1990 68236 2042
rect 68180 1978 68236 1990
rect 68404 800 68460 2772
rect 68516 1260 68572 4228
rect 68628 2604 68684 2614
rect 68628 2042 68684 2548
rect 68740 2380 68796 5796
rect 68964 5124 69020 7700
rect 68740 2314 68796 2324
rect 68852 5068 69020 5124
rect 68628 1990 68630 2042
rect 68682 1990 68684 2042
rect 68628 1978 68684 1990
rect 68516 1194 68572 1204
rect 66836 198 66838 250
rect 66890 198 66892 250
rect 66836 186 66892 198
rect 67144 0 67256 800
rect 67816 0 67928 800
rect 68376 0 68488 800
rect 68740 588 68796 598
rect 68740 474 68796 532
rect 68740 422 68742 474
rect 68794 422 68796 474
rect 68740 410 68796 422
rect 68852 250 68908 5068
rect 68964 4956 69020 4966
rect 68964 3274 69020 4900
rect 69076 4508 69132 8260
rect 69300 6870 69356 9604
rect 69412 8204 69468 11398
rect 69412 8138 69468 8148
rect 69524 7756 69580 7766
rect 69524 7308 69580 7700
rect 69524 7242 69580 7252
rect 69300 6858 69412 6870
rect 69300 6806 69358 6858
rect 69410 6806 69412 6858
rect 69300 6804 69412 6806
rect 69356 6794 69412 6804
rect 69468 6580 69524 6590
rect 69468 6578 69580 6580
rect 69468 6526 69470 6578
rect 69522 6526 69580 6578
rect 69468 6514 69580 6526
rect 69356 5908 69412 5918
rect 69356 5906 69468 5908
rect 69356 5854 69358 5906
rect 69410 5854 69468 5906
rect 69356 5852 69468 5854
rect 69356 5842 69412 5852
rect 69244 5740 69300 5750
rect 69244 5646 69300 5684
rect 69076 4442 69132 4452
rect 69188 5010 69244 5022
rect 69188 4958 69190 5010
rect 69242 4958 69244 5010
rect 69188 3612 69244 4958
rect 69188 3546 69244 3556
rect 68964 3222 68966 3274
rect 69018 3222 69020 3274
rect 68964 3210 69020 3222
rect 69412 3274 69468 5796
rect 69524 4844 69580 6514
rect 69636 5852 69692 12182
rect 69860 12236 69916 12246
rect 69860 12142 69916 12180
rect 69972 9324 70028 12854
rect 70980 11900 71036 14200
rect 71652 14026 71708 14200
rect 71652 13974 71654 14026
rect 71706 13974 71708 14026
rect 71652 13962 71708 13974
rect 71764 14140 71820 14150
rect 71764 12682 71820 14084
rect 71876 13916 71932 14756
rect 72408 14200 72520 15000
rect 73080 14200 73192 15000
rect 73332 14922 73388 14934
rect 73332 14870 73334 14922
rect 73386 14870 73388 14922
rect 73332 14698 73388 14870
rect 73332 14646 73334 14698
rect 73386 14646 73388 14698
rect 73332 14634 73388 14646
rect 73556 14698 73612 14710
rect 73556 14646 73558 14698
rect 73610 14646 73612 14698
rect 73556 14250 73612 14646
rect 71876 13850 71932 13860
rect 72436 13132 72492 14200
rect 71764 12630 71766 12682
rect 71818 12630 71820 12682
rect 71764 12618 71820 12630
rect 71876 13076 72492 13132
rect 71764 12124 71820 12134
rect 70980 11834 71036 11844
rect 71204 11900 71260 11910
rect 70980 10668 71036 10678
rect 70980 9894 71036 10612
rect 70924 9884 71036 9894
rect 70756 9882 71036 9884
rect 70756 9830 70926 9882
rect 70978 9830 71036 9882
rect 70756 9828 71036 9830
rect 69972 9258 70028 9268
rect 70196 9324 70252 9334
rect 70196 9210 70252 9268
rect 70196 9158 70198 9210
rect 70250 9158 70252 9210
rect 70196 9146 70252 9158
rect 69860 9098 69916 9110
rect 69860 9046 69862 9098
rect 69914 9046 69916 9098
rect 69860 8988 69916 9046
rect 70588 8988 70644 8998
rect 69860 8986 70644 8988
rect 69860 8934 70590 8986
rect 70642 8934 70644 8986
rect 69860 8932 70644 8934
rect 70588 8876 70644 8932
rect 70588 8810 70644 8820
rect 70196 8652 70252 8662
rect 69748 8428 69804 8438
rect 69748 6300 69804 8372
rect 70196 8426 70252 8596
rect 70196 8374 70198 8426
rect 70250 8374 70252 8426
rect 70196 8362 70252 8374
rect 70756 8258 70812 9828
rect 70924 9818 70980 9828
rect 71204 9324 71260 11844
rect 71204 9258 71260 9268
rect 71316 10778 71372 10790
rect 71316 10726 71318 10778
rect 71370 10726 71372 10778
rect 71316 9110 71372 10726
rect 71260 9100 71372 9110
rect 70644 8204 70700 8214
rect 70756 8206 70758 8258
rect 70810 8206 70812 8258
rect 70756 8194 70812 8206
rect 71204 9098 71372 9100
rect 71204 9046 71262 9098
rect 71314 9046 71372 9098
rect 71204 9044 71372 9046
rect 71204 9034 71316 9044
rect 71204 8204 71260 9034
rect 71764 8426 71820 12068
rect 71876 11450 71932 13076
rect 71876 11398 71878 11450
rect 71930 11398 71932 11450
rect 71876 11386 71932 11398
rect 71988 12682 72044 12694
rect 71988 12630 71990 12682
rect 72042 12630 72044 12682
rect 71764 8374 71766 8426
rect 71818 8374 71820 8426
rect 71764 8362 71820 8374
rect 71988 8998 72044 12630
rect 73108 12012 73164 14200
rect 73556 14198 73558 14250
rect 73610 14198 73612 14250
rect 73864 14200 73976 15000
rect 74536 14200 74648 15000
rect 74788 14644 75180 14700
rect 73556 14186 73612 14198
rect 73892 14140 73948 14200
rect 74004 14140 74060 14150
rect 73892 14138 74060 14140
rect 73892 14086 74006 14138
rect 74058 14086 74060 14138
rect 73892 14084 74060 14086
rect 74004 14074 74060 14084
rect 74004 13468 74060 13478
rect 74004 13244 74060 13412
rect 74004 13178 74060 13188
rect 74228 13468 74284 13478
rect 74228 13132 74284 13412
rect 74228 13066 74284 13076
rect 74452 13132 74508 13142
rect 73780 13020 73836 13030
rect 73780 13018 74060 13020
rect 73780 12966 73782 13018
rect 73834 12966 74060 13018
rect 73780 12964 74060 12966
rect 73780 12954 73836 12964
rect 73556 12908 73612 12918
rect 73556 12684 73612 12852
rect 74004 12906 74060 12964
rect 74452 13018 74508 13076
rect 74452 12966 74454 13018
rect 74506 12966 74508 13018
rect 74452 12954 74508 12966
rect 74004 12854 74006 12906
rect 74058 12854 74060 12906
rect 74004 12842 74060 12854
rect 73556 12618 73612 12628
rect 73108 11946 73164 11956
rect 74116 12124 74172 12134
rect 73220 11898 73276 11910
rect 73220 11846 73222 11898
rect 73274 11846 73276 11898
rect 72100 11450 72156 11462
rect 72100 11398 72102 11450
rect 72154 11398 72156 11450
rect 72100 9996 72156 11398
rect 72100 9930 72156 9940
rect 72660 11228 72716 11238
rect 72660 9884 72716 11172
rect 72660 9818 72716 9828
rect 72772 9772 72828 9782
rect 71988 8986 72100 8998
rect 71988 8934 72046 8986
rect 72098 8934 72100 8986
rect 71988 8922 72100 8934
rect 70644 8146 70700 8148
rect 70644 8094 70646 8146
rect 70698 8094 70700 8146
rect 71204 8138 71260 8148
rect 71428 8204 71484 8214
rect 71428 8110 71484 8148
rect 71988 8204 72044 8922
rect 72772 8540 72828 9716
rect 73220 9660 73276 11846
rect 74116 11898 74172 12068
rect 74116 11846 74118 11898
rect 74170 11846 74172 11898
rect 74116 11834 74172 11846
rect 74340 12124 74396 12134
rect 73556 11786 73612 11798
rect 73556 11734 73558 11786
rect 73610 11734 73612 11786
rect 73444 11228 73500 11238
rect 73444 10778 73500 11172
rect 73444 10726 73446 10778
rect 73498 10726 73500 10778
rect 73444 10714 73500 10726
rect 73220 9594 73276 9604
rect 73276 8988 73332 8998
rect 73276 8986 73388 8988
rect 73276 8934 73278 8986
rect 73330 8934 73388 8986
rect 73276 8922 73388 8934
rect 72772 8474 72828 8484
rect 71988 8138 72044 8148
rect 72100 8428 72156 8438
rect 70644 8082 70700 8094
rect 71764 7644 71820 7654
rect 70868 7474 70924 7486
rect 70868 7422 70870 7474
rect 70922 7422 70924 7474
rect 70868 7420 70924 7422
rect 70868 7354 70924 7364
rect 71428 7420 71484 7430
rect 70532 7306 70588 7318
rect 70532 7254 70534 7306
rect 70586 7254 70588 7306
rect 69860 7196 69916 7206
rect 69860 6748 69916 7140
rect 70532 6972 70588 7254
rect 70532 6906 70588 6916
rect 70140 6860 70196 6870
rect 70028 6748 70084 6758
rect 69860 6746 70084 6748
rect 69860 6694 70030 6746
rect 70082 6694 70084 6746
rect 69860 6692 70084 6694
rect 70028 6682 70084 6692
rect 70140 6690 70196 6804
rect 70140 6638 70142 6690
rect 70194 6638 70196 6690
rect 70140 6626 70196 6638
rect 70588 6412 70644 6422
rect 69748 6244 70084 6300
rect 70028 6020 70084 6244
rect 70588 6074 70644 6356
rect 70588 6022 70590 6074
rect 70642 6022 70644 6074
rect 70028 6018 70364 6020
rect 69916 5964 69972 5974
rect 70028 5966 70030 6018
rect 70082 5966 70364 6018
rect 70588 6010 70644 6022
rect 70700 6300 70756 6310
rect 70028 5964 70364 5966
rect 70028 5954 70084 5964
rect 69916 5870 69972 5908
rect 69636 5786 69692 5796
rect 70308 5852 70364 5964
rect 70700 5908 70756 6244
rect 71428 6188 71484 7364
rect 71428 6030 71484 6132
rect 71372 6018 71484 6030
rect 71372 5966 71374 6018
rect 71426 5966 71484 6018
rect 71372 5964 71484 5966
rect 71372 5954 71428 5964
rect 70700 5906 70812 5908
rect 70700 5854 70702 5906
rect 70754 5854 70812 5906
rect 70700 5842 70812 5854
rect 70308 5786 70364 5796
rect 69524 3948 69580 4788
rect 70420 5122 70476 5134
rect 70420 5070 70422 5122
rect 70474 5070 70476 5122
rect 70420 4506 70476 5070
rect 70420 4454 70422 4506
rect 70474 4454 70476 4506
rect 69636 3948 69692 3958
rect 69524 3892 69636 3948
rect 69636 3882 69692 3892
rect 69412 3222 69414 3274
rect 69466 3222 69468 3274
rect 69412 3210 69468 3222
rect 70196 3276 70252 3286
rect 69076 2604 69132 2614
rect 69076 1820 69132 2548
rect 69076 1754 69132 1764
rect 69636 2156 69692 2166
rect 68964 1036 69020 1046
rect 68964 922 69020 980
rect 68964 870 68966 922
rect 69018 870 69020 922
rect 68964 858 69020 870
rect 69076 868 69356 924
rect 69076 800 69132 868
rect 68852 198 68854 250
rect 68906 198 68908 250
rect 68852 186 68908 198
rect 69048 0 69160 800
rect 69300 474 69356 868
rect 69636 800 69692 2100
rect 69972 1258 70028 1270
rect 69972 1206 69974 1258
rect 70026 1206 70028 1258
rect 69972 810 70028 1206
rect 69300 422 69302 474
rect 69354 422 69356 474
rect 69300 410 69356 422
rect 69608 0 69720 800
rect 69972 758 69974 810
rect 70026 758 70028 810
rect 70196 800 70252 3220
rect 70308 2716 70364 2726
rect 70308 2378 70364 2660
rect 70308 2326 70310 2378
rect 70362 2326 70364 2378
rect 70308 2314 70364 2326
rect 69972 746 70028 758
rect 70168 0 70280 800
rect 70420 698 70476 4454
rect 70644 4394 70700 4406
rect 70644 4342 70646 4394
rect 70698 4342 70700 4394
rect 70644 3387 70700 4342
rect 70756 4060 70812 5842
rect 71260 5738 71316 5750
rect 71260 5686 71262 5738
rect 71314 5686 71316 5738
rect 71260 5078 71316 5686
rect 71764 5292 71820 7588
rect 72100 6412 72156 8372
rect 72380 8092 72436 8102
rect 72324 8090 72436 8092
rect 72324 8038 72382 8090
rect 72434 8038 72436 8090
rect 72324 8026 72436 8038
rect 72212 7980 72268 7990
rect 72212 6858 72268 7924
rect 72212 6806 72214 6858
rect 72266 6806 72268 6858
rect 72212 6794 72268 6806
rect 72324 7196 72380 8026
rect 72548 7476 72604 7486
rect 73332 7476 73388 8922
rect 72548 7474 73388 7476
rect 72548 7422 72550 7474
rect 72602 7422 73388 7474
rect 72548 7420 73388 7422
rect 72548 7410 72604 7420
rect 72100 6346 72156 6356
rect 71932 6076 71988 6086
rect 71932 5982 71988 6020
rect 72044 5908 72100 5918
rect 72044 5906 72156 5908
rect 72044 5854 72046 5906
rect 72098 5854 72156 5906
rect 72044 5842 72156 5854
rect 71764 5226 71820 5236
rect 71204 5068 71316 5078
rect 71260 5012 71316 5068
rect 71204 5002 71260 5012
rect 70868 4956 70924 4966
rect 70868 4394 70924 4900
rect 71596 4954 71652 4966
rect 71596 4902 71598 4954
rect 71650 4902 71652 4954
rect 71596 4506 71652 4902
rect 71596 4454 71598 4506
rect 71650 4454 71652 4506
rect 71596 4442 71652 4454
rect 72100 4506 72156 5842
rect 72100 4454 72102 4506
rect 72154 4454 72156 4506
rect 72100 4442 72156 4454
rect 70868 4342 70870 4394
rect 70922 4342 70924 4394
rect 70868 4330 70924 4342
rect 70756 3994 70812 4004
rect 72100 4284 72156 4294
rect 71876 3388 71932 3398
rect 70644 3331 70812 3387
rect 70532 3164 70588 3174
rect 70532 2378 70588 3108
rect 70756 3164 70812 3331
rect 70756 3098 70812 3108
rect 70532 2326 70534 2378
rect 70586 2326 70588 2378
rect 70532 2314 70588 2326
rect 70868 1820 70924 1830
rect 70532 1484 70588 1494
rect 70532 1258 70588 1428
rect 70532 1206 70534 1258
rect 70586 1206 70588 1258
rect 70532 1194 70588 1206
rect 70868 800 70924 1764
rect 71428 922 71484 934
rect 71428 870 71430 922
rect 71482 870 71484 922
rect 71428 800 71484 870
rect 70420 646 70422 698
rect 70474 646 70476 698
rect 70420 634 70476 646
rect 70840 0 70952 800
rect 71400 0 71512 800
rect 71876 252 71932 3332
rect 71988 1484 72044 1494
rect 71988 1146 72044 1428
rect 71988 1094 71990 1146
rect 72042 1094 72044 1146
rect 71988 1082 72044 1094
rect 72100 800 72156 4228
rect 72324 2940 72380 7140
rect 72548 6692 72604 6702
rect 72324 2874 72380 2884
rect 72436 6690 72604 6692
rect 72436 6638 72550 6690
rect 72602 6638 72604 6690
rect 72436 6636 72604 6638
rect 72436 2380 72492 6636
rect 72548 6626 72604 6636
rect 73332 6076 73388 7420
rect 73332 6010 73388 6020
rect 73388 5908 73444 5918
rect 72604 5906 73500 5908
rect 72604 5854 73390 5906
rect 73442 5854 73500 5906
rect 72604 5852 73500 5854
rect 72604 5850 72660 5852
rect 72604 5798 72606 5850
rect 72658 5798 72660 5850
rect 73388 5842 73500 5852
rect 72604 5786 72660 5798
rect 73276 5738 73332 5750
rect 73276 5686 73278 5738
rect 73330 5686 73332 5738
rect 73276 5628 73332 5686
rect 73276 5562 73332 5572
rect 72548 5292 72604 5302
rect 72548 5234 72604 5236
rect 72548 5182 72550 5234
rect 72602 5182 72604 5234
rect 72548 5170 72604 5182
rect 72436 2314 72492 2324
rect 72548 4844 72604 4854
rect 72548 1372 72604 4788
rect 73332 4060 73388 4070
rect 73220 3724 73276 3734
rect 72884 3668 73220 3724
rect 72772 3612 72828 3622
rect 72772 3388 72828 3556
rect 72884 3500 72940 3668
rect 73220 3658 73276 3668
rect 72884 3434 72940 3444
rect 72772 3322 72828 3332
rect 72884 3276 72940 3286
rect 72940 3220 73164 3276
rect 72884 3210 72940 3220
rect 73108 2492 73164 3220
rect 73108 2426 73164 2436
rect 72548 1306 72604 1316
rect 72660 2380 72716 2390
rect 72660 800 72716 2324
rect 73332 800 73388 4004
rect 73444 2940 73500 5842
rect 73556 4060 73612 11734
rect 73892 11228 73948 11238
rect 73780 10778 73836 10790
rect 73780 10726 73782 10778
rect 73834 10726 73836 10778
rect 73668 9212 73724 9222
rect 73668 4956 73724 9156
rect 73780 8314 73836 10726
rect 73780 8262 73782 8314
rect 73834 8262 73836 8314
rect 73780 8250 73836 8262
rect 73892 7532 73948 11172
rect 74116 9212 74172 9222
rect 74116 9118 74172 9156
rect 73892 7466 73948 7476
rect 74116 7644 74172 7654
rect 74116 7308 74172 7588
rect 74228 7308 74284 7318
rect 74116 7306 74284 7308
rect 74116 7254 74230 7306
rect 74282 7254 74284 7306
rect 74116 7252 74284 7254
rect 74228 7242 74284 7252
rect 74228 6690 74284 6702
rect 74228 6638 74230 6690
rect 74282 6638 74284 6690
rect 74228 6086 74284 6638
rect 74340 6636 74396 12068
rect 74564 11900 74620 14200
rect 74676 14026 74732 14038
rect 74676 13974 74678 14026
rect 74730 13974 74732 14026
rect 74676 13916 74732 13974
rect 74676 13850 74732 13860
rect 74788 12012 74844 14644
rect 74900 14474 74956 14486
rect 74900 14422 74902 14474
rect 74954 14422 74956 14474
rect 74900 13916 74956 14422
rect 75124 14140 75180 14644
rect 75320 14200 75432 15000
rect 75572 14474 75628 14486
rect 75572 14422 75574 14474
rect 75626 14422 75628 14474
rect 75348 14140 75404 14200
rect 75124 14084 75404 14140
rect 75572 14138 75628 14422
rect 75992 14200 76104 15000
rect 76776 14200 76888 15000
rect 77448 14200 77560 15000
rect 77700 14588 77756 14598
rect 77756 14532 77980 14588
rect 77700 14522 77756 14532
rect 75572 14086 75574 14138
rect 75626 14086 75628 14138
rect 75572 14074 75628 14086
rect 74900 13850 74956 13860
rect 75012 14026 75068 14038
rect 75012 13974 75014 14026
rect 75066 13974 75068 14026
rect 75012 12908 75068 13974
rect 75124 13914 75180 13926
rect 75124 13862 75126 13914
rect 75178 13862 75180 13914
rect 75124 13018 75180 13862
rect 75460 13804 75516 13814
rect 75684 13804 75740 13814
rect 75460 13802 75740 13804
rect 75460 13750 75462 13802
rect 75514 13750 75686 13802
rect 75738 13750 75740 13802
rect 75460 13748 75740 13750
rect 75460 13738 75516 13748
rect 75684 13738 75740 13748
rect 75796 13690 75852 13702
rect 75796 13638 75798 13690
rect 75850 13638 75852 13690
rect 75796 13466 75852 13638
rect 75796 13414 75798 13466
rect 75850 13414 75852 13466
rect 75796 13402 75852 13414
rect 76020 13466 76076 14200
rect 76804 14028 76860 14200
rect 76020 13414 76022 13466
rect 76074 13414 76076 13466
rect 76020 13402 76076 13414
rect 76468 13972 76860 14028
rect 76916 14138 76972 14150
rect 76916 14086 76918 14138
rect 76970 14086 76972 14138
rect 75124 12966 75126 13018
rect 75178 12966 75180 13018
rect 75124 12954 75180 12966
rect 75012 12842 75068 12852
rect 74788 11946 74844 11956
rect 75236 12346 75292 12358
rect 75236 12294 75238 12346
rect 75290 12294 75292 12346
rect 74564 11834 74620 11844
rect 74676 11898 74732 11910
rect 74676 11846 74678 11898
rect 74730 11846 74732 11898
rect 74452 11788 74508 11798
rect 74452 9210 74508 11732
rect 74452 9158 74454 9210
rect 74506 9158 74508 9210
rect 74452 9146 74508 9158
rect 74676 8428 74732 11846
rect 75236 10108 75292 12294
rect 76468 12236 76524 13972
rect 76916 13804 76972 14086
rect 77252 14140 77308 14150
rect 77252 13916 77308 14084
rect 77364 14140 77420 14150
rect 77476 14140 77532 14200
rect 77364 14138 77532 14140
rect 77364 14086 77366 14138
rect 77418 14086 77532 14138
rect 77364 14084 77532 14086
rect 77588 14138 77644 14150
rect 77588 14086 77590 14138
rect 77642 14086 77644 14138
rect 77364 14074 77420 14084
rect 77588 13916 77644 14086
rect 77252 13860 77644 13916
rect 77924 13916 77980 14532
rect 78232 14200 78344 15000
rect 78708 14698 78764 14710
rect 78708 14646 78710 14698
rect 78762 14646 78764 14698
rect 78036 14140 78092 14150
rect 78036 14046 78092 14084
rect 78260 13916 78316 14200
rect 77924 13860 78316 13916
rect 78372 14138 78428 14150
rect 78372 14086 78374 14138
rect 78426 14086 78428 14138
rect 77140 13804 77196 13814
rect 76916 13738 76972 13748
rect 77028 13748 77140 13804
rect 76916 13468 76972 13478
rect 76804 12682 76860 12694
rect 76804 12630 76806 12682
rect 76858 12630 76860 12682
rect 76468 12180 76636 12236
rect 76580 11788 76636 12180
rect 76580 11722 76636 11732
rect 76692 12234 76748 12246
rect 76692 12182 76694 12234
rect 76746 12182 76748 12234
rect 75236 10042 75292 10052
rect 76580 9996 76636 10006
rect 76692 9996 76748 12182
rect 76804 10332 76860 12630
rect 76916 11564 76972 13412
rect 77028 12908 77084 13748
rect 77140 13738 77196 13748
rect 77140 13468 77196 13478
rect 77140 13132 77196 13412
rect 77252 13244 77308 13254
rect 77308 13188 77532 13244
rect 77252 13178 77308 13188
rect 77476 13132 77532 13188
rect 77476 13076 77980 13132
rect 77140 13066 77196 13076
rect 77028 12842 77084 12852
rect 77364 13020 77420 13030
rect 77364 12906 77420 12964
rect 77364 12854 77366 12906
rect 77418 12854 77420 12906
rect 77364 12842 77420 12854
rect 77812 12906 77868 12918
rect 77812 12854 77814 12906
rect 77866 12854 77868 12906
rect 77812 12236 77868 12854
rect 77924 12796 77980 13076
rect 78036 12796 78092 12806
rect 77924 12740 78036 12796
rect 78036 12730 78092 12740
rect 77924 12460 77980 12470
rect 77924 12366 77980 12404
rect 78260 12348 78316 12358
rect 78260 12254 78316 12292
rect 77812 12180 78092 12236
rect 77812 12010 77868 12022
rect 77812 11958 77814 12010
rect 77866 11958 77868 12010
rect 77588 11900 77644 11910
rect 77812 11900 77868 11958
rect 77588 11898 77868 11900
rect 77588 11846 77590 11898
rect 77642 11846 77868 11898
rect 77588 11844 77868 11846
rect 77588 11834 77644 11844
rect 76916 11508 77756 11564
rect 77252 10780 77308 10790
rect 77700 10780 77756 11508
rect 78036 11004 78092 12180
rect 78372 12234 78428 14086
rect 78484 14028 78540 14038
rect 78708 14028 78764 14646
rect 78904 14200 79016 15000
rect 79156 14868 79436 14924
rect 79156 14700 79212 14868
rect 79156 14634 79212 14644
rect 79268 14698 79324 14710
rect 79268 14646 79270 14698
rect 79322 14646 79324 14698
rect 79268 14364 79324 14646
rect 79380 14474 79436 14868
rect 79492 14922 79548 14934
rect 79492 14870 79494 14922
rect 79546 14870 79548 14922
rect 79492 14586 79548 14870
rect 79492 14534 79494 14586
rect 79546 14534 79548 14586
rect 79492 14522 79548 14534
rect 79380 14422 79382 14474
rect 79434 14422 79436 14474
rect 79380 14410 79436 14422
rect 79156 14308 79324 14364
rect 78820 14140 78876 14150
rect 78932 14140 78988 14200
rect 78820 14138 78988 14140
rect 78820 14086 78822 14138
rect 78874 14086 78988 14138
rect 78820 14084 78988 14086
rect 79044 14138 79100 14150
rect 79044 14086 79046 14138
rect 79098 14086 79100 14138
rect 78820 14074 78876 14084
rect 78540 13972 78652 14028
rect 78484 13962 78540 13972
rect 78372 12182 78374 12234
rect 78426 12182 78428 12234
rect 78372 12170 78428 12182
rect 78484 13132 78540 13142
rect 78484 12012 78540 13076
rect 78596 12346 78652 13972
rect 78708 13962 78764 13972
rect 79044 13580 79100 14086
rect 79156 14028 79212 14308
rect 79688 14200 79800 15000
rect 79940 14700 79996 14710
rect 80164 14700 80220 14710
rect 79940 14698 80220 14700
rect 79940 14646 79942 14698
rect 79994 14646 80166 14698
rect 80218 14646 80220 14698
rect 79940 14644 80220 14646
rect 79940 14634 79996 14644
rect 80164 14634 80220 14644
rect 80360 14200 80472 15000
rect 80724 14922 80780 14934
rect 80724 14870 80726 14922
rect 80778 14870 80780 14922
rect 80724 14698 80780 14870
rect 80948 14700 81004 14710
rect 80724 14646 80726 14698
rect 80778 14646 80780 14698
rect 80724 14634 80780 14646
rect 80836 14698 81004 14700
rect 80836 14646 80950 14698
rect 81002 14646 81004 14698
rect 80836 14644 81004 14646
rect 80724 14252 80780 14262
rect 80836 14252 80892 14644
rect 80948 14634 81004 14644
rect 80724 14250 80892 14252
rect 79716 14140 79772 14200
rect 79156 13962 79212 13972
rect 79380 14084 79772 14140
rect 78708 13524 79100 13580
rect 78708 13018 78764 13524
rect 78708 12966 78710 13018
rect 78762 12966 78764 13018
rect 78708 12954 78764 12966
rect 78820 13412 79212 13468
rect 78708 12682 78764 12694
rect 78708 12630 78710 12682
rect 78762 12630 78764 12682
rect 78708 12460 78764 12630
rect 78708 12394 78764 12404
rect 78596 12294 78598 12346
rect 78650 12294 78652 12346
rect 78596 12282 78652 12294
rect 78820 12348 78876 13412
rect 79156 13356 79212 13412
rect 79156 13300 79324 13356
rect 79044 13242 79100 13254
rect 79044 13190 79046 13242
rect 79098 13190 79100 13242
rect 78932 13018 78988 13030
rect 78932 12966 78934 13018
rect 78986 12966 78988 13018
rect 78932 12684 78988 12966
rect 79044 12796 79100 13190
rect 79268 13020 79324 13300
rect 79268 12954 79324 12964
rect 79044 12740 79324 12796
rect 78932 12628 79100 12684
rect 78820 12282 78876 12292
rect 78932 12460 78988 12470
rect 78260 11956 78540 12012
rect 78036 10938 78092 10948
rect 78148 11116 78204 11126
rect 78148 10780 78204 11060
rect 77700 10724 78204 10780
rect 76804 10276 77084 10332
rect 76580 9994 76748 9996
rect 76580 9942 76582 9994
rect 76634 9942 76748 9994
rect 76580 9940 76748 9942
rect 76804 10108 76860 10118
rect 76580 9930 76636 9940
rect 76804 9828 76860 10052
rect 76020 9772 76860 9828
rect 76020 9660 76076 9772
rect 76020 9594 76076 9604
rect 76244 9658 76300 9670
rect 76244 9606 76246 9658
rect 76298 9606 76300 9658
rect 74844 9212 74900 9222
rect 76244 9212 76300 9606
rect 76748 9212 76804 9222
rect 76244 9210 76804 9212
rect 76244 9158 76750 9210
rect 76802 9158 76804 9210
rect 76244 9156 76804 9158
rect 74844 8988 74900 9156
rect 74844 8986 74956 8988
rect 74844 8934 74846 8986
rect 74898 8934 74956 8986
rect 74844 8922 74956 8934
rect 74676 8362 74732 8372
rect 74900 8316 74956 8922
rect 74788 8258 74844 8270
rect 74788 8206 74790 8258
rect 74842 8206 74844 8258
rect 74900 8250 74956 8260
rect 76468 8258 76524 8270
rect 74676 7586 74732 7598
rect 74676 7534 74678 7586
rect 74730 7534 74732 7586
rect 74564 7474 74620 7486
rect 74564 7422 74566 7474
rect 74618 7422 74620 7474
rect 74564 7308 74620 7422
rect 74676 7420 74732 7534
rect 74676 7354 74732 7364
rect 74564 7242 74620 7252
rect 74788 7196 74844 8206
rect 76468 8206 76470 8258
rect 76522 8206 76524 8258
rect 75012 7420 75068 7430
rect 75180 7420 75236 7430
rect 75068 7418 75236 7420
rect 75068 7366 75182 7418
rect 75234 7366 75236 7418
rect 75068 7364 75236 7366
rect 75012 7354 75068 7364
rect 74788 7130 74844 7140
rect 75068 6860 75124 6870
rect 75180 6860 75236 7364
rect 75628 7418 75684 7430
rect 75628 7366 75630 7418
rect 75682 7366 75684 7418
rect 75628 7308 75684 7366
rect 75628 6972 75684 7252
rect 75628 6906 75684 6916
rect 76076 7420 76132 7430
rect 76076 6870 76132 7364
rect 76020 6860 76132 6870
rect 75180 6804 75404 6860
rect 75068 6690 75124 6804
rect 75068 6638 75070 6690
rect 75122 6638 75124 6690
rect 74340 6580 74452 6636
rect 75068 6626 75124 6638
rect 75180 6636 75236 6646
rect 74228 6074 74340 6086
rect 74228 6022 74286 6074
rect 74338 6022 74340 6074
rect 74228 6020 74340 6022
rect 74284 6010 74340 6020
rect 74396 6020 74452 6580
rect 75180 6542 75236 6580
rect 74396 6018 74620 6020
rect 74396 5966 74398 6018
rect 74450 5966 74620 6018
rect 74396 5964 74620 5966
rect 74396 5954 74452 5964
rect 74564 5190 74620 5964
rect 75348 5852 75404 6804
rect 76076 6804 76132 6860
rect 76300 7196 76356 7206
rect 76020 6794 76076 6804
rect 76300 6748 76356 7140
rect 76132 6746 76356 6748
rect 75852 6696 75908 6702
rect 76132 6696 76302 6746
rect 75852 6694 76302 6696
rect 76354 6694 76356 6746
rect 75852 6692 76356 6694
rect 75852 6690 76188 6692
rect 75852 6638 75854 6690
rect 75906 6640 76188 6690
rect 76300 6682 76356 6692
rect 75906 6638 75908 6640
rect 75852 6626 75908 6638
rect 75740 6524 75796 6534
rect 75740 6430 75796 6468
rect 76020 6412 76076 6422
rect 75572 6300 75628 6310
rect 75572 6018 75628 6244
rect 75572 5966 75574 6018
rect 75626 5966 75628 6018
rect 75572 5954 75628 5966
rect 75348 5796 75852 5852
rect 75572 5628 75628 5638
rect 75180 5516 75236 5526
rect 74564 5178 74676 5190
rect 73892 5122 73948 5134
rect 74564 5126 74622 5178
rect 74674 5126 74676 5178
rect 74564 5124 74676 5126
rect 73892 5070 73894 5122
rect 73946 5070 73948 5122
rect 74620 5114 74676 5124
rect 75180 5178 75236 5460
rect 75180 5126 75182 5178
rect 75234 5126 75236 5178
rect 73892 5068 73948 5070
rect 73892 5002 73948 5012
rect 75180 5068 75236 5126
rect 75180 5002 75236 5012
rect 73668 4890 73724 4900
rect 73556 3994 73612 4004
rect 74004 4844 74060 4854
rect 74004 4060 74060 4788
rect 74116 4620 74172 4630
rect 74172 4564 74508 4620
rect 74116 4554 74172 4564
rect 74452 4284 74508 4564
rect 74452 4218 74508 4228
rect 74004 3994 74060 4004
rect 75572 4058 75628 5572
rect 75572 4006 75574 4058
rect 75626 4006 75628 4058
rect 75572 3994 75628 4006
rect 75684 4506 75740 4518
rect 75684 4454 75686 4506
rect 75738 4454 75740 4506
rect 75348 3946 75404 3958
rect 75348 3894 75350 3946
rect 75402 3894 75404 3946
rect 74676 3836 74732 3846
rect 73444 2874 73500 2884
rect 73668 3388 73724 3398
rect 74676 3388 74732 3780
rect 75348 3836 75404 3894
rect 75348 3770 75404 3780
rect 75012 3612 75068 3622
rect 74676 3332 74956 3388
rect 73556 2716 73612 2726
rect 73444 2378 73500 2390
rect 73444 2326 73446 2378
rect 73498 2326 73500 2378
rect 73444 2156 73500 2326
rect 73444 2090 73500 2100
rect 71876 186 71932 196
rect 72072 0 72184 800
rect 72632 0 72744 800
rect 73304 0 73416 800
rect 73556 362 73612 2660
rect 73668 2492 73724 3332
rect 73668 2426 73724 2436
rect 74004 2268 74060 2278
rect 73892 2266 74060 2268
rect 73892 2214 74006 2266
rect 74058 2214 74060 2266
rect 73892 2212 74060 2214
rect 73892 800 73948 2212
rect 74004 2202 74060 2212
rect 74564 1932 74620 1942
rect 74564 800 74620 1876
rect 74788 1482 74844 1494
rect 74788 1430 74790 1482
rect 74842 1430 74844 1482
rect 73556 310 73558 362
rect 73610 310 73612 362
rect 73556 298 73612 310
rect 73864 0 73976 800
rect 74536 0 74648 800
rect 74788 700 74844 1430
rect 74900 1260 74956 3332
rect 75012 3052 75068 3556
rect 75348 3276 75404 3286
rect 75012 2986 75068 2996
rect 75124 3220 75348 3276
rect 75124 2266 75180 3220
rect 75348 3210 75404 3220
rect 75684 2828 75740 4454
rect 75796 3276 75852 5796
rect 75908 4506 75964 4518
rect 75908 4454 75910 4506
rect 75962 4454 75964 4506
rect 75908 4284 75964 4454
rect 75908 4218 75964 4228
rect 75796 3210 75852 3220
rect 75684 2762 75740 2772
rect 75908 2604 75964 2614
rect 75684 2548 75908 2604
rect 75124 2214 75126 2266
rect 75178 2214 75180 2266
rect 75124 2202 75180 2214
rect 75236 2268 75292 2278
rect 75292 2212 75628 2268
rect 75236 2202 75292 2212
rect 75012 2156 75068 2166
rect 75012 2044 75068 2100
rect 75012 1988 75292 2044
rect 74900 1194 74956 1204
rect 75124 1146 75180 1158
rect 75124 1094 75126 1146
rect 75178 1094 75180 1146
rect 74788 634 74844 644
rect 74900 1034 74956 1046
rect 74900 982 74902 1034
rect 74954 982 74956 1034
rect 74900 362 74956 982
rect 75124 800 75180 1094
rect 75236 1034 75292 1988
rect 75460 1932 75516 1942
rect 75460 1594 75516 1876
rect 75460 1542 75462 1594
rect 75514 1542 75516 1594
rect 75460 1530 75516 1542
rect 75572 1482 75628 2212
rect 75572 1430 75574 1482
rect 75626 1430 75628 1482
rect 75572 1418 75628 1430
rect 75236 982 75238 1034
rect 75290 982 75292 1034
rect 75236 970 75292 982
rect 75348 1372 75404 1382
rect 75348 812 75404 1316
rect 74900 310 74902 362
rect 74954 310 74956 362
rect 74900 298 74956 310
rect 75096 0 75208 800
rect 75684 800 75740 2548
rect 75908 2538 75964 2548
rect 75908 2266 75964 2278
rect 75908 2214 75910 2266
rect 75962 2214 75964 2266
rect 75908 2042 75964 2214
rect 75908 1990 75910 2042
rect 75962 1990 75964 2042
rect 75908 1978 75964 1990
rect 76020 1036 76076 6356
rect 76468 6076 76524 8206
rect 76580 6747 76636 9156
rect 76748 9146 76804 9156
rect 76804 8316 76860 8326
rect 76580 6691 76748 6747
rect 76468 6010 76524 6020
rect 76692 4620 76748 6691
rect 76692 4554 76748 4564
rect 76468 4396 76524 4406
rect 76244 2378 76300 2390
rect 76244 2326 76246 2378
rect 76298 2326 76300 2378
rect 76244 2156 76300 2326
rect 76468 2378 76524 4340
rect 76468 2326 76470 2378
rect 76522 2326 76524 2378
rect 76468 2314 76524 2326
rect 76692 3052 76748 3062
rect 76356 2156 76412 2166
rect 76244 2154 76412 2156
rect 76244 2102 76358 2154
rect 76410 2102 76412 2154
rect 76244 2100 76412 2102
rect 76356 2090 76412 2100
rect 76468 2044 76524 2054
rect 76468 1820 76524 1988
rect 76692 2044 76748 2996
rect 76692 1978 76748 1988
rect 76468 1764 76636 1820
rect 76468 1484 76524 1494
rect 76020 970 76076 980
rect 76356 1428 76468 1484
rect 76244 924 76300 934
rect 76132 868 76244 924
rect 76132 810 76188 868
rect 76244 858 76300 868
rect 75348 746 75404 756
rect 75656 0 75768 800
rect 76132 758 76134 810
rect 76186 758 76188 810
rect 76356 800 76412 1428
rect 76468 1418 76524 1428
rect 76580 924 76636 1764
rect 76804 1594 76860 8260
rect 76916 6524 76972 6534
rect 76916 5906 76972 6468
rect 76916 5854 76918 5906
rect 76970 5854 76972 5906
rect 76916 5842 76972 5854
rect 77028 3948 77084 10276
rect 77140 9772 77196 9782
rect 77140 8316 77196 9716
rect 77140 8250 77196 8260
rect 77252 9658 77308 10724
rect 77588 9996 77644 10006
rect 77588 9902 77644 9940
rect 78260 9996 78316 11956
rect 78372 11844 78764 11900
rect 78372 10332 78428 11844
rect 78596 11676 78652 11686
rect 78708 11676 78764 11844
rect 78820 11676 78876 11686
rect 78708 11620 78820 11676
rect 78596 11564 78652 11620
rect 78820 11610 78876 11620
rect 78596 11508 78764 11564
rect 78708 11452 78764 11508
rect 78932 11452 78988 12404
rect 78708 11396 78988 11452
rect 79044 11340 79100 12628
rect 78372 10266 78428 10276
rect 78484 11284 79100 11340
rect 79156 12572 79212 12582
rect 78372 10108 78428 10118
rect 78372 10050 78428 10052
rect 78372 9998 78374 10050
rect 78426 9998 78428 10050
rect 78372 9986 78428 9998
rect 78260 9930 78316 9940
rect 78484 9828 78540 11284
rect 79156 11226 79212 12516
rect 79156 11174 79158 11226
rect 79210 11174 79212 11226
rect 79156 11162 79212 11174
rect 78820 11116 78876 11126
rect 79268 11116 79324 12740
rect 79380 12572 79436 14084
rect 80388 14028 80444 14200
rect 80724 14198 80726 14250
rect 80778 14198 80892 14250
rect 80724 14196 80892 14198
rect 80948 14362 81004 14374
rect 80948 14310 80950 14362
rect 81002 14310 81004 14362
rect 80724 14186 80780 14196
rect 79380 12506 79436 12516
rect 79492 13972 80444 14028
rect 80500 14138 80556 14150
rect 80500 14086 80502 14138
rect 80554 14086 80556 14138
rect 79492 11452 79548 13972
rect 79604 13802 79660 13814
rect 80500 13804 80556 14086
rect 79604 13750 79606 13802
rect 79658 13750 79660 13802
rect 79604 13242 79660 13750
rect 79604 13190 79606 13242
rect 79658 13190 79660 13242
rect 79604 13178 79660 13190
rect 80052 13748 80556 13804
rect 80836 14026 80892 14038
rect 80836 13974 80838 14026
rect 80890 13974 80892 14026
rect 80836 13804 80892 13974
rect 80948 14028 81004 14310
rect 81144 14200 81256 15000
rect 81508 14586 81564 14598
rect 81508 14534 81510 14586
rect 81562 14534 81564 14586
rect 80948 13962 81004 13972
rect 81060 14026 81116 14038
rect 81060 13974 81062 14026
rect 81114 13974 81116 14026
rect 81060 13804 81116 13974
rect 80836 13748 81116 13804
rect 79604 12796 79660 12806
rect 79604 12010 79660 12740
rect 79940 12458 79996 12470
rect 79940 12406 79942 12458
rect 79994 12406 79996 12458
rect 79716 12236 79772 12246
rect 79772 12180 79884 12236
rect 79716 12170 79772 12180
rect 79604 11958 79606 12010
rect 79658 11958 79660 12010
rect 79604 11946 79660 11958
rect 79380 11396 79548 11452
rect 79604 11674 79660 11686
rect 79604 11622 79606 11674
rect 79658 11622 79660 11674
rect 79380 11340 79436 11396
rect 79380 11274 79436 11284
rect 79604 11340 79660 11622
rect 79604 11274 79660 11284
rect 79492 11226 79548 11238
rect 79492 11174 79494 11226
rect 79546 11174 79548 11226
rect 79492 11116 79548 11174
rect 79268 11060 79548 11116
rect 78820 10892 78876 11060
rect 78820 10836 79772 10892
rect 78820 10388 79548 10444
rect 77252 9606 77254 9658
rect 77306 9606 77308 9658
rect 77252 7868 77308 9606
rect 78036 9772 78540 9828
rect 78596 10108 78652 10118
rect 78036 9324 78092 9772
rect 78260 9658 78316 9670
rect 78260 9606 78262 9658
rect 78314 9606 78316 9658
rect 78260 9436 78316 9606
rect 78428 9660 78484 9670
rect 78596 9660 78652 10052
rect 78428 9658 78652 9660
rect 78428 9606 78430 9658
rect 78482 9606 78652 9658
rect 78428 9604 78652 9606
rect 78428 9594 78484 9604
rect 78260 9380 78708 9436
rect 77476 9268 78092 9324
rect 78652 9324 78708 9380
rect 77476 8092 77532 9268
rect 78652 9210 78708 9268
rect 78652 9158 78654 9210
rect 78706 9158 78708 9210
rect 77588 9100 78428 9156
rect 78652 9146 78708 9158
rect 77588 8764 77644 9100
rect 78372 9055 78428 9100
rect 78820 9055 78876 10388
rect 79044 10220 79100 10230
rect 78932 10108 78988 10118
rect 78932 9770 78988 10052
rect 78932 9718 78934 9770
rect 78986 9718 78988 9770
rect 78932 9706 78988 9718
rect 78372 8999 78876 9055
rect 77588 8698 77644 8708
rect 77756 8986 77812 8998
rect 77756 8934 77758 8986
rect 77810 8934 77812 8986
rect 77756 8428 77812 8934
rect 78204 8988 78260 8998
rect 78204 8894 78260 8932
rect 77476 8026 77532 8036
rect 77588 8372 77812 8428
rect 77980 8652 78036 8662
rect 77588 7980 77644 8372
rect 77980 8314 78036 8596
rect 77980 8262 77982 8314
rect 78034 8262 78036 8314
rect 77980 8250 78036 8262
rect 77924 8092 77980 8102
rect 78316 8092 78372 8102
rect 77812 7980 77868 7990
rect 77588 7868 77644 7924
rect 77252 7812 77644 7868
rect 77700 7924 77812 7980
rect 77700 6860 77756 7924
rect 77812 7914 77868 7924
rect 77924 7457 77980 8036
rect 78148 8090 78372 8092
rect 78148 8038 78318 8090
rect 78370 8038 78372 8090
rect 78148 8036 78372 8038
rect 77196 6804 77756 6860
rect 77812 7401 77980 7457
rect 78036 7474 78092 7486
rect 78036 7422 78038 7474
rect 78090 7422 78092 7474
rect 77196 6690 77252 6804
rect 77196 6638 77198 6690
rect 77250 6638 77252 6690
rect 77196 6626 77252 6638
rect 77308 6524 77364 6534
rect 77308 6522 77420 6524
rect 77308 6470 77310 6522
rect 77362 6470 77420 6522
rect 77308 6458 77420 6470
rect 77364 5068 77420 6458
rect 77476 6086 77532 6804
rect 77476 6074 77588 6086
rect 77476 6022 77534 6074
rect 77586 6022 77588 6074
rect 77476 6020 77588 6022
rect 77532 6010 77588 6020
rect 77812 5964 77868 7401
rect 77924 7308 77980 7318
rect 77924 7214 77980 7252
rect 78036 6692 78092 7422
rect 77812 5898 77868 5908
rect 77980 6636 78092 6692
rect 78148 6681 78204 8036
rect 78316 8026 78372 8036
rect 78876 8092 78932 8102
rect 78876 7998 78932 8036
rect 79044 7868 79100 10164
rect 79268 10108 79324 10118
rect 79268 9994 79324 10052
rect 79268 9942 79270 9994
rect 79322 9942 79324 9994
rect 79268 9930 79324 9942
rect 78372 7812 79100 7868
rect 79156 9212 79212 9222
rect 78372 7586 78428 7812
rect 79156 7588 79212 9156
rect 79268 9098 79324 9110
rect 79268 9046 79270 9098
rect 79322 9046 79324 9098
rect 79268 8988 79324 9046
rect 79268 8316 79324 8932
rect 79492 8988 79548 10388
rect 79604 10220 79660 10230
rect 79604 9210 79660 10164
rect 79604 9158 79606 9210
rect 79658 9158 79660 9210
rect 79604 9146 79660 9158
rect 79492 8922 79548 8932
rect 79268 8250 79324 8260
rect 79436 8652 79492 8662
rect 79436 8146 79492 8596
rect 79716 8652 79772 10836
rect 79828 9660 79884 12180
rect 79940 12124 79996 12406
rect 80052 12460 80108 13748
rect 81172 13692 81228 14200
rect 80164 13636 81228 13692
rect 80164 12572 80220 13636
rect 80836 13242 80892 13254
rect 81172 13244 81228 13254
rect 80836 13190 80838 13242
rect 80890 13190 80892 13242
rect 80724 13130 80780 13142
rect 80724 13078 80726 13130
rect 80778 13078 80780 13130
rect 80164 12506 80220 12516
rect 80612 12682 80668 12694
rect 80612 12630 80614 12682
rect 80666 12630 80668 12682
rect 80052 12394 80108 12404
rect 80612 12458 80668 12630
rect 80612 12406 80614 12458
rect 80666 12406 80668 12458
rect 80612 12394 80668 12406
rect 80276 12346 80332 12358
rect 80276 12294 80278 12346
rect 80330 12294 80332 12346
rect 80276 12236 80332 12294
rect 80276 12180 80556 12236
rect 79940 12068 80444 12124
rect 80276 11898 80332 11910
rect 80276 11846 80278 11898
rect 80330 11846 80332 11898
rect 80164 11562 80220 11574
rect 80164 11510 80166 11562
rect 80218 11510 80220 11562
rect 80164 10780 80220 11510
rect 80276 11004 80332 11846
rect 80388 11674 80444 12068
rect 80500 11786 80556 12180
rect 80724 12234 80780 13078
rect 80836 12682 80892 13190
rect 80836 12630 80838 12682
rect 80890 12630 80892 12682
rect 80836 12618 80892 12630
rect 80948 13242 81228 13244
rect 80948 13190 81174 13242
rect 81226 13190 81228 13242
rect 80948 13188 81228 13190
rect 80948 12572 81004 13188
rect 81172 13178 81228 13188
rect 81508 13020 81564 14534
rect 81816 14200 81928 15000
rect 82068 14308 82348 14364
rect 81732 14140 81788 14150
rect 81844 14140 81900 14200
rect 82068 14140 82124 14308
rect 81732 14138 81900 14140
rect 81732 14086 81734 14138
rect 81786 14086 81900 14138
rect 81732 14084 81900 14086
rect 81956 14084 82124 14140
rect 82180 14138 82236 14150
rect 82180 14086 82182 14138
rect 82234 14086 82236 14138
rect 81732 14074 81788 14084
rect 81956 13804 82012 14084
rect 81732 13748 82012 13804
rect 82068 13916 82124 13926
rect 81732 13242 81788 13748
rect 82068 13690 82124 13860
rect 82068 13638 82070 13690
rect 82122 13638 82124 13690
rect 82068 13626 82124 13638
rect 81732 13190 81734 13242
rect 81786 13190 81788 13242
rect 81732 13178 81788 13190
rect 82180 13130 82236 14086
rect 82292 14140 82348 14308
rect 82600 14200 82712 15000
rect 82852 14812 82908 14822
rect 82852 14698 82908 14756
rect 82852 14646 82854 14698
rect 82906 14646 82908 14698
rect 82852 14634 82908 14646
rect 83076 14698 83132 14710
rect 83076 14646 83078 14698
rect 83130 14646 83132 14698
rect 82852 14476 82908 14486
rect 82628 14140 82684 14200
rect 82852 14140 82908 14420
rect 83076 14362 83132 14646
rect 83076 14310 83078 14362
rect 83130 14310 83132 14362
rect 83076 14298 83132 14310
rect 83272 14200 83384 15000
rect 83524 14924 83580 14934
rect 83748 14924 83804 14934
rect 83580 14868 83692 14924
rect 83524 14858 83580 14868
rect 82292 14084 82684 14140
rect 82740 14084 82908 14140
rect 82740 14028 82796 14084
rect 82292 13972 82796 14028
rect 82852 13972 83132 14028
rect 82292 13468 82348 13972
rect 82516 13802 82572 13814
rect 82516 13750 82518 13802
rect 82570 13750 82572 13802
rect 82292 13402 82348 13412
rect 82404 13690 82460 13702
rect 82404 13638 82406 13690
rect 82458 13638 82460 13690
rect 82404 13356 82460 13638
rect 82516 13692 82572 13750
rect 82740 13804 82796 13814
rect 82852 13804 82908 13972
rect 83076 13916 83132 13972
rect 83076 13850 83132 13860
rect 82740 13802 82908 13804
rect 82740 13750 82742 13802
rect 82794 13750 82908 13802
rect 82740 13748 82908 13750
rect 82964 13802 83020 13814
rect 82964 13750 82966 13802
rect 83018 13750 83020 13802
rect 82740 13738 82796 13748
rect 82516 13636 82684 13692
rect 82628 13580 82684 13636
rect 82852 13580 82908 13590
rect 82628 13578 82908 13580
rect 82628 13526 82854 13578
rect 82906 13526 82908 13578
rect 82628 13524 82908 13526
rect 82852 13514 82908 13524
rect 82404 13290 82460 13300
rect 82516 13468 82572 13478
rect 82180 13078 82182 13130
rect 82234 13078 82236 13130
rect 82180 13066 82236 13078
rect 82516 13020 82572 13412
rect 82740 13356 82796 13394
rect 82740 13290 82796 13300
rect 81508 12964 81788 13020
rect 81732 12908 81788 12964
rect 82292 12964 82572 13020
rect 82740 13130 82796 13142
rect 82740 13078 82742 13130
rect 82794 13078 82796 13130
rect 81732 12852 81900 12908
rect 81396 12684 81452 12694
rect 80948 12506 81004 12516
rect 81060 12682 81452 12684
rect 81060 12630 81398 12682
rect 81450 12630 81452 12682
rect 81060 12628 81452 12630
rect 81060 12458 81116 12628
rect 81396 12618 81452 12628
rect 81060 12406 81062 12458
rect 81114 12406 81116 12458
rect 81060 12394 81116 12406
rect 81732 12460 81788 12470
rect 81844 12460 81900 12852
rect 81956 12906 82012 12918
rect 82292 12908 82348 12964
rect 81956 12854 81958 12906
rect 82010 12854 82012 12906
rect 81956 12796 82012 12854
rect 82291 12852 82348 12908
rect 82291 12796 82347 12852
rect 81956 12740 82347 12796
rect 82404 12794 82460 12806
rect 82404 12742 82406 12794
rect 82458 12742 82460 12794
rect 82404 12684 82460 12742
rect 82292 12628 82460 12684
rect 82292 12570 82348 12628
rect 82292 12518 82294 12570
rect 82346 12518 82348 12570
rect 82292 12506 82348 12518
rect 82740 12460 82796 13078
rect 81732 12458 81900 12460
rect 81732 12406 81734 12458
rect 81786 12406 81900 12458
rect 81732 12404 81900 12406
rect 82516 12404 82796 12460
rect 81732 12394 81788 12404
rect 82516 12348 82572 12404
rect 80724 12182 80726 12234
rect 80778 12182 80780 12234
rect 80724 12170 80780 12182
rect 81956 12292 82572 12348
rect 81956 12234 82012 12292
rect 81956 12182 81958 12234
rect 82010 12182 82012 12234
rect 81956 12170 82012 12182
rect 82068 12180 82572 12236
rect 80836 12122 80892 12134
rect 81732 12124 81788 12134
rect 80836 12070 80838 12122
rect 80890 12070 80892 12122
rect 80500 11734 80502 11786
rect 80554 11734 80556 11786
rect 80500 11722 80556 11734
rect 80612 12010 80668 12022
rect 80612 11958 80614 12010
rect 80666 11958 80668 12010
rect 80388 11622 80390 11674
rect 80442 11622 80444 11674
rect 80388 11610 80444 11622
rect 80612 11226 80668 11958
rect 80612 11174 80614 11226
rect 80666 11174 80668 11226
rect 80612 11162 80668 11174
rect 80836 11226 80892 12070
rect 81396 12068 81732 12124
rect 80836 11174 80838 11226
rect 80890 11174 80892 11226
rect 80836 11162 80892 11174
rect 81060 12010 81116 12022
rect 81060 11958 81062 12010
rect 81114 11958 81116 12010
rect 81060 11004 81116 11958
rect 81284 11898 81340 11910
rect 81284 11846 81286 11898
rect 81338 11846 81340 11898
rect 81284 11452 81340 11846
rect 81396 11674 81452 12068
rect 81732 12058 81788 12068
rect 82068 12122 82124 12180
rect 82068 12070 82070 12122
rect 82122 12070 82124 12122
rect 82068 12058 82124 12070
rect 81956 12010 82012 12022
rect 81956 11958 81958 12010
rect 82010 11958 82012 12010
rect 81508 11900 81564 11910
rect 81508 11788 81564 11844
rect 81844 11898 81900 11910
rect 81844 11846 81846 11898
rect 81898 11846 81900 11898
rect 81508 11732 81788 11788
rect 81396 11622 81398 11674
rect 81450 11622 81452 11674
rect 81396 11610 81452 11622
rect 81732 11674 81788 11732
rect 81732 11622 81734 11674
rect 81786 11622 81788 11674
rect 81732 11610 81788 11622
rect 81844 11452 81900 11846
rect 81956 11900 82012 11958
rect 82516 12010 82572 12180
rect 82516 11958 82518 12010
rect 82570 11958 82572 12010
rect 82516 11946 82572 11958
rect 82740 12122 82796 12134
rect 82740 12070 82742 12122
rect 82794 12070 82796 12122
rect 82404 11900 82460 11910
rect 81956 11898 82460 11900
rect 81956 11846 82406 11898
rect 82458 11846 82460 11898
rect 81956 11844 82460 11846
rect 82404 11834 82460 11844
rect 82740 11900 82796 12070
rect 82852 12124 82908 12134
rect 82964 12124 83020 13750
rect 83188 13466 83244 13478
rect 83188 13414 83190 13466
rect 83242 13414 83244 13466
rect 83076 12572 83132 12582
rect 83076 12478 83132 12516
rect 83188 12348 83244 13414
rect 83188 12282 83244 12292
rect 82908 12068 83020 12124
rect 83076 12124 83132 12134
rect 82852 12058 82908 12068
rect 82740 11834 82796 11844
rect 81284 11396 81900 11452
rect 81956 11732 82236 11788
rect 81956 11340 82012 11732
rect 82180 11676 82236 11732
rect 83076 11676 83132 12068
rect 83300 12122 83356 14200
rect 83524 14026 83580 14038
rect 83524 13974 83526 14026
rect 83578 13974 83580 14026
rect 83412 12796 83468 12806
rect 83412 12572 83468 12740
rect 83412 12506 83468 12516
rect 83300 12070 83302 12122
rect 83354 12070 83356 12122
rect 83300 12058 83356 12070
rect 82180 11620 83132 11676
rect 83412 12012 83468 12022
rect 82068 11564 82124 11574
rect 82068 11562 82908 11564
rect 82068 11510 82070 11562
rect 82122 11510 82908 11562
rect 82068 11508 82908 11510
rect 82068 11498 82124 11508
rect 80276 10948 81116 11004
rect 81732 11284 82012 11340
rect 82404 11396 82796 11452
rect 81732 11004 81788 11284
rect 81732 10948 81900 11004
rect 81732 10780 81788 10790
rect 80164 10724 81732 10780
rect 81732 10714 81788 10724
rect 81844 10556 81900 10948
rect 82404 10892 82460 11396
rect 82516 11226 82572 11238
rect 82516 11174 82518 11226
rect 82570 11174 82572 11226
rect 82516 11004 82572 11174
rect 82740 11226 82796 11396
rect 82852 11450 82908 11508
rect 83188 11452 83244 11462
rect 82852 11398 82854 11450
rect 82906 11398 82908 11450
rect 82852 11386 82908 11398
rect 82964 11396 83188 11452
rect 82740 11174 82742 11226
rect 82794 11174 82796 11226
rect 82740 11162 82796 11174
rect 82964 11228 83020 11396
rect 83188 11386 83244 11396
rect 83412 11450 83468 11956
rect 83412 11398 83414 11450
rect 83466 11398 83468 11450
rect 83412 11386 83468 11398
rect 82964 11162 83020 11172
rect 82516 10948 82908 11004
rect 80948 10500 81900 10556
rect 82068 10836 82460 10892
rect 80948 9994 81004 10500
rect 82068 10444 82124 10836
rect 82852 10668 82908 10948
rect 83524 10780 83580 13974
rect 83636 13804 83692 14868
rect 83748 14138 83804 14868
rect 84056 14200 84168 15000
rect 84420 14698 84476 14710
rect 84420 14646 84422 14698
rect 84474 14646 84476 14698
rect 83748 14086 83750 14138
rect 83802 14086 83804 14138
rect 83748 14074 83804 14086
rect 83636 13748 83916 13804
rect 83748 13580 83804 13590
rect 83636 13356 83692 13366
rect 83636 12460 83692 13300
rect 83636 12394 83692 12404
rect 83748 12122 83804 13524
rect 83860 13356 83916 13748
rect 83860 13290 83916 13300
rect 83748 12070 83750 12122
rect 83802 12070 83804 12122
rect 83748 12058 83804 12070
rect 83860 12796 83916 12806
rect 83860 11452 83916 12740
rect 84084 12012 84140 14200
rect 84308 14138 84364 14150
rect 84308 14086 84310 14138
rect 84362 14086 84364 14138
rect 84308 13802 84364 14086
rect 84308 13750 84310 13802
rect 84362 13750 84364 13802
rect 84308 13738 84364 13750
rect 84196 13354 84252 13366
rect 84196 13302 84198 13354
rect 84250 13302 84252 13354
rect 84196 12460 84252 13302
rect 84420 13354 84476 14646
rect 84532 14362 84588 14374
rect 84532 14310 84534 14362
rect 84586 14310 84588 14362
rect 84532 14028 84588 14310
rect 84728 14200 84840 15000
rect 84980 14698 85036 14710
rect 84980 14646 84982 14698
rect 85034 14646 85036 14698
rect 84532 13972 84700 14028
rect 84420 13302 84422 13354
rect 84474 13302 84476 13354
rect 84420 13290 84476 13302
rect 84532 13802 84588 13814
rect 84532 13750 84534 13802
rect 84586 13750 84588 13802
rect 84532 12682 84588 13750
rect 84532 12630 84534 12682
rect 84586 12630 84588 12682
rect 84532 12618 84588 12630
rect 84644 12460 84700 13972
rect 84756 12572 84812 14200
rect 84980 13580 85036 14646
rect 85512 14200 85624 15000
rect 86184 14200 86296 15000
rect 86968 14200 87080 15000
rect 87640 14200 87752 15000
rect 88228 14250 88284 14262
rect 84980 13514 85036 13524
rect 84868 13132 84924 13142
rect 84868 12682 84924 13076
rect 84868 12630 84870 12682
rect 84922 12630 84924 12682
rect 84868 12618 84924 12630
rect 84756 12506 84812 12516
rect 84980 12572 85036 12582
rect 84196 12404 84700 12460
rect 83972 11956 84140 12012
rect 83972 11788 84028 11956
rect 83972 11722 84028 11732
rect 83860 11386 83916 11396
rect 83972 11562 84028 11574
rect 83972 11510 83974 11562
rect 84026 11510 84028 11562
rect 83972 11228 84028 11510
rect 84196 11340 84252 11350
rect 84420 11340 84476 11350
rect 84252 11284 84364 11340
rect 84196 11274 84252 11284
rect 83636 11172 84028 11228
rect 83636 11002 83692 11172
rect 83636 10950 83638 11002
rect 83690 10950 83692 11002
rect 83636 10938 83692 10950
rect 84308 11002 84364 11284
rect 84308 10950 84310 11002
rect 84362 10950 84364 11002
rect 84308 10938 84364 10950
rect 83524 10724 84140 10780
rect 82852 10612 84028 10668
rect 80948 9942 80950 9994
rect 81002 9942 81004 9994
rect 80948 9930 81004 9942
rect 81060 10388 82124 10444
rect 82180 10500 82460 10556
rect 81060 9828 81116 10388
rect 82180 10220 82236 10500
rect 82404 10444 82460 10500
rect 82404 10388 83356 10444
rect 82292 10332 82348 10342
rect 82348 10276 82572 10332
rect 82292 10266 82348 10276
rect 80108 9772 80164 9782
rect 80612 9772 80668 9782
rect 80108 9770 80668 9772
rect 80108 9718 80110 9770
rect 80162 9718 80614 9770
rect 80666 9718 80668 9770
rect 80108 9716 80668 9718
rect 80108 9706 80164 9716
rect 80612 9660 80668 9716
rect 80948 9772 81116 9828
rect 81172 10164 81452 10220
rect 80612 9604 80892 9660
rect 79828 9594 79884 9604
rect 80500 9212 80556 9222
rect 80612 9212 80668 9222
rect 80500 9210 80612 9212
rect 80500 9158 80502 9210
rect 80554 9158 80612 9210
rect 80500 9156 80612 9158
rect 80500 9146 80556 9156
rect 80612 9146 80668 9156
rect 80164 9100 80220 9110
rect 79716 8586 79772 8596
rect 79940 9098 80220 9100
rect 79940 9046 80166 9098
rect 80218 9046 80220 9098
rect 79940 9044 80220 9046
rect 79940 8764 79996 9044
rect 80164 9034 80220 9044
rect 80724 8988 80780 8998
rect 79324 8092 79380 8102
rect 78372 7534 78374 7586
rect 78426 7534 78428 7586
rect 78372 6758 78428 7534
rect 78708 7532 79212 7588
rect 79268 8090 79380 8092
rect 79268 8038 79326 8090
rect 79378 8038 79380 8090
rect 79268 8026 79380 8038
rect 79436 8094 79438 8146
rect 79490 8094 79492 8146
rect 78708 7308 78764 7532
rect 78708 7242 78764 7252
rect 78876 7418 78932 7430
rect 78876 7366 78878 7418
rect 78930 7366 78932 7418
rect 78876 7308 78932 7366
rect 78876 7242 78932 7252
rect 79268 7084 79324 8026
rect 79436 7868 79492 8094
rect 79436 7812 79884 7868
rect 79436 7644 79492 7654
rect 79436 7550 79492 7588
rect 78316 6746 78428 6758
rect 78316 6694 78318 6746
rect 78370 6694 78428 6746
rect 78316 6692 78428 6694
rect 78484 7028 79100 7084
rect 78316 6682 78372 6692
rect 77980 6522 78036 6636
rect 78148 6625 78260 6681
rect 78204 6580 78260 6625
rect 77980 6470 77982 6522
rect 78034 6470 78036 6522
rect 77980 5908 78036 6470
rect 78092 6524 78148 6534
rect 78204 6524 78428 6580
rect 78092 6074 78148 6468
rect 78092 6022 78094 6074
rect 78146 6022 78148 6074
rect 78092 6010 78148 6022
rect 77980 5852 78204 5908
rect 77364 5002 77420 5012
rect 77700 4620 77756 4630
rect 77028 3882 77084 3892
rect 77140 4116 77644 4172
rect 77140 3722 77196 4116
rect 77364 3948 77420 3986
rect 77364 3882 77420 3892
rect 77588 3946 77644 4116
rect 77588 3894 77590 3946
rect 77642 3894 77644 3946
rect 77588 3882 77644 3894
rect 77140 3670 77142 3722
rect 77194 3670 77196 3722
rect 77140 3658 77196 3670
rect 77364 3722 77420 3734
rect 77364 3670 77366 3722
rect 77418 3670 77420 3722
rect 77364 3498 77420 3670
rect 77700 3724 77756 4564
rect 78036 3946 78092 3958
rect 78036 3894 78038 3946
rect 78090 3894 78092 3946
rect 77700 3668 77980 3724
rect 77812 3500 77868 3510
rect 77364 3446 77366 3498
rect 77418 3446 77420 3498
rect 77364 3434 77420 3446
rect 77700 3444 77812 3500
rect 76804 1542 76806 1594
rect 76858 1542 76860 1594
rect 76804 1530 76860 1542
rect 76916 3052 76972 3062
rect 76692 1372 76748 1382
rect 76692 1036 76748 1316
rect 76692 970 76748 980
rect 76580 858 76636 868
rect 76692 812 76748 822
rect 76132 746 76188 758
rect 76328 0 76440 800
rect 76916 800 76972 2996
rect 77700 1148 77756 3444
rect 77812 3434 77868 3444
rect 77588 1092 77756 1148
rect 77812 2378 77868 2390
rect 77812 2326 77814 2378
rect 77866 2326 77868 2378
rect 77252 1034 77308 1046
rect 77252 982 77254 1034
rect 77306 982 77308 1034
rect 77140 810 77196 822
rect 76692 718 76748 756
rect 76888 0 77000 800
rect 77140 758 77142 810
rect 77194 758 77196 810
rect 77140 588 77196 758
rect 77252 812 77308 982
rect 77252 746 77308 756
rect 77364 810 77420 822
rect 77364 758 77366 810
rect 77418 758 77420 810
rect 77588 800 77644 1092
rect 77140 522 77196 532
rect 77364 250 77420 758
rect 77364 198 77366 250
rect 77418 198 77420 250
rect 77364 186 77420 198
rect 77560 0 77672 800
rect 77812 250 77868 2326
rect 77924 2156 77980 3668
rect 78036 3500 78092 3894
rect 78036 3434 78092 3444
rect 78148 2828 78204 5852
rect 78260 4620 78316 4630
rect 78260 4396 78316 4564
rect 78260 4330 78316 4340
rect 78260 4172 78316 4182
rect 78260 3946 78316 4116
rect 78260 3894 78262 3946
rect 78314 3894 78316 3946
rect 78260 3882 78316 3894
rect 78260 3612 78316 3622
rect 78372 3612 78428 6524
rect 78484 6412 78540 7028
rect 78484 6346 78540 6356
rect 78596 6860 78652 6870
rect 78596 5862 78652 6804
rect 79044 6748 79100 7028
rect 79548 7474 79604 7486
rect 79548 7422 79550 7474
rect 79602 7422 79604 7474
rect 79548 7084 79604 7422
rect 79828 7084 79884 7812
rect 79548 7028 79660 7084
rect 79268 7018 79324 7028
rect 79268 6748 79324 6758
rect 78820 6690 78876 6702
rect 79044 6692 79268 6748
rect 78820 6638 78822 6690
rect 78874 6638 78876 6690
rect 79268 6682 79324 6692
rect 78820 6636 78876 6638
rect 78820 6570 78876 6580
rect 78540 5852 78652 5862
rect 78484 5850 78652 5852
rect 78484 5798 78542 5850
rect 78594 5798 78652 5850
rect 78484 5796 78652 5798
rect 79604 5852 79660 7028
rect 79828 7018 79884 7028
rect 79828 6860 79884 6870
rect 79828 6690 79884 6804
rect 79828 6638 79830 6690
rect 79882 6638 79884 6690
rect 79828 6626 79884 6638
rect 79772 5852 79828 5862
rect 79604 5850 79884 5852
rect 79604 5798 79774 5850
rect 79826 5798 79884 5850
rect 79604 5796 79884 5798
rect 78484 5786 78596 5796
rect 79772 5786 79884 5796
rect 78484 4956 78540 5786
rect 79268 5122 79324 5134
rect 79268 5070 79270 5122
rect 79322 5070 79324 5122
rect 78484 4890 78540 4900
rect 79044 5010 79100 5022
rect 79044 4958 79046 5010
rect 79098 4958 79100 5010
rect 79044 4396 79100 4958
rect 79268 4956 79324 5070
rect 79828 5067 79884 5786
rect 79268 4890 79324 4900
rect 79604 5011 79884 5067
rect 79604 4732 79660 5011
rect 79604 4676 79772 4732
rect 79044 4330 79100 4340
rect 79492 4508 79548 4518
rect 78596 4060 78652 4070
rect 79380 4060 79436 4070
rect 78652 4004 79100 4060
rect 78596 3994 78652 4004
rect 79044 3948 79100 4004
rect 79268 4004 79380 4060
rect 79268 3948 79324 4004
rect 79380 3994 79436 4004
rect 78708 3892 78988 3948
rect 79044 3892 79324 3948
rect 78708 3834 78764 3892
rect 78708 3782 78710 3834
rect 78762 3782 78764 3834
rect 78708 3770 78764 3782
rect 78596 3722 78652 3734
rect 78596 3670 78598 3722
rect 78650 3670 78652 3722
rect 78316 3556 78540 3612
rect 78260 3546 78316 3556
rect 78484 3276 78540 3556
rect 78596 3500 78652 3670
rect 78596 3434 78652 3444
rect 78820 3722 78876 3734
rect 78820 3670 78822 3722
rect 78874 3670 78876 3722
rect 78820 3386 78876 3670
rect 78932 3724 78988 3892
rect 78932 3668 79324 3724
rect 79268 3610 79324 3668
rect 79268 3558 79270 3610
rect 79322 3558 79324 3610
rect 79268 3546 79324 3558
rect 79380 3612 79436 3622
rect 79044 3500 79100 3510
rect 79156 3500 79212 3510
rect 79044 3498 79156 3500
rect 79044 3446 79046 3498
rect 79098 3446 79156 3498
rect 79044 3444 79156 3446
rect 79044 3434 79100 3444
rect 79156 3434 79212 3444
rect 78820 3334 78822 3386
rect 78874 3334 78876 3386
rect 78820 3322 78876 3334
rect 78708 3276 78764 3286
rect 79380 3276 79436 3556
rect 78484 3210 78540 3220
rect 78596 3274 78764 3276
rect 78596 3222 78710 3274
rect 78762 3222 78764 3274
rect 78596 3220 78764 3222
rect 78484 3052 78540 3062
rect 78596 3052 78652 3220
rect 78708 3210 78764 3220
rect 79044 3220 79436 3276
rect 79492 3276 79548 4452
rect 79604 4506 79660 4518
rect 79604 4454 79606 4506
rect 79658 4454 79660 4506
rect 79604 4284 79660 4454
rect 79716 4508 79772 4676
rect 79716 4442 79772 4452
rect 79828 4394 79884 4406
rect 79828 4342 79830 4394
rect 79882 4342 79884 4394
rect 79828 4284 79884 4342
rect 79604 4228 79884 4284
rect 79940 3948 79996 8708
rect 80612 8932 80724 8988
rect 80052 8092 80108 8102
rect 80052 6972 80108 8036
rect 80388 8092 80444 8102
rect 80388 7998 80444 8036
rect 80052 5180 80108 6916
rect 80164 7530 80220 7542
rect 80164 7478 80166 7530
rect 80218 7478 80220 7530
rect 80164 7308 80220 7478
rect 80164 6188 80220 7252
rect 80276 7420 80332 7430
rect 80276 6412 80332 7364
rect 80500 7308 80556 7318
rect 80500 7214 80556 7252
rect 80276 6346 80332 6356
rect 80500 6412 80556 6422
rect 80500 6188 80556 6356
rect 80164 6132 80556 6188
rect 80500 5628 80556 5638
rect 80052 5114 80108 5124
rect 80276 5572 80500 5628
rect 80108 4956 80164 4966
rect 80276 4956 80332 5572
rect 80500 5562 80556 5572
rect 80164 4900 80332 4956
rect 80108 4824 80164 4900
rect 80052 4394 80108 4406
rect 80052 4342 80054 4394
rect 80106 4342 80108 4394
rect 80052 4172 80108 4342
rect 80052 4106 80108 4116
rect 80276 4394 80332 4406
rect 80276 4342 80278 4394
rect 80330 4342 80332 4394
rect 79940 3892 80108 3948
rect 79828 3834 79884 3846
rect 79828 3782 79830 3834
rect 79882 3782 79884 3834
rect 79716 3386 79772 3398
rect 79716 3334 79718 3386
rect 79770 3334 79772 3386
rect 79492 3220 79660 3276
rect 78932 3162 78988 3174
rect 78932 3110 78934 3162
rect 78986 3110 78988 3162
rect 78484 3050 78652 3052
rect 78484 2998 78486 3050
rect 78538 2998 78652 3050
rect 78484 2996 78652 2998
rect 78708 3050 78764 3062
rect 78708 2998 78710 3050
rect 78762 2998 78764 3050
rect 78484 2986 78540 2996
rect 78148 2772 78540 2828
rect 77924 2100 78092 2156
rect 78036 1036 78092 2100
rect 78260 1596 78316 1606
rect 78260 1594 78428 1596
rect 78260 1542 78262 1594
rect 78314 1542 78428 1594
rect 78260 1540 78428 1542
rect 78260 1530 78316 1540
rect 78036 980 78204 1036
rect 77924 922 77980 934
rect 77924 870 77926 922
rect 77978 870 77980 922
rect 77924 698 77980 870
rect 78148 800 78204 980
rect 77924 646 77926 698
rect 77978 646 77980 698
rect 77924 634 77980 646
rect 77812 198 77814 250
rect 77866 198 77868 250
rect 77812 186 77868 198
rect 78120 0 78232 800
rect 78372 698 78428 1540
rect 78484 1594 78540 2772
rect 78708 1708 78764 2998
rect 78932 2378 78988 3110
rect 79044 3050 79100 3220
rect 79604 3162 79660 3220
rect 79604 3110 79606 3162
rect 79658 3110 79660 3162
rect 79604 3098 79660 3110
rect 79044 2998 79046 3050
rect 79098 2998 79100 3050
rect 79044 2986 79100 2998
rect 79716 3050 79772 3334
rect 79716 2998 79718 3050
rect 79770 2998 79772 3050
rect 79716 2986 79772 2998
rect 79604 2938 79660 2950
rect 79604 2886 79606 2938
rect 79658 2886 79660 2938
rect 79044 2716 79100 2726
rect 79492 2716 79548 2726
rect 79044 2714 79548 2716
rect 79044 2662 79046 2714
rect 79098 2662 79494 2714
rect 79546 2662 79548 2714
rect 79044 2660 79548 2662
rect 79044 2650 79100 2660
rect 79492 2650 79548 2660
rect 79604 2602 79660 2886
rect 79604 2550 79606 2602
rect 79658 2550 79660 2602
rect 79604 2538 79660 2550
rect 78932 2326 78934 2378
rect 78986 2326 78988 2378
rect 78932 2314 78988 2326
rect 79828 2380 79884 3782
rect 79940 3612 79996 3622
rect 79940 3052 79996 3556
rect 79940 2986 79996 2996
rect 79828 2314 79884 2324
rect 78484 1542 78486 1594
rect 78538 1542 78540 1594
rect 78484 1530 78540 1542
rect 78596 1652 78764 1708
rect 78372 646 78374 698
rect 78426 646 78428 698
rect 78372 634 78428 646
rect 78596 700 78652 1652
rect 78932 1540 79212 1596
rect 78708 1372 78764 1382
rect 78764 1316 78876 1372
rect 78708 1306 78764 1316
rect 78820 800 78876 1316
rect 78932 1148 78988 1540
rect 79156 1484 79212 1540
rect 79492 1484 79548 1494
rect 79156 1428 79492 1484
rect 79492 1418 79548 1428
rect 79044 1372 79100 1382
rect 79100 1316 79436 1372
rect 79044 1306 79100 1316
rect 78932 1092 79100 1148
rect 78596 634 78652 644
rect 78792 0 78904 800
rect 79044 476 79100 1092
rect 79380 800 79436 1316
rect 80052 800 80108 3892
rect 80276 3836 80332 4342
rect 80276 3770 80332 3780
rect 80388 3610 80444 3622
rect 80388 3558 80390 3610
rect 80442 3558 80444 3610
rect 80388 3500 80444 3558
rect 80388 3434 80444 3444
rect 80164 3050 80220 3062
rect 80164 2998 80166 3050
rect 80218 2998 80220 3050
rect 80164 2602 80220 2998
rect 80164 2550 80166 2602
rect 80218 2550 80220 2602
rect 80164 2538 80220 2550
rect 80164 1372 80220 1382
rect 80164 924 80220 1316
rect 80164 858 80220 868
rect 80612 800 80668 8932
rect 80724 8922 80780 8932
rect 80836 6412 80892 9604
rect 80948 8764 81004 9772
rect 81060 9660 81116 9670
rect 81060 8988 81116 9604
rect 81172 9324 81228 10164
rect 81284 9996 81340 10006
rect 81396 9996 81452 10164
rect 82180 10154 82236 10164
rect 81844 9996 81900 10006
rect 81396 9994 81900 9996
rect 81396 9942 81846 9994
rect 81898 9942 81900 9994
rect 81396 9940 81900 9942
rect 82516 9996 82572 10276
rect 82704 10220 82968 10230
rect 82760 10164 82808 10220
rect 82864 10164 82912 10220
rect 82704 10154 82968 10164
rect 83188 10220 83244 10230
rect 83188 10052 83244 10164
rect 83300 10108 83356 10388
rect 83748 10442 83804 10454
rect 83748 10390 83750 10442
rect 83802 10390 83804 10442
rect 83748 10332 83804 10390
rect 83972 10442 84028 10612
rect 83972 10390 83974 10442
rect 84026 10390 84028 10442
rect 83972 10378 84028 10390
rect 83748 10266 83804 10276
rect 84084 10108 84140 10724
rect 83300 10052 84140 10108
rect 82908 9996 83244 10052
rect 84308 9996 84364 10006
rect 82516 9940 82964 9996
rect 83860 9940 84308 9996
rect 81284 9436 81340 9940
rect 81844 9930 81900 9940
rect 83860 9884 83916 9940
rect 84308 9930 84364 9940
rect 83412 9828 83916 9884
rect 81396 9772 82460 9828
rect 82628 9772 83020 9828
rect 83132 9772 83188 9782
rect 81396 9660 81452 9772
rect 82404 9770 82684 9772
rect 82404 9718 82406 9770
rect 82458 9718 82684 9770
rect 82404 9716 82684 9718
rect 82964 9770 83188 9772
rect 82964 9718 83134 9770
rect 83186 9718 83188 9770
rect 82964 9716 83188 9718
rect 82404 9706 82460 9716
rect 83132 9706 83188 9716
rect 81396 9594 81452 9604
rect 81508 9660 81564 9670
rect 81620 9660 81676 9670
rect 81508 9658 81620 9660
rect 81508 9606 81510 9658
rect 81562 9606 81620 9658
rect 81508 9604 81620 9606
rect 81508 9594 81564 9604
rect 81620 9594 81676 9604
rect 82740 9658 82796 9670
rect 82740 9606 82742 9658
rect 82794 9606 82796 9658
rect 82740 9548 82796 9606
rect 83412 9548 83468 9828
rect 83916 9660 83972 9670
rect 83916 9566 83972 9604
rect 84084 9660 84140 9670
rect 82740 9492 83468 9548
rect 84084 9436 84140 9604
rect 81284 9380 84140 9436
rect 84420 9324 84476 11284
rect 84644 10780 84700 10790
rect 84644 9436 84700 10724
rect 84644 9370 84700 9380
rect 81172 9268 82348 9324
rect 82292 9212 82348 9268
rect 82628 9268 84476 9324
rect 82292 9146 82348 9156
rect 82516 9212 82572 9250
rect 82516 9146 82572 9156
rect 81284 9098 81340 9110
rect 81284 9046 81286 9098
rect 81338 9046 81340 9098
rect 81284 8988 81340 9046
rect 82180 9098 82236 9110
rect 82180 9046 82182 9098
rect 82234 9046 82236 9098
rect 82180 8988 82236 9046
rect 82628 9044 82684 9268
rect 84980 9212 85036 12516
rect 85092 11002 85148 11014
rect 85092 10950 85094 11002
rect 85146 10950 85148 11002
rect 85092 10892 85148 10950
rect 85092 10826 85148 10836
rect 85316 11002 85372 11014
rect 85316 10950 85318 11002
rect 85370 10950 85372 11002
rect 81284 8932 81564 8988
rect 81060 8922 81116 8932
rect 81508 8876 81564 8932
rect 82180 8922 82236 8932
rect 82404 8988 82684 9044
rect 82740 9156 85036 9212
rect 80948 8708 81452 8764
rect 81396 8428 81452 8708
rect 81508 8540 81564 8820
rect 81620 8874 81676 8886
rect 81620 8822 81622 8874
rect 81674 8822 81676 8874
rect 81620 8764 81676 8822
rect 82404 8764 82460 8988
rect 82740 8876 82796 9156
rect 81620 8708 82460 8764
rect 82516 8820 82796 8876
rect 83076 9042 83132 9054
rect 83076 8990 83078 9042
rect 83130 8990 83132 9042
rect 82516 8652 82572 8820
rect 82516 8586 82572 8596
rect 82704 8652 82968 8662
rect 82760 8596 82808 8652
rect 82864 8596 82912 8652
rect 82704 8586 82968 8596
rect 83076 8652 83132 8990
rect 83076 8586 83132 8596
rect 83188 8988 83580 9044
rect 83804 8988 83860 8998
rect 81508 8484 81676 8540
rect 81396 8372 81564 8428
rect 81284 8204 81340 8214
rect 81284 7756 81340 8148
rect 81284 7700 81452 7756
rect 81284 7474 81340 7486
rect 81284 7422 81286 7474
rect 81338 7422 81340 7474
rect 81172 7362 81228 7374
rect 81172 7310 81174 7362
rect 81226 7310 81228 7362
rect 81172 7308 81228 7310
rect 81172 7242 81228 7252
rect 80836 6356 81116 6412
rect 80836 4956 80892 4966
rect 80836 4284 80892 4900
rect 80724 4228 80892 4284
rect 80724 3836 80780 4228
rect 80724 3770 80780 3780
rect 80836 3946 80892 3958
rect 80836 3894 80838 3946
rect 80890 3894 80892 3946
rect 80836 2380 80892 3894
rect 80948 3724 81004 3734
rect 80948 3050 81004 3668
rect 80948 2998 80950 3050
rect 81002 2998 81004 3050
rect 80948 2986 81004 2998
rect 80836 2314 80892 2324
rect 80948 1932 81004 1942
rect 80724 1876 80948 1932
rect 80724 1036 80780 1876
rect 80948 1866 81004 1876
rect 81060 1484 81116 6356
rect 81284 5180 81340 7422
rect 81396 6020 81452 7700
rect 81508 6746 81564 8372
rect 81508 6694 81510 6746
rect 81562 6694 81564 6746
rect 81508 6682 81564 6694
rect 81508 6020 81564 6030
rect 81396 6018 81564 6020
rect 81396 5966 81510 6018
rect 81562 5966 81564 6018
rect 81396 5964 81564 5966
rect 81508 5954 81564 5964
rect 81620 5852 81676 8484
rect 83188 8428 83244 8988
rect 82180 8372 83244 8428
rect 83412 8874 83468 8886
rect 83412 8822 83414 8874
rect 83466 8822 83468 8874
rect 81844 8316 81900 8326
rect 81508 5796 81676 5852
rect 81732 8204 81788 8214
rect 81396 5180 81452 5190
rect 81284 5178 81452 5180
rect 81284 5126 81398 5178
rect 81450 5126 81452 5178
rect 81284 5124 81452 5126
rect 81396 5114 81452 5124
rect 81284 4956 81340 4966
rect 81284 3276 81340 4900
rect 81396 4394 81452 4406
rect 81396 4342 81398 4394
rect 81450 4342 81452 4394
rect 81396 3946 81452 4342
rect 81396 3894 81398 3946
rect 81450 3894 81452 3946
rect 81396 3882 81452 3894
rect 81284 3210 81340 3220
rect 81396 3500 81452 3510
rect 81396 2940 81452 3444
rect 81508 3162 81564 5796
rect 81620 5516 81676 5526
rect 81620 5010 81676 5460
rect 81620 4958 81622 5010
rect 81674 4958 81676 5010
rect 81620 4946 81676 4958
rect 81732 3834 81788 8148
rect 81844 7644 81900 8260
rect 82068 8316 82124 8326
rect 81956 8092 82012 8102
rect 82068 8092 82124 8260
rect 81956 8090 82124 8092
rect 81956 8038 81958 8090
rect 82010 8038 82124 8090
rect 81956 8036 82124 8038
rect 82180 8092 82236 8372
rect 83412 8316 83468 8822
rect 83524 8428 83580 8988
rect 83748 8986 83860 8988
rect 83748 8934 83806 8986
rect 83858 8934 83860 8986
rect 83748 8922 83860 8934
rect 84252 8988 84308 8998
rect 83748 8652 83804 8922
rect 84252 8894 84308 8932
rect 84700 8986 84756 8998
rect 84700 8934 84702 8986
rect 84754 8934 84756 8986
rect 84700 8764 84756 8934
rect 84700 8698 84756 8708
rect 84868 8764 84924 8774
rect 83748 8586 83804 8596
rect 84868 8540 84924 8708
rect 84084 8484 84924 8540
rect 84084 8428 84140 8484
rect 83524 8372 84140 8428
rect 85316 8316 85372 10950
rect 85540 9212 85596 14200
rect 85988 10892 86044 10902
rect 85988 10108 86044 10836
rect 86212 10892 86268 14200
rect 86660 13132 86716 13142
rect 86212 10826 86268 10836
rect 86436 11226 86492 11238
rect 86436 11174 86438 11226
rect 86490 11174 86492 11226
rect 86436 10892 86492 11174
rect 86660 11226 86716 13076
rect 86996 11564 87052 14200
rect 86996 11498 87052 11508
rect 87220 14026 87276 14038
rect 87220 13974 87222 14026
rect 87274 13974 87276 14026
rect 87220 11564 87276 13974
rect 87220 11498 87276 11508
rect 86660 11174 86662 11226
rect 86714 11174 86716 11226
rect 86660 11162 86716 11174
rect 86436 10826 86492 10836
rect 86548 10780 86604 10790
rect 86100 10108 86156 10118
rect 85988 10052 86100 10108
rect 86100 10042 86156 10052
rect 85540 9146 85596 9156
rect 85932 9660 85988 9670
rect 85932 9044 85988 9604
rect 86436 9660 86492 9670
rect 86436 9566 86492 9604
rect 86548 9222 86604 10724
rect 86772 10108 86828 10118
rect 86772 9994 86828 10052
rect 86772 9942 86774 9994
rect 86826 9942 86828 9994
rect 86772 9930 86828 9942
rect 87668 9996 87724 14200
rect 88228 14198 88230 14250
rect 88282 14198 88284 14250
rect 88424 14200 88536 15000
rect 88676 14250 88732 14262
rect 88228 14026 88284 14198
rect 88228 13974 88230 14026
rect 88282 13974 88284 14026
rect 88228 13962 88284 13974
rect 88452 12906 88508 14200
rect 88676 14198 88678 14250
rect 88730 14198 88732 14250
rect 89096 14200 89208 15000
rect 89880 14200 89992 15000
rect 90552 14200 90664 15000
rect 90804 14698 90860 14710
rect 90804 14646 90806 14698
rect 90858 14646 90860 14698
rect 88676 13132 88732 14198
rect 88676 13066 88732 13076
rect 88452 12854 88454 12906
rect 88506 12854 88508 12906
rect 88452 12842 88508 12854
rect 88676 12906 88732 12918
rect 88676 12854 88678 12906
rect 88730 12854 88732 12906
rect 87668 9930 87724 9940
rect 87780 12572 87836 12582
rect 87332 9660 87388 9670
rect 86492 9212 86604 9222
rect 86044 9210 86604 9212
rect 86044 9158 86494 9210
rect 86546 9158 86604 9210
rect 86044 9156 86604 9158
rect 87220 9212 87276 9222
rect 86044 9154 86100 9156
rect 86044 9102 86046 9154
rect 86098 9102 86100 9154
rect 86492 9146 86548 9156
rect 86044 9090 86100 9102
rect 85652 8988 85708 8998
rect 85652 8652 85708 8932
rect 85652 8586 85708 8596
rect 85764 8988 85988 9044
rect 87052 8988 87108 8998
rect 85764 8316 85820 8988
rect 86548 8986 87108 8988
rect 86548 8934 87054 8986
rect 87106 8934 87108 8986
rect 86548 8932 87108 8934
rect 85932 8874 85988 8886
rect 85932 8822 85934 8874
rect 85986 8822 85988 8874
rect 85932 8428 85988 8822
rect 86212 8764 86268 8774
rect 86268 8708 86380 8764
rect 86212 8698 86268 8708
rect 85932 8362 85988 8372
rect 86100 8428 86156 8438
rect 81956 8026 82012 8036
rect 82180 8026 82236 8036
rect 83300 8258 83356 8270
rect 83412 8260 84252 8316
rect 83300 8206 83302 8258
rect 83354 8206 83356 8258
rect 83300 7868 83356 8206
rect 84084 7980 84140 7990
rect 83300 7812 83468 7868
rect 83300 7644 83356 7654
rect 81844 7588 83300 7644
rect 83300 7578 83356 7588
rect 81844 7474 81900 7486
rect 81844 7422 81846 7474
rect 81898 7422 81900 7474
rect 81844 6524 81900 7422
rect 83412 7420 83468 7812
rect 84084 7756 84140 7924
rect 84196 7868 84252 8260
rect 84420 8258 84476 8270
rect 84420 8206 84422 8258
rect 84474 8206 84476 8258
rect 85316 8250 85372 8260
rect 85540 8260 85820 8316
rect 84420 8092 84476 8206
rect 84420 8026 84476 8036
rect 85260 8090 85316 8102
rect 85260 8038 85262 8090
rect 85314 8038 85316 8090
rect 85260 7980 85316 8038
rect 85260 7914 85316 7924
rect 84196 7812 84476 7868
rect 84084 7700 84364 7756
rect 81844 6458 81900 6468
rect 81956 7364 83468 7420
rect 81844 5010 81900 5022
rect 81844 4958 81846 5010
rect 81898 4958 81900 5010
rect 81844 4058 81900 4958
rect 81956 4956 82012 7364
rect 82516 7252 83692 7308
rect 82292 7196 82348 7206
rect 82516 7196 82572 7252
rect 82348 7140 82572 7196
rect 83636 7196 83692 7252
rect 82292 7130 82348 7140
rect 83636 7130 83692 7140
rect 82704 7084 82968 7094
rect 82760 7028 82808 7084
rect 82864 7028 82912 7084
rect 82704 7018 82968 7028
rect 83412 6972 83468 6982
rect 83020 6916 83412 6972
rect 82628 6860 82684 6870
rect 83020 6860 83076 6916
rect 83412 6906 83468 6916
rect 84308 6972 84364 7700
rect 84420 7644 84476 7812
rect 85540 7756 85596 8260
rect 85820 8146 85876 8158
rect 84420 7578 84476 7588
rect 84756 7700 85596 7756
rect 85708 8090 85764 8102
rect 85708 8038 85710 8090
rect 85762 8038 85764 8090
rect 85708 7756 85764 8038
rect 85820 8094 85822 8146
rect 85874 8094 85876 8146
rect 85820 7980 85876 8094
rect 85820 7914 85876 7924
rect 84420 7308 84476 7318
rect 84420 7214 84476 7252
rect 84308 6906 84364 6916
rect 82516 6804 82628 6860
rect 82516 6636 82572 6804
rect 82628 6794 82684 6804
rect 82908 6804 83076 6860
rect 84196 6860 84252 6870
rect 82516 6570 82572 6580
rect 82740 6748 82796 6758
rect 82292 6524 82348 6534
rect 82348 6468 82460 6524
rect 82292 6458 82348 6468
rect 82180 6412 82236 6422
rect 82404 6412 82460 6468
rect 82740 6412 82796 6692
rect 82908 6690 82964 6804
rect 82908 6638 82910 6690
rect 82962 6638 82964 6690
rect 83468 6748 83524 6758
rect 83748 6748 83804 6758
rect 84028 6748 84084 6758
rect 83468 6746 83692 6748
rect 83468 6694 83470 6746
rect 83522 6694 83692 6746
rect 83468 6692 83692 6694
rect 83468 6682 83524 6692
rect 82908 6626 82964 6638
rect 83020 6522 83076 6534
rect 83020 6470 83022 6522
rect 83074 6470 83076 6522
rect 83020 6468 83076 6470
rect 83020 6412 83244 6468
rect 82404 6356 82796 6412
rect 82180 5740 82236 6356
rect 83188 6076 83244 6412
rect 82180 5674 82236 5684
rect 82516 6020 83132 6076
rect 82516 5516 82572 6020
rect 82740 5906 82796 5918
rect 82740 5854 82742 5906
rect 82794 5854 82796 5906
rect 82740 5740 82796 5854
rect 83076 5908 83132 6020
rect 83188 6010 83244 6020
rect 83636 5908 83692 6692
rect 83804 6746 84084 6748
rect 83804 6694 84030 6746
rect 84082 6694 84084 6746
rect 83804 6692 84084 6694
rect 83748 6682 83804 6692
rect 83076 5852 83692 5908
rect 82740 5674 82796 5684
rect 82516 5450 82572 5460
rect 82704 5516 82968 5526
rect 82760 5460 82808 5516
rect 82864 5460 82912 5516
rect 82704 5450 82968 5460
rect 83076 5348 83468 5404
rect 82292 5180 82348 5190
rect 83076 5180 83132 5348
rect 82348 5124 83132 5180
rect 83188 5180 83244 5190
rect 82292 5114 82348 5124
rect 83188 5122 83244 5124
rect 83188 5070 83190 5122
rect 83242 5070 83244 5122
rect 83188 5058 83244 5070
rect 81956 4890 82012 4900
rect 82964 4900 83356 4956
rect 81844 4006 81846 4058
rect 81898 4006 81900 4058
rect 81844 3994 81900 4006
rect 82068 4844 82124 4854
rect 82068 4058 82124 4788
rect 82292 4732 82348 4742
rect 82292 4394 82348 4676
rect 82292 4342 82294 4394
rect 82346 4342 82348 4394
rect 82292 4330 82348 4342
rect 82068 4006 82070 4058
rect 82122 4006 82124 4058
rect 82068 3994 82124 4006
rect 82180 4284 82236 4294
rect 81732 3782 81734 3834
rect 81786 3782 81788 3834
rect 81732 3770 81788 3782
rect 82180 3724 82236 4228
rect 82068 3668 82236 3724
rect 82292 3834 82348 3846
rect 82292 3782 82294 3834
rect 82346 3782 82348 3834
rect 82068 3388 82124 3668
rect 81508 3110 81510 3162
rect 81562 3110 81564 3162
rect 81508 3098 81564 3110
rect 81620 3332 82124 3388
rect 81620 2940 81676 3332
rect 81396 2884 81676 2940
rect 81956 3162 82012 3174
rect 82292 3164 82348 3782
rect 82516 3724 82572 3734
rect 81956 3110 81958 3162
rect 82010 3110 82012 3162
rect 81956 2604 82012 3110
rect 81844 2548 82012 2604
rect 82068 3108 82348 3164
rect 82404 3162 82460 3174
rect 82404 3110 82406 3162
rect 82458 3110 82460 3162
rect 81172 2380 81228 2390
rect 81172 1708 81228 2324
rect 81620 2380 81676 2390
rect 81620 2156 81676 2324
rect 81172 1642 81228 1652
rect 81284 2100 81676 2156
rect 81060 1428 81228 1484
rect 80724 970 80780 980
rect 81172 924 81228 1428
rect 81284 1034 81340 2100
rect 81732 2044 81788 2054
rect 81620 1988 81732 2044
rect 81508 1036 81564 1046
rect 81284 982 81286 1034
rect 81338 982 81340 1034
rect 81284 970 81340 982
rect 81396 1034 81564 1036
rect 81396 982 81510 1034
rect 81562 982 81564 1034
rect 81396 980 81564 982
rect 81172 800 81228 868
rect 81396 924 81452 980
rect 81508 970 81564 980
rect 81396 858 81452 868
rect 81508 812 81564 822
rect 79044 410 79100 420
rect 79352 0 79464 800
rect 80024 0 80136 800
rect 80584 0 80696 800
rect 81144 0 81256 800
rect 81508 718 81564 756
rect 81620 588 81676 1988
rect 81732 1978 81788 1988
rect 81732 1146 81788 1158
rect 81732 1094 81734 1146
rect 81786 1094 81788 1146
rect 81732 924 81788 1094
rect 81732 858 81788 868
rect 81844 800 81900 2548
rect 82068 2492 82124 3108
rect 81956 2436 82124 2492
rect 82292 2938 82348 2950
rect 82292 2886 82294 2938
rect 82346 2886 82348 2938
rect 81956 2378 82012 2436
rect 82180 2380 82236 2390
rect 81956 2326 81958 2378
rect 82010 2326 82012 2378
rect 81956 2314 82012 2326
rect 82068 2378 82236 2380
rect 82068 2326 82182 2378
rect 82234 2326 82236 2378
rect 82068 2324 82236 2326
rect 82068 2268 82124 2324
rect 82180 2314 82236 2324
rect 82068 2202 82124 2212
rect 81956 1932 82012 1942
rect 81956 1146 82012 1876
rect 82292 1932 82348 2886
rect 82404 2828 82460 3110
rect 82516 2938 82572 3668
rect 82628 3500 82684 3510
rect 82628 3050 82684 3444
rect 82628 2998 82630 3050
rect 82682 2998 82684 3050
rect 82628 2986 82684 2998
rect 82740 3276 82796 3286
rect 82516 2886 82518 2938
rect 82570 2886 82572 2938
rect 82516 2874 82572 2886
rect 82404 2762 82460 2772
rect 82628 2828 82684 2838
rect 82292 1866 82348 1876
rect 82516 2156 82572 2166
rect 82516 1708 82572 2100
rect 82068 1652 82572 1708
rect 82068 1370 82124 1652
rect 82068 1318 82070 1370
rect 82122 1318 82124 1370
rect 82068 1306 82124 1318
rect 82404 1370 82460 1382
rect 82404 1318 82406 1370
rect 82458 1318 82460 1370
rect 81956 1094 81958 1146
rect 82010 1094 82012 1146
rect 81956 1082 82012 1094
rect 82068 810 82124 822
rect 81396 532 81676 588
rect 81396 474 81452 532
rect 81396 422 81398 474
rect 81450 422 81452 474
rect 81396 410 81452 422
rect 81816 0 81928 800
rect 82068 758 82070 810
rect 82122 758 82124 810
rect 82404 800 82460 1318
rect 82628 1372 82684 2772
rect 82628 1306 82684 1316
rect 82740 1370 82796 3220
rect 82964 3162 83020 4900
rect 82964 3110 82966 3162
rect 83018 3110 83020 3162
rect 82964 3098 83020 3110
rect 83076 4732 83132 4742
rect 83076 3722 83132 4676
rect 83300 4732 83356 4900
rect 83300 4666 83356 4676
rect 83412 4060 83468 5348
rect 83636 5292 83692 5852
rect 83524 5236 83692 5292
rect 83748 5852 83804 5862
rect 83860 5852 83916 6692
rect 84028 6682 84084 6692
rect 84084 6524 84140 6534
rect 84196 6524 84252 6804
rect 84140 6468 84252 6524
rect 84308 6636 84364 6646
rect 84084 6458 84140 6468
rect 83972 6188 84028 6198
rect 83972 6018 84028 6132
rect 83972 5966 83974 6018
rect 84026 5966 84028 6018
rect 83972 5954 84028 5966
rect 83860 5796 84140 5852
rect 83524 4284 83580 5236
rect 83524 4218 83580 4228
rect 83636 4956 83692 4966
rect 83412 4004 83580 4060
rect 83076 3670 83078 3722
rect 83130 3670 83132 3722
rect 82852 3050 82908 3062
rect 82852 2998 82854 3050
rect 82906 2998 82908 3050
rect 82852 1594 82908 2998
rect 82852 1542 82854 1594
rect 82906 1542 82908 1594
rect 82852 1530 82908 1542
rect 82740 1318 82742 1370
rect 82794 1318 82796 1370
rect 82740 1306 82796 1318
rect 82740 1034 82796 1046
rect 82740 982 82742 1034
rect 82794 982 82796 1034
rect 82740 810 82796 982
rect 82068 586 82124 758
rect 82068 534 82070 586
rect 82122 534 82124 586
rect 82068 522 82124 534
rect 82376 0 82488 800
rect 82740 758 82742 810
rect 82794 758 82796 810
rect 83076 800 83132 3670
rect 83188 3724 83244 3734
rect 83188 3162 83244 3668
rect 83188 3110 83190 3162
rect 83242 3110 83244 3162
rect 83188 3098 83244 3110
rect 83412 3722 83468 3734
rect 83412 3670 83414 3722
rect 83466 3670 83468 3722
rect 83412 1482 83468 3670
rect 83412 1430 83414 1482
rect 83466 1430 83468 1482
rect 83412 1418 83468 1430
rect 83524 1034 83580 4004
rect 83524 982 83526 1034
rect 83578 982 83580 1034
rect 83524 970 83580 982
rect 83636 800 83692 4900
rect 83748 3946 83804 5796
rect 83916 5516 83972 5526
rect 83916 4956 83972 5460
rect 83916 4954 84028 4956
rect 83916 4902 83918 4954
rect 83970 4902 84028 4954
rect 83916 4890 84028 4902
rect 83748 3894 83750 3946
rect 83802 3894 83804 3946
rect 83748 3882 83804 3894
rect 83972 2828 84028 4890
rect 84084 3946 84140 5796
rect 84084 3894 84086 3946
rect 84138 3894 84140 3946
rect 84084 3882 84140 3894
rect 84196 4060 84252 4070
rect 84308 4060 84364 6580
rect 84476 6522 84532 6534
rect 84476 6470 84478 6522
rect 84530 6470 84532 6522
rect 84476 6468 84532 6470
rect 84476 6412 84700 6468
rect 84476 5740 84532 5750
rect 84476 5516 84532 5684
rect 84476 4954 84532 5460
rect 84476 4902 84478 4954
rect 84530 4902 84532 4954
rect 84476 4890 84532 4902
rect 84644 4732 84700 6412
rect 84532 4676 84700 4732
rect 84420 4060 84476 4070
rect 84308 4004 84420 4060
rect 83972 2762 84028 2772
rect 83860 2268 83916 2278
rect 83860 2174 83916 2212
rect 84196 2266 84252 4004
rect 84420 3994 84476 4004
rect 84420 3498 84476 3510
rect 84420 3446 84422 3498
rect 84474 3446 84476 3498
rect 84196 2214 84198 2266
rect 84250 2214 84252 2266
rect 84196 2202 84252 2214
rect 84308 2938 84364 2950
rect 84308 2886 84310 2938
rect 84362 2886 84364 2938
rect 83748 2154 83804 2166
rect 83748 2102 83750 2154
rect 83802 2102 83804 2154
rect 83748 1596 83804 2102
rect 83972 2154 84028 2166
rect 83972 2102 83974 2154
rect 84026 2102 84028 2154
rect 83972 1820 84028 2102
rect 83972 1754 84028 1764
rect 83748 1540 84028 1596
rect 83972 1482 84028 1540
rect 83972 1430 83974 1482
rect 84026 1430 84028 1482
rect 83972 1418 84028 1430
rect 84084 1146 84140 1158
rect 84084 1094 84086 1146
rect 84138 1094 84140 1146
rect 83860 810 83916 822
rect 82740 746 82796 758
rect 83048 0 83160 800
rect 83608 0 83720 800
rect 83860 758 83862 810
rect 83914 758 83916 810
rect 83860 250 83916 758
rect 83860 198 83862 250
rect 83914 198 83916 250
rect 83860 186 83916 198
rect 84084 250 84140 1094
rect 84308 800 84364 2886
rect 84420 1932 84476 3446
rect 84532 3050 84588 4676
rect 84644 4396 84700 4406
rect 84644 3498 84700 4340
rect 84644 3446 84646 3498
rect 84698 3446 84700 3498
rect 84644 3434 84700 3446
rect 84532 2998 84534 3050
rect 84586 2998 84588 3050
rect 84532 2986 84588 2998
rect 84420 1866 84476 1876
rect 84756 1594 84812 7700
rect 85708 7690 85764 7700
rect 86100 7644 86156 8372
rect 84868 7586 84924 7598
rect 84868 7534 84870 7586
rect 84922 7534 84924 7586
rect 86100 7578 86156 7588
rect 84868 7308 84924 7534
rect 84868 7242 84924 7252
rect 84980 7474 85036 7486
rect 84980 7422 84982 7474
rect 85034 7422 85036 7474
rect 84980 7084 85036 7422
rect 85372 7418 85428 7430
rect 85372 7366 85374 7418
rect 85426 7366 85428 7418
rect 85372 7308 85428 7366
rect 85372 7242 85428 7252
rect 85988 7362 86044 7374
rect 85988 7310 85990 7362
rect 86042 7310 86044 7362
rect 84980 7018 85036 7028
rect 85764 7084 85820 7094
rect 85764 6747 85820 7028
rect 85764 6691 85876 6747
rect 85148 6580 85204 6590
rect 85092 6578 85204 6580
rect 85092 6526 85150 6578
rect 85202 6526 85204 6578
rect 85092 6514 85204 6526
rect 85260 6522 85316 6534
rect 84868 6188 84924 6198
rect 84868 5964 84924 6132
rect 84868 5898 84924 5908
rect 84924 5180 84980 5190
rect 84924 4956 84980 5124
rect 84924 4862 84980 4900
rect 85092 3050 85148 6514
rect 85260 6470 85262 6522
rect 85314 6470 85316 6522
rect 85260 6076 85316 6470
rect 85820 6522 85876 6691
rect 85820 6470 85822 6522
rect 85874 6470 85876 6522
rect 85820 6188 85876 6470
rect 85988 6300 86044 7310
rect 86212 6636 86268 6646
rect 86212 6534 86268 6580
rect 86156 6522 86268 6534
rect 86156 6470 86158 6522
rect 86210 6470 86268 6522
rect 86156 6458 86268 6470
rect 86212 6412 86268 6458
rect 86212 6346 86268 6356
rect 85988 6244 86156 6300
rect 85820 6132 86044 6188
rect 85204 6020 85316 6076
rect 85204 5628 85260 6020
rect 85540 5964 85596 5974
rect 85316 5908 85372 5918
rect 85316 5906 85484 5908
rect 85316 5854 85318 5906
rect 85370 5854 85484 5906
rect 85316 5852 85484 5854
rect 85316 5842 85372 5852
rect 85428 5786 85484 5796
rect 85204 5572 85484 5628
rect 85204 5404 85260 5414
rect 85204 5067 85260 5348
rect 85428 5404 85484 5572
rect 85428 5338 85484 5348
rect 85540 5067 85596 5908
rect 85820 5852 85876 5862
rect 85820 5758 85876 5796
rect 85204 5011 85372 5067
rect 85092 2998 85094 3050
rect 85146 2998 85148 3050
rect 84868 2604 84924 2614
rect 84868 2156 84924 2548
rect 84868 2090 84924 2100
rect 84756 1542 84758 1594
rect 84810 1542 84812 1594
rect 84756 1530 84812 1542
rect 85092 1594 85148 2998
rect 85204 3274 85260 3286
rect 85204 3222 85206 3274
rect 85258 3222 85260 3274
rect 85204 2828 85260 3222
rect 85316 3050 85372 5011
rect 85428 5011 85596 5067
rect 85652 5124 85932 5180
rect 85428 4732 85484 5011
rect 85428 4666 85484 4676
rect 85652 4620 85708 5124
rect 85652 4554 85708 4564
rect 85764 5010 85820 5022
rect 85764 4958 85766 5010
rect 85818 4958 85820 5010
rect 85652 4058 85708 4070
rect 85652 4006 85654 4058
rect 85706 4006 85708 4058
rect 85652 3836 85708 4006
rect 85652 3770 85708 3780
rect 85428 3610 85484 3622
rect 85428 3558 85430 3610
rect 85482 3558 85484 3610
rect 85428 3274 85484 3558
rect 85428 3222 85430 3274
rect 85482 3222 85484 3274
rect 85428 3210 85484 3222
rect 85316 2998 85318 3050
rect 85370 2998 85372 3050
rect 85316 2986 85372 2998
rect 85652 3052 85708 3062
rect 85652 2828 85708 2996
rect 85204 2772 85708 2828
rect 85764 2716 85820 4958
rect 85876 4732 85932 5124
rect 85988 4956 86044 6132
rect 85988 4890 86044 4900
rect 86100 4732 86156 6244
rect 86324 6188 86380 8708
rect 86436 8540 86492 8550
rect 86436 7644 86492 8484
rect 86548 8204 86604 8932
rect 87052 8922 87108 8932
rect 87220 8204 87276 9156
rect 86548 8202 86828 8204
rect 86548 8150 86550 8202
rect 86602 8150 86828 8202
rect 86548 8148 86828 8150
rect 86548 8138 86604 8148
rect 86436 7578 86492 7588
rect 86548 7980 86604 7990
rect 86212 6132 86380 6188
rect 86212 4844 86268 6132
rect 86212 4788 86492 4844
rect 85876 4676 86156 4732
rect 86212 4620 86268 4630
rect 85988 4396 86044 4406
rect 85876 4060 85932 4070
rect 85876 3966 85932 4004
rect 85764 2650 85820 2660
rect 85988 2716 86044 4340
rect 86212 3610 86268 4564
rect 86436 4060 86492 4788
rect 86548 4620 86604 7924
rect 86660 6690 86716 6702
rect 86660 6638 86662 6690
rect 86714 6638 86716 6690
rect 86660 5068 86716 6638
rect 86660 5002 86716 5012
rect 86548 4554 86604 4564
rect 86436 3994 86492 4004
rect 86548 4396 86604 4406
rect 86548 3836 86604 4340
rect 86548 3770 86604 3780
rect 86212 3558 86214 3610
rect 86266 3558 86268 3610
rect 86212 3546 86268 3558
rect 85988 2650 86044 2660
rect 85988 2268 86044 2278
rect 85988 2156 86044 2212
rect 85540 2100 86044 2156
rect 86100 2156 86156 2166
rect 85540 1932 85596 2100
rect 85092 1542 85094 1594
rect 85146 1542 85148 1594
rect 85092 1530 85148 1542
rect 85316 1876 85596 1932
rect 84420 1370 84476 1382
rect 84420 1318 84422 1370
rect 84474 1318 84476 1370
rect 84420 1036 84476 1318
rect 84420 970 84476 980
rect 84868 1034 84924 1046
rect 84868 982 84870 1034
rect 84922 982 84924 1034
rect 84868 800 84924 982
rect 84084 198 84086 250
rect 84138 198 84140 250
rect 84084 186 84140 198
rect 84280 0 84392 800
rect 84840 0 84952 800
rect 85316 698 85372 1876
rect 85428 1708 85484 1718
rect 85428 1146 85484 1652
rect 85652 1708 85708 1718
rect 85652 1372 85708 1652
rect 85652 1306 85708 1316
rect 85428 1094 85430 1146
rect 85482 1094 85484 1146
rect 85428 1082 85484 1094
rect 85540 1036 85596 1046
rect 85540 800 85596 980
rect 85764 810 85820 822
rect 85316 646 85318 698
rect 85370 646 85372 698
rect 85316 634 85372 646
rect 85512 0 85624 800
rect 85764 758 85766 810
rect 85818 758 85820 810
rect 86100 800 86156 2100
rect 86772 1148 86828 8148
rect 87108 8148 87276 8204
rect 86884 8092 86940 8102
rect 86884 8090 87052 8092
rect 86884 8038 86886 8090
rect 86938 8038 87052 8090
rect 86884 8036 87052 8038
rect 86884 8026 86940 8036
rect 86996 6860 87052 8036
rect 86884 6804 87052 6860
rect 86884 4060 86940 6804
rect 86996 6188 87052 6198
rect 86996 5852 87052 6132
rect 86996 5786 87052 5796
rect 87108 5628 87164 8148
rect 87220 7586 87276 7598
rect 87220 7534 87222 7586
rect 87274 7534 87276 7586
rect 87220 5852 87276 7534
rect 87332 6188 87388 9604
rect 87556 9548 87612 9558
rect 87444 9212 87500 9222
rect 87444 7474 87500 9156
rect 87556 8428 87612 9492
rect 87780 9222 87836 12516
rect 87892 12570 87948 12582
rect 87892 12518 87894 12570
rect 87946 12518 87948 12570
rect 87892 9548 87948 12518
rect 88676 9660 88732 12854
rect 89124 12348 89180 14200
rect 89460 13020 89516 13030
rect 89460 12906 89516 12964
rect 89460 12854 89462 12906
rect 89514 12854 89516 12906
rect 89460 12842 89516 12854
rect 89796 12906 89852 12918
rect 89796 12854 89798 12906
rect 89850 12854 89852 12906
rect 89796 12458 89852 12854
rect 89796 12406 89798 12458
rect 89850 12406 89852 12458
rect 89796 12394 89852 12406
rect 89124 12282 89180 12292
rect 88788 12236 88844 12246
rect 88844 12180 88956 12236
rect 88788 12170 88844 12180
rect 88788 11452 88844 11462
rect 88788 11226 88844 11396
rect 88788 11174 88790 11226
rect 88842 11174 88844 11226
rect 88788 11162 88844 11174
rect 88900 10332 88956 12180
rect 89908 12124 89964 14200
rect 89908 12058 89964 12068
rect 90020 14026 90076 14038
rect 90020 13974 90022 14026
rect 90074 13974 90076 14026
rect 89012 12012 89068 12022
rect 89012 11226 89068 11956
rect 89012 11174 89014 11226
rect 89066 11174 89068 11226
rect 89012 11162 89068 11174
rect 89348 11340 89404 11350
rect 89348 10442 89404 11284
rect 89348 10390 89350 10442
rect 89402 10390 89404 10442
rect 89348 10378 89404 10390
rect 89572 11002 89628 11014
rect 89572 10950 89574 11002
rect 89626 10950 89628 11002
rect 89572 10442 89628 10950
rect 90020 11002 90076 13974
rect 90132 13578 90188 13590
rect 90132 13526 90134 13578
rect 90186 13526 90188 13578
rect 90132 12234 90188 13526
rect 90356 13578 90412 13590
rect 90356 13526 90358 13578
rect 90410 13526 90412 13578
rect 90244 13466 90300 13478
rect 90244 13414 90246 13466
rect 90298 13414 90300 13466
rect 90244 12346 90300 13414
rect 90356 13468 90412 13526
rect 90356 13402 90412 13412
rect 90244 12294 90246 12346
rect 90298 12294 90300 12346
rect 90244 12282 90300 12294
rect 90132 12182 90134 12234
rect 90186 12182 90188 12234
rect 90132 12170 90188 12182
rect 90580 11562 90636 14200
rect 90804 13466 90860 14646
rect 91028 14698 91084 14710
rect 91028 14646 91030 14698
rect 91082 14646 91084 14698
rect 91028 14138 91084 14646
rect 91336 14200 91448 15000
rect 91588 14362 91644 14374
rect 91588 14310 91590 14362
rect 91642 14310 91644 14362
rect 91364 14140 91420 14200
rect 91028 14086 91030 14138
rect 91082 14086 91084 14138
rect 91028 14074 91084 14086
rect 91308 14084 91420 14140
rect 91308 14028 91364 14084
rect 91140 13972 91364 14028
rect 91588 14026 91644 14310
rect 92008 14200 92120 15000
rect 92792 14200 92904 15000
rect 93464 14200 93576 15000
rect 94248 14200 94360 15000
rect 94920 14200 95032 15000
rect 95704 14200 95816 15000
rect 96376 14200 96488 15000
rect 97160 14200 97272 15000
rect 97832 14200 97944 15000
rect 98084 14812 98140 14822
rect 91588 13974 91590 14026
rect 91642 13974 91644 14026
rect 91028 13804 91084 13814
rect 91028 13578 91084 13748
rect 91028 13526 91030 13578
rect 91082 13526 91084 13578
rect 91028 13514 91084 13526
rect 90804 13414 90806 13466
rect 90858 13414 90860 13466
rect 90804 13402 90860 13414
rect 90580 11510 90582 11562
rect 90634 11510 90636 11562
rect 90580 11498 90636 11510
rect 90804 11562 90860 11574
rect 90804 11510 90806 11562
rect 90858 11510 90860 11562
rect 90020 10950 90022 11002
rect 90074 10950 90076 11002
rect 90020 10938 90076 10950
rect 89572 10390 89574 10442
rect 89626 10390 89628 10442
rect 89572 10378 89628 10390
rect 88900 10276 89292 10332
rect 88676 9594 88732 9604
rect 88900 9996 88956 10006
rect 88900 9660 88956 9940
rect 88900 9594 88956 9604
rect 87892 9482 87948 9492
rect 87724 9212 87836 9222
rect 87780 9156 87836 9212
rect 87724 9080 87780 9156
rect 88396 9042 88452 9054
rect 88396 8990 88398 9042
rect 88450 8990 88452 9042
rect 88396 8988 88452 8990
rect 89068 8988 89124 8998
rect 88396 8986 89124 8988
rect 88396 8934 89070 8986
rect 89122 8934 89124 8986
rect 88396 8932 89124 8934
rect 89236 8988 89292 10276
rect 90692 9884 90748 9894
rect 90692 9210 90748 9828
rect 90692 9158 90694 9210
rect 90746 9158 90748 9210
rect 90692 9146 90748 9158
rect 90356 9098 90412 9110
rect 90356 9046 90358 9098
rect 90410 9046 90412 9098
rect 89740 8988 89796 8998
rect 90356 8988 90412 9046
rect 89236 8986 90412 8988
rect 89236 8934 89742 8986
rect 89794 8934 90412 8986
rect 89236 8932 90412 8934
rect 88116 8876 88172 8886
rect 88284 8876 88340 8886
rect 88172 8874 88340 8876
rect 88172 8822 88286 8874
rect 88338 8822 88340 8874
rect 88172 8820 88340 8822
rect 88116 8810 88172 8820
rect 88284 8810 88340 8820
rect 88900 8652 88956 8662
rect 88452 8596 88900 8652
rect 88452 8540 88508 8596
rect 88900 8586 88956 8596
rect 88452 8474 88508 8484
rect 87724 8428 87780 8438
rect 87556 8426 87780 8428
rect 87556 8374 87726 8426
rect 87778 8374 87780 8426
rect 87556 8372 87780 8374
rect 87724 8362 87780 8372
rect 89068 8372 89124 8932
rect 89684 8922 89796 8932
rect 88508 8316 88564 8326
rect 89068 8316 89404 8372
rect 88508 8258 88564 8260
rect 87444 7422 87446 7474
rect 87498 7422 87500 7474
rect 87444 7410 87500 7422
rect 87556 8204 87612 8214
rect 88508 8206 88510 8258
rect 88562 8206 88564 8258
rect 87556 7980 87612 8148
rect 87836 8146 87892 8158
rect 87332 6122 87388 6132
rect 87556 5908 87612 7924
rect 87668 8092 87724 8102
rect 87668 6972 87724 8036
rect 87836 8094 87838 8146
rect 87890 8094 87892 8146
rect 87836 7644 87892 8094
rect 88396 8090 88452 8102
rect 88396 8038 88398 8090
rect 88450 8038 88452 8090
rect 88396 7868 88452 8038
rect 88396 7802 88452 7812
rect 88004 7756 88060 7766
rect 88060 7700 88172 7756
rect 88004 7690 88060 7700
rect 87836 7588 87948 7644
rect 87892 7430 87948 7588
rect 88116 7532 88172 7700
rect 88508 7642 88564 8206
rect 89068 8090 89124 8102
rect 89068 8038 89070 8090
rect 89122 8038 89124 8090
rect 89068 7980 89124 8038
rect 89068 7914 89124 7924
rect 89236 8092 89292 8102
rect 88508 7590 88510 7642
rect 88562 7590 88564 7642
rect 88508 7578 88564 7590
rect 88676 7644 88732 7654
rect 88116 7466 88172 7476
rect 87892 7420 88004 7430
rect 87892 7418 88060 7420
rect 87892 7366 87950 7418
rect 88002 7366 88060 7418
rect 87892 7364 88060 7366
rect 87948 7354 88060 7364
rect 87668 6906 87724 6916
rect 87780 7084 87836 7094
rect 87780 6748 87836 7028
rect 87668 6690 87724 6702
rect 87668 6638 87670 6690
rect 87722 6638 87724 6690
rect 87780 6682 87836 6692
rect 87668 6636 87724 6638
rect 87668 6570 87724 6580
rect 88004 6636 88060 7354
rect 88676 7308 88732 7588
rect 89236 7532 89292 8036
rect 88004 6570 88060 6580
rect 88116 7252 88732 7308
rect 88788 7476 89292 7532
rect 87220 5786 87276 5796
rect 87332 5852 87612 5908
rect 87948 5852 88004 5862
rect 87108 5572 87276 5628
rect 87108 5122 87164 5134
rect 87108 5070 87110 5122
rect 87162 5070 87164 5122
rect 87108 5068 87164 5070
rect 87108 5002 87164 5012
rect 86884 3994 86940 4004
rect 86996 4620 87052 4630
rect 86884 3836 86940 3846
rect 86884 1708 86940 3780
rect 86884 1642 86940 1652
rect 86660 1146 86828 1148
rect 86660 1094 86774 1146
rect 86826 1094 86828 1146
rect 86660 1092 86828 1094
rect 86660 800 86716 1092
rect 86772 1082 86828 1092
rect 86996 1034 87052 4564
rect 87108 2716 87164 2726
rect 87108 2492 87164 2660
rect 87108 2426 87164 2436
rect 87220 1146 87276 5572
rect 87220 1094 87222 1146
rect 87274 1094 87276 1146
rect 87220 1082 87276 1094
rect 86996 982 86998 1034
rect 87050 982 87052 1034
rect 86996 970 87052 982
rect 87332 800 87388 5852
rect 87948 5758 88004 5796
rect 87780 5740 87836 5750
rect 87780 2940 87836 5684
rect 87948 5068 88004 5078
rect 87948 4956 88004 5012
rect 88116 4956 88172 7252
rect 88340 6972 88396 6982
rect 88788 6972 88844 7476
rect 88396 6916 88844 6972
rect 89124 7362 89180 7374
rect 89124 7310 89126 7362
rect 89178 7310 89180 7362
rect 89124 6972 89180 7310
rect 88340 6906 88396 6916
rect 89124 6906 89180 6916
rect 88564 5852 88620 5862
rect 88788 5852 88844 5862
rect 88564 5404 88620 5796
rect 88564 5338 88620 5348
rect 88676 5796 88788 5852
rect 87948 4954 88172 4956
rect 87948 4902 87950 4954
rect 88002 4902 88172 4954
rect 87948 4900 88172 4902
rect 88228 5068 88284 5078
rect 87948 4890 88004 4900
rect 87892 2940 87948 2950
rect 87780 2884 87892 2940
rect 87892 2874 87948 2884
rect 87444 1148 87500 1158
rect 87444 1054 87500 1092
rect 87892 1146 87948 1158
rect 87892 1094 87894 1146
rect 87946 1094 87948 1146
rect 87892 800 87948 1094
rect 88228 922 88284 5012
rect 88340 4060 88396 4070
rect 88676 4060 88732 5796
rect 88788 5786 88844 5796
rect 88340 1708 88396 4004
rect 88452 4004 88732 4060
rect 89236 5010 89292 5022
rect 89236 4958 89238 5010
rect 89290 4958 89292 5010
rect 89236 4058 89292 4958
rect 89236 4006 89238 4058
rect 89290 4006 89292 4058
rect 88452 1820 88508 4004
rect 89236 3994 89292 4006
rect 89348 4060 89404 8316
rect 89572 8090 89628 8102
rect 89572 8038 89574 8090
rect 89626 8038 89628 8090
rect 89572 7980 89628 8038
rect 89572 7914 89628 7924
rect 89460 6522 89516 6534
rect 89460 6470 89462 6522
rect 89514 6470 89516 6522
rect 89460 5852 89516 6470
rect 89460 5786 89516 5796
rect 89572 4956 89628 4966
rect 89460 4060 89516 4070
rect 89348 4058 89516 4060
rect 89348 4006 89462 4058
rect 89514 4006 89516 4058
rect 89348 4004 89516 4006
rect 89460 3994 89516 4004
rect 88452 1754 88508 1764
rect 88564 3836 88620 3846
rect 88340 1642 88396 1652
rect 88228 870 88230 922
rect 88282 870 88284 922
rect 88228 858 88284 870
rect 88452 1594 88508 1606
rect 88452 1542 88454 1594
rect 88506 1542 88508 1594
rect 88452 922 88508 1542
rect 88452 870 88454 922
rect 88506 870 88508 922
rect 88452 858 88508 870
rect 88564 800 88620 3780
rect 89236 3610 89292 3622
rect 89236 3558 89238 3610
rect 89290 3558 89292 3610
rect 88676 2828 88732 2838
rect 88732 2772 89068 2828
rect 88676 2762 88732 2772
rect 88788 2268 88844 2278
rect 88788 1594 88844 2212
rect 88788 1542 88790 1594
rect 88842 1542 88844 1594
rect 88788 1530 88844 1542
rect 88900 2042 88956 2054
rect 88900 1990 88902 2042
rect 88954 1990 88956 2042
rect 88900 1484 88956 1990
rect 88900 1418 88956 1428
rect 89012 1372 89068 2772
rect 89236 2268 89292 3558
rect 89572 3610 89628 4900
rect 89572 3558 89574 3610
rect 89626 3558 89628 3610
rect 89572 3546 89628 3558
rect 89236 2202 89292 2212
rect 89012 1306 89068 1316
rect 89124 2042 89180 2054
rect 89124 1990 89126 2042
rect 89178 1990 89180 2042
rect 89124 800 89180 1990
rect 89684 1146 89740 8922
rect 90412 8764 90468 8774
rect 90412 8426 90468 8708
rect 90412 8374 90414 8426
rect 90466 8374 90468 8426
rect 90412 8362 90468 8374
rect 89908 8316 89964 8326
rect 89908 8222 89964 8260
rect 90356 8204 90412 8214
rect 90244 8092 90412 8148
rect 90524 8146 90580 8158
rect 90524 8094 90526 8146
rect 90578 8094 90580 8146
rect 90244 6412 90300 8092
rect 90356 7756 90412 7766
rect 90356 7586 90412 7700
rect 90524 7644 90580 8094
rect 90804 7980 90860 11510
rect 91140 10668 91196 13972
rect 91588 13962 91644 13974
rect 91476 13020 91532 13030
rect 91476 12796 91532 12964
rect 91476 12730 91532 12740
rect 91924 12572 91980 12582
rect 91364 12122 91420 12134
rect 91364 12070 91366 12122
rect 91418 12070 91420 12122
rect 91364 11900 91420 12070
rect 91700 11900 91756 11910
rect 91364 11898 91756 11900
rect 91364 11846 91702 11898
rect 91754 11846 91756 11898
rect 91364 11844 91756 11846
rect 91700 11834 91756 11844
rect 91924 11562 91980 12516
rect 91924 11510 91926 11562
rect 91978 11510 91980 11562
rect 91924 11498 91980 11510
rect 92036 11452 92092 14200
rect 92708 14138 92764 14150
rect 92708 14086 92710 14138
rect 92762 14086 92764 14138
rect 92708 13916 92764 14086
rect 92708 13850 92764 13860
rect 92036 11386 92092 11396
rect 91476 11340 91532 11350
rect 91140 10602 91196 10612
rect 91364 10892 91420 10902
rect 91364 10668 91420 10836
rect 91364 10602 91420 10612
rect 91476 10220 91532 11284
rect 92820 11116 92876 14200
rect 92932 14138 92988 14150
rect 92932 14086 92934 14138
rect 92986 14086 92988 14138
rect 92932 12572 92988 14086
rect 92932 12506 92988 12516
rect 93492 12348 93548 14200
rect 93492 12282 93548 12292
rect 94164 12348 94220 12358
rect 93828 11900 93884 11910
rect 92932 11786 92988 11798
rect 92932 11734 92934 11786
rect 92986 11734 92988 11786
rect 92932 11562 92988 11734
rect 92932 11510 92934 11562
rect 92986 11510 92988 11562
rect 92932 11498 92988 11510
rect 93156 11786 93212 11798
rect 93156 11734 93158 11786
rect 93210 11734 93212 11786
rect 92820 11050 92876 11060
rect 93044 11116 93100 11126
rect 91812 10780 91868 10790
rect 93044 10780 93100 11060
rect 91868 10724 93100 10780
rect 91812 10714 91868 10724
rect 91476 10154 91532 10164
rect 91252 9772 91308 9782
rect 91252 9548 91308 9716
rect 91252 9482 91308 9492
rect 91700 9548 91756 9558
rect 91700 9436 91756 9492
rect 91700 9380 92260 9436
rect 92204 9212 92260 9380
rect 92820 9212 92876 9222
rect 92204 9210 92876 9212
rect 92204 9158 92206 9210
rect 92258 9158 92822 9210
rect 92874 9158 92876 9210
rect 92204 9156 92876 9158
rect 92204 9146 92260 9156
rect 92820 9146 92876 9156
rect 91308 9042 91364 9054
rect 91308 8990 91310 9042
rect 91362 8990 91364 9042
rect 91308 8988 91364 8990
rect 91756 8988 91812 8998
rect 91308 8986 91812 8988
rect 91308 8934 91758 8986
rect 91810 8934 91812 8986
rect 91308 8932 91812 8934
rect 91196 8874 91252 8886
rect 91196 8822 91198 8874
rect 91250 8822 91252 8874
rect 91196 8540 91252 8822
rect 91196 8474 91252 8484
rect 91756 8427 91812 8932
rect 91756 8371 92204 8427
rect 91196 8204 91252 8214
rect 91644 8204 91700 8214
rect 91196 8202 91868 8204
rect 91196 8150 91198 8202
rect 91250 8150 91646 8202
rect 91698 8150 91868 8202
rect 91196 8148 91868 8150
rect 91196 8138 91252 8148
rect 91644 8138 91700 8148
rect 91084 8092 91140 8102
rect 91084 7998 91140 8036
rect 90804 7914 90860 7924
rect 91532 7756 91588 7766
rect 91812 7756 91868 8148
rect 91812 7700 91980 7756
rect 90524 7588 90748 7644
rect 90356 7534 90358 7586
rect 90410 7534 90412 7586
rect 90356 7522 90412 7534
rect 90580 7474 90636 7486
rect 90580 7422 90582 7474
rect 90634 7422 90636 7474
rect 90468 7308 90524 7318
rect 90468 6524 90524 7252
rect 90468 6458 90524 6468
rect 90244 6346 90300 6356
rect 90580 6412 90636 7422
rect 90692 7420 90748 7588
rect 91252 7532 91308 7542
rect 91084 7420 91140 7430
rect 90692 7418 91140 7420
rect 90692 7366 91086 7418
rect 91138 7366 91140 7418
rect 90692 7364 91140 7366
rect 91028 7354 91140 7364
rect 90580 6346 90636 6356
rect 90748 6972 90804 6982
rect 90748 6690 90804 6916
rect 90748 6638 90750 6690
rect 90802 6638 90804 6690
rect 90748 5964 90804 6638
rect 90860 6636 90916 6646
rect 90860 6542 90916 6580
rect 90748 5908 90972 5964
rect 89908 5180 89964 5190
rect 89908 4956 89964 5124
rect 90580 5180 90636 5190
rect 90580 5122 90636 5124
rect 90580 5070 90582 5122
rect 90634 5070 90636 5122
rect 90580 5058 90636 5070
rect 89684 1094 89686 1146
rect 89738 1094 89740 1146
rect 89684 1082 89740 1094
rect 89796 3276 89852 3286
rect 89796 1372 89852 3220
rect 89908 2042 89964 4900
rect 90916 4508 90972 5908
rect 91028 4732 91084 7354
rect 91252 7196 91308 7476
rect 91532 7420 91588 7700
rect 91532 7418 91644 7420
rect 91532 7366 91534 7418
rect 91586 7366 91644 7418
rect 91532 7354 91644 7366
rect 91476 7196 91532 7206
rect 91252 7130 91308 7140
rect 91364 7140 91476 7196
rect 91252 6972 91308 6982
rect 91364 6972 91420 7140
rect 91476 7130 91532 7140
rect 91308 6916 91420 6972
rect 91476 6972 91532 6982
rect 91252 6906 91308 6916
rect 91364 6748 91420 6758
rect 91476 6748 91532 6916
rect 91420 6692 91532 6748
rect 91364 6682 91420 6692
rect 91420 6522 91476 6534
rect 91420 6470 91422 6522
rect 91474 6470 91476 6522
rect 91420 6412 91476 6470
rect 91420 6346 91476 6356
rect 91196 5740 91252 5750
rect 91196 5180 91252 5684
rect 91196 5048 91252 5124
rect 91364 5180 91420 5190
rect 91028 4666 91084 4676
rect 91252 4508 91308 4518
rect 91364 4508 91420 5124
rect 90916 4452 91084 4508
rect 90020 4396 90076 4406
rect 90020 4172 90076 4340
rect 90020 4106 90076 4116
rect 90916 3162 90972 3174
rect 90916 3110 90918 3162
rect 90970 3110 90972 3162
rect 90580 3052 90636 3062
rect 90132 2996 90580 3052
rect 90132 2380 90188 2996
rect 90580 2986 90636 2996
rect 90132 2314 90188 2324
rect 90692 2938 90748 2950
rect 90692 2886 90694 2938
rect 90746 2886 90748 2938
rect 89908 1990 89910 2042
rect 89962 1990 89964 2042
rect 89908 1978 89964 1990
rect 90692 2042 90748 2886
rect 90916 2938 90972 3110
rect 90916 2886 90918 2938
rect 90970 2886 90972 2938
rect 90916 2874 90972 2886
rect 90692 1990 90694 2042
rect 90746 1990 90748 2042
rect 90692 1978 90748 1990
rect 89796 800 89852 1316
rect 90580 1372 90636 1382
rect 90580 1278 90636 1316
rect 89908 1260 89964 1270
rect 89908 1146 89964 1204
rect 89908 1094 89910 1146
rect 89962 1094 89964 1146
rect 89908 1082 89964 1094
rect 90356 922 90412 934
rect 90356 870 90358 922
rect 90410 870 90412 922
rect 90356 800 90412 870
rect 91028 800 91084 4452
rect 91308 4452 91420 4508
rect 91252 4442 91308 4452
rect 91588 4396 91644 7354
rect 91756 7196 91812 7206
rect 91756 6746 91812 7140
rect 91756 6694 91758 6746
rect 91810 6694 91812 6746
rect 91756 6682 91812 6694
rect 91924 4956 91980 7700
rect 91924 4890 91980 4900
rect 91700 4396 91756 4406
rect 91588 4340 91700 4396
rect 91700 4330 91756 4340
rect 92148 4284 92204 8371
rect 92820 7470 92876 7482
rect 92428 7420 92484 7430
rect 92372 7418 92484 7420
rect 92372 7366 92430 7418
rect 92482 7366 92484 7418
rect 92372 7354 92484 7366
rect 92820 7418 92822 7470
rect 92874 7418 92876 7470
rect 92372 6188 92428 7354
rect 92820 6524 92876 7418
rect 92820 6458 92876 6468
rect 92372 6122 92428 6132
rect 92148 4218 92204 4228
rect 92820 5010 92876 5022
rect 92820 4958 92822 5010
rect 92874 4958 92876 5010
rect 91364 4116 91980 4172
rect 91252 4058 91308 4070
rect 91252 4006 91254 4058
rect 91306 4006 91308 4058
rect 91252 1370 91308 4006
rect 91364 3500 91420 4116
rect 91700 3946 91756 3958
rect 91700 3894 91702 3946
rect 91754 3894 91756 3946
rect 91364 3434 91420 3444
rect 91588 3836 91644 3846
rect 91476 3164 91532 3174
rect 91476 3070 91532 3108
rect 91252 1318 91254 1370
rect 91306 1318 91308 1370
rect 91252 1306 91308 1318
rect 91588 800 91644 3780
rect 91700 3386 91756 3894
rect 91700 3334 91702 3386
rect 91754 3334 91756 3386
rect 91700 3322 91756 3334
rect 91924 3386 91980 4116
rect 92820 3498 92876 4958
rect 92820 3446 92822 3498
rect 92874 3446 92876 3498
rect 92820 3434 92876 3446
rect 91924 3334 91926 3386
rect 91978 3334 91980 3386
rect 91924 3322 91980 3334
rect 92036 3388 92092 3398
rect 92092 3332 92204 3387
rect 92036 3331 92204 3332
rect 92036 3322 92092 3331
rect 91924 3052 91980 3062
rect 91924 2958 91980 2996
rect 92148 3050 92204 3331
rect 93044 3276 93100 10724
rect 93156 9210 93212 11734
rect 93156 9158 93158 9210
rect 93210 9158 93212 9210
rect 93156 9146 93212 9158
rect 93268 8540 93324 8550
rect 93268 8092 93324 8484
rect 93828 8372 93884 11844
rect 93940 8876 93996 8886
rect 94164 8876 94220 12292
rect 94276 10108 94332 14200
rect 94948 11788 95004 14200
rect 94836 11732 95004 11788
rect 94276 10042 94332 10052
rect 94724 11562 94780 11574
rect 94724 11510 94726 11562
rect 94778 11510 94780 11562
rect 93996 8820 94220 8876
rect 93940 8810 93996 8820
rect 93940 8372 93996 8382
rect 93828 8370 93996 8372
rect 93828 8318 93942 8370
rect 93994 8318 93996 8370
rect 93828 8316 93996 8318
rect 93940 8306 93996 8316
rect 92148 2998 92150 3050
rect 92202 2998 92204 3050
rect 92148 2986 92204 2998
rect 92820 3220 93100 3276
rect 93156 3498 93212 3510
rect 93156 3446 93158 3498
rect 93210 3446 93212 3498
rect 93156 3274 93212 3446
rect 93156 3222 93158 3274
rect 93210 3222 93212 3274
rect 92148 2156 92204 2166
rect 92148 1594 92204 2100
rect 92148 1542 92150 1594
rect 92202 1542 92204 1594
rect 92148 1530 92204 1542
rect 92372 1594 92428 1606
rect 92372 1542 92374 1594
rect 92426 1542 92428 1594
rect 92372 1148 92428 1542
rect 92372 1082 92428 1092
rect 92148 1034 92204 1046
rect 92148 982 92150 1034
rect 92202 982 92204 1034
rect 92148 800 92204 982
rect 92820 800 92876 3220
rect 93156 3210 93212 3222
rect 93268 1596 93324 8036
rect 93828 7474 93884 7486
rect 93828 7422 93830 7474
rect 93882 7422 93884 7474
rect 93828 6188 93884 7422
rect 93828 6122 93884 6132
rect 93940 5404 93996 5414
rect 93940 5122 93996 5348
rect 93940 5070 93942 5122
rect 93994 5070 93996 5122
rect 93940 5058 93996 5070
rect 93380 4620 93436 4630
rect 93380 1820 93436 4564
rect 94164 3836 94220 8820
rect 94724 8204 94780 11510
rect 94836 10332 94892 11732
rect 94836 10266 94892 10276
rect 94948 11562 95004 11574
rect 94948 11510 94950 11562
rect 95002 11510 95004 11562
rect 94948 9222 95004 11510
rect 94892 9212 95004 9222
rect 94836 9210 95004 9212
rect 94836 9158 94894 9210
rect 94946 9158 95004 9210
rect 94836 9156 95004 9158
rect 94836 9146 94948 9156
rect 94836 8258 94892 9146
rect 95340 8988 95396 8998
rect 94836 8206 94838 8258
rect 94890 8206 94892 8258
rect 94836 8194 94892 8206
rect 95284 8932 95340 8988
rect 95284 8856 95396 8932
rect 94724 8138 94780 8148
rect 95172 5628 95228 5638
rect 94780 5404 94836 5414
rect 94780 5178 94836 5348
rect 94780 5126 94782 5178
rect 94834 5126 94836 5178
rect 94780 5114 94836 5126
rect 95172 4060 95228 5572
rect 95284 5292 95340 8856
rect 95732 8316 95788 14200
rect 96012 9660 96068 9670
rect 96012 9658 96124 9660
rect 96012 9606 96014 9658
rect 96066 9606 96124 9658
rect 96012 9594 96124 9606
rect 95956 9098 96012 9110
rect 95956 9046 95958 9098
rect 96010 9046 96012 9098
rect 95956 8988 96012 9046
rect 95956 8922 96012 8932
rect 95732 8260 95900 8316
rect 95396 8146 95452 8158
rect 95396 8094 95398 8146
rect 95450 8094 95452 8146
rect 95396 7980 95452 8094
rect 95396 7914 95452 7924
rect 95732 8092 95788 8102
rect 95620 7644 95676 7654
rect 95620 7550 95676 7588
rect 95284 5226 95340 5236
rect 95172 3994 95228 4004
rect 95284 4284 95340 4294
rect 94052 3780 94220 3836
rect 94052 2492 94108 3780
rect 94388 3386 94444 3398
rect 94388 3334 94390 3386
rect 94442 3334 94444 3386
rect 94164 3274 94220 3286
rect 94164 3222 94166 3274
rect 94218 3222 94220 3274
rect 94164 3052 94220 3222
rect 94164 2986 94220 2996
rect 94388 3052 94444 3334
rect 94388 2986 94444 2996
rect 93828 2436 94108 2492
rect 93828 1932 93884 2436
rect 94164 2380 94220 2390
rect 94164 2286 94220 2324
rect 93940 2266 93996 2278
rect 93940 2214 93942 2266
rect 93994 2214 93996 2266
rect 93940 2044 93996 2214
rect 94612 2156 94668 2166
rect 94500 2044 94556 2054
rect 93940 2042 94556 2044
rect 93940 1990 94502 2042
rect 94554 1990 94556 2042
rect 93940 1988 94556 1990
rect 94500 1978 94556 1988
rect 93828 1876 94108 1932
rect 93380 1754 93436 1764
rect 93268 1540 93436 1596
rect 93380 800 93436 1540
rect 94052 800 94108 1876
rect 94612 1370 94668 2100
rect 94612 1318 94614 1370
rect 94666 1318 94668 1370
rect 94612 800 94668 1318
rect 95284 800 95340 4228
rect 95732 3274 95788 8036
rect 95732 3222 95734 3274
rect 95786 3222 95788 3274
rect 95732 3210 95788 3222
rect 95732 2268 95788 2278
rect 95732 2174 95788 2212
rect 95844 2154 95900 8260
rect 96068 7980 96124 9594
rect 96292 8874 96348 8886
rect 96292 8822 96294 8874
rect 96346 8822 96348 8874
rect 96292 8540 96348 8822
rect 96292 8474 96348 8484
rect 96236 8092 96292 8102
rect 96068 7914 96124 7924
rect 96180 8090 96292 8092
rect 96180 8038 96238 8090
rect 96290 8038 96292 8090
rect 96180 8026 96292 8038
rect 96404 8092 96460 14200
rect 97076 12572 97132 12582
rect 96628 12516 97076 12572
rect 96628 10780 96684 12516
rect 97076 12506 97132 12516
rect 97188 12348 97244 14200
rect 97524 14138 97580 14150
rect 97524 14086 97526 14138
rect 97578 14086 97580 14138
rect 97524 14028 97580 14086
rect 97524 13962 97580 13972
rect 97860 13692 97916 14200
rect 98084 14138 98140 14756
rect 98084 14086 98086 14138
rect 98138 14086 98140 14138
rect 98084 14074 98140 14086
rect 98308 14474 98364 14486
rect 98308 14422 98310 14474
rect 98362 14422 98364 14474
rect 98308 13916 98364 14422
rect 98616 14200 98728 15000
rect 99288 14200 99400 15000
rect 100072 14200 100184 15000
rect 100436 14812 100492 14822
rect 100436 14700 100492 14756
rect 100436 14644 100604 14700
rect 98308 13860 98476 13916
rect 97860 13636 98028 13692
rect 96740 12292 97244 12348
rect 97412 12460 97468 12470
rect 96740 11004 96796 12292
rect 96740 10938 96796 10948
rect 96852 11452 96908 11462
rect 96628 10714 96684 10724
rect 96852 10780 96908 11396
rect 96852 10714 96908 10724
rect 97300 11452 97356 11462
rect 97300 10108 97356 11396
rect 97300 10042 97356 10052
rect 97412 9660 97468 12404
rect 97412 9594 97468 9604
rect 97748 11898 97804 11910
rect 97748 11846 97750 11898
rect 97802 11846 97804 11898
rect 97748 9266 97804 11846
rect 97748 9214 97750 9266
rect 97802 9214 97804 9266
rect 97748 9202 97804 9214
rect 97972 8427 98028 13636
rect 98196 12234 98252 12246
rect 98196 12182 98198 12234
rect 98250 12182 98252 12234
rect 98084 12012 98140 12022
rect 98084 11562 98140 11956
rect 98084 11510 98086 11562
rect 98138 11510 98140 11562
rect 98084 11498 98140 11510
rect 98196 11116 98252 12182
rect 98308 11898 98364 11910
rect 98308 11846 98310 11898
rect 98362 11846 98364 11898
rect 98308 11788 98364 11846
rect 98308 11722 98364 11732
rect 98196 11050 98252 11060
rect 98308 11450 98364 11462
rect 98308 11398 98310 11450
rect 98362 11398 98364 11450
rect 97972 8371 98252 8427
rect 96404 8026 96460 8036
rect 96068 6524 96124 6534
rect 96180 6524 96236 8026
rect 97636 7980 97692 7990
rect 97524 7924 97636 7980
rect 97524 7420 97580 7924
rect 97636 7914 97692 7924
rect 98084 7470 98140 7482
rect 97524 7354 97580 7364
rect 97692 7420 97748 7430
rect 97692 7326 97748 7364
rect 98084 7418 98086 7470
rect 98138 7418 98140 7470
rect 95956 6466 96012 6478
rect 95956 6414 95958 6466
rect 96010 6414 96012 6466
rect 95956 2938 96012 6414
rect 96124 6468 96236 6524
rect 96852 7196 96908 7206
rect 96068 5180 96124 6468
rect 96068 5114 96124 5124
rect 96068 5010 96124 5022
rect 96068 4958 96070 5010
rect 96122 4958 96124 5010
rect 96068 4506 96124 4958
rect 96068 4454 96070 4506
rect 96122 4454 96124 4506
rect 96068 4442 96124 4454
rect 96180 4732 96236 4742
rect 95956 2886 95958 2938
rect 96010 2886 96012 2938
rect 95956 2874 96012 2886
rect 96068 3274 96124 3286
rect 96068 3222 96070 3274
rect 96122 3222 96124 3274
rect 96068 2492 96124 3222
rect 96068 2426 96124 2436
rect 96180 2938 96236 4676
rect 96404 4732 96460 4742
rect 96292 4506 96348 4518
rect 96292 4454 96294 4506
rect 96346 4454 96348 4506
rect 96292 3276 96348 4454
rect 96404 4284 96460 4676
rect 96404 4218 96460 4228
rect 96292 3210 96348 3220
rect 96740 4060 96796 4070
rect 96180 2886 96182 2938
rect 96234 2886 96236 2938
rect 95844 2102 95846 2154
rect 95898 2102 95900 2154
rect 95844 2090 95900 2102
rect 95956 2268 96012 2278
rect 95956 1708 96012 2212
rect 95956 1642 96012 1652
rect 96180 1484 96236 2886
rect 95844 1428 96236 1484
rect 96292 2154 96348 2166
rect 96292 2102 96294 2154
rect 96346 2102 96348 2154
rect 95844 800 95900 1428
rect 96292 1036 96348 2102
rect 96292 970 96348 980
rect 96516 2156 96572 2166
rect 96516 800 96572 2100
rect 96628 1820 96684 1830
rect 96628 1034 96684 1764
rect 96628 982 96630 1034
rect 96682 982 96684 1034
rect 96628 970 96684 982
rect 96740 1036 96796 4004
rect 96852 3386 96908 7140
rect 97412 6690 97468 6702
rect 97412 6638 97414 6690
rect 97466 6638 97468 6690
rect 97300 6578 97356 6590
rect 97300 6526 97302 6578
rect 97354 6526 97356 6578
rect 97300 6020 97356 6526
rect 97412 6188 97468 6638
rect 97916 6524 97972 6534
rect 97412 6122 97468 6132
rect 97860 6522 97972 6524
rect 97860 6470 97918 6522
rect 97970 6470 97972 6522
rect 97860 6458 97972 6470
rect 97860 6020 97916 6458
rect 97300 5964 97916 6020
rect 97412 5180 97468 5190
rect 97412 5122 97468 5124
rect 96964 5068 97020 5078
rect 97412 5070 97414 5122
rect 97466 5070 97468 5122
rect 97412 5058 97468 5070
rect 96964 3836 97020 5012
rect 96964 3770 97020 3780
rect 97076 4956 97132 4966
rect 96852 3334 96854 3386
rect 96906 3334 96908 3386
rect 96852 3322 96908 3334
rect 97076 2156 97132 4900
rect 97860 3276 97916 5964
rect 97972 5516 98028 5526
rect 98084 5516 98140 7418
rect 98028 5460 98140 5516
rect 97972 5450 98028 5460
rect 98028 5180 98084 5190
rect 98028 5086 98084 5124
rect 98196 4058 98252 8371
rect 98308 8426 98364 11398
rect 98420 11004 98476 13860
rect 98420 10938 98476 10948
rect 98532 12234 98588 12246
rect 98532 12182 98534 12234
rect 98586 12182 98588 12234
rect 98532 10108 98588 12182
rect 98644 12236 98700 14200
rect 99204 14138 99260 14150
rect 99204 14086 99206 14138
rect 99258 14086 99260 14138
rect 98644 12170 98700 12180
rect 98980 13580 99036 13590
rect 98532 10042 98588 10052
rect 98756 11002 98812 11014
rect 98756 10950 98758 11002
rect 98810 10950 98812 11002
rect 98308 8374 98310 8426
rect 98362 8374 98364 8426
rect 98308 8362 98364 8374
rect 98532 8988 98588 8998
rect 98364 6522 98420 6534
rect 98364 6470 98366 6522
rect 98418 6470 98420 6522
rect 98364 6412 98420 6470
rect 98364 6188 98420 6356
rect 98364 6122 98420 6132
rect 98196 4006 98198 4058
rect 98250 4006 98252 4058
rect 98196 3994 98252 4006
rect 98420 4058 98476 4070
rect 98420 4006 98422 4058
rect 98474 4006 98476 4058
rect 97860 3210 97916 3220
rect 97972 3724 98028 3734
rect 97636 2156 97692 2166
rect 97076 2100 97636 2156
rect 96852 1036 96908 1046
rect 96740 1034 96908 1036
rect 96740 982 96854 1034
rect 96906 982 96908 1034
rect 96740 980 96908 982
rect 96852 970 96908 980
rect 97076 800 97132 2100
rect 97636 2090 97692 2100
rect 97412 1820 97468 1830
rect 97412 1370 97468 1764
rect 97636 1820 97692 1830
rect 97636 1594 97692 1764
rect 97636 1542 97638 1594
rect 97690 1542 97692 1594
rect 97636 1530 97692 1542
rect 97412 1318 97414 1370
rect 97466 1318 97468 1370
rect 97412 1306 97468 1318
rect 97972 1146 98028 3668
rect 98420 3610 98476 4006
rect 98420 3558 98422 3610
rect 98474 3558 98476 3610
rect 98420 3546 98476 3558
rect 97972 1094 97974 1146
rect 98026 1094 98028 1146
rect 97972 1082 98028 1094
rect 98308 1594 98364 1606
rect 98308 1542 98310 1594
rect 98362 1542 98364 1594
rect 97412 1036 97468 1046
rect 85764 364 85820 758
rect 85764 298 85820 308
rect 86072 0 86184 800
rect 86632 0 86744 800
rect 87304 0 87416 800
rect 87864 0 87976 800
rect 88536 0 88648 800
rect 89096 0 89208 800
rect 89768 0 89880 800
rect 90328 0 90440 800
rect 91000 0 91112 800
rect 91560 0 91672 800
rect 92120 0 92232 800
rect 92792 0 92904 800
rect 93352 0 93464 800
rect 94024 0 94136 800
rect 94584 0 94696 800
rect 95256 0 95368 800
rect 95816 0 95928 800
rect 96488 0 96600 800
rect 97048 0 97160 800
rect 97412 588 97468 980
rect 97636 868 98028 924
rect 97636 800 97692 868
rect 97300 532 97468 588
rect 97300 364 97356 532
rect 97300 298 97356 308
rect 97608 0 97720 800
rect 97972 700 98028 868
rect 98308 800 98364 1542
rect 98532 922 98588 8932
rect 98644 8258 98700 8270
rect 98644 8206 98646 8258
rect 98698 8206 98700 8258
rect 98644 6524 98700 8206
rect 98756 6802 98812 10950
rect 98980 11002 99036 13524
rect 99204 13580 99260 14086
rect 99204 13514 99260 13524
rect 99204 12124 99260 12134
rect 99204 11898 99260 12068
rect 99204 11846 99206 11898
rect 99258 11846 99260 11898
rect 99204 11834 99260 11846
rect 99316 11676 99372 14200
rect 99428 14138 99484 14150
rect 99428 14086 99430 14138
rect 99482 14086 99484 14138
rect 99428 13018 99484 14086
rect 99428 12966 99430 13018
rect 99482 12966 99484 13018
rect 99428 12954 99484 12966
rect 99652 13916 99708 13926
rect 99652 12906 99708 13860
rect 99652 12854 99654 12906
rect 99706 12854 99708 12906
rect 99652 12842 99708 12854
rect 100100 12572 100156 14200
rect 100548 14140 100604 14644
rect 100744 14200 100856 15000
rect 101332 14812 101388 14822
rect 101108 14588 101164 14598
rect 100996 14250 101052 14262
rect 100772 14140 100828 14200
rect 100548 14084 100828 14140
rect 100996 14198 100998 14250
rect 101050 14198 101052 14250
rect 100996 13802 101052 14198
rect 100996 13750 100998 13802
rect 101050 13750 101052 13802
rect 100996 13738 101052 13750
rect 99316 11610 99372 11620
rect 99428 12516 100156 12572
rect 100548 13690 100604 13702
rect 100548 13638 100550 13690
rect 100602 13638 100604 13690
rect 99428 11340 99484 12516
rect 100436 12460 100492 12470
rect 100324 12124 100380 12134
rect 100212 11788 100268 11798
rect 99316 11284 99484 11340
rect 99540 11676 99596 11686
rect 98980 10950 98982 11002
rect 99034 10950 99036 11002
rect 98980 10938 99036 10950
rect 99204 11004 99260 11014
rect 98924 10108 98980 10118
rect 98924 9660 98980 10052
rect 98924 9658 99036 9660
rect 98924 9606 98926 9658
rect 98978 9606 99036 9658
rect 98924 9594 99036 9606
rect 98980 9042 99036 9594
rect 99092 9436 99148 9446
rect 99092 9154 99148 9380
rect 99092 9102 99094 9154
rect 99146 9102 99148 9154
rect 99092 9090 99148 9102
rect 98980 8990 98982 9042
rect 99034 8990 99036 9042
rect 98980 8978 99036 8990
rect 99204 7868 99260 10948
rect 99204 7802 99260 7812
rect 99092 7474 99148 7486
rect 99092 7422 99094 7474
rect 99146 7422 99148 7474
rect 99092 7420 99148 7422
rect 99092 7354 99148 7364
rect 99316 7196 99372 11284
rect 99540 8316 99596 11620
rect 99652 11562 99708 11574
rect 99652 11510 99654 11562
rect 99706 11510 99708 11562
rect 99652 10668 99708 11510
rect 100212 11452 100268 11732
rect 100324 11564 100380 12068
rect 100436 11786 100492 12404
rect 100548 12124 100604 13638
rect 101108 13130 101164 14532
rect 101332 13802 101388 14756
rect 101528 14200 101640 15000
rect 102004 14362 102060 14374
rect 102004 14310 102006 14362
rect 102058 14310 102060 14362
rect 101332 13750 101334 13802
rect 101386 13750 101388 13802
rect 101332 13738 101388 13750
rect 101108 13078 101110 13130
rect 101162 13078 101164 13130
rect 101108 13066 101164 13078
rect 101556 12460 101612 14200
rect 101780 13802 101836 13814
rect 101780 13750 101782 13802
rect 101834 13750 101836 13802
rect 101780 12796 101836 13750
rect 101780 12730 101836 12740
rect 102004 12796 102060 14310
rect 102200 14200 102312 15000
rect 102676 14924 102732 14934
rect 102676 14698 102732 14868
rect 102676 14646 102678 14698
rect 102730 14646 102732 14698
rect 102676 14634 102732 14646
rect 102564 14588 102620 14598
rect 102564 14474 102620 14532
rect 102564 14422 102566 14474
rect 102618 14422 102620 14474
rect 102564 14410 102620 14422
rect 102452 14362 102508 14374
rect 102452 14310 102454 14362
rect 102506 14310 102508 14362
rect 102228 13916 102284 14200
rect 102116 13860 102284 13916
rect 102116 13802 102172 13860
rect 102116 13750 102118 13802
rect 102170 13750 102172 13802
rect 102116 13738 102172 13750
rect 102452 13690 102508 14310
rect 102676 14250 102732 14262
rect 102676 14198 102678 14250
rect 102730 14198 102732 14250
rect 102984 14200 103096 15000
rect 103236 14922 103292 14934
rect 103236 14870 103238 14922
rect 103290 14870 103292 14922
rect 102676 14140 102732 14198
rect 103012 14140 103068 14200
rect 102676 14084 103068 14140
rect 102452 13638 102454 13690
rect 102506 13638 102508 13690
rect 102452 13626 102508 13638
rect 102564 14026 102620 14038
rect 102564 13974 102566 14026
rect 102618 13974 102620 14026
rect 102564 13130 102620 13974
rect 103236 13916 103292 14870
rect 103656 14200 103768 15000
rect 104020 14812 104076 14822
rect 104020 14810 104188 14812
rect 104020 14758 104022 14810
rect 104074 14758 104188 14810
rect 104020 14756 104188 14758
rect 104020 14746 104076 14756
rect 103908 14586 103964 14598
rect 103908 14534 103910 14586
rect 103962 14534 103964 14586
rect 103684 13916 103740 14200
rect 103908 14026 103964 14534
rect 103908 13974 103910 14026
rect 103962 13974 103964 14026
rect 103908 13962 103964 13974
rect 104020 14252 104076 14262
rect 102564 13078 102566 13130
rect 102618 13078 102620 13130
rect 102564 13066 102620 13078
rect 102788 13860 103292 13916
rect 103348 13860 103740 13916
rect 102788 13018 102844 13860
rect 103348 13804 103404 13860
rect 102788 12966 102790 13018
rect 102842 12966 102844 13018
rect 102788 12954 102844 12966
rect 102900 13748 103404 13804
rect 102004 12730 102060 12740
rect 102340 12906 102396 12918
rect 102340 12854 102342 12906
rect 102394 12854 102396 12906
rect 101556 12394 101612 12404
rect 100548 12058 100604 12068
rect 100436 11734 100438 11786
rect 100490 11734 100492 11786
rect 100436 11722 100492 11734
rect 100996 11898 101052 11910
rect 100996 11846 100998 11898
rect 101050 11846 101052 11898
rect 100996 11674 101052 11846
rect 101892 11788 101948 11798
rect 101948 11732 102060 11788
rect 101892 11722 101948 11732
rect 100996 11622 100998 11674
rect 101050 11622 101052 11674
rect 100996 11610 101052 11622
rect 101556 11674 101612 11686
rect 101556 11622 101558 11674
rect 101610 11622 101612 11674
rect 100324 11508 100492 11564
rect 100436 11452 100492 11508
rect 100212 11396 100380 11452
rect 100436 11396 100940 11452
rect 100212 11228 100268 11238
rect 100324 11228 100380 11396
rect 100436 11228 100492 11238
rect 100324 11172 100436 11228
rect 100212 10780 100268 11172
rect 100436 11162 100492 11172
rect 100548 11116 100604 11126
rect 100548 10892 100604 11060
rect 100772 10892 100828 10902
rect 100548 10836 100772 10892
rect 100772 10826 100828 10836
rect 100884 10780 100940 11396
rect 101444 10780 101500 10790
rect 100884 10724 101444 10780
rect 100212 10714 100268 10724
rect 101444 10714 101500 10724
rect 99652 10602 99708 10612
rect 100436 10668 100492 10678
rect 100436 10556 100492 10612
rect 101556 10556 101612 11622
rect 100436 10500 101612 10556
rect 99876 10220 99932 10230
rect 99876 10108 99932 10164
rect 99876 10052 100268 10108
rect 99708 9658 99764 9670
rect 100044 9660 100100 9670
rect 99708 9606 99710 9658
rect 99762 9606 99764 9658
rect 99708 9436 99764 9606
rect 99708 9370 99764 9380
rect 99876 9658 100100 9660
rect 99876 9606 100046 9658
rect 100098 9606 100100 9658
rect 99876 9604 100100 9606
rect 99540 8250 99596 8260
rect 99764 9212 99820 9222
rect 99876 9212 99932 9604
rect 100044 9594 100100 9604
rect 100212 9548 100268 10052
rect 100884 9548 100940 9558
rect 100212 9492 100884 9548
rect 100884 9482 100940 9492
rect 101220 9436 101276 9446
rect 101276 9380 101948 9436
rect 101220 9370 101276 9380
rect 99764 9210 99932 9212
rect 99764 9158 99766 9210
rect 99818 9158 99932 9210
rect 99764 9156 99932 9158
rect 99316 7140 99484 7196
rect 98756 6750 98758 6802
rect 98810 6750 98812 6802
rect 98756 6738 98812 6750
rect 99316 6972 99372 6982
rect 98644 6458 98700 6468
rect 99316 6018 99372 6916
rect 99316 5966 99318 6018
rect 99370 5966 99372 6018
rect 99316 5954 99372 5966
rect 99204 5068 99260 5078
rect 99204 3724 99260 5012
rect 99428 4732 99484 7140
rect 99316 4676 99484 4732
rect 99316 4058 99372 4676
rect 99316 4006 99318 4058
rect 99370 4006 99372 4058
rect 99316 3994 99372 4006
rect 99428 4508 99484 4518
rect 99204 3658 99260 3668
rect 99428 3722 99484 4452
rect 99764 4506 99820 9156
rect 101668 9100 101724 9110
rect 100828 9042 100884 9054
rect 100828 8990 100830 9042
rect 100882 8990 100884 9042
rect 100100 8874 100156 8886
rect 100716 8876 100772 8886
rect 100100 8822 100102 8874
rect 100154 8822 100156 8874
rect 99876 8652 99932 8662
rect 99876 7868 99932 8596
rect 100100 8316 100156 8822
rect 100100 8250 100156 8260
rect 100324 8874 100772 8876
rect 100324 8822 100718 8874
rect 100770 8822 100772 8874
rect 100324 8820 100772 8822
rect 100324 8262 100380 8820
rect 100716 8810 100772 8820
rect 100324 8210 100326 8262
rect 100378 8210 100380 8262
rect 100324 8198 100380 8210
rect 100436 8652 100492 8662
rect 100828 8652 100884 8990
rect 101276 8988 101332 8998
rect 99876 7802 99932 7812
rect 100100 7532 100156 7542
rect 100100 6972 100156 7476
rect 100100 6906 100156 6916
rect 100324 6690 100380 6702
rect 100324 6638 100326 6690
rect 100378 6638 100380 6690
rect 100212 6578 100268 6590
rect 100212 6526 100214 6578
rect 100266 6526 100268 6578
rect 100212 6524 100268 6526
rect 100212 6458 100268 6468
rect 99764 4454 99766 4506
rect 99818 4454 99820 4506
rect 99764 4442 99820 4454
rect 100100 4956 100156 4966
rect 100100 4506 100156 4900
rect 100324 4956 100380 6638
rect 100436 5852 100492 8596
rect 100772 8596 100884 8652
rect 101220 8986 101332 8988
rect 101220 8934 101278 8986
rect 101330 8934 101332 8986
rect 101220 8922 101332 8934
rect 100436 5786 100492 5796
rect 100548 8316 100604 8326
rect 100324 4890 100380 4900
rect 100436 5628 100492 5638
rect 100100 4454 100102 4506
rect 100154 4454 100156 4506
rect 100100 4442 100156 4454
rect 100212 4396 100268 4406
rect 99540 4060 99596 4070
rect 99540 3966 99596 4004
rect 99988 4060 100044 4070
rect 99428 3670 99430 3722
rect 99482 3670 99484 3722
rect 99428 3658 99484 3670
rect 98644 3610 98700 3622
rect 98644 3558 98646 3610
rect 98698 3558 98700 3610
rect 98644 2604 98700 3558
rect 99092 3612 99148 3622
rect 99092 2826 99148 3556
rect 99876 3612 99932 3622
rect 99876 3050 99932 3556
rect 99876 2998 99878 3050
rect 99930 2998 99932 3050
rect 99876 2986 99932 2998
rect 99092 2774 99094 2826
rect 99146 2774 99148 2826
rect 99092 2762 99148 2774
rect 99316 2938 99372 2950
rect 99316 2886 99318 2938
rect 99370 2886 99372 2938
rect 98644 2538 98700 2548
rect 99316 2604 99372 2886
rect 99316 2538 99372 2548
rect 99764 2714 99820 2726
rect 99764 2662 99766 2714
rect 99818 2662 99820 2714
rect 99764 2604 99820 2662
rect 99764 2538 99820 2548
rect 99540 2268 99596 2278
rect 98532 870 98534 922
rect 98586 870 98588 922
rect 98532 858 98588 870
rect 98868 2044 98924 2054
rect 98868 800 98924 1988
rect 99428 1372 99484 1382
rect 99428 1034 99484 1316
rect 99428 982 99430 1034
rect 99482 982 99484 1034
rect 99428 970 99484 982
rect 99540 800 99596 2212
rect 99876 1820 99932 1830
rect 99876 922 99932 1764
rect 99988 1260 100044 4004
rect 100212 3050 100268 4340
rect 100212 2998 100214 3050
rect 100266 2998 100268 3050
rect 100212 2986 100268 2998
rect 100324 2826 100380 2838
rect 100324 2774 100326 2826
rect 100378 2774 100380 2826
rect 100212 2602 100268 2614
rect 100212 2550 100214 2602
rect 100266 2550 100268 2602
rect 99988 1194 100044 1204
rect 100100 1708 100156 1718
rect 99876 870 99878 922
rect 99930 870 99932 922
rect 99876 858 99932 870
rect 100100 800 100156 1652
rect 100212 1260 100268 2550
rect 100324 1594 100380 2774
rect 100436 2378 100492 5572
rect 100548 2604 100604 8260
rect 100772 8316 100828 8596
rect 100660 7418 100716 7430
rect 100660 7366 100662 7418
rect 100714 7366 100716 7418
rect 100660 6188 100716 7366
rect 100772 7196 100828 8260
rect 101220 8316 101276 8922
rect 101668 8370 101724 9044
rect 101892 9100 101948 9380
rect 101892 9034 101948 9044
rect 101220 8250 101276 8260
rect 101444 8316 101500 8326
rect 101668 8318 101670 8370
rect 101722 8318 101724 8370
rect 101668 8306 101724 8318
rect 101444 7980 101500 8260
rect 101444 7914 101500 7924
rect 101780 8092 101836 8102
rect 100772 7130 100828 7140
rect 101052 6524 101108 6534
rect 101052 6430 101108 6468
rect 101612 6524 101668 6534
rect 101612 6430 101668 6468
rect 100660 6122 100716 6132
rect 101780 6020 101836 8036
rect 101556 5964 101836 6020
rect 100660 5906 100716 5918
rect 100660 5854 100662 5906
rect 100714 5854 100716 5906
rect 100660 5852 100716 5854
rect 100660 5786 100716 5796
rect 101276 5852 101332 5862
rect 101276 5850 101388 5852
rect 101276 5798 101278 5850
rect 101330 5798 101388 5850
rect 101276 5786 101388 5798
rect 100996 5292 101052 5302
rect 100772 3836 100828 3846
rect 100660 3164 100716 3174
rect 100772 3164 100828 3780
rect 100996 3610 101052 5236
rect 101332 4956 101388 5786
rect 101556 5068 101612 5964
rect 101724 5852 101780 5862
rect 101780 5796 101836 5852
rect 101724 5720 101836 5796
rect 101556 5002 101612 5012
rect 101780 5068 101836 5720
rect 102004 5068 102060 11732
rect 102228 11786 102284 11798
rect 102228 11734 102230 11786
rect 102282 11734 102284 11786
rect 102228 11340 102284 11734
rect 102340 11788 102396 12854
rect 102564 12906 102620 12918
rect 102564 12854 102566 12906
rect 102618 12854 102620 12906
rect 102564 11898 102620 12854
rect 102900 12906 102956 13748
rect 103460 13692 103516 13702
rect 103236 13690 103516 13692
rect 103236 13638 103462 13690
rect 103514 13638 103516 13690
rect 103236 13636 103516 13638
rect 103012 13356 103068 13366
rect 103012 13018 103068 13300
rect 103236 13242 103292 13636
rect 103460 13626 103516 13636
rect 103236 13190 103238 13242
rect 103290 13190 103292 13242
rect 103236 13178 103292 13190
rect 103348 13466 103404 13478
rect 103348 13414 103350 13466
rect 103402 13414 103404 13466
rect 103348 13132 103404 13414
rect 104020 13356 104076 14196
rect 104132 13466 104188 14756
rect 104132 13414 104134 13466
rect 104186 13414 104188 13466
rect 104132 13402 104188 13414
rect 104244 14362 104300 14374
rect 104244 14310 104246 14362
rect 104298 14310 104300 14362
rect 103796 13300 104076 13356
rect 103348 13066 103404 13076
rect 103460 13130 103516 13142
rect 103460 13078 103462 13130
rect 103514 13078 103516 13130
rect 103012 12966 103014 13018
rect 103066 12966 103068 13018
rect 103012 12954 103068 12966
rect 102900 12854 102902 12906
rect 102954 12854 102956 12906
rect 102900 12842 102956 12854
rect 103124 12796 103180 12806
rect 103012 12794 103180 12796
rect 103012 12742 103126 12794
rect 103178 12742 103180 12794
rect 103012 12740 103180 12742
rect 102676 12682 102732 12694
rect 102676 12630 102678 12682
rect 102730 12630 102732 12682
rect 102676 12572 102732 12630
rect 102900 12572 102956 12582
rect 102676 12570 102956 12572
rect 102676 12518 102902 12570
rect 102954 12518 102956 12570
rect 102676 12516 102956 12518
rect 102900 12506 102956 12516
rect 102900 12124 102956 12134
rect 103012 12124 103068 12740
rect 103124 12730 103180 12740
rect 103460 12460 103516 13078
rect 103796 13018 103852 13300
rect 103796 12966 103798 13018
rect 103850 12966 103852 13018
rect 103796 12954 103852 12966
rect 104020 13018 104076 13030
rect 104020 12966 104022 13018
rect 104074 12966 104076 13018
rect 103572 12684 103628 12694
rect 104020 12684 104076 12966
rect 104244 12908 104300 14310
rect 104440 14200 104552 15000
rect 104804 14922 104860 14934
rect 104804 14870 104806 14922
rect 104858 14870 104860 14922
rect 104692 14586 104748 14598
rect 104692 14534 104694 14586
rect 104746 14534 104748 14586
rect 104244 12842 104300 12852
rect 104356 13020 104412 13030
rect 103572 12682 104076 12684
rect 103572 12630 103574 12682
rect 103626 12630 104076 12682
rect 103572 12628 104076 12630
rect 103572 12618 103628 12628
rect 103348 12404 103516 12460
rect 104132 12570 104188 12582
rect 104132 12518 104134 12570
rect 104186 12518 104188 12570
rect 102900 12122 103068 12124
rect 102900 12070 102902 12122
rect 102954 12070 103068 12122
rect 102900 12068 103068 12070
rect 103124 12348 103180 12358
rect 103124 12122 103180 12292
rect 103348 12346 103404 12404
rect 103348 12294 103350 12346
rect 103402 12294 103404 12346
rect 103348 12282 103404 12294
rect 103684 12346 103740 12358
rect 103684 12294 103686 12346
rect 103738 12294 103740 12346
rect 103124 12070 103126 12122
rect 103178 12070 103180 12122
rect 102900 12058 102956 12068
rect 103124 12058 103180 12070
rect 103236 12234 103292 12246
rect 103236 12182 103238 12234
rect 103290 12182 103292 12234
rect 102564 11846 102566 11898
rect 102618 11846 102620 11898
rect 102564 11834 102620 11846
rect 103012 11898 103068 11910
rect 103012 11846 103014 11898
rect 103066 11846 103068 11898
rect 102452 11788 102508 11798
rect 102340 11786 102508 11788
rect 102340 11734 102454 11786
rect 102506 11734 102508 11786
rect 102340 11732 102508 11734
rect 102452 11722 102508 11732
rect 102900 11340 102956 11350
rect 102228 11284 102900 11340
rect 102900 11274 102956 11284
rect 103012 11002 103068 11846
rect 103236 11788 103292 12182
rect 103460 12234 103516 12246
rect 103460 12182 103462 12234
rect 103514 12182 103516 12234
rect 103460 12124 103516 12182
rect 103460 12058 103516 12068
rect 103236 11732 103628 11788
rect 103012 10950 103014 11002
rect 103066 10950 103068 11002
rect 103012 10938 103068 10950
rect 103348 11450 103404 11462
rect 103348 11398 103350 11450
rect 103402 11398 103404 11450
rect 103348 11002 103404 11398
rect 103572 11450 103628 11732
rect 103684 11786 103740 12294
rect 104132 12348 104188 12518
rect 104132 12282 104188 12292
rect 104244 12572 104300 12582
rect 104132 12124 104188 12134
rect 104020 11900 104076 11910
rect 104020 11806 104076 11844
rect 103684 11734 103686 11786
rect 103738 11734 103740 11786
rect 103684 11722 103740 11734
rect 103572 11398 103574 11450
rect 103626 11398 103628 11450
rect 103572 11386 103628 11398
rect 103348 10950 103350 11002
rect 103402 10950 103404 11002
rect 103348 10938 103404 10950
rect 103796 10108 103852 10118
rect 103460 9996 103516 10006
rect 102956 9772 103012 9782
rect 102900 9716 102956 9772
rect 102900 9678 103012 9716
rect 102228 9548 102284 9558
rect 102228 9436 102284 9492
rect 102228 9380 102732 9436
rect 102452 8540 102508 8550
rect 102116 6690 102172 6702
rect 102116 6638 102118 6690
rect 102170 6638 102172 6690
rect 102116 6636 102172 6638
rect 102116 6570 102172 6580
rect 102452 5234 102508 8484
rect 102452 5182 102454 5234
rect 102506 5182 102508 5234
rect 102452 5170 102508 5182
rect 102564 8258 102620 8270
rect 102564 8206 102566 8258
rect 102618 8206 102620 8258
rect 102564 8092 102620 8206
rect 102004 5012 102508 5068
rect 101780 5002 101836 5012
rect 101332 4890 101388 4900
rect 101780 4732 101836 4742
rect 101108 4564 101612 4620
rect 101108 3948 101164 4564
rect 101444 4396 101500 4406
rect 101108 3882 101164 3892
rect 101220 4060 101276 4070
rect 100996 3558 100998 3610
rect 101050 3558 101052 3610
rect 100996 3546 101052 3558
rect 100660 3162 100828 3164
rect 100660 3110 100662 3162
rect 100714 3110 100828 3162
rect 100660 3108 100828 3110
rect 100884 3500 100940 3510
rect 100660 3098 100716 3108
rect 100660 2828 100716 2838
rect 100884 2828 100940 3444
rect 100660 2826 100940 2828
rect 100660 2774 100662 2826
rect 100714 2774 100940 2826
rect 100660 2772 100940 2774
rect 100996 3388 101052 3398
rect 100660 2762 100716 2772
rect 100548 2548 100828 2604
rect 100436 2326 100438 2378
rect 100490 2326 100492 2378
rect 100436 2314 100492 2326
rect 100660 1818 100716 1830
rect 100660 1766 100662 1818
rect 100714 1766 100716 1818
rect 100324 1542 100326 1594
rect 100378 1542 100380 1594
rect 100324 1530 100380 1542
rect 100548 1706 100604 1718
rect 100548 1654 100550 1706
rect 100602 1654 100604 1706
rect 100548 1372 100604 1654
rect 100660 1596 100716 1766
rect 100660 1530 100716 1540
rect 100772 1594 100828 2548
rect 100996 1818 101052 3332
rect 101108 3386 101164 3398
rect 101108 3334 101110 3386
rect 101162 3334 101164 3386
rect 101108 3164 101164 3334
rect 101108 3098 101164 3108
rect 101108 2938 101164 2950
rect 101108 2886 101110 2938
rect 101162 2886 101164 2938
rect 101108 1930 101164 2886
rect 101108 1878 101110 1930
rect 101162 1878 101164 1930
rect 101108 1866 101164 1878
rect 100996 1766 100998 1818
rect 101050 1766 101052 1818
rect 100996 1754 101052 1766
rect 101220 1708 101276 4004
rect 101220 1642 101276 1652
rect 101332 3948 101388 3958
rect 100772 1542 100774 1594
rect 100826 1542 100828 1594
rect 100772 1530 100828 1542
rect 100884 1372 100940 1382
rect 100548 1370 100940 1372
rect 100548 1318 100886 1370
rect 100938 1318 100940 1370
rect 100548 1316 100940 1318
rect 100884 1306 100940 1316
rect 100996 1372 101052 1382
rect 100212 1194 100268 1204
rect 100772 1146 100828 1158
rect 100772 1094 100774 1146
rect 100826 1094 100828 1146
rect 100772 800 100828 1094
rect 100996 922 101052 1316
rect 100996 870 100998 922
rect 101050 870 101052 922
rect 100996 858 101052 870
rect 101332 800 101388 3892
rect 101444 1146 101500 4340
rect 101556 3164 101612 4564
rect 101556 3098 101612 3108
rect 101780 3162 101836 4676
rect 102004 4732 102060 4742
rect 101780 3110 101782 3162
rect 101834 3110 101836 3162
rect 101780 3098 101836 3110
rect 101892 4620 101948 4630
rect 101892 2826 101948 4564
rect 102004 4506 102060 4676
rect 102004 4454 102006 4506
rect 102058 4454 102060 4506
rect 102004 4442 102060 4454
rect 102340 4506 102396 4518
rect 102340 4454 102342 4506
rect 102394 4454 102396 4506
rect 102004 3836 102060 3846
rect 102340 3836 102396 4454
rect 102004 3834 102396 3836
rect 102004 3782 102006 3834
rect 102058 3782 102396 3834
rect 102004 3780 102396 3782
rect 102452 3836 102508 5012
rect 102564 4058 102620 8036
rect 102676 7420 102732 9380
rect 102900 8988 102956 9678
rect 102900 8922 102956 8932
rect 103460 8988 103516 9940
rect 103684 9772 103740 9782
rect 103684 9678 103740 9716
rect 103460 8922 103516 8932
rect 103012 8146 103068 8158
rect 103012 8094 103014 8146
rect 103066 8094 103068 8146
rect 103012 8092 103068 8094
rect 103628 8092 103684 8102
rect 103012 8090 103684 8092
rect 103012 8038 103630 8090
rect 103682 8038 103684 8090
rect 103012 8036 103684 8038
rect 103348 7868 103404 7878
rect 102676 7354 102732 7364
rect 102788 7362 102844 7374
rect 102788 7310 102790 7362
rect 102842 7310 102844 7362
rect 102788 6972 102844 7310
rect 103348 7308 103404 7812
rect 103628 7532 103684 8036
rect 103796 7868 103852 10052
rect 104020 10108 104076 10118
rect 104020 9994 104076 10052
rect 104020 9942 104022 9994
rect 104074 9942 104076 9994
rect 104020 9930 104076 9942
rect 104132 8372 104188 12068
rect 104244 9222 104300 12516
rect 104356 9436 104412 12964
rect 104468 11004 104524 14200
rect 104580 13802 104636 13814
rect 104580 13750 104582 13802
rect 104634 13750 104636 13802
rect 104580 11786 104636 13750
rect 104692 12908 104748 14534
rect 104692 12842 104748 12852
rect 104804 12906 104860 14870
rect 105112 14200 105224 15000
rect 105896 14200 106008 15000
rect 106568 14200 106680 15000
rect 107352 14200 107464 15000
rect 108024 14200 108136 15000
rect 108808 14200 108920 15000
rect 109480 14200 109592 15000
rect 110264 14200 110376 15000
rect 111048 14200 111160 15000
rect 111720 14200 111832 15000
rect 112504 14200 112616 15000
rect 113176 14200 113288 15000
rect 113652 14812 113708 14822
rect 113428 14586 113484 14598
rect 113428 14534 113430 14586
rect 113482 14534 113484 14586
rect 104804 12854 104806 12906
rect 104858 12854 104860 12906
rect 104804 12842 104860 12854
rect 104580 11734 104582 11786
rect 104634 11734 104636 11786
rect 104580 11722 104636 11734
rect 104468 10938 104524 10948
rect 105140 9772 105196 14200
rect 105364 12908 105420 12918
rect 105140 9706 105196 9716
rect 105252 12572 105308 12582
rect 104356 9370 104412 9380
rect 104244 9212 104356 9222
rect 105140 9212 105196 9222
rect 104244 9210 105196 9212
rect 104244 9158 104302 9210
rect 104354 9158 105142 9210
rect 105194 9158 105196 9210
rect 104244 9156 105196 9158
rect 104300 9146 104356 9156
rect 105140 9146 105196 9156
rect 103908 8316 104188 8372
rect 103908 8250 103964 8260
rect 104076 8092 104132 8102
rect 104076 7998 104132 8036
rect 104524 8090 104580 8102
rect 104524 8038 104526 8090
rect 104578 8038 104580 8090
rect 103796 7812 104076 7868
rect 103628 7476 103964 7532
rect 103348 7242 103404 7252
rect 102788 6906 102844 6916
rect 103012 7196 103068 7206
rect 103012 6972 103068 7140
rect 103012 6906 103068 6916
rect 103796 6860 103852 6870
rect 103124 6690 103180 6702
rect 103124 6638 103126 6690
rect 103178 6638 103180 6690
rect 103124 6524 103180 6638
rect 103124 6458 103180 6468
rect 103684 5852 103740 5862
rect 102564 4006 102566 4058
rect 102618 4006 102620 4058
rect 102564 3994 102620 4006
rect 102676 5516 102732 5526
rect 102452 3780 102620 3836
rect 102004 3770 102060 3780
rect 102340 3610 102396 3622
rect 102340 3558 102342 3610
rect 102394 3558 102396 3610
rect 102340 3386 102396 3558
rect 102340 3334 102342 3386
rect 102394 3334 102396 3386
rect 102340 3322 102396 3334
rect 101892 2774 101894 2826
rect 101946 2774 101948 2826
rect 101892 2762 101948 2774
rect 102004 3276 102060 3286
rect 101556 2378 101612 2390
rect 101556 2326 101558 2378
rect 101610 2326 101612 2378
rect 101556 2044 101612 2326
rect 101780 2268 101836 2278
rect 101780 2154 101836 2212
rect 101780 2102 101782 2154
rect 101834 2102 101836 2154
rect 101780 2090 101836 2102
rect 101556 1978 101612 1988
rect 102004 2044 102060 3220
rect 102452 3050 102508 3062
rect 102452 2998 102454 3050
rect 102506 2998 102508 3050
rect 102452 2492 102508 2998
rect 102452 2426 102508 2436
rect 102004 1978 102060 1988
rect 102340 2380 102396 2390
rect 102340 1930 102396 2324
rect 102564 2154 102620 3780
rect 102676 3722 102732 5460
rect 103684 5190 103740 5796
rect 103628 5180 103740 5190
rect 103460 5178 103740 5180
rect 102788 5124 102844 5134
rect 103460 5126 103630 5178
rect 103682 5126 103740 5178
rect 103460 5124 103740 5126
rect 102788 5122 103516 5124
rect 102788 5070 102790 5122
rect 102842 5070 103516 5122
rect 103628 5114 103684 5124
rect 102788 5068 103516 5070
rect 102788 5058 102844 5068
rect 103460 4058 103516 4070
rect 103460 4006 103462 4058
rect 103514 4006 103516 4058
rect 102676 3670 102678 3722
rect 102730 3670 102732 3722
rect 102676 3658 102732 3670
rect 102900 3946 102956 3958
rect 102900 3894 102902 3946
rect 102954 3894 102956 3946
rect 102676 3388 102732 3398
rect 102676 2828 102732 3332
rect 102900 3388 102956 3894
rect 103460 3498 103516 4006
rect 103460 3446 103462 3498
rect 103514 3446 103516 3498
rect 103460 3434 103516 3446
rect 102900 3322 102956 3332
rect 102676 2762 102732 2772
rect 102900 3050 102956 3062
rect 102900 2998 102902 3050
rect 102954 2998 102956 3050
rect 102900 2268 102956 2998
rect 103684 2604 103740 2614
rect 103684 2380 103740 2548
rect 103684 2314 103740 2324
rect 102900 2202 102956 2212
rect 102564 2102 102566 2154
rect 102618 2102 102620 2154
rect 102564 2090 102620 2102
rect 102340 1878 102342 1930
rect 102394 1878 102396 1930
rect 102340 1866 102396 1878
rect 102452 1818 102508 1830
rect 102452 1766 102454 1818
rect 102506 1766 102508 1818
rect 102452 1708 102508 1766
rect 103012 1820 103068 1830
rect 102900 1708 102956 1718
rect 102452 1706 102956 1708
rect 102452 1654 102902 1706
rect 102954 1654 102956 1706
rect 102452 1652 102956 1654
rect 102900 1642 102956 1652
rect 101444 1094 101446 1146
rect 101498 1094 101500 1146
rect 101444 1082 101500 1094
rect 101780 1594 101836 1606
rect 101780 1542 101782 1594
rect 101834 1542 101836 1594
rect 101780 1146 101836 1542
rect 101780 1094 101782 1146
rect 101834 1094 101836 1146
rect 101780 1082 101836 1094
rect 102004 1594 102060 1606
rect 102004 1542 102006 1594
rect 102058 1542 102060 1594
rect 102004 800 102060 1542
rect 103012 924 103068 1764
rect 102564 868 103068 924
rect 103124 1708 103180 1718
rect 102564 800 102620 868
rect 103124 800 103180 1652
rect 103796 800 103852 6804
rect 103908 2380 103964 7476
rect 104020 7084 104076 7812
rect 104132 7586 104188 7598
rect 104132 7534 104134 7586
rect 104186 7534 104188 7586
rect 104132 7532 104188 7534
rect 104524 7532 104580 8038
rect 104132 7466 104188 7476
rect 104244 7476 104580 7532
rect 104972 7532 105028 7542
rect 104244 7474 104300 7476
rect 104244 7422 104246 7474
rect 104298 7422 104300 7474
rect 104020 7018 104076 7028
rect 104132 7196 104188 7206
rect 104020 6748 104076 6758
rect 104020 5180 104076 6692
rect 104132 5852 104188 7140
rect 104132 5786 104188 5796
rect 104020 5114 104076 5124
rect 104132 4058 104188 4070
rect 104132 4006 104134 4058
rect 104186 4006 104188 4058
rect 104132 3722 104188 4006
rect 104132 3670 104134 3722
rect 104186 3670 104188 3722
rect 104132 3658 104188 3670
rect 104020 3610 104076 3622
rect 104020 3558 104022 3610
rect 104074 3558 104076 3610
rect 104020 3050 104076 3558
rect 104020 2998 104022 3050
rect 104074 2998 104076 3050
rect 104020 2986 104076 2998
rect 104244 3050 104300 7422
rect 104972 7418 105028 7476
rect 104972 7366 104974 7418
rect 105026 7366 105028 7418
rect 104972 6860 105028 7366
rect 104972 6804 105196 6860
rect 104916 6522 104972 6534
rect 104916 6470 104918 6522
rect 104970 6470 104972 6522
rect 104244 2998 104246 3050
rect 104298 2998 104300 3050
rect 104244 2986 104300 2998
rect 104356 5852 104412 5862
rect 103908 2314 103964 2324
rect 104356 800 104412 5796
rect 104916 5852 104972 6470
rect 104916 5786 104972 5796
rect 105028 6524 105084 6534
rect 104692 4282 104748 4294
rect 104692 4230 104694 4282
rect 104746 4230 104748 4282
rect 104692 3498 104748 4230
rect 104692 3446 104694 3498
rect 104746 3446 104748 3498
rect 104692 3434 104748 3446
rect 104916 4282 104972 4294
rect 104916 4230 104918 4282
rect 104970 4230 104972 4282
rect 104916 2602 104972 4230
rect 104916 2550 104918 2602
rect 104970 2550 104972 2602
rect 104916 2538 104972 2550
rect 105028 800 105084 6468
rect 105140 2602 105196 6804
rect 105140 2550 105142 2602
rect 105194 2550 105196 2602
rect 105140 2538 105196 2550
rect 105252 1594 105308 12516
rect 105364 6524 105420 12852
rect 105812 11786 105868 11798
rect 105812 11734 105814 11786
rect 105866 11734 105868 11786
rect 105588 11004 105644 11014
rect 105476 8874 105532 8886
rect 105476 8822 105478 8874
rect 105530 8822 105532 8874
rect 105476 6858 105532 8822
rect 105476 6806 105478 6858
rect 105530 6806 105532 6858
rect 105476 6794 105532 6806
rect 105364 6458 105420 6468
rect 105364 5740 105420 5750
rect 105364 5234 105420 5684
rect 105364 5182 105366 5234
rect 105418 5182 105420 5234
rect 105364 5170 105420 5182
rect 105252 1542 105254 1594
rect 105306 1542 105308 1594
rect 105252 1530 105308 1542
rect 105588 800 105644 10948
rect 105812 10444 105868 11734
rect 105924 11788 105980 14200
rect 105924 11722 105980 11732
rect 106372 12124 106428 12134
rect 105812 10378 105868 10388
rect 105700 8428 105756 8438
rect 105700 7362 105756 8372
rect 105700 7310 105702 7362
rect 105754 7310 105756 7362
rect 105700 7298 105756 7310
rect 105700 6860 105756 6870
rect 105700 6766 105756 6804
rect 105700 6412 105756 6422
rect 105700 5740 105756 6356
rect 105700 5674 105756 5684
rect 105812 4058 105868 4070
rect 105812 4006 105814 4058
rect 105866 4006 105868 4058
rect 105812 1260 105868 4006
rect 106372 3387 106428 12068
rect 106596 12012 106652 14200
rect 107380 12796 107436 14200
rect 107380 12730 107436 12740
rect 107940 12796 107996 12806
rect 106596 11946 106652 11956
rect 106484 11340 106540 11350
rect 106484 10332 106540 11284
rect 106484 10266 106540 10276
rect 106876 9660 106932 9670
rect 107828 9660 107884 9670
rect 106820 9658 107884 9660
rect 106820 9606 106878 9658
rect 106930 9606 107830 9658
rect 107882 9606 107884 9658
rect 106820 9604 107884 9606
rect 106820 9594 106932 9604
rect 107828 9594 107884 9604
rect 106708 5180 106764 5190
rect 106708 5122 106764 5124
rect 106708 5070 106710 5122
rect 106762 5070 106764 5122
rect 106708 5058 106764 5070
rect 106820 3387 106876 9594
rect 107940 8326 107996 12740
rect 108052 11450 108108 14200
rect 108052 11398 108054 11450
rect 108106 11398 108108 11450
rect 108052 11386 108108 11398
rect 108724 11898 108780 11910
rect 108724 11846 108726 11898
rect 108778 11846 108780 11898
rect 108724 9772 108780 11846
rect 108836 10780 108892 14200
rect 109172 12908 109228 12918
rect 109172 12814 109228 12852
rect 108948 12012 109004 12022
rect 108948 11898 109004 11956
rect 108948 11846 108950 11898
rect 109002 11846 109004 11898
rect 108948 11834 109004 11846
rect 109284 11674 109340 11686
rect 109284 11622 109286 11674
rect 109338 11622 109340 11674
rect 109284 11338 109340 11622
rect 109508 11564 109564 14200
rect 109844 12906 109900 12918
rect 109844 12854 109846 12906
rect 109898 12854 109900 12906
rect 109620 12460 109676 12470
rect 109620 12236 109676 12404
rect 109844 12460 109900 12854
rect 109844 12394 109900 12404
rect 109620 12170 109676 12180
rect 109508 11498 109564 11508
rect 109732 11674 109788 11686
rect 109732 11622 109734 11674
rect 109786 11622 109788 11674
rect 109284 11286 109286 11338
rect 109338 11286 109340 11338
rect 109284 11274 109340 11286
rect 108836 10714 108892 10724
rect 109396 10668 109452 10678
rect 108332 9770 108780 9772
rect 108332 9718 108726 9770
rect 108778 9718 108780 9770
rect 108332 9716 108780 9718
rect 108164 9660 108220 9670
rect 108164 9566 108220 9604
rect 108332 9210 108388 9716
rect 108724 9706 108780 9716
rect 108836 9884 108892 9894
rect 108836 9436 108892 9828
rect 109060 9884 109116 9894
rect 109060 9790 109116 9828
rect 109284 9436 109340 9446
rect 108836 9380 109284 9436
rect 109284 9370 109340 9380
rect 109396 9268 109452 10612
rect 109732 10666 109788 11622
rect 109732 10614 109734 10666
rect 109786 10614 109788 10666
rect 109732 10602 109788 10614
rect 109956 10666 110012 10678
rect 109956 10614 109958 10666
rect 110010 10614 110012 10666
rect 109956 9994 110012 10614
rect 110292 10107 110348 14200
rect 110852 12906 110908 12918
rect 110852 12854 110854 12906
rect 110906 12854 110908 12906
rect 110852 11340 110908 12854
rect 110964 11898 111020 11910
rect 110964 11846 110966 11898
rect 111018 11846 111020 11898
rect 110964 11564 111020 11846
rect 110964 11498 111020 11508
rect 110852 11274 110908 11284
rect 111076 10107 111132 14200
rect 111188 14026 111244 14038
rect 111188 13974 111190 14026
rect 111242 13974 111244 14026
rect 111188 11898 111244 13974
rect 111188 11846 111190 11898
rect 111242 11846 111244 11898
rect 111188 11834 111244 11846
rect 109956 9942 109958 9994
rect 110010 9942 110012 9994
rect 109956 9930 110012 9942
rect 110180 10051 110348 10107
rect 110628 10051 111132 10107
rect 111636 10444 111692 10454
rect 110180 9996 110236 10051
rect 110180 9930 110236 9940
rect 108332 9158 108334 9210
rect 108386 9158 108388 9210
rect 108332 9146 108388 9158
rect 109060 9212 109452 9268
rect 109620 9658 109676 9670
rect 109620 9606 109622 9658
rect 109674 9606 109676 9658
rect 107268 8316 107324 8326
rect 107156 7586 107212 7598
rect 107156 7534 107158 7586
rect 107210 7534 107212 7586
rect 107156 6524 107212 7534
rect 107268 7474 107324 8260
rect 107884 8316 107996 8326
rect 107940 8260 107996 8316
rect 107884 8184 107940 8260
rect 107548 8090 107604 8102
rect 107548 8038 107550 8090
rect 107602 8038 107604 8090
rect 107548 7644 107604 8038
rect 107548 7588 107996 7644
rect 107268 7422 107270 7474
rect 107322 7422 107324 7474
rect 107940 7532 107996 7588
rect 107940 7476 108780 7532
rect 107268 7410 107324 7422
rect 107828 7455 107884 7467
rect 107828 7403 107830 7455
rect 107882 7403 107884 7455
rect 107828 6972 107884 7403
rect 107828 6906 107884 6916
rect 107660 6524 107716 6534
rect 107156 6522 107772 6524
rect 107156 6470 107662 6522
rect 107714 6470 107772 6522
rect 107156 6468 107772 6470
rect 107660 6458 107772 6468
rect 107548 5180 107604 5190
rect 107548 4954 107604 5124
rect 107548 4902 107550 4954
rect 107602 4902 107604 4954
rect 107548 4890 107604 4902
rect 106260 3331 106428 3387
rect 106708 3331 106876 3387
rect 106932 3948 106988 3958
rect 105812 1194 105868 1204
rect 105924 1594 105980 1606
rect 105924 1542 105926 1594
rect 105978 1542 105980 1594
rect 105924 1036 105980 1542
rect 105924 970 105980 980
rect 106148 1036 106204 1046
rect 106148 942 106204 980
rect 106260 800 106316 3331
rect 106708 1482 106764 3331
rect 106708 1430 106710 1482
rect 106762 1430 106764 1482
rect 106708 1418 106764 1430
rect 106820 2492 106876 2502
rect 106372 1036 106428 1046
rect 106372 942 106428 980
rect 106820 800 106876 2436
rect 106932 1594 106988 3892
rect 107604 3276 107660 3286
rect 107492 3220 107604 3276
rect 107492 2716 107548 3220
rect 107604 3210 107660 3220
rect 107492 2650 107548 2660
rect 107716 2716 107772 6458
rect 107940 3387 107996 7476
rect 108724 7474 108780 7476
rect 108724 7422 108726 7474
rect 108778 7422 108780 7474
rect 108724 7410 108780 7422
rect 108500 6636 108556 6646
rect 108500 5964 108556 6580
rect 108500 5898 108556 5908
rect 107828 3331 107996 3387
rect 108948 5010 109004 5022
rect 108948 4958 108950 5010
rect 109002 4958 109004 5010
rect 107828 3162 107884 3331
rect 107828 3110 107830 3162
rect 107882 3110 107884 3162
rect 107828 3098 107884 3110
rect 108500 3162 108556 3174
rect 108500 3110 108502 3162
rect 108554 3110 108556 3162
rect 108500 2828 108556 3110
rect 107716 2650 107772 2660
rect 108164 2772 108556 2828
rect 106932 1542 106934 1594
rect 106986 1542 106988 1594
rect 106932 1530 106988 1542
rect 107492 1706 107548 1718
rect 107492 1654 107494 1706
rect 107546 1654 107548 1706
rect 107492 800 107548 1654
rect 108164 1706 108220 2772
rect 108948 2716 109004 4958
rect 109060 4282 109116 9212
rect 109228 8988 109284 8998
rect 109172 8986 109284 8988
rect 109172 8934 109230 8986
rect 109282 8934 109284 8986
rect 109172 8922 109284 8934
rect 109172 8316 109228 8922
rect 109172 8250 109228 8260
rect 109620 8316 109676 9606
rect 109868 9436 110132 9446
rect 109924 9380 109972 9436
rect 110028 9380 110076 9436
rect 109868 9370 110132 9380
rect 110628 9100 110684 10051
rect 111524 9772 111580 9782
rect 110852 9770 111580 9772
rect 110852 9718 111526 9770
rect 111578 9718 111580 9770
rect 110852 9716 111580 9718
rect 110852 9670 110908 9716
rect 111524 9706 111580 9716
rect 110796 9660 110908 9670
rect 110628 9034 110684 9044
rect 110740 9658 110908 9660
rect 110740 9606 110798 9658
rect 110850 9606 110908 9658
rect 110740 9604 110908 9606
rect 110740 9594 110852 9604
rect 109620 8250 109676 8260
rect 110460 8316 110516 8326
rect 110460 8258 110516 8260
rect 110460 8206 110462 8258
rect 110514 8206 110516 8258
rect 110348 8092 110404 8102
rect 109284 8090 110404 8092
rect 109284 8038 110350 8090
rect 110402 8038 110404 8090
rect 109284 8036 110404 8038
rect 109172 6972 109228 6982
rect 109284 6972 109340 8036
rect 110348 8026 110404 8036
rect 109868 7868 110132 7878
rect 109924 7812 109972 7868
rect 110028 7812 110076 7868
rect 110460 7868 110516 8206
rect 110740 8092 110796 9594
rect 110964 9548 111020 9558
rect 110964 9212 111020 9492
rect 110964 9146 111020 9156
rect 111188 9100 111244 9110
rect 110740 8026 110796 8036
rect 110908 8092 110964 8102
rect 110908 7868 110964 8036
rect 110460 7812 110964 7868
rect 109868 7802 110132 7812
rect 109508 7756 109564 7766
rect 111076 7756 111132 7766
rect 110180 7700 111076 7756
rect 109508 7644 110236 7700
rect 111076 7690 111132 7700
rect 111188 7588 111244 9044
rect 110964 7532 111244 7588
rect 110964 7306 111020 7532
rect 111636 7308 111692 10388
rect 111748 7980 111804 14200
rect 111972 14026 112028 14038
rect 111972 13974 111974 14026
rect 112026 13974 112028 14026
rect 111860 11564 111916 11574
rect 111860 9994 111916 11508
rect 111860 9942 111862 9994
rect 111914 9942 111916 9994
rect 111860 9930 111916 9942
rect 111748 7914 111804 7924
rect 110964 7254 110966 7306
rect 111018 7254 111020 7306
rect 110964 7242 111020 7254
rect 111524 7252 111692 7308
rect 109228 6916 109340 6972
rect 109172 6906 109228 6916
rect 110180 6860 110236 6870
rect 110068 6804 110180 6860
rect 110068 6636 110124 6804
rect 110180 6794 110236 6804
rect 110516 6692 110572 6702
rect 111524 6692 111580 7252
rect 110516 6690 111580 6692
rect 110516 6638 110518 6690
rect 110570 6638 111580 6690
rect 110516 6636 111580 6638
rect 110516 6626 110572 6636
rect 110068 6570 110124 6580
rect 110404 6578 110460 6590
rect 110404 6526 110406 6578
rect 110458 6526 110460 6578
rect 110404 6524 110460 6526
rect 111300 6524 111356 6534
rect 109060 4230 109062 4282
rect 109114 4230 109116 4282
rect 109060 4218 109116 4230
rect 109284 6466 109340 6478
rect 110404 6468 110684 6524
rect 109284 6414 109286 6466
rect 109338 6414 109340 6466
rect 109284 3387 109340 6414
rect 109868 6300 110132 6310
rect 109924 6244 109972 6300
rect 110028 6244 110076 6300
rect 109868 6234 110132 6244
rect 109732 6188 109788 6198
rect 109732 5964 109788 6132
rect 110516 6188 110572 6198
rect 109732 5898 109788 5908
rect 110068 5964 110124 5974
rect 109732 5628 109788 5638
rect 109396 4732 109452 4742
rect 109396 4282 109452 4676
rect 109396 4230 109398 4282
rect 109450 4230 109452 4282
rect 109396 4218 109452 4230
rect 109172 3331 109340 3387
rect 109732 3387 109788 5572
rect 110068 5068 110124 5908
rect 110068 5002 110124 5012
rect 110292 5122 110348 5134
rect 110292 5070 110294 5122
rect 110346 5070 110348 5122
rect 110292 5068 110348 5070
rect 110292 5002 110348 5012
rect 110516 4956 110572 6132
rect 110628 5852 110684 6468
rect 111300 6466 111356 6468
rect 111300 6414 111302 6466
rect 111354 6414 111356 6466
rect 111300 6402 111356 6414
rect 111524 6086 111580 6636
rect 111468 6074 111580 6086
rect 111468 6022 111470 6074
rect 111522 6022 111580 6074
rect 111468 6020 111580 6022
rect 111636 7084 111692 7094
rect 111468 6010 111524 6020
rect 110908 5852 110964 5862
rect 110628 5850 111020 5852
rect 110628 5798 110910 5850
rect 110962 5798 111020 5850
rect 110628 5796 111020 5798
rect 110908 5786 111020 5796
rect 110516 4890 110572 4900
rect 110964 4956 111020 5786
rect 110964 4890 111020 4900
rect 111468 5068 111524 5078
rect 111468 4956 111524 5012
rect 111636 4956 111692 7028
rect 111972 6188 112028 13974
rect 112532 13020 112588 14200
rect 112980 14026 113036 14038
rect 112980 13974 112982 14026
rect 113034 13974 113036 14026
rect 112980 13916 113036 13974
rect 113204 13916 113260 14200
rect 113428 14026 113484 14534
rect 113428 13974 113430 14026
rect 113482 13974 113484 14026
rect 113428 13962 113484 13974
rect 112980 13860 113260 13916
rect 113652 13804 113708 14756
rect 113764 14588 113820 14598
rect 113764 13804 113820 14532
rect 113960 14200 114072 15000
rect 114212 14250 114268 14262
rect 113876 13804 113932 13814
rect 113764 13748 113876 13804
rect 113652 13738 113708 13748
rect 113876 13738 113932 13748
rect 112308 12964 112588 13020
rect 112084 12572 112140 12582
rect 112084 11562 112140 12516
rect 112084 11510 112086 11562
rect 112138 11510 112140 11562
rect 112084 11498 112140 11510
rect 112308 11116 112364 12964
rect 113988 12572 114044 14200
rect 114212 14198 114214 14250
rect 114266 14198 114268 14250
rect 114632 14200 114744 15000
rect 115220 14924 115276 14934
rect 114884 14476 114940 14514
rect 114884 14410 114940 14420
rect 115220 14476 115276 14868
rect 115220 14410 115276 14420
rect 114996 14362 115052 14374
rect 114996 14310 114998 14362
rect 115050 14310 115052 14362
rect 114212 14026 114268 14198
rect 114212 13974 114214 14026
rect 114266 13974 114268 14026
rect 114212 13962 114268 13974
rect 114660 13468 114716 14200
rect 114996 14026 115052 14310
rect 115416 14200 115528 15000
rect 115892 14812 115948 14822
rect 115668 14810 115948 14812
rect 115668 14758 115894 14810
rect 115946 14758 115948 14810
rect 115668 14756 115948 14758
rect 115668 14698 115724 14756
rect 115892 14746 115948 14756
rect 115668 14646 115670 14698
rect 115722 14646 115724 14698
rect 115668 14634 115724 14646
rect 116088 14200 116200 15000
rect 116340 14698 116396 14710
rect 116340 14646 116342 14698
rect 116394 14646 116396 14698
rect 116340 14250 116396 14646
rect 114996 13974 114998 14026
rect 115050 13974 115052 14026
rect 114996 13962 115052 13974
rect 115444 14028 115500 14200
rect 116116 14028 116172 14200
rect 116340 14198 116342 14250
rect 116394 14198 116396 14250
rect 116340 14186 116396 14198
rect 116564 14586 116620 14598
rect 116564 14534 116566 14586
rect 116618 14534 116620 14586
rect 116564 14028 116620 14534
rect 116676 14474 116732 14486
rect 116676 14422 116678 14474
rect 116730 14422 116732 14474
rect 116676 14138 116732 14422
rect 116872 14200 116984 15000
rect 117124 14474 117180 14486
rect 117124 14422 117126 14474
rect 117178 14422 117180 14474
rect 116676 14086 116678 14138
rect 116730 14086 116732 14138
rect 116676 14074 116732 14086
rect 115444 13962 115500 13972
rect 115780 13972 116172 14028
rect 116228 13972 116620 14028
rect 113652 12516 114044 12572
rect 114212 13412 114716 13468
rect 114212 12572 114268 13412
rect 115220 13354 115276 13366
rect 115220 13302 115222 13354
rect 115274 13302 115276 13354
rect 114660 13242 114716 13254
rect 114660 13190 114662 13242
rect 114714 13190 114716 13242
rect 112308 11050 112364 11060
rect 112420 12236 112476 12246
rect 111972 6122 112028 6132
rect 112308 6578 112364 6590
rect 112308 6526 112310 6578
rect 112362 6526 112364 6578
rect 112308 6188 112364 6526
rect 112420 6412 112476 12180
rect 113652 11900 113708 12516
rect 114212 12506 114268 12516
rect 114436 12906 114492 12918
rect 114436 12854 114438 12906
rect 114490 12854 114492 12906
rect 114436 12460 114492 12854
rect 114660 12906 114716 13190
rect 114660 12854 114662 12906
rect 114714 12854 114716 12906
rect 114660 12842 114716 12854
rect 114548 12794 114604 12806
rect 114548 12742 114550 12794
rect 114602 12742 114604 12794
rect 114548 12684 114604 12742
rect 114772 12740 115052 12796
rect 114772 12684 114828 12740
rect 114548 12628 114828 12684
rect 114996 12682 115052 12740
rect 114996 12630 114998 12682
rect 115050 12630 115052 12682
rect 114996 12618 115052 12630
rect 114884 12570 114940 12582
rect 114884 12518 114886 12570
rect 114938 12518 114940 12570
rect 114436 12404 114828 12460
rect 114212 12236 114268 12246
rect 114212 12012 114268 12180
rect 114548 12124 114604 12134
rect 114548 12122 114716 12124
rect 114548 12070 114550 12122
rect 114602 12070 114716 12122
rect 114548 12068 114716 12070
rect 114548 12058 114604 12068
rect 113204 11844 113708 11900
rect 114156 11956 114268 12012
rect 113092 11788 113148 11798
rect 112756 11564 112812 11574
rect 112756 11228 112812 11508
rect 112756 11162 112812 11172
rect 112532 10108 112588 10118
rect 112532 8092 112588 10052
rect 112532 8026 112588 8036
rect 113092 8092 113148 11732
rect 113092 8026 113148 8036
rect 113204 7644 113260 11844
rect 114156 11788 114212 11956
rect 114156 11732 114268 11788
rect 113652 11452 113708 11462
rect 113876 11452 113932 11462
rect 113652 11450 113932 11452
rect 113652 11398 113654 11450
rect 113706 11398 113878 11450
rect 113930 11398 113932 11450
rect 113652 11396 113932 11398
rect 113652 11386 113708 11396
rect 113876 11386 113932 11396
rect 113428 11340 113484 11350
rect 113204 7578 113260 7588
rect 113316 11116 113372 11126
rect 113316 6758 113372 11060
rect 113428 11004 113484 11284
rect 113428 10938 113484 10948
rect 114100 11338 114156 11350
rect 114100 11286 114102 11338
rect 114154 11286 114156 11338
rect 114100 10444 114156 11286
rect 114212 10666 114268 11732
rect 114212 10614 114214 10666
rect 114266 10614 114268 10666
rect 114212 10602 114268 10614
rect 114324 11676 114380 11686
rect 113876 10388 114156 10444
rect 113652 8204 113708 8214
rect 113652 7868 113708 8148
rect 113652 7802 113708 7812
rect 113764 7644 113820 7654
rect 113260 6748 113372 6758
rect 112756 6746 113372 6748
rect 112756 6694 113262 6746
rect 113314 6694 113372 6746
rect 112756 6692 113372 6694
rect 113652 7588 113764 7644
rect 113652 6692 113708 7588
rect 113764 7578 113820 7588
rect 112756 6690 112812 6692
rect 112756 6638 112758 6690
rect 112810 6638 112812 6690
rect 113260 6682 113316 6692
rect 112756 6626 112812 6638
rect 113540 6636 113708 6692
rect 112420 6356 112812 6412
rect 112308 6122 112364 6132
rect 112644 5068 112700 5078
rect 112196 5012 112252 5022
rect 111468 4954 111692 4956
rect 111468 4902 111470 4954
rect 111522 4902 111692 4954
rect 111468 4900 111692 4902
rect 111860 5010 112252 5012
rect 111860 4958 112198 5010
rect 112250 4958 112252 5010
rect 111860 4956 112252 4958
rect 111468 4890 111524 4900
rect 109868 4732 110132 4742
rect 109924 4676 109972 4732
rect 110028 4676 110076 4732
rect 109868 4666 110132 4676
rect 110516 4732 110572 4742
rect 110516 4396 110572 4676
rect 110516 4330 110572 4340
rect 110628 4620 110684 4630
rect 110628 3948 110684 4564
rect 111860 4508 111916 4956
rect 112196 4946 112252 4956
rect 112532 4956 112588 4966
rect 110516 3892 110684 3948
rect 111636 4452 111916 4508
rect 112420 4844 112476 4854
rect 109732 3331 109900 3387
rect 109060 3276 109116 3286
rect 109060 2940 109116 3220
rect 109172 3164 109228 3331
rect 109172 3098 109228 3108
rect 109060 2874 109116 2884
rect 108164 1654 108166 1706
rect 108218 1654 108220 1706
rect 108164 1642 108220 1654
rect 108276 2660 109004 2716
rect 108276 1372 108332 2660
rect 109060 2604 109116 2614
rect 108388 2548 109060 2604
rect 108388 2044 108444 2548
rect 109060 2538 109116 2548
rect 108948 2380 109004 2390
rect 109004 2324 109116 2380
rect 108948 2314 109004 2324
rect 108388 1978 108444 1988
rect 108612 2044 108668 2054
rect 108388 1708 108444 1718
rect 108388 1594 108444 1652
rect 108388 1542 108390 1594
rect 108442 1542 108444 1594
rect 108388 1530 108444 1542
rect 108276 1306 108332 1316
rect 108052 980 108332 1036
rect 108052 800 108108 980
rect 108276 812 108332 980
rect 97972 644 98140 700
rect 98084 486 98140 644
rect 98084 476 98196 486
rect 98084 420 98140 476
rect 98140 410 98196 420
rect 98280 0 98392 800
rect 98840 0 98952 800
rect 99512 0 99624 800
rect 100072 0 100184 800
rect 100744 0 100856 800
rect 101304 0 101416 800
rect 101976 0 102088 800
rect 102536 0 102648 800
rect 103096 0 103208 800
rect 103768 0 103880 800
rect 104328 0 104440 800
rect 105000 0 105112 800
rect 105560 0 105672 800
rect 106232 0 106344 800
rect 106792 0 106904 800
rect 107464 0 107576 800
rect 108024 0 108136 800
rect 108612 800 108668 1988
rect 109060 1932 109116 2324
rect 109060 1876 109228 1932
rect 109172 1820 109228 1876
rect 109172 1754 109228 1764
rect 109732 1482 109788 1494
rect 109732 1430 109734 1482
rect 109786 1430 109788 1482
rect 109284 1372 109340 1382
rect 109284 800 109340 1316
rect 109732 922 109788 1430
rect 109732 870 109734 922
rect 109786 870 109788 922
rect 109732 858 109788 870
rect 109844 800 109900 3331
rect 110292 2828 110348 2838
rect 109956 2044 110012 2054
rect 109956 1594 110012 1988
rect 109956 1542 109958 1594
rect 110010 1542 110012 1594
rect 109956 1530 110012 1542
rect 110292 1146 110348 2772
rect 110292 1094 110294 1146
rect 110346 1094 110348 1146
rect 110292 1082 110348 1094
rect 110516 800 110572 3892
rect 110628 3722 110684 3734
rect 110628 3670 110630 3722
rect 110682 3670 110684 3722
rect 110628 3052 110684 3670
rect 111636 3386 111692 4452
rect 112420 4060 112476 4788
rect 111636 3334 111638 3386
rect 111690 3334 111692 3386
rect 111636 3322 111692 3334
rect 111748 4004 112476 4060
rect 110628 2986 110684 2996
rect 110852 2828 110908 2838
rect 110852 2826 111244 2828
rect 110852 2774 110854 2826
rect 110906 2774 111244 2826
rect 110852 2772 111244 2774
rect 110852 2762 110908 2772
rect 110740 2714 110796 2726
rect 110740 2662 110742 2714
rect 110794 2662 110796 2714
rect 110740 2604 110796 2662
rect 111188 2714 111244 2772
rect 111188 2662 111190 2714
rect 111242 2662 111244 2714
rect 111188 2650 111244 2662
rect 111076 2604 111132 2614
rect 110740 2602 111132 2604
rect 110740 2550 111078 2602
rect 111130 2550 111132 2602
rect 110740 2548 111132 2550
rect 111076 2538 111132 2548
rect 111412 1372 111468 1382
rect 111412 1278 111468 1316
rect 111636 1372 111692 1382
rect 110740 1148 110796 1158
rect 110740 1034 110796 1092
rect 110740 982 110742 1034
rect 110794 982 110796 1034
rect 110740 970 110796 982
rect 111076 1146 111132 1158
rect 111076 1094 111078 1146
rect 111130 1094 111132 1146
rect 111076 800 111132 1094
rect 111636 1034 111692 1316
rect 111636 982 111638 1034
rect 111690 982 111692 1034
rect 111636 970 111692 982
rect 111748 800 111804 4004
rect 112420 3612 112476 3622
rect 111860 3498 111916 3510
rect 111860 3446 111862 3498
rect 111914 3446 111916 3498
rect 111860 1146 111916 3446
rect 112308 3388 112364 3398
rect 111860 1094 111862 1146
rect 111914 1094 111916 1146
rect 111860 1082 111916 1094
rect 112084 1146 112140 1158
rect 112084 1094 112086 1146
rect 112138 1094 112140 1146
rect 112084 812 112140 1094
rect 108276 746 108332 756
rect 108584 0 108696 800
rect 109256 0 109368 800
rect 109816 0 109928 800
rect 110488 0 110600 800
rect 111048 0 111160 800
rect 111720 0 111832 800
rect 112308 800 112364 3332
rect 112420 3052 112476 3556
rect 112532 3164 112588 4900
rect 112644 4732 112700 5012
rect 112644 4666 112700 4676
rect 112756 3722 112812 6356
rect 113204 6188 113260 6198
rect 112756 3670 112758 3722
rect 112810 3670 112812 3722
rect 112756 3658 112812 3670
rect 112868 4732 112924 4742
rect 112644 3612 112700 3622
rect 112644 3518 112700 3556
rect 112868 3387 112924 4676
rect 113204 3722 113260 6132
rect 113428 5292 113484 5302
rect 113428 5122 113484 5236
rect 113428 5070 113430 5122
rect 113482 5070 113484 5122
rect 113428 5058 113484 5070
rect 113540 4284 113596 6636
rect 113708 6522 113764 6534
rect 113708 6470 113710 6522
rect 113762 6470 113764 6522
rect 113708 6188 113764 6470
rect 113708 6122 113764 6132
rect 113540 4218 113596 4228
rect 113876 3948 113932 10388
rect 113988 10220 114044 10230
rect 114044 10164 114156 10220
rect 113988 10154 114044 10164
rect 114100 7588 114156 10164
rect 114324 7756 114380 11620
rect 114436 11228 114492 11238
rect 114436 10666 114492 11172
rect 114436 10614 114438 10666
rect 114490 10614 114492 10666
rect 114436 10602 114492 10614
rect 114660 9894 114716 12068
rect 114772 12122 114828 12404
rect 114772 12070 114774 12122
rect 114826 12070 114828 12122
rect 114772 12058 114828 12070
rect 114884 12012 114940 12518
rect 115220 12234 115276 13302
rect 115556 13132 115612 13142
rect 115556 12794 115612 13076
rect 115556 12742 115558 12794
rect 115610 12742 115612 12794
rect 115556 12730 115612 12742
rect 115780 12460 115836 13972
rect 115892 13804 115948 13814
rect 115892 13132 115948 13748
rect 116228 13578 116284 13972
rect 116228 13526 116230 13578
rect 116282 13526 116284 13578
rect 116228 13514 116284 13526
rect 116340 13804 116396 13814
rect 116340 13580 116396 13748
rect 116564 13804 116620 13814
rect 116452 13580 116508 13590
rect 116340 13578 116508 13580
rect 116340 13526 116454 13578
rect 116506 13526 116508 13578
rect 116340 13524 116508 13526
rect 116452 13514 116508 13524
rect 115892 13066 115948 13076
rect 116564 12908 116620 13748
rect 116004 12852 116620 12908
rect 116004 12572 116060 12852
rect 116228 12572 116284 12582
rect 116004 12516 116172 12572
rect 115220 12182 115222 12234
rect 115274 12182 115276 12234
rect 115220 12170 115276 12182
rect 115332 12404 115836 12460
rect 114884 11956 115164 12012
rect 114996 11788 115052 11798
rect 115108 11788 115164 11956
rect 115220 11788 115276 11798
rect 115108 11786 115276 11788
rect 115108 11734 115222 11786
rect 115274 11734 115276 11786
rect 115108 11732 115276 11734
rect 114996 11694 115052 11732
rect 115220 11722 115276 11732
rect 115332 11452 115388 12404
rect 115668 12124 115724 12134
rect 115668 12030 115724 12068
rect 115892 12122 115948 12134
rect 115892 12070 115894 12122
rect 115946 12070 115948 12122
rect 115892 11900 115948 12070
rect 115892 11834 115948 11844
rect 115332 11386 115388 11396
rect 116004 11340 116060 11350
rect 116116 11340 116172 12516
rect 116228 12236 116284 12516
rect 116564 12570 116620 12582
rect 116564 12518 116566 12570
rect 116618 12518 116620 12570
rect 116564 12460 116620 12518
rect 116788 12460 116844 12470
rect 116564 12458 116844 12460
rect 116564 12406 116790 12458
rect 116842 12406 116844 12458
rect 116564 12404 116844 12406
rect 116788 12394 116844 12404
rect 116676 12236 116732 12246
rect 116228 12234 116732 12236
rect 116228 12182 116678 12234
rect 116730 12182 116732 12234
rect 116228 12180 116732 12182
rect 116676 12170 116732 12180
rect 116060 11284 116172 11340
rect 116228 12012 116284 12022
rect 116900 12012 116956 14200
rect 117124 13914 117180 14422
rect 117544 14200 117656 15000
rect 118020 14924 118076 14934
rect 117796 14476 117852 14486
rect 117124 13862 117126 13914
rect 117178 13862 117180 13914
rect 117124 13850 117180 13862
rect 117348 14138 117404 14150
rect 117348 14086 117350 14138
rect 117402 14086 117404 14138
rect 117348 13914 117404 14086
rect 117348 13862 117350 13914
rect 117402 13862 117404 13914
rect 117348 13850 117404 13862
rect 117236 13018 117292 13030
rect 117236 12966 117238 13018
rect 117290 12966 117292 13018
rect 117124 12572 117180 12582
rect 117012 12348 117068 12358
rect 117012 12234 117068 12292
rect 117012 12182 117014 12234
rect 117066 12182 117068 12234
rect 117012 12170 117068 12182
rect 116004 11274 116060 11284
rect 116228 10780 116284 11956
rect 116564 11956 116956 12012
rect 116564 11676 116620 11956
rect 117124 11900 117180 12516
rect 117236 12234 117292 12966
rect 117236 12182 117238 12234
rect 117290 12182 117292 12234
rect 117236 12170 117292 12182
rect 117460 13018 117516 13030
rect 117460 12966 117462 13018
rect 117514 12966 117516 13018
rect 117460 12010 117516 12966
rect 117460 11958 117462 12010
rect 117514 11958 117516 12010
rect 117460 11946 117516 11958
rect 116564 11610 116620 11620
rect 116900 11844 117180 11900
rect 116452 11338 116508 11350
rect 116452 11286 116454 11338
rect 116506 11286 116508 11338
rect 116452 11004 116508 11286
rect 116452 10948 116732 11004
rect 116228 10724 116620 10780
rect 115556 10276 116060 10332
rect 115556 10108 115612 10276
rect 115556 10042 115612 10052
rect 115780 10108 115836 10118
rect 115780 9994 115836 10052
rect 115780 9942 115782 9994
rect 115834 9942 115836 9994
rect 115780 9930 115836 9942
rect 116004 9996 116060 10276
rect 116564 10220 116620 10724
rect 116676 10444 116732 10948
rect 116676 10378 116732 10388
rect 116564 10164 116732 10220
rect 116004 9930 116060 9940
rect 114660 9884 114772 9894
rect 114660 9882 115500 9884
rect 114660 9830 114718 9882
rect 114770 9830 115500 9882
rect 114660 9828 115500 9830
rect 114716 9818 114772 9828
rect 115444 9770 115500 9828
rect 115444 9718 115446 9770
rect 115498 9718 115500 9770
rect 115444 9706 115500 9718
rect 114772 9604 115388 9660
rect 114772 9548 114828 9604
rect 114772 9482 114828 9492
rect 115332 9548 115388 9604
rect 115332 9482 115388 9492
rect 115220 9436 115276 9446
rect 115220 8652 115276 9380
rect 116676 9324 116732 10164
rect 116900 9996 116956 11844
rect 117572 11788 117628 14200
rect 117684 13916 117740 13926
rect 117684 13356 117740 13860
rect 117796 13468 117852 14420
rect 118020 14476 118076 14868
rect 118020 14410 118076 14420
rect 118132 14252 118188 14262
rect 118328 14200 118440 15000
rect 118580 14924 118636 14934
rect 118132 14140 118188 14196
rect 118356 14140 118412 14200
rect 118132 14084 118412 14140
rect 117908 13916 117964 13926
rect 117908 13692 117964 13860
rect 118580 13916 118636 14868
rect 118804 14362 118860 14374
rect 118804 14310 118806 14362
rect 118858 14310 118860 14362
rect 118580 13850 118636 13860
rect 118692 14250 118748 14262
rect 118692 14198 118694 14250
rect 118746 14198 118748 14250
rect 117908 13636 118412 13692
rect 118020 13468 118076 13478
rect 117796 13412 118020 13468
rect 118020 13402 118076 13412
rect 117684 13300 117852 13356
rect 116900 9930 116956 9940
rect 117012 11732 117628 11788
rect 117796 11788 117852 13300
rect 118356 12684 118412 13636
rect 118468 13690 118524 13702
rect 118468 13638 118470 13690
rect 118522 13638 118524 13690
rect 118468 13356 118524 13638
rect 118692 13690 118748 14198
rect 118692 13638 118694 13690
rect 118746 13638 118748 13690
rect 118692 13626 118748 13638
rect 118468 13300 118748 13356
rect 118356 12628 118636 12684
rect 118468 12458 118524 12470
rect 118468 12406 118470 12458
rect 118522 12406 118524 12458
rect 118020 12180 118412 12236
rect 118020 12012 118076 12180
rect 118020 11946 118076 11956
rect 118244 12012 118300 12022
rect 118244 11898 118300 11956
rect 118244 11846 118246 11898
rect 118298 11846 118300 11898
rect 118244 11834 118300 11846
rect 117796 11732 118188 11788
rect 116676 9258 116732 9268
rect 116228 9212 116284 9222
rect 115668 9156 116228 9212
rect 115668 8876 115724 9156
rect 116228 9146 116284 9156
rect 115220 8586 115276 8596
rect 115332 8820 115724 8876
rect 115332 7980 115388 8820
rect 114324 7690 114380 7700
rect 114660 7924 115388 7980
rect 115444 8652 115500 8662
rect 114100 7532 114380 7588
rect 113988 7362 114044 7374
rect 113988 7310 113990 7362
rect 114042 7310 114044 7362
rect 113988 4282 114044 7310
rect 114156 5292 114212 5302
rect 114156 5178 114212 5236
rect 114156 5126 114158 5178
rect 114210 5126 114212 5178
rect 114156 5114 114212 5126
rect 114324 4620 114380 7532
rect 114212 4564 114380 4620
rect 113988 4230 113990 4282
rect 114042 4230 114044 4282
rect 113988 4218 114044 4230
rect 114100 4284 114156 4294
rect 113204 3670 113206 3722
rect 113258 3670 113260 3722
rect 113204 3658 113260 3670
rect 113316 3892 113932 3948
rect 112644 3331 112924 3387
rect 112644 3276 112700 3331
rect 112644 3210 112700 3220
rect 112532 3098 112588 3108
rect 112420 2986 112476 2996
rect 113316 2044 113372 3892
rect 113652 3722 113708 3734
rect 113652 3670 113654 3722
rect 113706 3670 113708 3722
rect 113540 3498 113596 3510
rect 113540 3446 113542 3498
rect 113594 3446 113596 3498
rect 113540 3388 113596 3446
rect 113540 3322 113596 3332
rect 113428 3164 113484 3174
rect 113428 2156 113484 3108
rect 113652 2268 113708 3670
rect 113652 2202 113708 2212
rect 113876 3722 113932 3734
rect 113876 3670 113878 3722
rect 113930 3670 113932 3722
rect 113540 2156 113596 2166
rect 113428 2100 113540 2156
rect 113876 2156 113932 3670
rect 114100 3722 114156 4228
rect 114100 3670 114102 3722
rect 114154 3670 114156 3722
rect 114100 3658 114156 3670
rect 113988 3610 114044 3622
rect 113988 3558 113990 3610
rect 114042 3558 114044 3610
rect 113988 3386 114044 3558
rect 114212 3610 114268 4564
rect 114324 4396 114380 4406
rect 114324 4282 114380 4340
rect 114324 4230 114326 4282
rect 114378 4230 114380 4282
rect 114324 4218 114380 4230
rect 114660 4060 114716 7924
rect 114212 3558 114214 3610
rect 114266 3558 114268 3610
rect 114212 3546 114268 3558
rect 114436 4004 114716 4060
rect 114772 7756 114828 7766
rect 115444 7756 115500 8596
rect 114436 3498 114492 4004
rect 114772 3946 114828 7700
rect 115332 7700 115500 7756
rect 115780 8652 115836 8662
rect 117012 8652 117068 11732
rect 117460 11620 117964 11676
rect 117236 11450 117292 11462
rect 117236 11398 117238 11450
rect 117290 11398 117292 11450
rect 117236 11228 117292 11398
rect 117460 11450 117516 11620
rect 117460 11398 117462 11450
rect 117514 11398 117516 11450
rect 117460 11386 117516 11398
rect 117796 11450 117852 11462
rect 117796 11398 117798 11450
rect 117850 11398 117852 11450
rect 117684 11340 117740 11378
rect 117684 11274 117740 11284
rect 117236 11172 117628 11228
rect 117348 11004 117404 11014
rect 117348 10892 117404 10948
rect 117348 10836 117516 10892
rect 117124 10780 117180 10790
rect 117180 10724 117292 10780
rect 117124 10714 117180 10724
rect 114772 3894 114774 3946
rect 114826 3894 114828 3946
rect 114772 3882 114828 3894
rect 115108 6860 115164 6870
rect 115108 3948 115164 6804
rect 115108 3892 115276 3948
rect 114436 3446 114438 3498
rect 114490 3446 114492 3498
rect 114436 3434 114492 3446
rect 114548 3834 114604 3846
rect 114548 3782 114550 3834
rect 114602 3782 114604 3834
rect 113988 3334 113990 3386
rect 114042 3334 114044 3386
rect 113988 3322 114044 3334
rect 114548 2940 114604 3782
rect 115220 3836 115276 3892
rect 115332 3946 115388 7700
rect 115556 7644 115612 7654
rect 115444 7586 115500 7598
rect 115444 7534 115446 7586
rect 115498 7534 115500 7586
rect 115444 7308 115500 7534
rect 115556 7474 115612 7588
rect 115556 7422 115558 7474
rect 115610 7422 115612 7474
rect 115556 7410 115612 7422
rect 115780 7308 115836 8596
rect 116340 8596 117068 8652
rect 116004 8428 116060 8438
rect 116004 7980 116060 8372
rect 116228 8428 116284 8438
rect 116228 8214 116284 8372
rect 116172 8202 116284 8214
rect 116172 8150 116174 8202
rect 116226 8150 116284 8202
rect 116172 8148 116284 8150
rect 116172 8138 116228 8148
rect 116004 7924 116284 7980
rect 115948 7644 116004 7654
rect 115948 7550 116004 7588
rect 115444 7252 115836 7308
rect 115780 6804 115836 7252
rect 115780 6748 116004 6804
rect 115948 6746 116004 6748
rect 115948 6694 115950 6746
rect 116002 6694 116004 6746
rect 115948 6682 116004 6694
rect 115780 6636 115836 6646
rect 116228 6636 116284 7924
rect 116340 6748 116396 8596
rect 117012 8428 117068 8438
rect 116452 8316 116508 8326
rect 116508 8260 116620 8316
rect 116452 8250 116508 8260
rect 116340 6692 116508 6748
rect 116228 6580 116396 6636
rect 115780 6524 116060 6580
rect 115892 5068 115948 5078
rect 115668 5010 115724 5022
rect 115668 4958 115670 5010
rect 115722 4958 115724 5010
rect 115668 4506 115724 4958
rect 115668 4454 115670 4506
rect 115722 4454 115724 4506
rect 115668 4442 115724 4454
rect 115892 4394 115948 5012
rect 116004 4506 116060 6524
rect 116228 6300 116284 6310
rect 116004 4454 116006 4506
rect 116058 4454 116060 4506
rect 116004 4442 116060 4454
rect 116116 4620 116172 4630
rect 115892 4342 115894 4394
rect 115946 4342 115948 4394
rect 115892 4330 115948 4342
rect 116116 4394 116172 4564
rect 116116 4342 116118 4394
rect 116170 4342 116172 4394
rect 116116 4330 116172 4342
rect 115668 4172 115724 4182
rect 115332 3894 115334 3946
rect 115386 3894 115388 3946
rect 115332 3882 115388 3894
rect 115556 3948 115612 3958
rect 115668 3948 115724 4116
rect 115612 3892 115724 3948
rect 115556 3882 115612 3892
rect 115220 3770 115276 3780
rect 115444 3834 115500 3846
rect 115444 3782 115446 3834
rect 115498 3782 115500 3834
rect 115108 3724 115164 3734
rect 114996 3722 115164 3724
rect 114996 3670 115110 3722
rect 115162 3670 115164 3722
rect 114996 3668 115164 3670
rect 114884 3498 114940 3510
rect 114884 3446 114886 3498
rect 114938 3446 114940 3498
rect 114884 3276 114940 3446
rect 114884 3210 114940 3220
rect 114996 3052 115052 3668
rect 115108 3658 115164 3668
rect 115444 3612 115500 3782
rect 115332 3556 115500 3612
rect 115780 3834 115836 3846
rect 115780 3782 115782 3834
rect 115834 3782 115836 3834
rect 115220 3500 115276 3510
rect 115220 3406 115276 3444
rect 114548 2874 114604 2884
rect 114660 2996 115052 3052
rect 114324 2268 114380 2278
rect 113876 2100 114156 2156
rect 113540 2090 113596 2100
rect 113316 1978 113372 1988
rect 113652 2044 113708 2054
rect 113652 1932 113708 1988
rect 113540 1876 113708 1932
rect 112644 1594 112700 1606
rect 112644 1542 112646 1594
rect 112698 1542 112700 1594
rect 112644 1034 112700 1542
rect 112644 982 112646 1034
rect 112698 982 112700 1034
rect 112644 970 112700 982
rect 112868 1594 112924 1606
rect 112868 1542 112870 1594
rect 112922 1542 112924 1594
rect 112868 800 112924 1542
rect 113540 800 113596 1876
rect 114100 800 114156 2100
rect 114324 1932 114380 2212
rect 114324 1866 114380 1876
rect 114660 1146 114716 2996
rect 115108 2940 115164 2950
rect 114772 2884 115108 2940
rect 114772 2604 114828 2884
rect 115108 2874 115164 2884
rect 114772 2538 114828 2548
rect 114660 1094 114662 1146
rect 114714 1094 114716 1146
rect 114660 1082 114716 1094
rect 114884 1036 114940 1046
rect 114772 1034 114940 1036
rect 114772 982 114886 1034
rect 114938 982 114940 1034
rect 114772 980 114940 982
rect 114772 800 114828 980
rect 114884 970 114940 980
rect 115332 800 115388 3556
rect 115444 3388 115500 3398
rect 115444 2154 115500 3332
rect 115780 3386 115836 3782
rect 115780 3334 115782 3386
rect 115834 3334 115836 3386
rect 115780 3322 115836 3334
rect 116116 3836 116172 3846
rect 115444 2102 115446 2154
rect 115498 2102 115500 2154
rect 115444 2090 115500 2102
rect 115892 2826 115948 2838
rect 115892 2774 115894 2826
rect 115946 2774 115948 2826
rect 115668 1820 115724 1830
rect 115556 1596 115612 1606
rect 115668 1596 115724 1764
rect 115892 1820 115948 2774
rect 115892 1754 115948 1764
rect 116004 2154 116060 2166
rect 116004 2102 116006 2154
rect 116058 2102 116060 2154
rect 116004 1596 116060 2102
rect 115668 1540 116060 1596
rect 115556 1484 115612 1540
rect 115556 1428 116060 1484
rect 116004 800 116060 1428
rect 116116 922 116172 3780
rect 116228 3386 116284 6244
rect 116340 6188 116396 6580
rect 116340 6122 116396 6132
rect 116340 4620 116396 4630
rect 116340 4282 116396 4564
rect 116340 4230 116342 4282
rect 116394 4230 116396 4282
rect 116340 4218 116396 4230
rect 116228 3334 116230 3386
rect 116282 3334 116284 3386
rect 116228 3322 116284 3334
rect 116452 3050 116508 6692
rect 116564 6300 116620 8260
rect 117012 8277 117068 8372
rect 117012 8225 117014 8277
rect 117066 8225 117068 8277
rect 117012 8213 117068 8225
rect 116564 6234 116620 6244
rect 116900 7868 116956 7878
rect 116676 4956 116732 4966
rect 116452 2998 116454 3050
rect 116506 2998 116508 3050
rect 116452 2986 116508 2998
rect 116564 4620 116620 4630
rect 116452 1036 116508 1046
rect 116452 942 116508 980
rect 116116 870 116118 922
rect 116170 870 116172 922
rect 116116 858 116172 870
rect 116564 800 116620 4564
rect 116676 1370 116732 4900
rect 116900 3498 116956 7812
rect 117012 7362 117068 7374
rect 117012 7310 117014 7362
rect 117066 7310 117068 7362
rect 117012 6748 117068 7310
rect 117236 6972 117292 10724
rect 117348 10666 117404 10678
rect 117348 10614 117350 10666
rect 117402 10614 117404 10666
rect 117348 7980 117404 10614
rect 117460 9884 117516 10836
rect 117572 10444 117628 11172
rect 117684 10668 117740 10678
rect 117684 10574 117740 10612
rect 117572 10378 117628 10388
rect 117460 9818 117516 9828
rect 117796 8764 117852 11398
rect 117908 11338 117964 11620
rect 117908 11286 117910 11338
rect 117962 11286 117964 11338
rect 117908 11274 117964 11286
rect 118132 8988 118188 11732
rect 118356 11564 118412 12180
rect 118468 12124 118524 12406
rect 118580 12348 118636 12628
rect 118692 12458 118748 13300
rect 118804 13244 118860 14310
rect 119000 14200 119112 15000
rect 119784 14200 119896 15000
rect 120148 14924 120204 14934
rect 118804 13178 118860 13188
rect 118692 12406 118694 12458
rect 118746 12406 118748 12458
rect 118692 12394 118748 12406
rect 118580 12282 118636 12292
rect 118468 12058 118524 12068
rect 119028 12012 119084 14200
rect 119252 14138 119308 14150
rect 119252 14086 119254 14138
rect 119306 14086 119308 14138
rect 119252 13580 119308 14086
rect 119252 13514 119308 13524
rect 119364 13802 119420 13814
rect 119364 13750 119366 13802
rect 119418 13750 119420 13802
rect 119364 13020 119420 13750
rect 119364 12954 119420 12964
rect 119588 13802 119644 13814
rect 119588 13750 119590 13802
rect 119642 13750 119644 13802
rect 119588 12570 119644 13750
rect 119588 12518 119590 12570
rect 119642 12518 119644 12570
rect 119588 12506 119644 12518
rect 119700 13132 119756 13142
rect 119140 12404 119532 12460
rect 119140 12236 119196 12404
rect 119140 12170 119196 12180
rect 119364 12236 119420 12246
rect 118804 11956 119084 12012
rect 118468 11900 118524 11910
rect 118468 11806 118524 11844
rect 118804 11788 118860 11956
rect 118804 11722 118860 11732
rect 119028 11788 119084 11798
rect 118356 11508 118636 11564
rect 118356 11226 118412 11238
rect 118356 11174 118358 11226
rect 118410 11174 118412 11226
rect 118356 10892 118412 11174
rect 118580 11226 118636 11508
rect 119028 11562 119084 11732
rect 119028 11510 119030 11562
rect 119082 11510 119084 11562
rect 119028 11498 119084 11510
rect 119252 11786 119308 11798
rect 119252 11734 119254 11786
rect 119306 11734 119308 11786
rect 119252 11340 119308 11734
rect 119252 11274 119308 11284
rect 118580 11174 118582 11226
rect 118634 11174 118636 11226
rect 118580 11162 118636 11174
rect 118356 10836 118860 10892
rect 118580 10108 118636 10118
rect 118580 9772 118636 10052
rect 118580 9706 118636 9716
rect 118804 9772 118860 10836
rect 118804 9706 118860 9716
rect 118356 9436 118412 9446
rect 118412 9380 118468 9436
rect 118356 9370 118468 9380
rect 118412 9210 118468 9370
rect 118412 9158 118414 9210
rect 118466 9158 118468 9210
rect 118412 9146 118468 9158
rect 118524 9154 118580 9166
rect 118524 9102 118526 9154
rect 118578 9102 118580 9154
rect 118524 9100 118580 9102
rect 118524 9044 118972 9100
rect 118916 8998 118972 9044
rect 118132 8932 118860 8988
rect 118916 8986 119028 8998
rect 118916 8934 118974 8986
rect 119026 8934 119028 8986
rect 118916 8932 119028 8934
rect 117460 8708 117852 8764
rect 117460 8316 117516 8708
rect 117572 8540 117628 8550
rect 117628 8484 118636 8540
rect 117572 8474 117628 8484
rect 117460 8250 117516 8260
rect 117908 8258 117964 8270
rect 117908 8206 117910 8258
rect 117962 8206 117964 8258
rect 117908 8204 117964 8206
rect 117908 8138 117964 8148
rect 118132 8204 118188 8214
rect 118132 7980 118188 8148
rect 118468 8092 118524 8102
rect 117348 7924 118188 7980
rect 118244 8036 118468 8092
rect 118244 7756 118300 8036
rect 118468 8026 118524 8036
rect 118580 7980 118636 8484
rect 118580 7914 118636 7924
rect 117460 7700 118300 7756
rect 117460 7196 117516 7700
rect 118804 7698 118860 8932
rect 118972 8652 119028 8932
rect 119252 8988 119308 8998
rect 118972 8596 119196 8652
rect 118804 7646 118806 7698
rect 118858 7646 118860 7698
rect 117460 7130 117516 7140
rect 117796 7586 117852 7598
rect 117796 7534 117798 7586
rect 117850 7534 117852 7586
rect 117796 7084 117852 7534
rect 118020 7588 118412 7644
rect 118804 7634 118860 7646
rect 118916 8426 118972 8438
rect 118916 8374 118918 8426
rect 118970 8374 118972 8426
rect 118020 7532 118076 7588
rect 118020 7466 118076 7476
rect 118132 7474 118188 7486
rect 118132 7422 118134 7474
rect 118186 7422 118188 7474
rect 117796 7028 118076 7084
rect 117236 6916 117964 6972
rect 117012 6682 117068 6692
rect 117124 6860 117180 6870
rect 117124 6636 117180 6804
rect 117796 6748 117852 6758
rect 117684 6636 117740 6646
rect 117124 6580 117684 6636
rect 117684 6570 117740 6580
rect 117684 5964 117740 5974
rect 117684 5516 117740 5908
rect 117012 5460 117740 5516
rect 117012 5122 117068 5460
rect 117012 5070 117014 5122
rect 117066 5070 117068 5122
rect 117012 5058 117068 5070
rect 117348 5292 117404 5302
rect 116900 3446 116902 3498
rect 116954 3446 116956 3498
rect 116900 3434 116956 3446
rect 117012 4282 117068 4294
rect 117012 4230 117014 4282
rect 117066 4230 117068 4282
rect 116900 2828 116956 2838
rect 116900 2734 116956 2772
rect 117012 2154 117068 4230
rect 117124 3498 117180 3510
rect 117124 3446 117126 3498
rect 117178 3446 117180 3498
rect 117124 3164 117180 3446
rect 117124 3098 117180 3108
rect 117236 3276 117292 3286
rect 117236 2828 117292 3220
rect 117348 3274 117404 5236
rect 117684 5190 117740 5460
rect 117628 5178 117740 5190
rect 117628 5126 117630 5178
rect 117682 5126 117740 5178
rect 117628 5124 117740 5126
rect 117628 5114 117684 5124
rect 117796 5067 117852 6692
rect 117908 6018 117964 6916
rect 118020 6468 118076 7028
rect 118132 6748 118188 7422
rect 118356 7196 118412 7588
rect 118916 7420 118972 8374
rect 118916 7354 118972 7364
rect 119028 7644 119084 7654
rect 119028 7196 119084 7588
rect 118356 7140 119084 7196
rect 118132 6682 118188 6692
rect 118412 6748 118468 6758
rect 118412 6634 118468 6692
rect 118412 6582 118414 6634
rect 118466 6582 118468 6634
rect 118412 6570 118468 6582
rect 118748 6522 118804 6534
rect 118748 6470 118750 6522
rect 118802 6470 118804 6522
rect 118748 6468 118804 6470
rect 118020 6412 118860 6468
rect 117908 5966 117910 6018
rect 117962 5966 117964 6018
rect 117908 5954 117964 5966
rect 117796 5011 118076 5067
rect 117460 4508 117516 4518
rect 117460 4172 117516 4452
rect 117796 4508 117852 4518
rect 117908 4508 117964 4518
rect 117796 4506 117908 4508
rect 117796 4454 117798 4506
rect 117850 4454 117908 4506
rect 117796 4452 117908 4454
rect 117796 4442 117852 4452
rect 117908 4442 117964 4452
rect 118020 4506 118076 5011
rect 118020 4454 118022 4506
rect 118074 4454 118076 4506
rect 118020 4442 118076 4454
rect 117460 4116 117740 4172
rect 117684 3386 117740 4116
rect 118468 4060 118524 4070
rect 118244 3724 118300 3734
rect 117684 3334 117686 3386
rect 117738 3334 117740 3386
rect 117684 3322 117740 3334
rect 118020 3500 118076 3510
rect 117348 3222 117350 3274
rect 117402 3222 117404 3274
rect 117348 3210 117404 3222
rect 117572 3276 117628 3286
rect 117572 3162 117628 3220
rect 117572 3110 117574 3162
rect 117626 3110 117628 3162
rect 117572 3098 117628 3110
rect 117796 3162 117852 3174
rect 117796 3110 117798 3162
rect 117850 3110 117852 3162
rect 117236 2762 117292 2772
rect 117348 3050 117404 3062
rect 117348 2998 117350 3050
rect 117402 2998 117404 3050
rect 117012 2102 117014 2154
rect 117066 2102 117068 2154
rect 117012 2090 117068 2102
rect 117236 2156 117292 2166
rect 117236 2062 117292 2100
rect 117348 1482 117404 2998
rect 117796 2826 117852 3110
rect 117796 2774 117798 2826
rect 117850 2774 117852 2826
rect 117796 2762 117852 2774
rect 117460 2714 117516 2726
rect 117460 2662 117462 2714
rect 117514 2662 117516 2714
rect 117460 2380 117516 2662
rect 117684 2714 117740 2726
rect 117684 2662 117686 2714
rect 117738 2662 117740 2714
rect 117684 2604 117740 2662
rect 117684 2538 117740 2548
rect 117908 2604 117964 2614
rect 117460 2314 117516 2324
rect 117348 1430 117350 1482
rect 117402 1430 117404 1482
rect 117348 1418 117404 1430
rect 117796 1596 117852 1606
rect 116676 1318 116678 1370
rect 116730 1318 116732 1370
rect 116676 1306 116732 1318
rect 117012 1370 117068 1382
rect 117012 1318 117014 1370
rect 117066 1318 117068 1370
rect 116788 1260 116844 1270
rect 116788 1034 116844 1204
rect 117012 1260 117068 1318
rect 117012 1194 117068 1204
rect 116788 982 116790 1034
rect 116842 982 116844 1034
rect 116788 970 116844 982
rect 117012 868 117292 924
rect 112084 746 112140 756
rect 112280 0 112392 800
rect 112840 0 112952 800
rect 113512 0 113624 800
rect 114072 0 114184 800
rect 114744 0 114856 800
rect 115304 0 115416 800
rect 115976 0 116088 800
rect 116536 0 116648 800
rect 117012 700 117068 868
rect 117236 800 117292 868
rect 117796 800 117852 1540
rect 117908 1146 117964 2548
rect 118020 1594 118076 3444
rect 118020 1542 118022 1594
rect 118074 1542 118076 1594
rect 118020 1530 118076 1542
rect 118132 2604 118188 2614
rect 118132 1482 118188 2548
rect 118132 1430 118134 1482
rect 118186 1430 118188 1482
rect 118132 1418 118188 1430
rect 117908 1094 117910 1146
rect 117962 1094 117964 1146
rect 117908 1082 117964 1094
rect 118244 922 118300 3668
rect 118356 3500 118412 3510
rect 118468 3500 118524 4004
rect 118692 3836 118748 3846
rect 118580 3780 118692 3836
rect 118580 3722 118636 3780
rect 118692 3770 118748 3780
rect 118804 3834 118860 6412
rect 119028 5964 119084 5974
rect 118804 3782 118806 3834
rect 118858 3782 118860 3834
rect 118804 3770 118860 3782
rect 118916 5908 119028 5964
rect 118580 3670 118582 3722
rect 118634 3670 118636 3722
rect 118580 3658 118636 3670
rect 118468 3444 118748 3500
rect 118356 2380 118412 3444
rect 118468 3052 118524 3062
rect 118468 2826 118524 2996
rect 118468 2774 118470 2826
rect 118522 2774 118524 2826
rect 118468 2762 118524 2774
rect 118356 2314 118412 2324
rect 118244 870 118246 922
rect 118298 870 118300 922
rect 118244 858 118300 870
rect 118356 1932 118412 1942
rect 118356 800 118412 1876
rect 118692 1708 118748 3444
rect 118916 2604 118972 5908
rect 119028 5898 119084 5908
rect 119140 3162 119196 8596
rect 119252 7588 119308 8932
rect 119364 8092 119420 12180
rect 119476 11340 119532 12404
rect 119476 11274 119532 11284
rect 119588 11562 119644 11574
rect 119588 11510 119590 11562
rect 119642 11510 119644 11562
rect 119588 9324 119644 11510
rect 119588 9258 119644 9268
rect 119364 8026 119420 8036
rect 119700 7644 119756 13076
rect 119812 12796 119868 14200
rect 120036 14026 120092 14038
rect 120036 13974 120038 14026
rect 120090 13974 120092 14026
rect 119812 12730 119868 12740
rect 119924 13914 119980 13926
rect 119924 13862 119926 13914
rect 119978 13862 119980 13914
rect 119924 12570 119980 13862
rect 120036 12796 120092 13974
rect 120148 13916 120204 14868
rect 120148 13850 120204 13860
rect 120260 14810 120316 14822
rect 120260 14758 120262 14810
rect 120314 14758 120316 14810
rect 120260 13802 120316 14758
rect 120456 14200 120568 15000
rect 121044 14922 121100 14934
rect 121044 14870 121046 14922
rect 121098 14870 121100 14922
rect 120708 14588 120764 14598
rect 120708 14362 120764 14532
rect 121044 14476 121100 14870
rect 121044 14410 121100 14420
rect 120708 14310 120710 14362
rect 120762 14310 120764 14362
rect 120708 14298 120764 14310
rect 121240 14200 121352 15000
rect 121492 14810 121548 14822
rect 121492 14758 121494 14810
rect 121546 14758 121548 14810
rect 121492 14476 121548 14758
rect 121492 14410 121548 14420
rect 121604 14362 121660 14374
rect 121604 14310 121606 14362
rect 121658 14310 121660 14362
rect 120260 13750 120262 13802
rect 120314 13750 120316 13802
rect 120260 13738 120316 13750
rect 120036 12730 120092 12740
rect 119924 12518 119926 12570
rect 119978 12518 119980 12570
rect 119924 12506 119980 12518
rect 120484 12572 120540 14200
rect 120596 13972 121100 14028
rect 120596 13130 120652 13972
rect 121044 13914 121100 13972
rect 121044 13862 121046 13914
rect 121098 13862 121100 13914
rect 121044 13850 121100 13862
rect 120596 13078 120598 13130
rect 120650 13078 120652 13130
rect 120596 13066 120652 13078
rect 120820 13130 120876 13142
rect 120820 13078 120822 13130
rect 120874 13078 120876 13130
rect 120708 12796 120764 12806
rect 120820 12796 120876 13078
rect 120764 12740 120876 12796
rect 120708 12730 120764 12740
rect 120484 12506 120540 12516
rect 120820 12572 120876 12582
rect 120820 12570 120988 12572
rect 120820 12518 120822 12570
rect 120874 12518 120988 12570
rect 120820 12516 120988 12518
rect 120820 12506 120876 12516
rect 120932 12460 120988 12516
rect 121044 12460 121100 12470
rect 120932 12458 121100 12460
rect 120932 12406 121046 12458
rect 121098 12406 121100 12458
rect 120932 12404 121100 12406
rect 121044 12394 121100 12404
rect 121268 12460 121324 14200
rect 121604 12906 121660 14310
rect 121912 14200 122024 15000
rect 122500 14810 122556 14822
rect 122500 14758 122502 14810
rect 122554 14758 122556 14810
rect 121604 12854 121606 12906
rect 121658 12854 121660 12906
rect 121604 12842 121660 12854
rect 121268 12394 121324 12404
rect 120820 12348 120876 12358
rect 120372 12236 120428 12246
rect 119812 12124 119868 12134
rect 119868 12068 119980 12124
rect 119812 12058 119868 12068
rect 119812 10220 119868 10230
rect 119812 9212 119868 10164
rect 119812 9146 119868 9156
rect 119924 7868 119980 12068
rect 119924 7802 119980 7812
rect 120148 12012 120204 12022
rect 120148 7756 120204 11956
rect 120372 12012 120428 12180
rect 120372 11946 120428 11956
rect 120372 11788 120428 11798
rect 120596 11788 120652 11798
rect 120372 11694 120428 11732
rect 120484 11786 120652 11788
rect 120484 11734 120598 11786
rect 120650 11734 120652 11786
rect 120484 11732 120652 11734
rect 120484 10892 120540 11732
rect 120596 11722 120652 11732
rect 120372 10836 120540 10892
rect 120708 10892 120764 10902
rect 120260 10668 120316 10678
rect 120260 9548 120316 10612
rect 120260 9482 120316 9492
rect 120372 8652 120428 10836
rect 120484 10666 120540 10678
rect 120484 10614 120486 10666
rect 120538 10614 120540 10666
rect 120484 9782 120540 10614
rect 120484 9772 120596 9782
rect 120484 9716 120540 9772
rect 120540 9678 120596 9716
rect 120372 8586 120428 8596
rect 120708 8652 120764 10836
rect 120820 9996 120876 12292
rect 121940 12236 121996 14200
rect 122500 13914 122556 14758
rect 122696 14200 122808 15000
rect 122948 14476 123004 14486
rect 122500 13862 122502 13914
rect 122554 13862 122556 13914
rect 122500 13850 122556 13862
rect 122276 13018 122332 13030
rect 122276 12966 122278 13018
rect 122330 12966 122332 13018
rect 122164 12236 122220 12246
rect 121940 12170 121996 12180
rect 122052 12180 122164 12236
rect 121380 11788 121436 11798
rect 121044 11338 121100 11350
rect 121044 11286 121046 11338
rect 121098 11286 121100 11338
rect 120932 11004 120988 11014
rect 120932 10668 120988 10948
rect 121044 10892 121100 11286
rect 121044 10826 121100 10836
rect 120932 10602 120988 10612
rect 120820 9940 121324 9996
rect 121044 9772 121100 9782
rect 121044 9678 121100 9716
rect 121268 9772 121324 9940
rect 121380 9994 121436 11732
rect 122052 11564 122108 12180
rect 122164 12170 122220 12180
rect 122276 11900 122332 12966
rect 122500 13018 122556 13030
rect 122500 12966 122502 13018
rect 122554 12966 122556 13018
rect 122500 12122 122556 12966
rect 122724 12348 122780 14200
rect 122948 13914 123004 14420
rect 123368 14200 123480 15000
rect 124152 14200 124264 15000
rect 124404 14476 124460 14486
rect 124460 14420 124572 14476
rect 124404 14410 124460 14420
rect 122948 13862 122950 13914
rect 123002 13862 123004 13914
rect 122948 13850 123004 13862
rect 122724 12282 122780 12292
rect 122948 13020 123004 13030
rect 122500 12070 122502 12122
rect 122554 12070 122556 12122
rect 122500 12058 122556 12070
rect 122724 12122 122780 12134
rect 122724 12070 122726 12122
rect 122778 12070 122780 12122
rect 122724 11900 122780 12070
rect 122276 11844 122780 11900
rect 121716 11508 122108 11564
rect 121380 9942 121382 9994
rect 121434 9942 121436 9994
rect 121380 9930 121436 9942
rect 121604 10666 121660 10678
rect 121604 10614 121606 10666
rect 121658 10614 121660 10666
rect 121268 9706 121324 9716
rect 120708 8586 120764 8596
rect 120932 9324 120988 9334
rect 120260 7756 120316 7766
rect 120148 7700 120260 7756
rect 120260 7690 120316 7700
rect 120932 7654 120988 9268
rect 120876 7644 120988 7654
rect 120372 7642 120988 7644
rect 119252 7532 119532 7588
rect 119700 7578 119756 7588
rect 119924 7586 119980 7598
rect 119364 6300 119420 6310
rect 119252 5964 119308 5974
rect 119252 5906 119308 5908
rect 119252 5854 119254 5906
rect 119306 5854 119308 5906
rect 119252 5842 119308 5854
rect 119364 4060 119420 6244
rect 119364 3994 119420 4004
rect 119140 3110 119142 3162
rect 119194 3110 119196 3162
rect 119140 3098 119196 3110
rect 118916 2538 118972 2548
rect 119028 2828 119084 2838
rect 118916 1708 118972 1718
rect 118692 1652 118916 1708
rect 118916 1642 118972 1652
rect 118468 1596 118524 1606
rect 118468 1146 118524 1540
rect 118468 1094 118470 1146
rect 118522 1094 118524 1146
rect 118468 1082 118524 1094
rect 119028 800 119084 2772
rect 119140 2268 119196 2278
rect 119140 1820 119196 2212
rect 119364 2268 119420 2278
rect 119364 2154 119420 2212
rect 119364 2102 119366 2154
rect 119418 2102 119420 2154
rect 119364 2090 119420 2102
rect 119476 1932 119532 7532
rect 119924 7534 119926 7586
rect 119978 7534 119980 7586
rect 119700 7420 119756 7430
rect 119700 6300 119756 7364
rect 119924 7420 119980 7534
rect 120372 7590 120878 7642
rect 120930 7590 120988 7642
rect 120372 7588 120988 7590
rect 121156 8540 121212 8550
rect 120260 7476 120316 7486
rect 120372 7476 120428 7588
rect 120876 7578 120932 7588
rect 120260 7474 120428 7476
rect 120260 7422 120262 7474
rect 120314 7422 120428 7474
rect 120260 7420 120428 7422
rect 120260 7410 120316 7420
rect 119924 7354 119980 7364
rect 121044 7308 121100 7318
rect 120372 6972 120428 6982
rect 120372 6804 120428 6916
rect 120372 6748 120876 6804
rect 119700 6234 119756 6244
rect 120708 6076 120764 6086
rect 119756 5964 119812 5974
rect 119756 5870 119812 5908
rect 120372 5852 120428 5862
rect 119700 4676 120316 4732
rect 119700 3498 119756 4676
rect 119924 4564 120204 4620
rect 119700 3446 119702 3498
rect 119754 3446 119756 3498
rect 119700 3434 119756 3446
rect 119812 4396 119868 4406
rect 119588 3162 119644 3174
rect 119588 3110 119590 3162
rect 119642 3110 119644 3162
rect 119588 2154 119644 3110
rect 119588 2102 119590 2154
rect 119642 2102 119644 2154
rect 119588 2090 119644 2102
rect 119476 1876 119756 1932
rect 119140 1764 119644 1820
rect 119476 1370 119532 1382
rect 119476 1318 119478 1370
rect 119530 1318 119532 1370
rect 119476 1036 119532 1318
rect 119476 970 119532 980
rect 119588 800 119644 1764
rect 119700 1370 119756 1876
rect 119812 1482 119868 4340
rect 119924 4282 119980 4564
rect 119924 4230 119926 4282
rect 119978 4230 119980 4282
rect 119924 4218 119980 4230
rect 120036 4394 120092 4406
rect 120036 4342 120038 4394
rect 120090 4342 120092 4394
rect 119924 4060 119980 4070
rect 119924 2604 119980 4004
rect 120036 3162 120092 4342
rect 120148 4396 120204 4564
rect 120148 4330 120204 4340
rect 120260 4282 120316 4676
rect 120372 4394 120428 5796
rect 120708 5068 120764 6020
rect 120820 5234 120876 6748
rect 121044 6802 121100 7252
rect 121044 6750 121046 6802
rect 121098 6750 121100 6802
rect 121044 6738 121100 6750
rect 120820 5182 120822 5234
rect 120874 5182 120876 5234
rect 120820 5170 120876 5182
rect 120708 5012 120988 5068
rect 120372 4342 120374 4394
rect 120426 4342 120428 4394
rect 120372 4330 120428 4342
rect 120260 4230 120262 4282
rect 120314 4230 120316 4282
rect 120260 4218 120316 4230
rect 120148 4172 120204 4182
rect 120148 4058 120204 4116
rect 120372 4172 120428 4182
rect 120932 4172 120988 5012
rect 121156 4956 121212 8484
rect 121604 8427 121660 10614
rect 121492 8371 121660 8427
rect 121324 7420 121380 7430
rect 121324 7084 121380 7364
rect 121324 7018 121380 7028
rect 121380 4956 121436 4966
rect 121156 4900 121380 4956
rect 121380 4890 121436 4900
rect 120372 4170 120652 4172
rect 120372 4118 120374 4170
rect 120426 4118 120652 4170
rect 120372 4116 120652 4118
rect 120932 4116 121100 4172
rect 120372 4106 120428 4116
rect 120148 4006 120150 4058
rect 120202 4006 120204 4058
rect 120148 3994 120204 4006
rect 120260 4060 120316 4070
rect 120260 3500 120316 4004
rect 120596 3722 120652 4116
rect 121044 3836 121100 4116
rect 121156 4060 121212 4070
rect 121380 4060 121436 4070
rect 121156 3966 121212 4004
rect 121268 4004 121380 4060
rect 121268 3836 121324 4004
rect 121380 3994 121436 4004
rect 121044 3780 121324 3836
rect 120596 3670 120598 3722
rect 120650 3670 120652 3722
rect 120596 3658 120652 3670
rect 121156 3612 121212 3622
rect 120820 3610 121212 3612
rect 120820 3558 121158 3610
rect 121210 3558 121212 3610
rect 120820 3556 121212 3558
rect 120036 3110 120038 3162
rect 120090 3110 120092 3162
rect 120036 3098 120092 3110
rect 120148 3444 120316 3500
rect 120372 3498 120428 3510
rect 120372 3446 120374 3498
rect 120426 3446 120428 3498
rect 119924 2538 119980 2548
rect 119812 1430 119814 1482
rect 119866 1430 119868 1482
rect 119812 1418 119868 1430
rect 119700 1318 119702 1370
rect 119754 1318 119756 1370
rect 119700 1306 119756 1318
rect 119700 1036 119756 1046
rect 120148 1036 120204 3444
rect 120372 3388 120428 3446
rect 120820 3388 120876 3556
rect 121156 3546 121212 3556
rect 121492 3498 121548 8371
rect 121716 8316 121772 11508
rect 121716 8250 121772 8260
rect 121828 11338 121884 11350
rect 121828 11286 121830 11338
rect 121882 11286 121884 11338
rect 121660 8092 121716 8102
rect 121660 8090 121772 8092
rect 121660 8038 121662 8090
rect 121714 8038 121772 8090
rect 121660 8026 121772 8038
rect 121716 7420 121772 8026
rect 121716 7354 121772 7364
rect 121604 5964 121660 5974
rect 121828 5964 121884 11286
rect 122164 8652 122220 8662
rect 122052 8092 122108 8102
rect 121940 8036 122052 8092
rect 121940 7485 121996 8036
rect 122052 8026 122108 8036
rect 122164 7756 122220 8596
rect 121940 7433 121942 7485
rect 121994 7433 121996 7485
rect 121940 7421 121996 7433
rect 122052 7700 122220 7756
rect 122388 8652 122444 8662
rect 121660 5908 121884 5964
rect 121940 7308 121996 7318
rect 121604 5898 121660 5908
rect 121828 5740 121884 5750
rect 121716 5292 121772 5302
rect 121604 4956 121660 4966
rect 121604 4396 121660 4900
rect 121716 4620 121772 5236
rect 121828 4956 121884 5684
rect 121828 4890 121884 4900
rect 121940 4732 121996 7252
rect 122052 4956 122108 7700
rect 122276 7308 122332 7318
rect 122276 6748 122332 7252
rect 122276 6682 122332 6692
rect 122164 6524 122220 6534
rect 122164 6300 122220 6468
rect 122164 6234 122220 6244
rect 122388 6086 122444 8596
rect 122500 8540 122556 8550
rect 122500 6748 122556 8484
rect 122836 7474 122892 7486
rect 122836 7422 122838 7474
rect 122890 7422 122892 7474
rect 122836 7420 122892 7422
rect 122836 7354 122892 7364
rect 122948 7084 123004 12964
rect 123396 9100 123452 14200
rect 124180 11116 124236 14200
rect 124516 14140 124572 14420
rect 124824 14200 124936 15000
rect 125608 14200 125720 15000
rect 126280 14200 126392 15000
rect 127064 14200 127176 15000
rect 127428 14922 127484 14934
rect 127428 14870 127430 14922
rect 127482 14870 127484 14922
rect 124852 14140 124908 14200
rect 124516 14084 124908 14140
rect 124516 13804 124572 13814
rect 124516 12908 124572 13748
rect 124516 12842 124572 12852
rect 124964 13020 125020 13030
rect 124180 11050 124236 11060
rect 124404 11450 124460 11462
rect 124404 11398 124406 11450
rect 124458 11398 124460 11450
rect 124292 10892 124348 10902
rect 123396 9034 123452 9044
rect 123732 9324 123788 9334
rect 123732 8652 123788 9268
rect 123732 8586 123788 8596
rect 123956 9324 124012 9334
rect 123340 8204 123396 8224
rect 123340 8146 123396 8148
rect 123228 8092 123284 8102
rect 123340 8094 123342 8146
rect 123394 8094 123396 8146
rect 123340 8092 123396 8094
rect 123788 8092 123844 8102
rect 123340 8090 123844 8092
rect 123340 8038 123790 8090
rect 123842 8038 123844 8090
rect 123340 8036 123844 8038
rect 123228 7998 123284 8036
rect 123732 8026 123844 8036
rect 122948 7018 123004 7028
rect 123284 7084 123340 7094
rect 122500 6682 122556 6692
rect 122612 6690 122668 6702
rect 122612 6638 122614 6690
rect 122666 6638 122668 6690
rect 122500 6578 122556 6590
rect 122500 6526 122502 6578
rect 122554 6526 122556 6578
rect 122500 6524 122556 6526
rect 122612 6524 122668 6638
rect 123116 6524 123172 6534
rect 122612 6522 123228 6524
rect 122612 6470 123118 6522
rect 123170 6470 123228 6522
rect 122612 6468 123228 6470
rect 122500 6458 122556 6468
rect 123116 6458 123228 6468
rect 122388 6076 122500 6086
rect 122276 6074 122500 6076
rect 122276 6022 122446 6074
rect 122498 6022 122500 6074
rect 122276 6020 122500 6022
rect 122164 5124 122220 5134
rect 122276 5124 122332 6020
rect 122444 6010 122500 6020
rect 122948 6076 123004 6086
rect 122612 5964 122668 5974
rect 122612 5292 122668 5908
rect 122612 5226 122668 5236
rect 122836 5964 122892 5974
rect 122164 5122 122332 5124
rect 122164 5070 122166 5122
rect 122218 5070 122332 5122
rect 122164 5068 122332 5070
rect 122164 5058 122220 5068
rect 122052 4900 122780 4956
rect 121940 4676 122220 4732
rect 121716 4564 122108 4620
rect 121828 4396 121884 4406
rect 121604 4394 121884 4396
rect 121604 4342 121830 4394
rect 121882 4342 121884 4394
rect 121604 4340 121884 4342
rect 121828 4330 121884 4340
rect 121940 4282 121996 4294
rect 121940 4230 121942 4282
rect 121994 4230 121996 4282
rect 121604 4170 121660 4182
rect 121604 4118 121606 4170
rect 121658 4118 121660 4170
rect 121604 4060 121660 4118
rect 121940 4060 121996 4230
rect 121604 4004 121996 4060
rect 121492 3446 121494 3498
rect 121546 3446 121548 3498
rect 121492 3434 121548 3446
rect 120372 3332 120876 3388
rect 120260 3276 120316 3286
rect 120316 3220 121548 3276
rect 120260 3210 120316 3220
rect 121268 2940 121324 2950
rect 121268 2492 121324 2884
rect 121492 2716 121548 3220
rect 121492 2650 121548 2660
rect 120932 2436 121324 2492
rect 120372 2380 120428 2390
rect 120820 2380 120876 2390
rect 120428 2324 120652 2380
rect 120372 2314 120428 2324
rect 119756 980 120204 1036
rect 120260 1594 120316 1606
rect 120260 1542 120262 1594
rect 120314 1542 120316 1594
rect 119700 970 119756 980
rect 120260 800 120316 1542
rect 120484 1594 120540 1606
rect 120484 1542 120486 1594
rect 120538 1542 120540 1594
rect 120484 1370 120540 1542
rect 120596 1596 120652 2324
rect 120820 1708 120876 2324
rect 120932 2268 120988 2436
rect 121604 2380 121660 2390
rect 121156 2268 121212 2278
rect 120932 2202 120988 2212
rect 121044 2212 121156 2268
rect 120932 2044 120988 2054
rect 121044 2044 121100 2212
rect 121156 2202 121212 2212
rect 120988 1988 121100 2044
rect 121156 2044 121212 2054
rect 120932 1978 120988 1988
rect 121044 1820 121100 1830
rect 121156 1820 121212 1988
rect 121100 1764 121212 1820
rect 121044 1754 121100 1764
rect 120820 1652 120988 1708
rect 120708 1596 120764 1606
rect 120596 1540 120708 1596
rect 120708 1530 120764 1540
rect 120820 1484 120876 1494
rect 120932 1484 120988 1652
rect 120932 1428 121548 1484
rect 120484 1318 120486 1370
rect 120538 1318 120540 1370
rect 120484 1306 120540 1318
rect 120708 1372 120764 1382
rect 120708 1278 120764 1316
rect 120820 800 120876 1428
rect 121268 1146 121324 1158
rect 121268 1094 121270 1146
rect 121322 1094 121324 1146
rect 117012 634 117068 644
rect 117208 0 117320 800
rect 117768 0 117880 800
rect 118328 0 118440 800
rect 119000 0 119112 800
rect 119560 0 119672 800
rect 120232 0 120344 800
rect 120792 0 120904 800
rect 121268 364 121324 1094
rect 121492 800 121548 1428
rect 121604 1370 121660 2324
rect 121604 1318 121606 1370
rect 121658 1318 121660 1370
rect 121604 1306 121660 1318
rect 121716 1146 121772 1158
rect 121716 1094 121718 1146
rect 121770 1094 121772 1146
rect 121268 298 121324 308
rect 121464 0 121576 800
rect 121716 700 121772 1094
rect 122052 800 122108 4564
rect 122164 3498 122220 4676
rect 122164 3446 122166 3498
rect 122218 3446 122220 3498
rect 122164 3434 122220 3446
rect 122612 4394 122668 4406
rect 122612 4342 122614 4394
rect 122666 4342 122668 4394
rect 122612 3500 122668 4342
rect 122612 3434 122668 3444
rect 122164 2828 122220 2838
rect 122164 2604 122220 2772
rect 122164 2538 122220 2548
rect 122724 800 122780 4900
rect 122836 4282 122892 5908
rect 122836 4230 122838 4282
rect 122890 4230 122892 4282
rect 122836 4218 122892 4230
rect 122948 1370 123004 6020
rect 123172 5516 123228 6458
rect 123284 5852 123340 7028
rect 123564 6524 123620 6534
rect 123620 6468 123676 6524
rect 123564 6392 123676 6468
rect 123284 5786 123340 5796
rect 123172 5450 123228 5460
rect 123508 5010 123564 5022
rect 123284 4956 123340 4966
rect 123060 3724 123116 3734
rect 123284 3724 123340 4900
rect 123508 4958 123510 5010
rect 123562 4958 123564 5010
rect 123508 4506 123564 4958
rect 123508 4454 123510 4506
rect 123562 4454 123564 4506
rect 123508 4442 123564 4454
rect 123116 3668 123340 3724
rect 123060 3658 123116 3668
rect 122948 1318 122950 1370
rect 123002 1318 123004 1370
rect 122948 1306 123004 1318
rect 123284 3276 123340 3286
rect 123284 800 123340 3220
rect 123396 1596 123452 1606
rect 123396 1594 123564 1596
rect 123396 1542 123398 1594
rect 123450 1542 123564 1594
rect 123396 1540 123564 1542
rect 123396 1530 123452 1540
rect 121716 634 121772 644
rect 122024 0 122136 800
rect 122696 0 122808 800
rect 123256 0 123368 800
rect 123508 700 123564 1540
rect 123620 1594 123676 6392
rect 123732 5628 123788 8026
rect 123844 7306 123900 7318
rect 123844 7254 123846 7306
rect 123898 7254 123900 7306
rect 123844 6524 123900 7254
rect 123844 6458 123900 6468
rect 123732 5562 123788 5572
rect 123956 5122 124012 9268
rect 123956 5070 123958 5122
rect 124010 5070 124012 5122
rect 123956 4506 124012 5070
rect 123956 4454 123958 4506
rect 124010 4454 124012 4506
rect 123956 4442 124012 4454
rect 124068 8540 124124 8550
rect 123956 4172 124012 4182
rect 124068 4172 124124 8484
rect 124292 4394 124348 10836
rect 124404 6188 124460 11398
rect 124964 11226 125020 12964
rect 124964 11174 124966 11226
rect 125018 11174 125020 11226
rect 124964 11162 125020 11174
rect 125636 11004 125692 14200
rect 125972 13914 126028 13926
rect 125972 13862 125974 13914
rect 126026 13862 126028 13914
rect 125860 12906 125916 12918
rect 125860 12854 125862 12906
rect 125914 12854 125916 12906
rect 125860 11786 125916 12854
rect 125972 11900 126028 13862
rect 126196 13914 126252 13926
rect 126196 13862 126198 13914
rect 126250 13862 126252 13914
rect 126196 13130 126252 13862
rect 126196 13078 126198 13130
rect 126250 13078 126252 13130
rect 126196 13066 126252 13078
rect 126084 11900 126140 11910
rect 125972 11898 126140 11900
rect 125972 11846 126086 11898
rect 126138 11846 126140 11898
rect 125972 11844 126140 11846
rect 126084 11834 126140 11844
rect 125860 11734 125862 11786
rect 125914 11734 125916 11786
rect 125860 11722 125916 11734
rect 126308 11562 126364 14200
rect 126756 13916 126812 13926
rect 126756 13468 126812 13860
rect 126756 13402 126812 13412
rect 126980 13244 127036 13254
rect 126756 13130 126812 13142
rect 126756 13078 126758 13130
rect 126810 13078 126812 13130
rect 126756 12906 126812 13078
rect 126756 12854 126758 12906
rect 126810 12854 126812 12906
rect 126756 12842 126812 12854
rect 126980 12572 127036 13188
rect 126980 12506 127036 12516
rect 127092 11900 127148 14200
rect 127428 12906 127484 14870
rect 127736 14200 127848 15000
rect 128520 14200 128632 15000
rect 129192 14200 129304 15000
rect 129976 14200 130088 15000
rect 130648 14200 130760 15000
rect 131124 14922 131180 14934
rect 131124 14870 131126 14922
rect 131178 14870 131180 14922
rect 127428 12854 127430 12906
rect 127482 12854 127484 12906
rect 127428 12842 127484 12854
rect 127092 11834 127148 11844
rect 127316 12796 127372 12806
rect 126308 11510 126310 11562
rect 126362 11510 126364 11562
rect 126308 11498 126364 11510
rect 126532 11562 126588 11574
rect 126532 11510 126534 11562
rect 126586 11510 126588 11562
rect 125524 10948 125692 11004
rect 125524 10890 125580 10948
rect 125524 10838 125526 10890
rect 125578 10838 125580 10890
rect 125524 10826 125580 10838
rect 125748 10890 125804 10902
rect 125748 10838 125750 10890
rect 125802 10838 125804 10890
rect 125636 10778 125692 10790
rect 125636 10726 125638 10778
rect 125690 10726 125692 10778
rect 125636 9884 125692 10726
rect 125636 9818 125692 9828
rect 125748 9548 125804 10838
rect 125860 10778 125916 10790
rect 125860 10726 125862 10778
rect 125914 10726 125916 10778
rect 125860 10332 125916 10726
rect 126532 10444 126588 11510
rect 126532 10378 126588 10388
rect 125860 10266 125916 10276
rect 125748 9482 125804 9492
rect 127316 10220 127372 12740
rect 127764 11674 127820 14200
rect 127764 11622 127766 11674
rect 127818 11622 127820 11674
rect 127764 11610 127820 11622
rect 127988 11900 128044 11910
rect 124796 8988 124852 8998
rect 124740 8986 124852 8988
rect 124740 8934 124798 8986
rect 124850 8934 124852 8986
rect 124740 8922 124852 8934
rect 124740 8316 124796 8922
rect 124740 6636 124796 8260
rect 124852 8764 124908 8774
rect 127092 8764 127148 8774
rect 124852 6802 124908 8708
rect 126532 8708 127092 8764
rect 126532 8540 126588 8708
rect 127092 8698 127148 8708
rect 126532 8474 126588 8484
rect 125076 8428 125132 8438
rect 125076 8277 125132 8372
rect 125076 8225 125078 8277
rect 125130 8225 125132 8277
rect 125076 8213 125132 8225
rect 125972 8316 126028 8326
rect 125972 8258 126028 8260
rect 125972 8206 125974 8258
rect 126026 8206 126028 8258
rect 126644 8316 126700 8326
rect 125972 8194 126028 8206
rect 126420 8204 126476 8214
rect 125412 7532 125468 7542
rect 125412 7308 125468 7476
rect 125412 7242 125468 7252
rect 124852 6750 124854 6802
rect 124906 6750 124908 6802
rect 124852 6738 124908 6750
rect 126420 6748 126476 8148
rect 126644 7654 126700 8260
rect 127316 7654 127372 10164
rect 127764 11226 127820 11238
rect 127764 11174 127766 11226
rect 127818 11174 127820 11226
rect 127652 8316 127708 8326
rect 127540 8092 127596 8102
rect 127540 7998 127596 8036
rect 126644 7642 126756 7654
rect 127260 7644 127372 7654
rect 126644 7590 126702 7642
rect 126754 7590 126756 7642
rect 126644 7588 126756 7590
rect 126700 7578 126756 7588
rect 126812 7642 127372 7644
rect 126812 7590 127262 7642
rect 127314 7590 127372 7642
rect 126812 7588 127372 7590
rect 126812 7586 126868 7588
rect 126812 7534 126814 7586
rect 126866 7534 126868 7586
rect 127260 7578 127316 7588
rect 126812 7522 126868 7534
rect 124740 6570 124796 6580
rect 126196 6692 126476 6748
rect 126196 6300 126252 6692
rect 126420 6690 126476 6692
rect 126420 6638 126422 6690
rect 126474 6638 126476 6690
rect 126420 6626 126476 6638
rect 126308 6578 126364 6590
rect 126308 6526 126310 6578
rect 126362 6526 126364 6578
rect 126308 6412 126364 6526
rect 127652 6412 127708 8260
rect 126308 6356 127708 6412
rect 126196 6244 126756 6300
rect 124404 6122 124460 6132
rect 126700 6074 126756 6244
rect 126700 6022 126702 6074
rect 126754 6022 126756 6074
rect 126700 6010 126756 6022
rect 127036 6074 127092 6356
rect 127036 6022 127038 6074
rect 127090 6022 127092 6074
rect 127036 6010 127092 6022
rect 127428 5010 127484 5022
rect 125468 4954 125524 4966
rect 125468 4902 125470 4954
rect 125522 4902 125524 4954
rect 125468 4506 125524 4902
rect 125468 4454 125470 4506
rect 125522 4454 125524 4506
rect 125468 4442 125524 4454
rect 126532 4956 126588 4966
rect 124292 4342 124294 4394
rect 124346 4342 124348 4394
rect 124292 4330 124348 4342
rect 125636 4396 125692 4406
rect 124012 4116 124124 4172
rect 124180 4282 124236 4294
rect 124180 4230 124182 4282
rect 124234 4230 124236 4282
rect 124180 4172 124236 4230
rect 123956 4106 124012 4116
rect 124180 4106 124236 4116
rect 125636 3836 125692 4340
rect 126532 4060 126588 4900
rect 126756 4956 126812 4966
rect 126756 4732 126812 4900
rect 126756 4666 126812 4676
rect 127428 4958 127430 5010
rect 127482 4958 127484 5010
rect 127428 4170 127484 4958
rect 127428 4118 127430 4170
rect 127482 4118 127484 4170
rect 127428 4106 127484 4118
rect 127204 4060 127260 4070
rect 126532 4004 127204 4060
rect 127204 3994 127260 4004
rect 125636 3770 125692 3780
rect 127764 3387 127820 11174
rect 127988 8652 128044 11844
rect 128548 11900 128604 14200
rect 129220 11900 129276 14200
rect 128548 11834 128604 11844
rect 129108 11844 129276 11900
rect 129108 11228 129164 11844
rect 129556 11676 129612 11686
rect 129108 11162 129164 11172
rect 129220 11450 129276 11462
rect 129220 11398 129222 11450
rect 129274 11398 129276 11450
rect 129108 10668 129164 10678
rect 129220 10668 129276 11398
rect 129108 10666 129276 10668
rect 129108 10614 129110 10666
rect 129162 10614 129276 10666
rect 129108 10612 129276 10614
rect 129108 10602 129164 10612
rect 129220 10444 129276 10454
rect 129108 10108 129164 10118
rect 129108 9772 129164 10052
rect 129220 9994 129276 10388
rect 129556 10444 129612 11620
rect 130004 11114 130060 14200
rect 130004 11062 130006 11114
rect 130058 11062 130060 11114
rect 130004 11050 130060 11062
rect 130452 11114 130508 11126
rect 130452 11062 130454 11114
rect 130506 11062 130508 11114
rect 130452 10668 130508 11062
rect 129556 10378 129612 10388
rect 130004 10556 130060 10566
rect 129220 9942 129222 9994
rect 129274 9942 129276 9994
rect 129220 9930 129276 9942
rect 130004 9772 130060 10500
rect 129108 9716 129276 9772
rect 128380 9660 128436 9670
rect 128884 9660 128940 9670
rect 128380 9658 128940 9660
rect 128380 9606 128382 9658
rect 128434 9606 128886 9658
rect 128938 9606 128940 9658
rect 128380 9604 128940 9606
rect 128380 9436 128436 9604
rect 128884 9594 128940 9604
rect 128380 9370 128436 9380
rect 127876 8596 128044 8652
rect 127876 7420 127932 8596
rect 127876 7354 127932 7364
rect 127988 8428 128044 8438
rect 127988 6858 128044 8372
rect 129052 8090 129108 8102
rect 129052 8038 129054 8090
rect 129106 8038 129108 8090
rect 128436 7868 128492 7878
rect 128268 7420 128324 7430
rect 127988 6806 127990 6858
rect 128042 6806 128044 6858
rect 127988 6794 128044 6806
rect 128100 7364 128268 7420
rect 127876 4170 127932 4182
rect 127876 4118 127878 4170
rect 127930 4118 127932 4170
rect 127876 3498 127932 4118
rect 128100 4172 128156 7364
rect 128268 7288 128324 7364
rect 128268 6636 128324 6646
rect 128268 6074 128324 6580
rect 128268 6022 128270 6074
rect 128322 6022 128324 6074
rect 128268 6010 128324 6022
rect 128436 6578 128492 7812
rect 129052 7868 129108 8038
rect 129052 7802 129108 7812
rect 129220 7308 129276 9716
rect 129612 9770 130060 9772
rect 129612 9718 130006 9770
rect 130058 9718 130060 9770
rect 129612 9716 130060 9718
rect 129612 9210 129668 9716
rect 130004 9706 130060 9716
rect 130340 9658 130396 9670
rect 130340 9606 130342 9658
rect 130394 9606 130396 9658
rect 129612 9158 129614 9210
rect 129666 9158 129668 9210
rect 129612 9146 129668 9158
rect 130004 9212 130060 9222
rect 129444 7756 129500 7766
rect 129444 7532 129500 7700
rect 129388 7476 129500 7532
rect 129388 7474 129444 7476
rect 129388 7422 129390 7474
rect 129442 7422 129444 7474
rect 129388 7410 129444 7422
rect 129220 7252 129388 7308
rect 129332 6802 129388 7252
rect 129332 6750 129334 6802
rect 129386 6750 129388 6802
rect 129332 6738 129388 6750
rect 128436 6526 128438 6578
rect 128490 6526 128492 6578
rect 128548 6690 128604 6702
rect 128548 6638 128550 6690
rect 128602 6638 128604 6690
rect 128548 6636 128604 6638
rect 128548 6570 128604 6580
rect 128436 4506 128492 6526
rect 129220 6188 129276 6198
rect 129220 6018 129276 6132
rect 129220 5966 129222 6018
rect 129274 5966 129276 6018
rect 129220 5954 129276 5966
rect 129444 6188 129500 6198
rect 128772 5292 128828 5302
rect 128772 5122 128828 5236
rect 128772 5070 128774 5122
rect 128826 5070 128828 5122
rect 128772 5058 128828 5070
rect 129444 5292 129500 6132
rect 129444 4966 129500 5236
rect 129388 4954 129500 4966
rect 129388 4902 129390 4954
rect 129442 4902 129500 4954
rect 129388 4900 129500 4902
rect 129388 4890 129444 4900
rect 130004 4844 130060 9156
rect 130340 9212 130396 9606
rect 130340 9146 130396 9156
rect 130452 8270 130508 10612
rect 130676 8652 130732 14200
rect 131012 12348 131068 12358
rect 130900 10668 130956 10678
rect 130900 10574 130956 10612
rect 130900 10220 130956 10230
rect 131012 10220 131068 12292
rect 131124 12122 131180 14870
rect 131432 14200 131544 15000
rect 132104 14200 132216 15000
rect 132888 14200 133000 15000
rect 133560 14200 133672 15000
rect 134148 14364 134204 14374
rect 131124 12070 131126 12122
rect 131178 12070 131180 12122
rect 131124 12058 131180 12070
rect 130956 10164 131068 10220
rect 131236 11900 131292 11910
rect 130900 10154 130956 10164
rect 131236 9772 131292 11844
rect 131460 11004 131516 14200
rect 131460 10948 131964 11004
rect 131348 10780 131404 10790
rect 131572 10780 131628 10790
rect 131404 10724 131516 10780
rect 131348 10714 131404 10724
rect 130844 9770 131292 9772
rect 130844 9718 131238 9770
rect 131290 9718 131292 9770
rect 130844 9716 131292 9718
rect 130844 9210 130900 9716
rect 131236 9706 131292 9716
rect 131348 10332 131404 10342
rect 131236 9436 131292 9446
rect 131348 9436 131404 10276
rect 131292 9380 131404 9436
rect 131460 10108 131516 10724
rect 131236 9370 131292 9380
rect 130844 9158 130846 9210
rect 130898 9158 130900 9210
rect 130844 9146 130900 9158
rect 131124 9324 131180 9334
rect 130676 8586 130732 8596
rect 130452 8260 130564 8270
rect 130452 8258 131012 8260
rect 130452 8206 130510 8258
rect 130562 8206 131012 8258
rect 130452 8204 131012 8206
rect 130508 8194 130564 8204
rect 130956 8202 131012 8204
rect 130956 8150 130958 8202
rect 131010 8150 131012 8202
rect 130956 8138 131012 8150
rect 130396 8090 130452 8102
rect 130396 8038 130398 8090
rect 130450 8038 130452 8090
rect 130396 7756 130452 8038
rect 130396 7690 130452 7700
rect 130228 7474 130284 7486
rect 130228 7422 130230 7474
rect 130282 7422 130284 7474
rect 130228 7420 130284 7422
rect 130228 7354 130284 7364
rect 130452 7420 130508 7430
rect 130452 6972 130508 7364
rect 130452 6906 130508 6916
rect 130900 6690 130956 6702
rect 130900 6638 130902 6690
rect 130954 6638 130956 6690
rect 130900 6636 130956 6638
rect 130788 6578 130844 6590
rect 130788 6526 130790 6578
rect 130842 6526 130844 6578
rect 130900 6570 130956 6580
rect 130788 6524 130844 6526
rect 130788 6458 130844 6468
rect 131124 6086 131180 9268
rect 131460 9222 131516 10052
rect 131572 9994 131628 10724
rect 131572 9942 131574 9994
rect 131626 9942 131628 9994
rect 131572 9930 131628 9942
rect 131684 10668 131740 10678
rect 131404 9210 131516 9222
rect 131404 9158 131406 9210
rect 131458 9158 131516 9210
rect 131404 9156 131516 9158
rect 131404 9146 131460 9156
rect 131684 8316 131740 10612
rect 131460 8260 131740 8316
rect 131796 9772 131852 9782
rect 131796 9042 131852 9716
rect 131796 8990 131798 9042
rect 131850 8990 131852 9042
rect 131460 6646 131516 8260
rect 131628 8092 131684 8102
rect 131796 8092 131852 8990
rect 131628 8090 131852 8092
rect 131628 8038 131630 8090
rect 131682 8038 131852 8090
rect 131628 8036 131852 8038
rect 131628 8026 131684 8036
rect 131908 6804 131964 10948
rect 132132 10332 132188 14200
rect 132132 10266 132188 10276
rect 132356 13132 132412 13142
rect 132020 10108 132076 10118
rect 132020 9826 132076 10052
rect 132020 9774 132022 9826
rect 132074 9774 132076 9826
rect 132020 9762 132076 9774
rect 132076 8316 132132 8326
rect 132356 8316 132412 13076
rect 132916 12012 132972 14200
rect 132916 11956 133084 12012
rect 132916 11788 132972 11798
rect 132692 11676 132748 11686
rect 132468 11452 132524 11462
rect 132692 11452 132748 11620
rect 132524 11396 132748 11452
rect 132468 11386 132524 11396
rect 132916 11114 132972 11732
rect 132916 11062 132918 11114
rect 132970 11062 132972 11114
rect 132916 11050 132972 11062
rect 132916 10220 132972 10230
rect 132076 8314 132412 8316
rect 132076 8262 132078 8314
rect 132130 8262 132412 8314
rect 132076 8260 132412 8262
rect 132076 8250 132132 8260
rect 132356 8204 132412 8260
rect 132356 8138 132412 8148
rect 132580 9994 132636 10006
rect 132580 9942 132582 9994
rect 132634 9942 132636 9994
rect 132468 7980 132524 7990
rect 132468 7306 132524 7924
rect 132468 7254 132470 7306
rect 132522 7254 132524 7306
rect 132468 7242 132524 7254
rect 132580 6972 132636 9942
rect 132916 9996 132972 10164
rect 132916 9930 132972 9940
rect 132916 8428 132972 8438
rect 132580 6906 132636 6916
rect 132804 7756 132860 7766
rect 131404 6636 131516 6646
rect 131460 6580 131516 6636
rect 131684 6748 131964 6804
rect 132804 6802 132860 7700
rect 132804 6750 132806 6802
rect 132858 6750 132860 6802
rect 131404 6504 131460 6580
rect 131684 6300 131740 6748
rect 132804 6738 132860 6750
rect 131852 6524 131908 6534
rect 131908 6468 131964 6524
rect 131852 6392 131964 6468
rect 131684 6244 131852 6300
rect 130900 6076 130956 6086
rect 130564 5964 130620 5974
rect 130564 5906 130620 5908
rect 130564 5854 130566 5906
rect 130618 5854 130620 5906
rect 130564 5842 130620 5854
rect 130004 4778 130060 4788
rect 128436 4454 128438 4506
rect 128490 4454 128492 4506
rect 128436 4442 128492 4454
rect 128100 4106 128156 4116
rect 127876 3446 127878 3498
rect 127930 3446 127932 3498
rect 127876 3434 127932 3446
rect 129556 3836 129612 3846
rect 127652 3331 127820 3387
rect 125860 3052 125916 3062
rect 125860 2716 125916 2996
rect 125860 2650 125916 2660
rect 126084 2716 126140 2726
rect 125412 2492 125468 2502
rect 125468 2436 125580 2492
rect 125412 2426 125468 2436
rect 123620 1542 123622 1594
rect 123674 1542 123676 1594
rect 123620 1530 123676 1542
rect 123844 1932 123900 1942
rect 123844 800 123900 1876
rect 124516 1820 124572 1830
rect 124516 800 124572 1764
rect 125300 1146 125356 1158
rect 125300 1094 125302 1146
rect 125354 1094 125356 1146
rect 124852 868 125132 924
rect 123508 634 123564 644
rect 123816 0 123928 800
rect 124488 0 124600 800
rect 124740 476 124796 486
rect 124852 476 124908 868
rect 125076 800 125132 868
rect 124796 420 124908 476
rect 124740 410 124796 420
rect 125048 0 125160 800
rect 125300 588 125356 1094
rect 125524 1146 125580 2436
rect 125860 2266 125916 2278
rect 125860 2214 125862 2266
rect 125914 2214 125916 2266
rect 125860 1932 125916 2214
rect 125860 1866 125916 1876
rect 126084 1372 126140 2660
rect 126756 2716 126812 2726
rect 127316 2716 127372 2726
rect 126756 2714 127372 2716
rect 126756 2662 126758 2714
rect 126810 2662 127318 2714
rect 127370 2662 127372 2714
rect 126756 2660 127372 2662
rect 126756 2650 126812 2660
rect 127316 2650 127372 2660
rect 127652 2716 127708 3331
rect 129332 2940 129388 2950
rect 127652 2650 127708 2660
rect 128772 2828 128828 2838
rect 127764 2492 127820 2502
rect 127820 2436 127932 2492
rect 127764 2426 127820 2436
rect 126420 2380 126476 2390
rect 126756 2380 126812 2390
rect 126420 2378 126812 2380
rect 126420 2326 126422 2378
rect 126474 2326 126758 2378
rect 126810 2326 126812 2378
rect 126420 2324 126812 2326
rect 126420 2314 126476 2324
rect 126756 2314 126812 2324
rect 126084 1306 126140 1316
rect 126308 2154 126364 2166
rect 126308 2102 126310 2154
rect 126362 2102 126364 2154
rect 126308 1372 126364 2102
rect 127652 2156 127708 2166
rect 127652 2062 127708 2100
rect 127876 2156 127932 2436
rect 127876 2090 127932 2100
rect 126308 1306 126364 1316
rect 128212 1820 128268 1830
rect 125524 1094 125526 1146
rect 125578 1094 125580 1146
rect 125524 1082 125580 1094
rect 125748 1260 125804 1270
rect 125748 800 125804 1204
rect 127540 1260 127596 1270
rect 126308 1146 126364 1158
rect 126308 1094 126310 1146
rect 126362 1094 126364 1146
rect 126308 800 126364 1094
rect 126980 1148 127036 1158
rect 126980 800 127036 1092
rect 127540 800 127596 1204
rect 128212 800 128268 1764
rect 128772 800 128828 2772
rect 129332 800 129388 2884
rect 129556 2380 129612 3780
rect 130900 3498 130956 6020
rect 131068 6074 131180 6086
rect 131068 6022 131070 6074
rect 131122 6022 131180 6074
rect 131068 6020 131180 6022
rect 131068 5964 131124 6020
rect 131068 5898 131124 5908
rect 131628 5852 131684 5862
rect 131628 5850 131740 5852
rect 131628 5798 131630 5850
rect 131682 5798 131740 5850
rect 131628 5786 131740 5798
rect 131460 5010 131516 5022
rect 131460 4958 131462 5010
rect 131514 4958 131516 5010
rect 130900 3446 130902 3498
rect 130954 3446 130956 3498
rect 130900 3434 130956 3446
rect 131236 3834 131292 3846
rect 131236 3782 131238 3834
rect 131290 3782 131292 3834
rect 129556 2314 129612 2324
rect 130900 2828 130956 2838
rect 130900 2266 130956 2772
rect 130900 2214 130902 2266
rect 130954 2214 130956 2266
rect 130900 2202 130956 2214
rect 130564 1148 130620 1158
rect 130004 1034 130060 1046
rect 130004 982 130006 1034
rect 130058 982 130060 1034
rect 130004 800 130060 982
rect 130564 800 130620 1092
rect 131236 800 131292 3782
rect 131460 3610 131516 4958
rect 131460 3558 131462 3610
rect 131514 3558 131516 3610
rect 131460 3546 131516 3558
rect 131684 3164 131740 5786
rect 131796 4170 131852 6244
rect 131796 4118 131798 4170
rect 131850 4118 131852 4170
rect 131796 4106 131852 4118
rect 131684 3098 131740 3108
rect 131908 2940 131964 6392
rect 132076 5852 132132 5862
rect 132076 5850 132188 5852
rect 132076 5798 132078 5850
rect 132130 5798 132188 5850
rect 132076 5786 132188 5798
rect 132020 4170 132076 4182
rect 132020 4118 132022 4170
rect 132074 4118 132076 4170
rect 132020 3836 132076 4118
rect 132020 3770 132076 3780
rect 131908 2874 131964 2884
rect 132020 3610 132076 3622
rect 132020 3558 132022 3610
rect 132074 3558 132076 3610
rect 131796 1708 131852 1718
rect 131796 800 131852 1652
rect 125300 522 125356 532
rect 125720 0 125832 800
rect 126280 0 126392 800
rect 126952 0 127064 800
rect 127512 0 127624 800
rect 128184 0 128296 800
rect 128744 0 128856 800
rect 129304 0 129416 800
rect 129976 0 130088 800
rect 130536 0 130648 800
rect 131208 0 131320 800
rect 131768 0 131880 800
rect 132020 588 132076 3558
rect 132132 2716 132188 5786
rect 132524 5850 132580 5862
rect 132524 5798 132526 5850
rect 132578 5798 132580 5850
rect 132524 5628 132580 5798
rect 132524 5562 132580 5572
rect 132356 5292 132412 5302
rect 132356 3722 132412 5236
rect 132580 5122 132636 5134
rect 132580 5070 132582 5122
rect 132634 5070 132636 5122
rect 132580 4844 132636 5070
rect 132580 4778 132636 4788
rect 132356 3670 132358 3722
rect 132410 3670 132412 3722
rect 132356 3658 132412 3670
rect 132692 3500 132748 3510
rect 132244 3276 132300 3286
rect 132692 3276 132748 3444
rect 132300 3220 132748 3276
rect 132804 3386 132860 3398
rect 132804 3334 132806 3386
rect 132858 3334 132860 3386
rect 132244 3210 132300 3220
rect 132691 3052 132747 3062
rect 132468 2996 132691 3052
rect 132468 2938 132524 2996
rect 132691 2986 132747 2996
rect 132468 2886 132470 2938
rect 132522 2886 132524 2938
rect 132468 2874 132524 2886
rect 132804 2938 132860 3334
rect 132916 3387 132972 8372
rect 133028 5516 133084 11956
rect 133588 11676 133644 14200
rect 134148 14026 134204 14308
rect 134344 14200 134456 15000
rect 134708 14364 134764 14374
rect 134148 13974 134150 14026
rect 134202 13974 134204 14026
rect 134148 13962 134204 13974
rect 134372 14028 134428 14200
rect 134372 13972 134540 14028
rect 134260 13916 134316 13926
rect 134260 13914 134428 13916
rect 134260 13862 134262 13914
rect 134314 13862 134428 13914
rect 134260 13860 134428 13862
rect 134260 13850 134316 13860
rect 134148 12124 134204 12134
rect 133588 11610 133644 11620
rect 134036 11674 134092 11686
rect 134036 11622 134038 11674
rect 134090 11622 134092 11674
rect 133588 11116 133644 11126
rect 133588 11022 133644 11060
rect 133924 10556 133980 10566
rect 133924 10462 133980 10500
rect 133140 10444 133196 10454
rect 133140 9996 133196 10388
rect 133140 9930 133196 9940
rect 133588 10444 133644 10454
rect 133476 9826 133532 9838
rect 133476 9774 133478 9826
rect 133530 9774 133532 9826
rect 133476 9100 133532 9774
rect 133252 9044 133476 9100
rect 133252 9042 133308 9044
rect 133252 8990 133254 9042
rect 133306 8990 133308 9042
rect 133476 9034 133532 9044
rect 133252 8978 133308 8990
rect 133140 8930 133196 8942
rect 133140 8878 133142 8930
rect 133194 8878 133196 8930
rect 133140 8092 133196 8878
rect 133588 8876 133644 10388
rect 134036 10444 134092 11622
rect 134148 10556 134204 12068
rect 134372 12124 134428 13860
rect 134484 13020 134540 13972
rect 134708 13914 134764 14308
rect 135016 14200 135128 15000
rect 135800 14200 135912 15000
rect 136276 14362 136332 14374
rect 136276 14310 136278 14362
rect 136330 14310 136332 14362
rect 134708 13862 134710 13914
rect 134762 13862 134764 13914
rect 134708 13850 134764 13862
rect 134484 12954 134540 12964
rect 134372 12058 134428 12068
rect 134932 12012 134988 12022
rect 134260 11900 134316 11910
rect 134260 11228 134316 11844
rect 134260 11162 134316 11172
rect 134148 10490 134204 10500
rect 134820 10778 134876 10790
rect 134820 10726 134822 10778
rect 134874 10726 134876 10778
rect 134036 10378 134092 10388
rect 134260 10444 134316 10454
rect 134260 10350 134316 10388
rect 134484 10444 134540 10454
rect 134372 10332 134428 10342
rect 134092 9658 134148 9670
rect 134092 9606 134094 9658
rect 134146 9606 134148 9658
rect 133476 8820 133644 8876
rect 133924 9100 133980 9110
rect 133364 8652 133420 8662
rect 133252 8204 133308 8214
rect 133252 8110 133308 8148
rect 133140 8026 133196 8036
rect 133364 7474 133420 8596
rect 133364 7422 133366 7474
rect 133418 7422 133420 7474
rect 133364 7410 133420 7422
rect 133140 5794 133196 5806
rect 133140 5742 133142 5794
rect 133194 5742 133196 5794
rect 133140 5740 133196 5742
rect 133140 5674 133196 5684
rect 133028 5450 133084 5460
rect 133476 5180 133532 8820
rect 133700 8764 133756 8774
rect 133588 8316 133644 8326
rect 133700 8316 133756 8708
rect 133588 8314 133756 8316
rect 133588 8262 133590 8314
rect 133642 8262 133756 8314
rect 133588 8260 133756 8262
rect 133924 8326 133980 9044
rect 134092 9100 134148 9606
rect 134092 9034 134148 9044
rect 134260 9042 134316 9054
rect 134260 8990 134262 9042
rect 134314 8990 134316 9042
rect 134260 8988 134316 8990
rect 134260 8922 134316 8932
rect 133924 8314 134036 8326
rect 133924 8262 133982 8314
rect 134034 8262 134036 8314
rect 133588 8250 133644 8260
rect 133924 8250 134036 8262
rect 133924 8204 133980 8250
rect 133812 8148 133980 8204
rect 133812 8092 133868 8148
rect 133588 8036 133868 8092
rect 133588 7586 133644 8036
rect 133588 7534 133590 7586
rect 133642 7534 133644 7586
rect 133588 7522 133644 7534
rect 133812 7532 133868 7542
rect 133812 7306 133868 7476
rect 133812 7254 133814 7306
rect 133866 7254 133868 7306
rect 133812 7242 133868 7254
rect 134372 6690 134428 10276
rect 134484 7980 134540 10388
rect 134820 8316 134876 10726
rect 134932 10668 134988 11956
rect 135044 11116 135100 14200
rect 135828 13804 135884 14200
rect 135492 13748 135884 13804
rect 135380 12124 135436 12134
rect 135380 11450 135436 12068
rect 135380 11398 135382 11450
rect 135434 11398 135436 11450
rect 135380 11386 135436 11398
rect 135044 11050 135100 11060
rect 135156 11116 135212 11126
rect 135268 11116 135324 11126
rect 135156 11114 135268 11116
rect 135156 11062 135158 11114
rect 135210 11062 135268 11114
rect 135156 11060 135268 11062
rect 135156 11050 135212 11060
rect 135268 11050 135324 11060
rect 135380 11114 135436 11126
rect 135380 11062 135382 11114
rect 135434 11062 135436 11114
rect 135380 10892 135436 11062
rect 135492 11004 135548 13748
rect 135492 10938 135548 10948
rect 135604 13580 135660 13590
rect 135380 10826 135436 10836
rect 135604 10892 135660 13524
rect 135828 13020 135884 13030
rect 135716 11562 135772 11574
rect 135716 11510 135718 11562
rect 135770 11510 135772 11562
rect 135716 11002 135772 11510
rect 135716 10950 135718 11002
rect 135770 10950 135772 11002
rect 135716 10938 135772 10950
rect 135604 10826 135660 10836
rect 135828 10780 135884 12964
rect 136276 12122 136332 14310
rect 136472 14200 136584 15000
rect 136724 14308 137116 14364
rect 136276 12070 136278 12122
rect 136330 12070 136332 12122
rect 136276 12058 136332 12070
rect 135940 11452 135996 11462
rect 135940 11002 135996 11396
rect 135940 10950 135942 11002
rect 135994 10950 135996 11002
rect 135940 10938 135996 10950
rect 135828 10714 135884 10724
rect 136388 10778 136444 10790
rect 136388 10726 136390 10778
rect 136442 10726 136444 10778
rect 134932 10612 135660 10668
rect 135492 9994 135548 10006
rect 135492 9942 135494 9994
rect 135546 9942 135548 9994
rect 134932 9884 134988 9894
rect 134932 9826 134988 9828
rect 134932 9774 134934 9826
rect 134986 9774 134988 9826
rect 134932 9762 134988 9774
rect 135492 9772 135548 9942
rect 135492 9706 135548 9716
rect 134484 7914 134540 7924
rect 134596 8247 134652 8259
rect 134820 8250 134876 8260
rect 134932 9436 134988 9446
rect 134596 8195 134598 8247
rect 134650 8195 134652 8247
rect 134596 7644 134652 8195
rect 134596 7578 134652 7588
rect 134820 6860 134876 6870
rect 134820 6802 134876 6804
rect 134820 6750 134822 6802
rect 134874 6750 134876 6802
rect 134820 6738 134876 6750
rect 134372 6638 134374 6690
rect 134426 6638 134428 6690
rect 133252 5124 133532 5180
rect 133812 6578 133868 6590
rect 133812 6526 133814 6578
rect 133866 6526 133868 6578
rect 133812 5190 133868 6526
rect 134148 6300 134204 6310
rect 134148 5292 134204 6244
rect 134260 5906 134316 5918
rect 134260 5854 134262 5906
rect 134314 5854 134316 5906
rect 134260 5628 134316 5854
rect 134260 5404 134316 5572
rect 134260 5338 134316 5348
rect 134148 5226 134204 5236
rect 134372 5190 134428 6638
rect 133812 5180 133924 5190
rect 133812 5178 133980 5180
rect 133812 5126 133870 5178
rect 133922 5126 133980 5178
rect 133812 5124 133980 5126
rect 133252 4394 133308 5124
rect 133868 5114 133980 5124
rect 134316 5178 134428 5190
rect 134316 5126 134318 5178
rect 134370 5126 134428 5178
rect 134316 5124 134428 5126
rect 134316 5114 134372 5124
rect 133420 4954 133476 4966
rect 133420 4902 133422 4954
rect 133474 4902 133476 4954
rect 133420 4844 133476 4902
rect 133420 4778 133476 4788
rect 133252 4342 133254 4394
rect 133306 4342 133308 4394
rect 133252 4330 133308 4342
rect 133588 4506 133644 4518
rect 133588 4454 133590 4506
rect 133642 4454 133644 4506
rect 133476 3498 133532 3510
rect 133476 3446 133478 3498
rect 133530 3446 133532 3498
rect 132916 3331 133084 3387
rect 132804 2886 132806 2938
rect 132858 2886 132860 2938
rect 132804 2874 132860 2886
rect 132692 2828 132748 2838
rect 132692 2716 132748 2772
rect 132916 2716 132972 2726
rect 132692 2660 132916 2716
rect 132132 2650 132188 2660
rect 132916 2650 132972 2660
rect 132804 1820 132860 1830
rect 132860 1764 132972 1820
rect 132804 1754 132860 1764
rect 132468 1594 132524 1606
rect 132468 1542 132470 1594
rect 132522 1542 132524 1594
rect 132468 800 132524 1542
rect 132916 1596 132972 1764
rect 132916 1530 132972 1540
rect 133028 800 133084 3331
rect 133476 3050 133532 3446
rect 133476 2998 133478 3050
rect 133530 2998 133532 3050
rect 133476 2986 133532 2998
rect 133364 2380 133420 2390
rect 133364 2044 133420 2324
rect 133364 1978 133420 1988
rect 133588 1596 133644 4454
rect 133700 4508 133756 4518
rect 133700 3276 133756 4452
rect 133700 3210 133756 3220
rect 133924 1708 133980 5114
rect 134148 4060 134204 4070
rect 134148 3966 134204 4004
rect 134820 4060 134876 4070
rect 134260 3946 134316 3958
rect 134260 3894 134262 3946
rect 134314 3894 134316 3946
rect 134036 3722 134092 3734
rect 134036 3670 134038 3722
rect 134090 3670 134092 3722
rect 134036 3500 134092 3670
rect 134036 3434 134092 3444
rect 134260 3500 134316 3894
rect 134260 3434 134316 3444
rect 134372 3834 134428 3846
rect 134372 3782 134374 3834
rect 134426 3782 134428 3834
rect 134148 3276 134204 3286
rect 134148 3164 134204 3220
rect 134036 3108 134204 3164
rect 134036 2828 134092 3108
rect 134036 2762 134092 2772
rect 134148 2940 134204 2950
rect 133924 1642 133980 1652
rect 133588 1540 133756 1596
rect 133700 800 133756 1540
rect 133924 1034 133980 1046
rect 133924 982 133926 1034
rect 133978 982 133980 1034
rect 133924 924 133980 982
rect 134148 924 134204 2884
rect 134260 2380 134316 2390
rect 134260 2286 134316 2324
rect 134372 1596 134428 3782
rect 134820 3722 134876 4004
rect 134820 3670 134822 3722
rect 134874 3670 134876 3722
rect 134820 3658 134876 3670
rect 134932 3724 134988 9380
rect 135268 9100 135324 9110
rect 135268 9042 135324 9044
rect 135268 8990 135270 9042
rect 135322 8990 135324 9042
rect 135268 8978 135324 8990
rect 135380 8930 135436 8942
rect 135380 8878 135382 8930
rect 135434 8878 135436 8930
rect 135156 8652 135212 8662
rect 135156 7654 135212 8596
rect 135380 8428 135436 8878
rect 135604 8428 135660 10612
rect 135940 9714 135996 9726
rect 135940 9662 135942 9714
rect 135994 9662 135996 9714
rect 135772 8988 135828 8998
rect 135772 8894 135828 8932
rect 135940 8988 135996 9662
rect 135604 8372 135772 8428
rect 135380 8362 135436 8372
rect 135492 8258 135548 8270
rect 135492 8206 135494 8258
rect 135546 8206 135548 8258
rect 135156 7642 135268 7654
rect 135156 7590 135214 7642
rect 135266 7590 135268 7642
rect 135156 7588 135268 7590
rect 135212 7578 135268 7588
rect 135492 6748 135548 8206
rect 135268 6692 135548 6748
rect 135268 6524 135324 6692
rect 135100 6468 135324 6524
rect 135380 6578 135436 6590
rect 135380 6526 135382 6578
rect 135434 6526 135436 6578
rect 135100 6074 135156 6468
rect 135100 6022 135102 6074
rect 135154 6022 135156 6074
rect 135100 5964 135156 6022
rect 135100 5898 135156 5908
rect 135268 5068 135324 5078
rect 135268 5010 135324 5012
rect 135268 4958 135270 5010
rect 135322 4958 135324 5010
rect 135268 4946 135324 4958
rect 135380 4956 135436 6526
rect 135548 5964 135604 6002
rect 135548 5898 135604 5908
rect 135604 5740 135660 5750
rect 135604 4956 135660 5684
rect 135380 4900 135548 4956
rect 135044 3724 135100 3734
rect 134932 3722 135100 3724
rect 134932 3670 135046 3722
rect 135098 3670 135100 3722
rect 134932 3668 135100 3670
rect 135044 3658 135100 3668
rect 134372 1530 134428 1540
rect 134484 3388 134540 3398
rect 134148 868 134316 924
rect 133924 858 133980 868
rect 134260 800 134316 868
rect 132020 522 132076 532
rect 132440 0 132552 800
rect 133000 0 133112 800
rect 133672 0 133784 800
rect 134232 0 134344 800
rect 134484 588 134540 3332
rect 134820 3276 134876 3286
rect 135380 3276 135436 3286
rect 134876 3220 135380 3276
rect 134820 3210 134876 3220
rect 135380 3210 135436 3220
rect 134596 3164 134652 3174
rect 134596 2940 134652 3108
rect 134596 2874 134652 2884
rect 135492 2940 135548 4900
rect 135604 4890 135660 4900
rect 135716 3388 135772 8372
rect 135940 7868 135996 8932
rect 135828 7812 135996 7868
rect 136276 8764 136332 8774
rect 135828 6860 135884 7812
rect 135996 7644 136052 7654
rect 135996 7550 136052 7588
rect 136108 7474 136164 7486
rect 136108 7422 136110 7474
rect 136162 7422 136164 7474
rect 136108 6972 136164 7422
rect 136108 6906 136164 6916
rect 135828 6804 135996 6860
rect 136276 6804 136332 8708
rect 135828 6690 135884 6702
rect 135828 6638 135830 6690
rect 135882 6638 135884 6690
rect 135828 4058 135884 6638
rect 135940 6086 135996 6804
rect 136164 6748 136332 6804
rect 135940 6074 136052 6086
rect 135940 6022 135998 6074
rect 136050 6022 136052 6074
rect 135940 6010 136052 6022
rect 135940 5964 135996 6010
rect 135940 5898 135996 5908
rect 136164 4170 136220 6748
rect 136164 4118 136166 4170
rect 136218 4118 136220 4170
rect 136164 4106 136220 4118
rect 136276 6636 136332 6646
rect 135828 4006 135830 4058
rect 135882 4006 135884 4058
rect 135828 3994 135884 4006
rect 135716 3322 135772 3332
rect 136164 3836 136220 3846
rect 134820 1708 134876 1718
rect 134820 800 134876 1652
rect 135044 1372 135100 1382
rect 135044 1278 135100 1316
rect 135492 800 135548 2884
rect 136052 3276 136108 3286
rect 136052 800 136108 3220
rect 136164 1708 136220 3780
rect 136276 2268 136332 6580
rect 136276 2202 136332 2212
rect 136388 2156 136444 10726
rect 136500 10220 136556 14200
rect 136500 10154 136556 10164
rect 136612 11338 136668 11350
rect 136612 11286 136614 11338
rect 136666 11286 136668 11338
rect 136500 6972 136556 6982
rect 136500 4732 136556 6916
rect 136612 5964 136668 11286
rect 136724 9996 136780 14308
rect 137060 14140 137116 14308
rect 137256 14200 137368 15000
rect 137928 14200 138040 15000
rect 138712 14200 138824 15000
rect 138964 14586 139020 14598
rect 138964 14534 138966 14586
rect 139018 14534 139020 14586
rect 137284 14140 137340 14200
rect 137060 14084 137340 14140
rect 137396 12908 137452 12918
rect 137396 12796 137452 12852
rect 137844 12796 137900 12806
rect 137396 12740 137844 12796
rect 137844 12730 137900 12740
rect 137620 12012 137676 12022
rect 136724 9930 136780 9940
rect 136836 10442 136892 10454
rect 136836 10390 136838 10442
rect 136890 10390 136892 10442
rect 136836 7644 136892 10390
rect 137032 10220 137296 10230
rect 137088 10164 137136 10220
rect 137192 10164 137240 10220
rect 137032 10154 137296 10164
rect 137620 10220 137676 11956
rect 137956 11900 138012 14200
rect 138516 14026 138572 14038
rect 138516 13974 138518 14026
rect 138570 13974 138572 14026
rect 138292 13916 138348 13926
rect 137956 11834 138012 11844
rect 138068 13860 138292 13916
rect 137732 11676 137788 11686
rect 137732 10554 137788 11620
rect 138068 11452 138124 13860
rect 138292 13850 138348 13860
rect 138516 13578 138572 13974
rect 138740 13916 138796 14200
rect 138740 13850 138796 13860
rect 138516 13526 138518 13578
rect 138570 13526 138572 13578
rect 138516 13514 138572 13526
rect 138740 13468 138796 13478
rect 138628 13466 138796 13468
rect 138628 13414 138742 13466
rect 138794 13414 138796 13466
rect 138628 13412 138796 13414
rect 138628 13356 138684 13412
rect 138740 13402 138796 13412
rect 138180 13300 138684 13356
rect 138180 13018 138236 13300
rect 138964 13242 139020 14534
rect 139384 14200 139496 15000
rect 140168 14200 140280 15000
rect 140840 14200 140952 15000
rect 141092 14362 141148 14374
rect 141092 14310 141094 14362
rect 141146 14310 141148 14362
rect 138964 13190 138966 13242
rect 139018 13190 139020 13242
rect 138964 13178 139020 13190
rect 139076 13578 139132 13590
rect 139076 13526 139078 13578
rect 139130 13526 139132 13578
rect 138180 12966 138182 13018
rect 138234 12966 138236 13018
rect 138180 12954 138236 12966
rect 138404 13018 138460 13030
rect 138404 12966 138406 13018
rect 138458 12966 138460 13018
rect 138404 12682 138460 12966
rect 138404 12630 138406 12682
rect 138458 12630 138460 12682
rect 138404 12618 138460 12630
rect 139076 12682 139132 13526
rect 139076 12630 139078 12682
rect 139130 12630 139132 12682
rect 139076 12618 139132 12630
rect 139188 12122 139244 12134
rect 139188 12070 139190 12122
rect 139242 12070 139244 12122
rect 138852 12010 138908 12022
rect 138852 11958 138854 12010
rect 138906 11958 138908 12010
rect 138852 11788 138908 11958
rect 138292 11676 138348 11686
rect 138292 11582 138348 11620
rect 138516 11674 138572 11686
rect 138516 11622 138518 11674
rect 138570 11622 138572 11674
rect 137732 10502 137734 10554
rect 137786 10502 137788 10554
rect 137732 10490 137788 10502
rect 137956 11396 138124 11452
rect 137060 9996 137116 10006
rect 137060 9770 137116 9940
rect 137396 9996 137452 10006
rect 137396 9902 137452 9940
rect 137060 9718 137062 9770
rect 137114 9718 137116 9770
rect 137060 9706 137116 9718
rect 137396 9212 137452 9222
rect 137396 8874 137452 9156
rect 137620 9042 137676 10164
rect 137788 9884 137844 9894
rect 137788 9790 137844 9828
rect 137956 9436 138012 11396
rect 137956 9370 138012 9380
rect 138068 11226 138124 11238
rect 138068 11174 138070 11226
rect 138122 11174 138124 11226
rect 137620 8990 137622 9042
rect 137674 8990 137676 9042
rect 137620 8978 137676 8990
rect 137396 8822 137398 8874
rect 137450 8822 137452 8874
rect 137396 8810 137452 8822
rect 137032 8652 137296 8662
rect 137088 8596 137136 8652
rect 137192 8596 137240 8652
rect 137032 8586 137296 8596
rect 137620 8316 137676 8326
rect 136724 7588 136892 7644
rect 136948 8092 137004 8102
rect 136724 6860 136780 7588
rect 136948 7474 137004 8036
rect 137284 8092 137340 8102
rect 137284 8090 137564 8092
rect 137284 8038 137286 8090
rect 137338 8038 137564 8090
rect 137284 8036 137564 8038
rect 137284 8026 137340 8036
rect 136948 7422 136950 7474
rect 137002 7422 137004 7474
rect 136948 7410 137004 7422
rect 137396 7306 137452 7318
rect 137396 7254 137398 7306
rect 137450 7254 137452 7306
rect 137032 7084 137296 7094
rect 137088 7028 137136 7084
rect 137192 7028 137240 7084
rect 137032 7018 137296 7028
rect 136724 6804 137228 6860
rect 136612 5898 136668 5908
rect 136948 6690 137004 6702
rect 136948 6638 136950 6690
rect 137002 6638 137004 6690
rect 136948 5740 137004 6638
rect 137172 6690 137228 6804
rect 137172 6638 137174 6690
rect 137226 6638 137228 6690
rect 137172 6626 137228 6638
rect 137396 5964 137452 7254
rect 137508 7084 137564 8036
rect 137508 7018 137564 7028
rect 137620 6018 137676 8260
rect 137844 6858 137900 6870
rect 137844 6806 137846 6858
rect 137898 6806 137900 6858
rect 137620 5966 137622 6018
rect 137674 5966 137676 6018
rect 137396 5908 137564 5964
rect 137620 5954 137676 5966
rect 137732 6076 137788 6086
rect 136836 5684 137004 5740
rect 136612 5180 136668 5190
rect 136612 5122 136668 5124
rect 136612 5070 136614 5122
rect 136666 5070 136668 5122
rect 136612 5058 136668 5070
rect 136500 4666 136556 4676
rect 136724 3724 136780 3734
rect 136500 3276 136556 3286
rect 136724 3276 136780 3668
rect 136556 3220 136668 3276
rect 136500 3210 136556 3220
rect 136612 3052 136668 3220
rect 136724 3210 136780 3220
rect 136836 3052 136892 5684
rect 137508 5628 137564 5908
rect 137508 5562 137564 5572
rect 137032 5516 137296 5526
rect 137088 5460 137136 5516
rect 137192 5460 137240 5516
rect 137032 5450 137296 5460
rect 137620 5516 137676 5526
rect 137620 5190 137676 5460
rect 137564 5178 137676 5190
rect 137564 5126 137566 5178
rect 137618 5126 137676 5178
rect 137564 5124 137676 5126
rect 137564 5114 137620 5124
rect 137116 4954 137172 4966
rect 137116 4902 137118 4954
rect 137170 4902 137172 4954
rect 137116 4732 137172 4902
rect 137116 4666 137172 4676
rect 137284 4732 137340 4742
rect 136612 2996 136892 3052
rect 136724 2268 136780 2278
rect 136388 2100 136556 2156
rect 136388 1932 136444 1942
rect 136388 1818 136444 1876
rect 136388 1766 136390 1818
rect 136442 1766 136444 1818
rect 136388 1754 136444 1766
rect 136164 1642 136220 1652
rect 136500 1482 136556 2100
rect 136500 1430 136502 1482
rect 136554 1430 136556 1482
rect 136500 1418 136556 1430
rect 136724 800 136780 2212
rect 137172 1372 137228 1382
rect 137172 1036 137228 1316
rect 137172 970 137228 980
rect 137284 800 137340 4676
rect 137732 4170 137788 6020
rect 137844 5852 137900 6806
rect 137844 5786 137900 5796
rect 138068 5740 138124 11174
rect 138516 10890 138572 11622
rect 138516 10838 138518 10890
rect 138570 10838 138572 10890
rect 138516 10826 138572 10838
rect 138628 11450 138684 11462
rect 138628 11398 138630 11450
rect 138682 11398 138684 11450
rect 138292 9042 138348 9054
rect 138292 8990 138294 9042
rect 138346 8990 138348 9042
rect 138292 8988 138348 8990
rect 138292 7474 138348 8932
rect 138628 8540 138684 11398
rect 138852 9042 138908 11732
rect 138964 11226 139020 11238
rect 138964 11174 138966 11226
rect 139018 11174 139020 11226
rect 138964 10890 139020 11174
rect 138964 10838 138966 10890
rect 139018 10838 139020 10890
rect 138964 10826 139020 10838
rect 138964 9660 139020 9670
rect 138964 9658 139132 9660
rect 138964 9606 138966 9658
rect 139018 9606 139132 9658
rect 138964 9604 139132 9606
rect 138964 9594 139020 9604
rect 138852 8990 138854 9042
rect 138906 8990 138908 9042
rect 138852 8978 138908 8990
rect 138852 8540 138908 8550
rect 138628 8484 138852 8540
rect 138852 8474 138908 8484
rect 138292 7422 138294 7474
rect 138346 7422 138348 7474
rect 138292 6860 138348 7422
rect 138964 8146 139020 8158
rect 138964 8094 138966 8146
rect 139018 8094 139020 8146
rect 138292 6804 138852 6860
rect 138796 6746 138852 6804
rect 138796 6694 138798 6746
rect 138850 6694 138852 6746
rect 138796 6682 138852 6694
rect 138068 5674 138124 5684
rect 138292 6412 138348 6422
rect 138124 4956 138180 4966
rect 138124 4954 138236 4956
rect 138124 4902 138126 4954
rect 138178 4902 138236 4954
rect 138124 4890 138236 4902
rect 137732 4118 137734 4170
rect 137786 4118 137788 4170
rect 137732 4106 137788 4118
rect 137956 4844 138012 4854
rect 137956 800 138012 4788
rect 138180 4058 138236 4890
rect 138292 4506 138348 6356
rect 138628 6412 138684 6422
rect 138628 5292 138684 6356
rect 138740 5906 138796 5918
rect 138740 5854 138742 5906
rect 138794 5854 138796 5906
rect 138740 5852 138796 5854
rect 138740 5786 138796 5796
rect 138628 5226 138684 5236
rect 138964 4732 139020 8094
rect 138964 4666 139020 4676
rect 139076 6524 139132 9604
rect 139188 8258 139244 12070
rect 139300 12124 139356 12134
rect 139300 9994 139356 12068
rect 139412 10668 139468 14200
rect 139524 13916 139580 13926
rect 139524 13578 139580 13860
rect 139524 13526 139526 13578
rect 139578 13526 139580 13578
rect 139524 13514 139580 13526
rect 140084 13804 140140 13814
rect 139748 12010 139804 12022
rect 139748 11958 139750 12010
rect 139802 11958 139804 12010
rect 139748 11900 139804 11958
rect 139524 11676 139580 11686
rect 139524 11226 139580 11620
rect 139524 11174 139526 11226
rect 139578 11174 139580 11226
rect 139524 11162 139580 11174
rect 139412 10602 139468 10612
rect 139300 9942 139302 9994
rect 139354 9942 139356 9994
rect 139300 9930 139356 9942
rect 139748 9826 139804 11844
rect 139748 9774 139750 9826
rect 139802 9774 139804 9826
rect 139748 9762 139804 9774
rect 139748 8988 139804 8998
rect 139524 8876 139580 8886
rect 139524 8426 139580 8820
rect 139524 8374 139526 8426
rect 139578 8374 139580 8426
rect 139524 8362 139580 8374
rect 139636 8652 139692 8662
rect 139188 8206 139190 8258
rect 139242 8206 139244 8258
rect 139188 8194 139244 8206
rect 139412 6860 139468 6870
rect 139636 6860 139692 8596
rect 139244 6524 139300 6534
rect 139076 6522 139300 6524
rect 139076 6470 139246 6522
rect 139298 6470 139300 6522
rect 139076 6468 139300 6470
rect 138292 4454 138294 4506
rect 138346 4454 138348 4506
rect 138292 4442 138348 4454
rect 138180 4006 138182 4058
rect 138234 4006 138236 4058
rect 138180 3994 138236 4006
rect 138516 3388 138572 3398
rect 138180 2604 138236 2614
rect 138180 1820 138236 2548
rect 138180 1754 138236 1764
rect 138516 800 138572 3332
rect 138628 3162 138684 3174
rect 138628 3110 138630 3162
rect 138682 3110 138684 3162
rect 138628 2490 138684 3110
rect 139076 2940 139132 6468
rect 139244 6458 139300 6468
rect 139412 6076 139468 6804
rect 139412 6010 139468 6020
rect 139524 6804 139692 6860
rect 139300 5964 139356 5974
rect 139300 5234 139356 5908
rect 139300 5182 139302 5234
rect 139354 5182 139356 5234
rect 139300 5170 139356 5182
rect 139412 5906 139468 5918
rect 139412 5854 139414 5906
rect 139466 5854 139468 5906
rect 139412 4844 139468 5854
rect 139412 4620 139468 4788
rect 139412 4554 139468 4564
rect 139412 4170 139468 4182
rect 139412 4118 139414 4170
rect 139466 4118 139468 4170
rect 139076 2874 139132 2884
rect 139188 3946 139244 3958
rect 139188 3894 139190 3946
rect 139242 3894 139244 3946
rect 138628 2438 138630 2490
rect 138682 2438 138684 2490
rect 138628 2426 138684 2438
rect 139188 800 139244 3894
rect 139412 2940 139468 4118
rect 139524 3724 139580 6804
rect 139748 6646 139804 8932
rect 139972 7586 140028 7598
rect 139972 7534 139974 7586
rect 140026 7534 140028 7586
rect 139860 7306 139916 7318
rect 139860 7254 139862 7306
rect 139914 7254 139916 7306
rect 139860 7196 139916 7254
rect 139860 7130 139916 7140
rect 139692 6634 139804 6646
rect 139692 6582 139694 6634
rect 139746 6582 139804 6634
rect 139692 6580 139804 6582
rect 139860 6860 139916 6870
rect 139692 6570 139748 6580
rect 139860 4508 139916 6804
rect 139860 4442 139916 4452
rect 139524 3658 139580 3668
rect 139636 4172 139692 4182
rect 139636 3500 139692 4116
rect 139636 3434 139692 3444
rect 139748 3724 139804 3734
rect 139412 2874 139468 2884
rect 139636 3164 139692 3174
rect 139636 2716 139692 3108
rect 139636 2650 139692 2660
rect 139748 800 139804 3668
rect 139972 3387 140028 7534
rect 140084 5794 140140 13748
rect 140196 13132 140252 14200
rect 140756 14140 140812 14150
rect 140196 13066 140252 13076
rect 140644 13466 140700 13478
rect 140644 13414 140646 13466
rect 140698 13414 140700 13466
rect 140308 9042 140364 9054
rect 140308 8990 140310 9042
rect 140362 8990 140364 9042
rect 140308 8988 140364 8990
rect 140308 8922 140364 8932
rect 140420 8930 140476 8942
rect 140420 8878 140422 8930
rect 140474 8878 140476 8930
rect 140084 5742 140086 5794
rect 140138 5742 140140 5794
rect 140084 5730 140140 5742
rect 140196 8764 140252 8774
rect 139860 3331 140028 3387
rect 140196 3386 140252 8708
rect 140308 7474 140364 7486
rect 140308 7422 140310 7474
rect 140362 7422 140364 7474
rect 140308 4394 140364 7422
rect 140420 7420 140476 8878
rect 140420 7354 140476 7364
rect 140644 6748 140700 13414
rect 140756 10108 140812 14084
rect 140868 11114 140924 14200
rect 141092 12010 141148 14310
rect 141624 14200 141736 15000
rect 142296 14200 142408 15000
rect 143080 14200 143192 15000
rect 143752 14200 143864 15000
rect 144536 14200 144648 15000
rect 145208 14200 145320 15000
rect 145992 14200 146104 15000
rect 146664 14200 146776 15000
rect 147448 14200 147560 15000
rect 147924 14362 147980 14374
rect 147924 14310 147926 14362
rect 147978 14310 147980 14362
rect 141652 13468 141708 14200
rect 141092 11958 141094 12010
rect 141146 11958 141148 12010
rect 141092 11946 141148 11958
rect 141204 13412 141708 13468
rect 141092 11786 141148 11798
rect 141092 11734 141094 11786
rect 141146 11734 141148 11786
rect 141092 11676 141148 11734
rect 141092 11610 141148 11620
rect 140868 11062 140870 11114
rect 140922 11062 140924 11114
rect 140868 11050 140924 11062
rect 141204 10332 141260 13412
rect 142324 13244 142380 14200
rect 142884 13914 142940 13926
rect 142884 13862 142886 13914
rect 142938 13862 142940 13914
rect 141204 10266 141260 10276
rect 141316 13188 142380 13244
rect 142660 13692 142716 13702
rect 140756 10042 140812 10052
rect 140756 9714 140812 9726
rect 140756 9662 140758 9714
rect 140810 9662 140812 9714
rect 140756 9212 140812 9662
rect 140980 9602 141036 9614
rect 140980 9550 140982 9602
rect 141034 9550 141036 9602
rect 140980 9436 141036 9550
rect 140980 9370 141036 9380
rect 140756 8988 140812 9156
rect 141316 9210 141372 13188
rect 142660 13130 142716 13636
rect 142660 13078 142662 13130
rect 142714 13078 142716 13130
rect 142660 13066 142716 13078
rect 142324 13018 142380 13030
rect 142324 12966 142326 13018
rect 142378 12966 142380 13018
rect 142324 10892 142380 12966
rect 142660 12908 142716 12918
rect 142660 12794 142716 12852
rect 142660 12742 142662 12794
rect 142714 12742 142716 12794
rect 142660 12730 142716 12742
rect 142884 12794 142940 13862
rect 142884 12742 142886 12794
rect 142938 12742 142940 12794
rect 142884 12730 142940 12742
rect 142996 13244 143052 13254
rect 141316 9158 141318 9210
rect 141370 9158 141372 9210
rect 141316 9146 141372 9158
rect 141540 10220 141596 10230
rect 141540 9212 141596 10164
rect 141708 9996 141764 10006
rect 141708 9882 141764 9940
rect 141708 9830 141710 9882
rect 141762 9830 141764 9882
rect 141708 9818 141764 9830
rect 141708 9212 141764 9222
rect 141540 9210 141764 9212
rect 141540 9158 141710 9210
rect 141762 9158 141764 9210
rect 141540 9156 141764 9158
rect 141708 9146 141764 9156
rect 140756 8922 140812 8932
rect 140980 9098 141036 9110
rect 140980 9046 140982 9098
rect 141034 9046 141036 9098
rect 140980 8764 141036 9046
rect 142324 9042 142380 10836
rect 142772 11788 142828 11798
rect 142324 8990 142326 9042
rect 142378 8990 142380 9042
rect 142324 8978 142380 8990
rect 142436 10220 142492 10230
rect 140980 8698 141036 8708
rect 141092 8540 141148 8550
rect 141092 8204 141148 8484
rect 141092 8138 141148 8148
rect 141876 8090 141932 8102
rect 141876 8038 141878 8090
rect 141930 8038 141932 8090
rect 141876 7980 141932 8038
rect 141876 7914 141932 7924
rect 140980 7474 141036 7486
rect 140980 7422 140982 7474
rect 141034 7422 141036 7474
rect 140980 6748 141036 7422
rect 142436 7474 142492 10164
rect 142772 7654 142828 11732
rect 142884 9772 142940 9782
rect 142884 9678 142940 9716
rect 142996 8540 143052 13188
rect 143108 12684 143164 14200
rect 143220 13914 143276 13926
rect 143220 13862 143222 13914
rect 143274 13862 143276 13914
rect 143220 13578 143276 13862
rect 143220 13526 143222 13578
rect 143274 13526 143276 13578
rect 143220 13514 143276 13526
rect 143108 12618 143164 12628
rect 143220 12236 143276 12246
rect 143220 9994 143276 12180
rect 143332 11900 143388 11910
rect 143332 11452 143388 11844
rect 143332 11386 143388 11396
rect 143220 9942 143222 9994
rect 143274 9942 143276 9994
rect 143220 9930 143276 9942
rect 143332 11226 143388 11238
rect 143332 11174 143334 11226
rect 143386 11174 143388 11226
rect 143332 10442 143388 11174
rect 143668 11116 143724 11126
rect 143332 10390 143334 10442
rect 143386 10390 143388 10442
rect 142996 8474 143052 8484
rect 143108 9772 143164 9782
rect 142772 7642 142884 7654
rect 142772 7590 142830 7642
rect 142882 7590 142884 7642
rect 142772 7588 142884 7590
rect 142828 7578 142884 7588
rect 142436 7422 142438 7474
rect 142490 7422 142492 7474
rect 142436 7410 142492 7422
rect 141876 7308 141932 7318
rect 141876 7214 141932 7252
rect 142660 6972 142716 6982
rect 142996 6972 143052 6982
rect 142716 6916 142828 6972
rect 142660 6906 142716 6916
rect 141764 6860 141820 6870
rect 141764 6766 141820 6804
rect 142772 6802 142828 6916
rect 140644 6682 140700 6692
rect 140868 6692 141036 6748
rect 142772 6750 142774 6802
rect 142826 6750 142828 6802
rect 142772 6738 142828 6750
rect 140868 6524 140924 6692
rect 142324 6690 142380 6702
rect 142324 6638 142326 6690
rect 142378 6638 142380 6690
rect 140308 4342 140310 4394
rect 140362 4342 140364 4394
rect 140308 4330 140364 4342
rect 140420 6468 140924 6524
rect 140980 6578 141036 6590
rect 140980 6526 140982 6578
rect 141034 6526 141036 6578
rect 140420 3946 140476 6468
rect 140868 5964 140924 5974
rect 140868 5906 140924 5908
rect 140868 5854 140870 5906
rect 140922 5854 140924 5906
rect 140868 5842 140924 5854
rect 140644 5122 140700 5134
rect 140644 5070 140646 5122
rect 140698 5070 140700 5122
rect 140644 5068 140700 5070
rect 140644 5002 140700 5012
rect 140420 3894 140422 3946
rect 140474 3894 140476 3946
rect 140420 3882 140476 3894
rect 140532 4956 140588 4966
rect 140196 3334 140198 3386
rect 140250 3334 140252 3386
rect 139860 3164 139916 3331
rect 140196 3322 140252 3334
rect 140308 3500 140364 3510
rect 139860 2268 139916 3108
rect 139860 2202 139916 2212
rect 140308 800 140364 3444
rect 140532 3164 140588 4900
rect 140980 4732 141036 6526
rect 142324 5964 142380 6638
rect 142996 6578 143052 6916
rect 142996 6526 142998 6578
rect 143050 6526 143052 6578
rect 141428 5906 141484 5918
rect 142324 5908 142492 5964
rect 141428 5854 141430 5906
rect 141482 5854 141484 5906
rect 141316 5794 141372 5806
rect 141316 5742 141318 5794
rect 141370 5742 141372 5794
rect 140644 4676 141036 4732
rect 141148 4954 141204 4966
rect 141148 4902 141150 4954
rect 141202 4902 141204 4954
rect 141148 4732 141204 4902
rect 140644 4170 140700 4676
rect 141148 4666 141204 4676
rect 140980 4508 141036 4518
rect 140868 4452 140980 4508
rect 140868 4396 140924 4452
rect 140980 4442 141036 4452
rect 140644 4118 140646 4170
rect 140698 4118 140700 4170
rect 140644 3388 140700 4118
rect 140756 4340 140924 4396
rect 140756 3500 140812 4340
rect 140980 4284 141036 4294
rect 140756 3434 140812 3444
rect 140868 4172 140924 4182
rect 140644 3322 140700 3332
rect 140532 3098 140588 3108
rect 140756 3164 140812 3174
rect 140756 2716 140812 3108
rect 140756 2650 140812 2660
rect 140868 1596 140924 4116
rect 140980 3498 141036 4228
rect 141204 4284 141260 4294
rect 141204 4170 141260 4228
rect 141204 4118 141206 4170
rect 141258 4118 141260 4170
rect 141204 4106 141260 4118
rect 140980 3446 140982 3498
rect 141034 3446 141036 3498
rect 140980 3434 141036 3446
rect 141092 3610 141148 3622
rect 141092 3558 141094 3610
rect 141146 3558 141148 3610
rect 140980 2380 141036 2390
rect 141092 2380 141148 3558
rect 141316 3500 141372 5742
rect 141428 5124 141484 5854
rect 142156 5516 142212 5526
rect 142156 5180 142212 5460
rect 141428 5068 141820 5124
rect 141428 3724 141484 5068
rect 141596 4956 141652 4966
rect 141596 4862 141652 4900
rect 141764 4956 141820 5068
rect 141764 4890 141820 4900
rect 142156 4954 142212 5124
rect 142156 4902 142158 4954
rect 142210 4902 142212 4954
rect 142156 4890 142212 4902
rect 141988 4506 142044 4518
rect 141988 4454 141990 4506
rect 142042 4454 142044 4506
rect 141540 3948 141596 3958
rect 141540 3854 141596 3892
rect 141428 3658 141484 3668
rect 141316 3434 141372 3444
rect 141764 3500 141820 3510
rect 141036 2324 141148 2380
rect 141540 3388 141596 3398
rect 141540 2380 141596 3332
rect 141764 3276 141820 3444
rect 141764 3210 141820 3220
rect 140980 2314 141036 2324
rect 141540 2314 141596 2324
rect 141540 2156 141596 2166
rect 140868 1540 141036 1596
rect 140980 800 141036 1540
rect 141540 800 141596 2100
rect 134484 522 134540 532
rect 134792 0 134904 800
rect 135464 0 135576 800
rect 136024 0 136136 800
rect 136696 0 136808 800
rect 137256 0 137368 800
rect 137928 0 138040 800
rect 138488 0 138600 800
rect 139160 0 139272 800
rect 139720 0 139832 800
rect 140280 0 140392 800
rect 140952 0 141064 800
rect 141512 0 141624 800
rect 141988 476 142044 4454
rect 142436 4506 142492 5908
rect 142660 5906 142716 5918
rect 142660 5854 142662 5906
rect 142714 5854 142716 5906
rect 142660 4732 142716 5854
rect 142828 4954 142884 4966
rect 142828 4902 142830 4954
rect 142882 4902 142884 4954
rect 142828 4844 142884 4902
rect 142828 4778 142884 4788
rect 142660 4666 142716 4676
rect 142436 4454 142438 4506
rect 142490 4454 142492 4506
rect 142436 4442 142492 4454
rect 142996 4508 143052 6526
rect 142996 4442 143052 4452
rect 142772 4396 142828 4406
rect 142548 3612 142604 3622
rect 142212 1484 142268 1494
rect 142212 800 142268 1428
rect 142548 812 142604 3556
rect 142772 3500 142828 4340
rect 142772 3434 142828 3444
rect 143108 3386 143164 9716
rect 143332 8428 143388 10390
rect 143556 10778 143612 10790
rect 143556 10726 143558 10778
rect 143610 10726 143612 10778
rect 143556 10442 143612 10726
rect 143556 10390 143558 10442
rect 143610 10390 143612 10442
rect 143556 10378 143612 10390
rect 143668 9660 143724 11060
rect 143780 9884 143836 14200
rect 144116 13916 144172 13926
rect 144116 9994 144172 13860
rect 144452 13242 144508 13254
rect 144452 13190 144454 13242
rect 144506 13190 144508 13242
rect 144228 12908 144284 12918
rect 144228 12122 144284 12852
rect 144452 12234 144508 13190
rect 144452 12182 144454 12234
rect 144506 12182 144508 12234
rect 144452 12170 144508 12182
rect 144228 12070 144230 12122
rect 144282 12070 144284 12122
rect 144228 12058 144284 12070
rect 144116 9942 144118 9994
rect 144170 9942 144172 9994
rect 144116 9930 144172 9942
rect 144452 11900 144508 11910
rect 144452 9894 144508 11844
rect 144564 11788 144620 14200
rect 144564 11722 144620 11732
rect 145124 12458 145180 12470
rect 145124 12406 145126 12458
rect 145178 12406 145180 12458
rect 143780 9828 144060 9884
rect 144452 9882 144564 9894
rect 144452 9830 144510 9882
rect 144562 9830 144564 9882
rect 144452 9828 144564 9830
rect 143780 9660 143836 9670
rect 143668 9658 143836 9660
rect 143668 9606 143782 9658
rect 143834 9606 143836 9658
rect 143668 9604 143836 9606
rect 143780 9594 143836 9604
rect 143780 9212 143836 9222
rect 143780 9042 143836 9156
rect 143780 8990 143782 9042
rect 143834 8990 143836 9042
rect 143780 8978 143836 8990
rect 143892 8988 143948 8998
rect 143892 8930 143948 8932
rect 143892 8878 143894 8930
rect 143946 8878 143948 8930
rect 143892 8866 143948 8878
rect 143220 8372 143388 8428
rect 143668 8428 143724 8438
rect 143220 6076 143276 8372
rect 143332 8258 143388 8270
rect 143332 8206 143334 8258
rect 143386 8206 143388 8258
rect 143332 6188 143388 8206
rect 143668 8204 143724 8372
rect 143612 8148 143724 8204
rect 143612 7474 143668 8148
rect 143724 7644 143780 7654
rect 143724 7550 143780 7588
rect 143612 7422 143614 7474
rect 143666 7422 143668 7474
rect 143612 6870 143668 7422
rect 143556 6860 143668 6870
rect 143612 6804 143668 6860
rect 143556 6794 143612 6804
rect 143332 6132 143780 6188
rect 143220 6020 143444 6076
rect 143388 5962 143444 6020
rect 143388 5910 143390 5962
rect 143442 5910 143444 5962
rect 143388 5898 143444 5910
rect 143556 5628 143612 6132
rect 143724 6074 143780 6132
rect 143724 6022 143726 6074
rect 143778 6022 143780 6074
rect 143724 6010 143780 6022
rect 143444 5572 143612 5628
rect 143276 4954 143332 4966
rect 143276 4902 143278 4954
rect 143330 4902 143332 4954
rect 143276 4396 143332 4902
rect 143276 4394 143388 4396
rect 143276 4342 143278 4394
rect 143330 4342 143388 4394
rect 143276 4330 143388 4342
rect 143332 4170 143388 4330
rect 143332 4118 143334 4170
rect 143386 4118 143388 4170
rect 143332 4106 143388 4118
rect 143108 3334 143110 3386
rect 143162 3334 143164 3386
rect 143108 3322 143164 3334
rect 141988 410 142044 420
rect 142184 0 142296 800
rect 142772 2828 142828 2838
rect 142772 800 142828 2772
rect 143444 1932 143500 5572
rect 143780 5404 143836 5414
rect 143612 4954 143668 4966
rect 143612 4902 143614 4954
rect 143666 4902 143668 4954
rect 143612 4620 143668 4902
rect 143612 4554 143668 4564
rect 143780 4620 143836 5348
rect 143780 4554 143836 4564
rect 143556 4394 143612 4406
rect 143556 4342 143558 4394
rect 143610 4342 143612 4394
rect 143556 3722 143612 4342
rect 144004 4058 144060 9828
rect 144508 9818 144564 9828
rect 144956 9772 145012 9782
rect 144956 9678 145012 9716
rect 144676 9212 144732 9222
rect 144452 8876 144508 8886
rect 144452 8316 144508 8820
rect 144228 8247 144284 8259
rect 144452 8250 144508 8260
rect 144676 8876 144732 9156
rect 144228 8195 144230 8247
rect 144282 8195 144284 8247
rect 144228 7644 144284 8195
rect 144228 7578 144284 7588
rect 144564 8092 144620 8102
rect 144564 7084 144620 8036
rect 144676 7430 144732 8820
rect 145012 9212 145068 9222
rect 144788 8204 144844 8214
rect 144788 7644 144844 8148
rect 144788 7578 144844 7588
rect 144676 7418 144788 7430
rect 144676 7366 144734 7418
rect 144786 7366 144788 7418
rect 144676 7364 144788 7366
rect 144732 7354 144788 7364
rect 144676 7084 144732 7094
rect 144564 7028 144676 7084
rect 144676 7018 144732 7028
rect 144564 6860 144620 6870
rect 144340 6690 144396 6702
rect 144340 6638 144342 6690
rect 144394 6638 144396 6690
rect 144228 5852 144284 5862
rect 144228 4620 144284 5796
rect 144340 4844 144396 6638
rect 144452 5852 144508 5862
rect 144452 5292 144508 5796
rect 144452 5226 144508 5236
rect 144564 5234 144620 6804
rect 145012 6524 145068 9156
rect 145124 9044 145180 12406
rect 145236 12012 145292 14200
rect 145236 11946 145292 11956
rect 145348 12908 145404 12918
rect 145348 12458 145404 12852
rect 145348 12406 145350 12458
rect 145402 12406 145404 12458
rect 145124 9042 145292 9044
rect 145124 8990 145126 9042
rect 145178 8990 145292 9042
rect 145124 8988 145292 8990
rect 145124 8978 145180 8988
rect 145236 8316 145292 8988
rect 145124 8258 145180 8270
rect 145124 8206 145126 8258
rect 145178 8206 145180 8258
rect 145236 8250 145292 8260
rect 145124 8204 145180 8206
rect 145124 8138 145180 8148
rect 145348 7654 145404 12406
rect 146020 11226 146076 14200
rect 146692 13020 146748 14200
rect 146692 12954 146748 12964
rect 147140 13244 147196 13254
rect 147028 12908 147084 12918
rect 146020 11174 146022 11226
rect 146074 11174 146076 11226
rect 146020 11162 146076 11174
rect 146132 11340 146188 11350
rect 145516 9660 145572 9670
rect 145964 9660 146020 9670
rect 145516 9658 146076 9660
rect 145516 9606 145518 9658
rect 145570 9606 145966 9658
rect 146018 9606 146076 9658
rect 145516 9604 146076 9606
rect 145516 9594 145572 9604
rect 145964 9594 146076 9604
rect 145292 7642 145404 7654
rect 145292 7590 145294 7642
rect 145346 7590 145404 7642
rect 145292 7588 145404 7590
rect 145572 8874 145628 8886
rect 145572 8822 145574 8874
rect 145626 8822 145628 8874
rect 145292 7578 145348 7588
rect 145572 7420 145628 8822
rect 146020 8876 146076 9594
rect 146020 8810 146076 8820
rect 145684 8428 145740 8438
rect 145684 8334 145740 8372
rect 145572 7354 145628 7364
rect 145796 6860 145852 6870
rect 145796 6766 145852 6804
rect 145012 6458 145068 6468
rect 145236 6636 145292 6646
rect 145236 6130 145292 6580
rect 144788 6076 144844 6086
rect 145124 6076 145180 6086
rect 145012 6020 145124 6076
rect 145236 6078 145238 6130
rect 145290 6078 145292 6130
rect 145236 6066 145292 6078
rect 145348 6578 145404 6590
rect 145348 6526 145350 6578
rect 145402 6526 145404 6578
rect 144676 5964 144732 5974
rect 144788 5964 145068 6020
rect 145124 6010 145180 6020
rect 145236 5964 145292 5974
rect 144676 5628 144732 5908
rect 145012 5628 145068 5638
rect 144676 5572 145012 5628
rect 145012 5562 145068 5572
rect 144564 5182 144566 5234
rect 144618 5182 144620 5234
rect 144564 5170 144620 5182
rect 145236 5068 145292 5908
rect 144676 5012 145292 5068
rect 144452 4844 144508 4854
rect 144340 4788 144452 4844
rect 144452 4778 144508 4788
rect 144676 4620 144732 5012
rect 144228 4564 144732 4620
rect 144900 4844 144956 4854
rect 144004 4006 144006 4058
rect 144058 4006 144060 4058
rect 144004 3994 144060 4006
rect 143556 3670 143558 3722
rect 143610 3670 143612 3722
rect 143556 3658 143612 3670
rect 144004 3724 144060 3734
rect 144004 3630 144060 3668
rect 144900 2156 144956 4788
rect 145348 4284 145404 6526
rect 146020 6018 146076 6030
rect 146020 5966 146022 6018
rect 146074 5966 146076 6018
rect 145684 5906 145740 5918
rect 145684 5854 145686 5906
rect 145738 5854 145740 5906
rect 145572 4620 145628 4630
rect 145348 3946 145404 4228
rect 145460 4506 145516 4518
rect 145460 4454 145462 4506
rect 145514 4454 145516 4506
rect 145460 4058 145516 4454
rect 145572 4284 145628 4564
rect 145684 4506 145740 5854
rect 145908 5292 145964 5302
rect 145908 5122 145964 5236
rect 145908 5070 145910 5122
rect 145962 5070 145964 5122
rect 145908 5058 145964 5070
rect 146020 4844 146076 5966
rect 146020 4778 146076 4788
rect 145684 4454 145686 4506
rect 145738 4454 145740 4506
rect 145684 4442 145740 4454
rect 145572 4218 145628 4228
rect 145460 4006 145462 4058
rect 145514 4006 145516 4058
rect 145460 3994 145516 4006
rect 145348 3894 145350 3946
rect 145402 3894 145404 3946
rect 145348 3882 145404 3894
rect 146132 3722 146188 11284
rect 146916 10892 146972 10902
rect 146804 10780 146860 10790
rect 146580 10444 146636 10454
rect 146580 10220 146636 10388
rect 146580 10154 146636 10164
rect 146804 10220 146860 10724
rect 146804 9770 146860 10164
rect 146804 9718 146806 9770
rect 146858 9718 146860 9770
rect 146804 9706 146860 9718
rect 146916 9222 146972 10836
rect 147028 9436 147084 12852
rect 147140 9994 147196 13188
rect 147476 11562 147532 14200
rect 147924 13692 147980 14310
rect 148120 14200 148232 15000
rect 148596 14922 148652 14934
rect 148596 14870 148598 14922
rect 148650 14870 148652 14922
rect 148372 14698 148428 14710
rect 148372 14646 148374 14698
rect 148426 14646 148428 14698
rect 147924 13626 147980 13636
rect 148148 12124 148204 14200
rect 148372 13804 148428 14646
rect 148372 13738 148428 13748
rect 148372 13468 148428 13478
rect 148372 13374 148428 13412
rect 148596 13018 148652 14870
rect 148708 14250 148764 14262
rect 148708 14198 148710 14250
rect 148762 14198 148764 14250
rect 148904 14200 149016 15000
rect 149156 14476 149212 14486
rect 148708 14028 148764 14198
rect 148708 13962 148764 13972
rect 148932 13132 148988 14200
rect 149156 13802 149212 14420
rect 149268 14252 149324 14262
rect 149576 14200 149688 15000
rect 149828 14474 149884 14486
rect 149828 14422 149830 14474
rect 149882 14422 149884 14474
rect 149828 14252 149884 14422
rect 149268 14158 149324 14196
rect 149156 13750 149158 13802
rect 149210 13750 149212 13802
rect 149156 13738 149212 13750
rect 149380 14138 149436 14150
rect 149380 14086 149382 14138
rect 149434 14086 149436 14138
rect 149380 13690 149436 14086
rect 149380 13638 149382 13690
rect 149434 13638 149436 13690
rect 149380 13626 149436 13638
rect 149268 13580 149324 13590
rect 148932 13066 148988 13076
rect 149156 13354 149212 13366
rect 149156 13302 149158 13354
rect 149210 13302 149212 13354
rect 148596 12966 148598 13018
rect 148650 12966 148652 13018
rect 148596 12954 148652 12966
rect 149156 13020 149212 13302
rect 149268 13130 149324 13524
rect 149492 13580 149548 13590
rect 149380 13356 149436 13366
rect 149380 13262 149436 13300
rect 149492 13242 149548 13524
rect 149492 13190 149494 13242
rect 149546 13190 149548 13242
rect 149492 13178 149548 13190
rect 149268 13078 149270 13130
rect 149322 13078 149324 13130
rect 149268 13066 149324 13078
rect 149156 12954 149212 12964
rect 149044 12906 149100 12918
rect 149044 12854 149046 12906
rect 149098 12854 149100 12906
rect 148708 12572 148764 12610
rect 148708 12506 148764 12516
rect 149044 12572 149100 12854
rect 149044 12506 149100 12516
rect 149268 12906 149324 12918
rect 149268 12854 149270 12906
rect 149322 12854 149324 12906
rect 149268 12570 149324 12854
rect 149268 12518 149270 12570
rect 149322 12518 149324 12570
rect 149268 12506 149324 12518
rect 148708 12348 148764 12358
rect 148596 12234 148652 12246
rect 148596 12182 148598 12234
rect 148650 12182 148652 12234
rect 148148 12068 148316 12124
rect 147812 11900 147868 11910
rect 147476 11510 147478 11562
rect 147530 11510 147532 11562
rect 147476 11498 147532 11510
rect 147700 11788 147756 11798
rect 147700 11004 147756 11732
rect 147700 10938 147756 10948
rect 147812 10556 147868 11844
rect 148148 11898 148204 11910
rect 148148 11846 148150 11898
rect 148202 11846 148204 11898
rect 147812 10490 147868 10500
rect 147924 11116 147980 11126
rect 147140 9942 147142 9994
rect 147194 9942 147196 9994
rect 147140 9930 147196 9942
rect 147252 10444 147308 10454
rect 147028 9380 147196 9436
rect 146916 9210 147028 9222
rect 146916 9158 146974 9210
rect 147026 9158 147028 9210
rect 146916 9156 147028 9158
rect 146972 9146 147028 9156
rect 146468 9042 146524 9054
rect 146468 8990 146470 9042
rect 146522 8990 146524 9042
rect 146468 8876 146524 8990
rect 147140 8988 147196 9380
rect 146916 8932 147196 8988
rect 146580 8876 146636 8886
rect 146468 8820 146580 8876
rect 146580 8258 146636 8820
rect 146356 8204 146412 8214
rect 146580 8206 146582 8258
rect 146634 8206 146636 8258
rect 146580 8194 146636 8206
rect 146244 7532 146300 7542
rect 146244 6300 146300 7476
rect 146356 6690 146412 8148
rect 146356 6638 146358 6690
rect 146410 6638 146412 6690
rect 146356 6626 146412 6638
rect 146748 6524 146804 6534
rect 146244 6234 146300 6244
rect 146580 6522 146804 6524
rect 146580 6470 146750 6522
rect 146802 6470 146804 6522
rect 146580 6468 146804 6470
rect 146132 3670 146134 3722
rect 146186 3670 146188 3722
rect 146132 3658 146188 3670
rect 146468 4172 146524 4182
rect 144900 2090 144956 2100
rect 143444 1866 143500 1876
rect 145796 1820 145852 1830
rect 143444 1596 143500 1606
rect 143444 800 143500 1540
rect 144004 1596 144060 1606
rect 144004 800 144060 1540
rect 144788 1594 144844 1606
rect 144788 1542 144790 1594
rect 144842 1542 144844 1594
rect 144788 1036 144844 1542
rect 144732 980 144844 1036
rect 145236 1596 145292 1606
rect 144732 924 144788 980
rect 144676 868 144788 924
rect 144676 800 144732 868
rect 145236 800 145292 1540
rect 145796 800 145852 1764
rect 146468 800 146524 4116
rect 146580 3948 146636 6468
rect 146748 6458 146804 6468
rect 146916 6188 146972 8932
rect 147252 8876 147308 10388
rect 147532 10108 147588 10118
rect 147532 9882 147588 10052
rect 147532 9830 147534 9882
rect 147586 9830 147588 9882
rect 147532 9818 147588 9830
rect 147924 9894 147980 11060
rect 147924 9882 148036 9894
rect 147924 9830 147982 9882
rect 148034 9830 148036 9882
rect 147924 9828 148036 9830
rect 147980 9818 148036 9828
rect 148148 9884 148204 11846
rect 148148 9042 148204 9828
rect 147084 8820 147308 8876
rect 147420 8986 147476 8998
rect 147420 8934 147422 8986
rect 147474 8934 147476 8986
rect 148148 8990 148150 9042
rect 148202 8990 148204 9042
rect 148148 8978 148204 8990
rect 147420 8876 147476 8934
rect 147084 8314 147140 8820
rect 147420 8810 147476 8820
rect 147084 8262 147086 8314
rect 147138 8262 147140 8314
rect 147084 8250 147140 8262
rect 147532 8316 147588 8326
rect 147532 8222 147588 8260
rect 147980 8092 148036 8102
rect 147812 8090 148036 8092
rect 147812 8038 147982 8090
rect 148034 8038 148036 8090
rect 147812 8036 148036 8038
rect 147588 7532 147644 7542
rect 147588 7306 147644 7476
rect 147588 7254 147590 7306
rect 147642 7254 147644 7306
rect 147588 7242 147644 7254
rect 147812 6972 147868 8036
rect 147980 8026 148036 8036
rect 147812 6906 147868 6916
rect 147924 7532 147980 7552
rect 147924 7474 147980 7476
rect 147924 7422 147926 7474
rect 147978 7422 147980 7474
rect 147644 6860 147700 6870
rect 147196 6524 147252 6534
rect 147644 6524 147700 6804
rect 147196 6522 147308 6524
rect 147196 6470 147198 6522
rect 147250 6470 147308 6522
rect 147196 6458 147308 6470
rect 146916 6076 146972 6132
rect 146804 6020 146972 6076
rect 146804 5190 146860 6020
rect 146748 5178 146860 5190
rect 146748 5126 146750 5178
rect 146802 5126 146860 5178
rect 146748 5124 146860 5126
rect 146916 5906 146972 5918
rect 146916 5854 146918 5906
rect 146970 5854 146972 5906
rect 146748 5114 146804 5124
rect 146580 3882 146636 3892
rect 146916 4732 146972 5854
rect 147084 4956 147140 4966
rect 147084 4862 147140 4900
rect 146916 3836 146972 4676
rect 147252 4396 147308 6458
rect 147644 6430 147700 6468
rect 147252 4330 147308 4340
rect 147476 5906 147532 5918
rect 147476 5854 147478 5906
rect 147530 5854 147532 5906
rect 147476 4396 147532 5854
rect 147812 5738 147868 5750
rect 147812 5686 147814 5738
rect 147866 5686 147868 5738
rect 147644 4956 147700 4966
rect 147644 4862 147700 4900
rect 147700 4508 147756 4518
rect 147812 4508 147868 5686
rect 147756 4452 147868 4508
rect 147700 4442 147756 4452
rect 147476 4330 147532 4340
rect 146916 3770 146972 3780
rect 147476 4060 147532 4070
rect 147364 1708 147420 1718
rect 147252 1652 147364 1708
rect 147252 1484 147308 1652
rect 147364 1642 147420 1652
rect 147476 1594 147532 4004
rect 147924 3834 147980 7422
rect 148092 4956 148148 4966
rect 148092 4954 148204 4956
rect 148092 4902 148094 4954
rect 148146 4902 148204 4954
rect 148092 4890 148204 4902
rect 148148 4058 148204 4890
rect 148260 4170 148316 12068
rect 148428 10220 148484 10230
rect 148428 9882 148484 10164
rect 148428 9830 148430 9882
rect 148482 9830 148484 9882
rect 148428 9818 148484 9830
rect 148596 9548 148652 12182
rect 148708 11116 148764 12292
rect 149492 12348 149548 12358
rect 148932 11900 148988 11910
rect 148932 11806 148988 11844
rect 148708 11050 148764 11060
rect 149380 9996 149436 10006
rect 149492 9996 149548 12292
rect 149436 9940 149548 9996
rect 149380 9930 149436 9940
rect 148876 9660 148932 9670
rect 148876 9566 148932 9604
rect 149436 9660 149492 9670
rect 149436 9658 149548 9660
rect 149436 9606 149438 9658
rect 149490 9606 149548 9658
rect 149436 9594 149548 9606
rect 148596 9492 148764 9548
rect 148596 8874 148652 8886
rect 148596 8822 148598 8874
rect 148650 8822 148652 8874
rect 148596 6300 148652 8822
rect 148708 8540 148764 9492
rect 149492 9042 149548 9594
rect 149492 8990 149494 9042
rect 149546 8990 149548 9042
rect 149604 9100 149660 14200
rect 150360 14200 150472 15000
rect 150724 14364 150780 14374
rect 150780 14308 150892 14364
rect 150724 14298 150780 14308
rect 149828 14186 149884 14196
rect 150164 13468 150220 13478
rect 149716 13132 149772 13142
rect 149716 10444 149772 13076
rect 150052 11450 150108 11462
rect 150052 11398 150054 11450
rect 150106 11398 150108 11450
rect 150052 11340 150108 11398
rect 150052 11274 150108 11284
rect 149716 10378 149772 10388
rect 149772 9884 149828 9894
rect 149772 9790 149828 9828
rect 149604 9034 149660 9044
rect 149492 8988 149548 8990
rect 148820 8932 149548 8988
rect 148820 8876 148876 8932
rect 148820 8810 148876 8820
rect 148708 8258 148764 8484
rect 149268 8764 149324 8774
rect 149268 8426 149324 8708
rect 149268 8374 149270 8426
rect 149322 8374 149324 8426
rect 149268 8362 149324 8374
rect 149492 8428 149548 8932
rect 149604 8428 149660 8438
rect 149492 8372 149604 8428
rect 149604 8362 149660 8372
rect 150052 8428 150108 8438
rect 148708 8206 148710 8258
rect 148762 8206 148764 8258
rect 148708 8194 148764 8206
rect 150052 8146 150108 8372
rect 150052 8094 150054 8146
rect 150106 8094 150108 8146
rect 150052 8082 150108 8094
rect 150164 8204 150220 13412
rect 150388 12458 150444 14200
rect 150836 14140 150892 14308
rect 151032 14200 151144 15000
rect 151396 14924 151452 14934
rect 151284 14588 151340 14598
rect 151060 14140 151116 14200
rect 150836 14084 151116 14140
rect 150388 12406 150390 12458
rect 150442 12406 150444 12458
rect 150388 12394 150444 12406
rect 150500 14028 150556 14038
rect 151284 14028 151340 14532
rect 150388 11340 150444 11350
rect 150388 11114 150444 11284
rect 150388 11062 150390 11114
rect 150442 11062 150444 11114
rect 150388 11050 150444 11062
rect 150276 11004 150332 11014
rect 150276 10910 150332 10948
rect 148708 7868 148764 7878
rect 148708 6802 148764 7812
rect 149996 7532 150052 7542
rect 149604 7470 149660 7482
rect 149604 7418 149606 7470
rect 149658 7418 149660 7470
rect 149996 7438 150052 7476
rect 150164 7532 150220 8148
rect 150164 7466 150220 7476
rect 150276 9884 150332 9894
rect 148708 6750 148710 6802
rect 148762 6750 148764 6802
rect 148708 6738 148764 6750
rect 148820 6972 148876 6982
rect 148596 6234 148652 6244
rect 148820 6086 148876 6916
rect 149604 6636 149660 7418
rect 150276 6860 150332 9828
rect 150388 9772 150444 9782
rect 150388 9100 150444 9716
rect 150388 9034 150444 9044
rect 150500 9044 150556 13972
rect 150948 13972 151340 14028
rect 150724 10108 150780 10118
rect 150724 9770 150780 10052
rect 150948 9884 151004 13972
rect 151060 13242 151116 13254
rect 151060 13190 151062 13242
rect 151114 13190 151116 13242
rect 151060 12684 151116 13190
rect 151060 12618 151116 12628
rect 151172 12796 151228 12806
rect 151060 11676 151116 11686
rect 151060 11002 151116 11620
rect 151172 11338 151228 12740
rect 151172 11286 151174 11338
rect 151226 11286 151228 11338
rect 151172 11274 151228 11286
rect 151284 11674 151340 11686
rect 151284 11622 151286 11674
rect 151338 11622 151340 11674
rect 151060 10950 151062 11002
rect 151114 10950 151116 11002
rect 151060 10938 151116 10950
rect 151172 11116 151228 11126
rect 151060 9996 151116 10006
rect 151060 9902 151116 9940
rect 150948 9818 151004 9828
rect 151172 9884 151228 11060
rect 151172 9818 151228 9828
rect 150724 9718 150726 9770
rect 150778 9718 150780 9770
rect 150724 9706 150780 9718
rect 150500 9042 150892 9044
rect 150500 8990 150502 9042
rect 150554 8990 150892 9042
rect 150500 8988 150892 8990
rect 150500 8978 150556 8988
rect 150500 8428 150556 8438
rect 150500 8204 150556 8372
rect 150668 8204 150724 8214
rect 150444 8148 150668 8204
rect 150444 7642 150500 8148
rect 150668 8110 150724 8148
rect 150444 7590 150446 7642
rect 150498 7590 150500 7642
rect 150444 7578 150500 7590
rect 150836 7644 150892 8988
rect 150948 8874 151004 8886
rect 150948 8822 150950 8874
rect 151002 8822 151004 8874
rect 150948 8428 151004 8822
rect 150948 8362 151004 8372
rect 151116 8540 151172 8550
rect 151116 8314 151172 8484
rect 151116 8262 151118 8314
rect 151170 8262 151172 8314
rect 151116 8250 151172 8262
rect 151284 8092 151340 11622
rect 151396 10890 151452 14868
rect 151508 14810 151564 14822
rect 151508 14758 151510 14810
rect 151562 14758 151564 14810
rect 151508 14476 151564 14758
rect 151508 14410 151564 14420
rect 151816 14200 151928 15000
rect 152488 14200 152600 15000
rect 152852 14252 152908 14262
rect 151844 13692 151900 14200
rect 151844 13626 151900 13636
rect 152068 13692 152124 13702
rect 152068 13468 152124 13636
rect 152068 13402 152124 13412
rect 152516 12908 152572 14200
rect 152516 12842 152572 12852
rect 153272 14200 153384 15000
rect 153944 14200 154056 15000
rect 154728 14200 154840 15000
rect 155204 14476 155260 14486
rect 152852 12570 152908 14196
rect 152852 12518 152854 12570
rect 152906 12518 152908 12570
rect 152852 12506 152908 12518
rect 152964 13804 153020 13814
rect 151508 11900 151564 11910
rect 151508 11806 151564 11844
rect 151396 10838 151398 10890
rect 151450 10838 151452 10890
rect 151396 10826 151452 10838
rect 151732 11564 151788 11574
rect 151732 10780 151788 11508
rect 151732 10714 151788 10724
rect 152068 10892 152124 10902
rect 151452 10108 151508 10118
rect 151452 9882 151508 10052
rect 151452 9830 151454 9882
rect 151506 9830 151508 9882
rect 151452 9818 151508 9830
rect 151844 9042 151900 9054
rect 151844 8990 151846 9042
rect 151898 8990 151900 9042
rect 151172 8036 151340 8092
rect 151396 8540 151452 8550
rect 151396 8204 151452 8484
rect 151844 8540 151900 8990
rect 151844 8474 151900 8484
rect 151900 8258 151956 8270
rect 151900 8249 151902 8258
rect 151004 7644 151060 7654
rect 150836 7642 151060 7644
rect 150836 7590 151006 7642
rect 151058 7590 151060 7642
rect 150836 7588 151060 7590
rect 151004 7578 151060 7588
rect 148764 6076 148876 6086
rect 148708 6074 148876 6076
rect 148708 6022 148766 6074
rect 148818 6022 148876 6074
rect 148708 6020 148876 6022
rect 149268 6578 149324 6590
rect 149268 6526 149270 6578
rect 149322 6526 149324 6578
rect 149604 6570 149660 6580
rect 150164 6804 150332 6860
rect 150724 7532 150780 7542
rect 149268 6524 149324 6526
rect 150164 6524 150220 6804
rect 150500 6748 150556 6758
rect 150276 6692 150500 6748
rect 150276 6690 150332 6692
rect 150276 6638 150278 6690
rect 150330 6638 150332 6690
rect 150500 6682 150556 6692
rect 150276 6626 150332 6638
rect 150724 6646 150780 7476
rect 151172 7196 151228 8036
rect 151396 7654 151452 8148
rect 151340 7642 151452 7654
rect 151340 7590 151342 7642
rect 151394 7590 151452 7642
rect 151340 7588 151452 7590
rect 151508 8206 151902 8249
rect 151954 8206 151956 8258
rect 151508 8204 151956 8206
rect 151508 8193 151900 8204
rect 151340 7578 151396 7588
rect 151508 7420 151564 8193
rect 151900 8117 151956 8148
rect 151788 8092 151844 8102
rect 151396 7364 151564 7420
rect 151620 8090 151844 8092
rect 151620 8038 151790 8090
rect 151842 8038 151844 8090
rect 151620 8036 151844 8038
rect 151172 7140 151340 7196
rect 150724 6634 150836 6646
rect 150724 6582 150782 6634
rect 150834 6582 150836 6634
rect 150724 6580 150836 6582
rect 150780 6570 150836 6580
rect 151116 6524 151172 6534
rect 150164 6468 150444 6524
rect 149268 6076 149324 6468
rect 149268 6020 149436 6076
rect 148708 6010 148820 6020
rect 148540 5068 148596 5078
rect 148540 4974 148596 5012
rect 148260 4118 148262 4170
rect 148314 4118 148316 4170
rect 148260 4106 148316 4118
rect 148148 4006 148150 4058
rect 148202 4006 148204 4058
rect 148148 3994 148204 4006
rect 147924 3782 147926 3834
rect 147978 3782 147980 3834
rect 147924 3770 147980 3782
rect 148708 3724 148764 6010
rect 149212 5852 149268 5862
rect 149156 5850 149268 5852
rect 149156 5798 149214 5850
rect 149266 5798 149268 5850
rect 149156 5786 149268 5798
rect 148876 4954 148932 4966
rect 148876 4902 148878 4954
rect 148930 4902 148932 4954
rect 148876 4844 148932 4902
rect 148876 4778 148932 4788
rect 149156 3946 149212 5786
rect 149380 5516 149436 6020
rect 149940 6018 149996 6030
rect 149940 5966 149942 6018
rect 149994 5966 149996 6018
rect 149156 3894 149158 3946
rect 149210 3894 149212 3946
rect 149156 3882 149212 3894
rect 149268 5460 149436 5516
rect 149716 5794 149772 5806
rect 149716 5742 149718 5794
rect 149770 5742 149772 5794
rect 148708 3658 148764 3668
rect 147812 3498 147868 3510
rect 147812 3446 147814 3498
rect 147866 3446 147868 3498
rect 147812 3276 147868 3446
rect 147812 3210 147868 3220
rect 149268 2828 149324 5460
rect 149716 5404 149772 5742
rect 149716 5338 149772 5348
rect 149436 5068 149492 5078
rect 149436 4956 149492 5012
rect 149436 4954 149548 4956
rect 149436 4902 149438 4954
rect 149490 4902 149548 4954
rect 149436 4890 149548 4902
rect 149492 4506 149548 4890
rect 149772 4954 149828 4966
rect 149772 4902 149774 4954
rect 149826 4902 149828 4954
rect 149772 4732 149828 4902
rect 149940 4844 149996 5966
rect 149940 4778 149996 4788
rect 149772 4666 149828 4676
rect 150052 4732 150108 4742
rect 149492 4454 149494 4506
rect 149546 4454 149548 4506
rect 149492 4442 149548 4454
rect 150052 4058 150108 4676
rect 150052 4006 150054 4058
rect 150106 4006 150108 4058
rect 150052 3994 150108 4006
rect 150164 3388 150220 3398
rect 149268 2762 149324 2772
rect 149492 3276 149548 3286
rect 148932 2156 148988 2166
rect 147476 1542 147478 1594
rect 147530 1542 147532 1594
rect 147476 1530 147532 1542
rect 148260 1932 148316 1942
rect 147028 1428 147308 1484
rect 147028 800 147084 1428
rect 147700 1036 147756 1046
rect 147700 800 147756 980
rect 148260 800 148316 1876
rect 148932 800 148988 2100
rect 149492 800 149548 3220
rect 150052 2940 150108 2950
rect 150052 2268 150108 2884
rect 150164 2716 150220 3332
rect 150388 3274 150444 6468
rect 151116 6430 151172 6468
rect 150948 5906 151004 5918
rect 150948 5854 150950 5906
rect 151002 5854 151004 5906
rect 150948 5852 151004 5854
rect 150948 5786 151004 5796
rect 151284 5234 151340 7140
rect 151284 5182 151286 5234
rect 151338 5182 151340 5234
rect 151284 5170 151340 5182
rect 151284 4620 151340 4630
rect 151396 4620 151452 7364
rect 151620 6860 151676 8036
rect 151788 8026 151844 8036
rect 152068 7980 152124 10836
rect 152404 10444 152460 10454
rect 152236 9660 152292 9670
rect 152236 9658 152348 9660
rect 152236 9606 152238 9658
rect 152290 9606 152348 9658
rect 152236 9594 152348 9606
rect 152292 8540 152348 9594
rect 152292 8474 152348 8484
rect 151956 7924 152124 7980
rect 151956 7868 152012 7924
rect 151788 7812 152012 7868
rect 151788 7642 151844 7812
rect 151788 7590 151790 7642
rect 151842 7590 151844 7642
rect 151788 7578 151844 7590
rect 151508 6804 151676 6860
rect 151508 6636 151564 6804
rect 151508 6570 151564 6580
rect 151732 6690 151788 6702
rect 151732 6638 151734 6690
rect 151786 6638 151788 6690
rect 151732 6636 151788 6638
rect 151732 6570 151788 6580
rect 151788 5852 151844 5862
rect 151788 5292 151844 5796
rect 151788 5226 151844 5236
rect 151340 4564 151452 4620
rect 151508 4620 151564 4630
rect 151284 4554 151340 4564
rect 151060 3612 151116 3622
rect 151060 3518 151116 3556
rect 150388 3222 150390 3274
rect 150442 3222 150444 3274
rect 150388 3210 150444 3222
rect 151508 3162 151564 4564
rect 151956 4396 152012 7812
rect 152180 6972 152236 6982
rect 152180 6858 152236 6916
rect 152180 6806 152182 6858
rect 152234 6806 152236 6858
rect 152180 6794 152236 6806
rect 152404 4620 152460 10388
rect 152964 9894 153020 13748
rect 153188 13804 153244 13814
rect 153188 13710 153244 13748
rect 153300 12124 153356 14200
rect 153860 14140 153916 14150
rect 153972 14140 154028 14200
rect 153916 14084 154028 14140
rect 153860 14074 153916 14084
rect 154756 13468 154812 14200
rect 154756 13402 154812 13412
rect 154980 13468 155036 13478
rect 154644 13132 154700 13142
rect 153300 12058 153356 12068
rect 153524 12124 153580 12134
rect 153524 11450 153580 12068
rect 153524 11398 153526 11450
rect 153578 11398 153580 11450
rect 153524 11386 153580 11398
rect 154532 12012 154588 12022
rect 154532 11228 154588 11956
rect 154532 11162 154588 11172
rect 154644 10892 154700 13076
rect 154756 12572 154812 12582
rect 154756 11676 154812 12516
rect 154868 11898 154924 11910
rect 154868 11846 154870 11898
rect 154922 11846 154924 11898
rect 154868 11788 154924 11846
rect 154868 11722 154924 11732
rect 154756 11610 154812 11620
rect 154644 10826 154700 10836
rect 153412 10444 153468 10454
rect 152964 9882 153076 9894
rect 152964 9830 153022 9882
rect 153074 9830 153076 9882
rect 152516 9772 152908 9828
rect 152516 9660 152572 9772
rect 152684 9660 152740 9670
rect 152516 9594 152572 9604
rect 152628 9658 152740 9660
rect 152628 9606 152686 9658
rect 152738 9606 152740 9658
rect 152628 9594 152740 9606
rect 152628 8204 152684 9594
rect 152852 8428 152908 9772
rect 152964 9818 153076 9830
rect 152964 9042 153020 9818
rect 152964 8990 152966 9042
rect 153018 8990 153020 9042
rect 152964 8978 153020 8990
rect 153076 9154 153132 9166
rect 153076 9102 153078 9154
rect 153130 9102 153132 9154
rect 153076 8540 153132 9102
rect 152964 8428 153020 8438
rect 152852 8372 152964 8428
rect 152964 8362 153020 8372
rect 152628 8138 152684 8148
rect 152964 7586 153020 7598
rect 152964 7534 152966 7586
rect 153018 7534 153020 7586
rect 152852 6130 152908 6142
rect 152852 6078 152854 6130
rect 152906 6078 152908 6130
rect 152852 6076 152908 6078
rect 152852 6010 152908 6020
rect 152852 5906 152908 5918
rect 152852 5854 152854 5906
rect 152906 5854 152908 5906
rect 152628 5404 152684 5414
rect 152628 5122 152684 5348
rect 152628 5070 152630 5122
rect 152682 5070 152684 5122
rect 152628 5058 152684 5070
rect 151956 4330 152012 4340
rect 152180 4564 152460 4620
rect 152852 4956 152908 5854
rect 152180 3948 152236 4564
rect 152852 4508 152908 4900
rect 152852 4442 152908 4452
rect 152180 3882 152236 3892
rect 152292 4396 152348 4406
rect 151508 3110 151510 3162
rect 151562 3110 151564 3162
rect 151508 3098 151564 3110
rect 150724 3050 150780 3062
rect 150724 2998 150726 3050
rect 150778 2998 150780 3050
rect 150164 2650 150220 2660
rect 150276 2828 150332 2838
rect 150052 2202 150108 2212
rect 150276 2154 150332 2772
rect 150276 2102 150278 2154
rect 150330 2102 150332 2154
rect 150276 2090 150332 2102
rect 150276 1708 150332 1718
rect 150276 1614 150332 1652
rect 150164 1372 150220 1382
rect 150164 800 150220 1316
rect 150724 800 150780 2998
rect 152292 2490 152348 4340
rect 152964 4172 153020 7534
rect 153076 6748 153132 8484
rect 153300 7644 153356 7654
rect 153300 7308 153356 7588
rect 153412 7474 153468 10388
rect 154644 9996 154700 10006
rect 154644 9770 154700 9940
rect 154980 9994 155036 13412
rect 155092 13356 155148 13366
rect 155092 12012 155148 13300
rect 155092 11946 155148 11956
rect 154980 9942 154982 9994
rect 155034 9942 155036 9994
rect 154980 9930 155036 9942
rect 154644 9718 154646 9770
rect 154698 9718 154700 9770
rect 154644 9706 154700 9718
rect 153580 9660 153636 9670
rect 153580 9658 153692 9660
rect 153580 9606 153582 9658
rect 153634 9606 153692 9658
rect 153580 9594 153692 9606
rect 153636 8876 153692 9594
rect 155204 9042 155260 14420
rect 155400 14200 155512 15000
rect 156184 14200 156296 15000
rect 156856 14200 156968 15000
rect 157108 14700 157164 14710
rect 157108 14364 157164 14644
rect 157108 14298 157164 14308
rect 157640 14200 157752 15000
rect 158312 14200 158424 15000
rect 158900 14252 158956 14262
rect 155316 13356 155372 13366
rect 155316 13242 155372 13300
rect 155316 13190 155318 13242
rect 155370 13190 155372 13242
rect 155316 13178 155372 13190
rect 155428 12236 155484 14200
rect 156212 14028 156268 14200
rect 156212 13962 156268 13972
rect 155428 12170 155484 12180
rect 155540 13804 155596 13814
rect 155372 9996 155428 10006
rect 155372 9882 155428 9940
rect 155372 9830 155374 9882
rect 155426 9830 155428 9882
rect 155372 9818 155428 9830
rect 155204 8990 155206 9042
rect 155258 8990 155260 9042
rect 154420 8930 154476 8942
rect 154420 8878 154422 8930
rect 154474 8878 154476 8930
rect 153636 8820 154364 8876
rect 153972 8428 154028 8438
rect 153972 8334 154028 8372
rect 153412 7422 153414 7474
rect 153466 7422 153468 7474
rect 153412 7410 153468 7422
rect 154308 8258 154364 8820
rect 154308 8206 154310 8258
rect 154362 8206 154364 8258
rect 153300 7252 153468 7308
rect 153076 6690 153132 6692
rect 153076 6638 153078 6690
rect 153130 6638 153132 6690
rect 153076 6626 153132 6638
rect 153132 4954 153188 4966
rect 153132 4902 153134 4954
rect 153186 4902 153188 4954
rect 153132 4844 153188 4902
rect 153132 4778 153188 4788
rect 153300 4508 153356 4518
rect 153076 4172 153132 4182
rect 152964 4116 153076 4172
rect 152628 4058 152684 4070
rect 152628 4006 152630 4058
rect 152682 4006 152684 4058
rect 152516 3948 152572 3958
rect 152292 2438 152294 2490
rect 152346 2438 152348 2490
rect 152292 2426 152348 2438
rect 152404 3610 152460 3622
rect 152404 3558 152406 3610
rect 152458 3558 152460 3610
rect 151284 2378 151340 2390
rect 151284 2326 151286 2378
rect 151338 2326 151340 2378
rect 151060 1932 151116 1942
rect 151060 1838 151116 1876
rect 151284 800 151340 2326
rect 152404 1820 152460 3558
rect 152516 3386 152572 3892
rect 152516 3334 152518 3386
rect 152570 3334 152572 3386
rect 152516 3322 152572 3334
rect 152628 3052 152684 4006
rect 153076 3948 153132 4116
rect 153076 3882 153132 3892
rect 153076 3722 153132 3734
rect 153076 3670 153078 3722
rect 153130 3670 153132 3722
rect 152628 2986 152684 2996
rect 152852 3386 152908 3398
rect 152852 3334 152854 3386
rect 152906 3334 152908 3386
rect 152628 2492 152684 2502
rect 152628 2398 152684 2436
rect 152404 1754 152460 1764
rect 152516 2380 152572 2390
rect 151956 924 152012 934
rect 151956 800 152012 868
rect 152516 800 152572 2324
rect 152852 2268 152908 3334
rect 153076 2938 153132 3670
rect 153188 3724 153244 3734
rect 153188 3500 153244 3668
rect 153300 3722 153356 4452
rect 153412 4170 153468 7252
rect 153748 7306 153804 7318
rect 153748 7254 153750 7306
rect 153802 7254 153804 7306
rect 153748 7196 153804 7254
rect 153748 7130 153804 7140
rect 154308 7084 154364 8206
rect 154420 7420 154476 8878
rect 154420 7354 154476 7364
rect 154196 7028 154364 7084
rect 153692 6636 153748 6646
rect 153692 6542 153748 6580
rect 153580 4954 153636 4966
rect 153580 4902 153582 4954
rect 153634 4902 153636 4954
rect 153580 4732 153636 4902
rect 153580 4666 153636 4676
rect 153412 4118 153414 4170
rect 153466 4118 153468 4170
rect 153412 4106 153468 4118
rect 153300 3670 153302 3722
rect 153354 3670 153356 3722
rect 153300 3658 153356 3670
rect 153188 3434 153244 3444
rect 153076 2886 153078 2938
rect 153130 2886 153132 2938
rect 153076 2874 153132 2886
rect 152852 2202 152908 2212
rect 153188 2604 153244 2614
rect 153188 800 153244 2548
rect 154196 2490 154252 7028
rect 154980 6636 155036 6646
rect 154308 6524 154364 6534
rect 154308 5906 154364 6468
rect 154532 6466 154588 6478
rect 154532 6414 154534 6466
rect 154586 6414 154588 6466
rect 154532 6412 154588 6414
rect 154532 6346 154588 6356
rect 154700 6412 154756 6422
rect 154700 6074 154756 6356
rect 154700 6022 154702 6074
rect 154754 6022 154756 6074
rect 154700 6010 154756 6022
rect 154980 6412 155036 6580
rect 154308 5854 154310 5906
rect 154362 5854 154364 5906
rect 154308 5842 154364 5854
rect 154980 4966 155036 6356
rect 155204 6086 155260 8990
rect 155428 8874 155484 8886
rect 155428 8822 155430 8874
rect 155482 8822 155484 8874
rect 155316 7306 155372 7318
rect 155316 7254 155318 7306
rect 155370 7254 155372 7306
rect 155316 6748 155372 7254
rect 155428 7308 155484 8822
rect 155428 7242 155484 7252
rect 155540 7474 155596 13748
rect 156884 12460 156940 14200
rect 157668 13916 157724 14200
rect 157668 13850 157724 13860
rect 158340 13916 158396 14200
rect 158340 13850 158396 13860
rect 159096 14200 159208 15000
rect 159768 14200 159880 15000
rect 160552 14200 160664 15000
rect 161224 14200 161336 15000
rect 161532 14924 161588 14934
rect 161476 14868 161532 14924
rect 161476 14858 161588 14868
rect 156884 12394 156940 12404
rect 157220 13580 157276 13590
rect 156436 11676 156492 11686
rect 156212 11620 156436 11676
rect 156212 10444 156268 11620
rect 156436 11610 156492 11620
rect 157108 11676 157164 11686
rect 156436 10444 156492 10454
rect 156212 10378 156268 10388
rect 156324 10388 156436 10444
rect 156324 9826 156380 10388
rect 156436 10378 156492 10388
rect 156324 9774 156326 9826
rect 156378 9774 156380 9826
rect 156324 9772 156380 9774
rect 156212 9716 156380 9772
rect 155988 8258 156044 8270
rect 155988 8206 155990 8258
rect 156042 8206 156044 8258
rect 155988 8204 156044 8206
rect 155988 8138 156044 8148
rect 156212 7868 156268 9716
rect 156324 9602 156380 9614
rect 156324 9550 156326 9602
rect 156378 9550 156380 9602
rect 156324 9436 156380 9550
rect 156324 9370 156380 9380
rect 156324 9042 156380 9054
rect 156324 8990 156326 9042
rect 156378 8990 156380 9042
rect 156324 8092 156380 8990
rect 156604 8092 156660 8102
rect 156324 8090 156660 8092
rect 156324 8038 156606 8090
rect 156658 8038 156660 8090
rect 156324 8036 156660 8038
rect 156548 8026 156660 8036
rect 156212 7812 156380 7868
rect 155540 7422 155542 7474
rect 155594 7422 155596 7474
rect 155316 6682 155372 6692
rect 155540 6636 155596 7422
rect 155428 6578 155484 6590
rect 155428 6526 155430 6578
rect 155482 6526 155484 6578
rect 155988 7644 156044 7654
rect 155988 6690 156044 7588
rect 155988 6638 155990 6690
rect 156042 6638 156044 6690
rect 155988 6626 156044 6638
rect 156100 7586 156156 7598
rect 156100 7534 156102 7586
rect 156154 7534 156156 7586
rect 155540 6570 155596 6580
rect 155204 6074 155316 6086
rect 155204 6022 155262 6074
rect 155314 6022 155316 6074
rect 155204 6020 155316 6022
rect 155260 6010 155316 6020
rect 155428 4966 155484 6526
rect 156100 6412 156156 7534
rect 156100 6346 156156 6356
rect 156100 5906 156156 5918
rect 156100 5854 156102 5906
rect 156154 5854 156156 5906
rect 154476 4956 154532 4966
rect 154476 4862 154532 4900
rect 154924 4954 155036 4966
rect 155372 4956 155484 4966
rect 154924 4902 154926 4954
rect 154978 4902 155036 4954
rect 154924 4900 155036 4902
rect 155316 4954 155484 4956
rect 155316 4902 155374 4954
rect 155426 4902 155484 4954
rect 155316 4900 155484 4902
rect 155652 5628 155708 5638
rect 154924 4890 154980 4900
rect 155316 4890 155428 4900
rect 154644 4732 154700 4742
rect 154420 4172 154476 4182
rect 154420 2826 154476 4116
rect 154644 3388 154700 4676
rect 155316 4060 155372 4890
rect 155652 4508 155708 5572
rect 156100 5292 156156 5854
rect 155652 4442 155708 4452
rect 155988 5236 156156 5292
rect 155988 4732 156044 5236
rect 155316 3994 155372 4004
rect 154644 3322 154700 3332
rect 154868 3498 154924 3510
rect 154868 3446 154870 3498
rect 154922 3446 154924 3498
rect 154532 3164 154588 3174
rect 154532 2940 154588 3108
rect 154532 2884 154812 2940
rect 154420 2774 154422 2826
rect 154474 2774 154476 2826
rect 154420 2762 154476 2774
rect 154196 2438 154198 2490
rect 154250 2438 154252 2490
rect 154196 2426 154252 2438
rect 154532 2492 154588 2502
rect 154532 2398 154588 2436
rect 154756 2492 154812 2884
rect 154756 2426 154812 2436
rect 153860 2268 153916 2278
rect 153860 2174 153916 2212
rect 154420 2154 154476 2166
rect 154420 2102 154422 2154
rect 154474 2102 154476 2154
rect 153748 1036 153804 1046
rect 153748 800 153804 980
rect 154420 800 154476 2102
rect 154868 1484 154924 3446
rect 154868 1418 154924 1428
rect 154980 3050 155036 3062
rect 154980 2998 154982 3050
rect 155034 2998 155036 3050
rect 154980 800 155036 2998
rect 155988 2716 156044 4676
rect 156100 5122 156156 5134
rect 156100 5070 156102 5122
rect 156154 5070 156156 5122
rect 156100 4508 156156 5070
rect 156100 4442 156156 4452
rect 156212 5010 156268 5022
rect 156212 4958 156214 5010
rect 156266 4958 156268 5010
rect 156100 4284 156156 4294
rect 156100 4190 156156 4228
rect 155988 2650 156044 2660
rect 155652 2266 155708 2278
rect 155652 2214 155654 2266
rect 155706 2214 155708 2266
rect 155652 800 155708 2214
rect 155988 1818 156044 1830
rect 155988 1766 155990 1818
rect 156042 1766 156044 1818
rect 155988 1708 156044 1766
rect 155988 1642 156044 1652
rect 156212 800 156268 4958
rect 156324 3610 156380 7812
rect 156548 6524 156604 8026
rect 157108 7654 157164 11620
rect 157220 9436 157276 13524
rect 158788 12234 158844 12246
rect 158788 12182 158790 12234
rect 158842 12182 158844 12234
rect 158788 10892 158844 12182
rect 158788 10826 158844 10836
rect 158900 10668 158956 14196
rect 159124 13356 159180 14200
rect 159572 14028 159628 14038
rect 159124 13290 159180 13300
rect 159236 13802 159292 13814
rect 159236 13750 159238 13802
rect 159290 13750 159292 13802
rect 159012 11900 159068 11910
rect 159012 10892 159068 11844
rect 159236 11564 159292 13750
rect 159236 11498 159292 11508
rect 159348 13020 159404 13030
rect 159012 10826 159068 10836
rect 159236 11116 159292 11126
rect 159236 10668 159292 11060
rect 158900 10612 159068 10668
rect 157780 10220 157836 10230
rect 157780 9826 157836 10164
rect 157780 9774 157782 9826
rect 157834 9774 157836 9826
rect 157780 9762 157836 9774
rect 158676 9772 158732 9782
rect 157220 9042 157276 9380
rect 157220 8990 157222 9042
rect 157274 8990 157276 9042
rect 157220 8978 157276 8990
rect 158564 9658 158620 9670
rect 158564 9606 158566 9658
rect 158618 9606 158620 9658
rect 158564 9100 158620 9606
rect 157780 8874 157836 8886
rect 157780 8822 157782 8874
rect 157834 8822 157836 8874
rect 157780 8540 157836 8822
rect 157780 8474 157836 8484
rect 158564 8428 158620 9044
rect 158564 8362 158620 8372
rect 158676 9042 158732 9716
rect 158900 9660 158956 9670
rect 158676 8990 158678 9042
rect 158730 8990 158732 9042
rect 158676 8260 158732 8990
rect 158228 8204 158732 8260
rect 158788 9658 158956 9660
rect 158788 9606 158902 9658
rect 158954 9606 158956 9658
rect 158788 9604 158956 9606
rect 157108 7642 157220 7654
rect 157108 7590 157166 7642
rect 157218 7590 157220 7642
rect 157108 7588 157220 7590
rect 157164 7578 157220 7588
rect 156716 7420 156772 7430
rect 157612 7420 157668 7430
rect 156548 6458 156604 6468
rect 156660 7418 156772 7420
rect 156660 7366 156718 7418
rect 156770 7366 156772 7418
rect 156660 7354 156772 7366
rect 157556 7418 157668 7420
rect 157556 7366 157614 7418
rect 157666 7366 157668 7418
rect 157556 7354 157668 7366
rect 156324 3558 156326 3610
rect 156378 3558 156380 3610
rect 156324 3546 156380 3558
rect 156436 4956 156492 4966
rect 156436 3498 156492 4900
rect 156660 4060 156716 7354
rect 157332 6860 157388 6870
rect 157332 6766 157388 6804
rect 156772 6690 156828 6702
rect 156772 6638 156774 6690
rect 156826 6638 156828 6690
rect 156772 6412 156828 6638
rect 157556 6636 157612 7354
rect 157556 6570 157612 6580
rect 158228 6690 158284 8204
rect 158564 8092 158620 8102
rect 158564 7644 158620 8036
rect 158228 6638 158230 6690
rect 158282 6638 158284 6690
rect 158228 6524 158284 6638
rect 158228 6458 158284 6468
rect 158452 7362 158508 7374
rect 158452 7310 158454 7362
rect 158506 7310 158508 7362
rect 156772 6346 156828 6356
rect 157556 6412 157612 6422
rect 157556 5906 157612 6356
rect 157556 5854 157558 5906
rect 157610 5854 157612 5906
rect 157556 5842 157612 5854
rect 158116 6188 158172 6198
rect 158116 5906 158172 6132
rect 158116 5854 158118 5906
rect 158170 5854 158172 5906
rect 158116 5842 158172 5854
rect 156996 5740 157052 5750
rect 156996 5646 157052 5684
rect 157444 5068 157500 5078
rect 156660 3994 156716 4004
rect 156772 4172 156828 4182
rect 156436 3446 156438 3498
rect 156490 3446 156492 3498
rect 156436 3434 156492 3446
rect 156436 1818 156492 1830
rect 156436 1766 156438 1818
rect 156490 1766 156492 1818
rect 156436 1708 156492 1766
rect 156436 1642 156492 1652
rect 156772 800 156828 4116
rect 157444 800 157500 5012
rect 158452 3387 158508 7310
rect 158564 5122 158620 7588
rect 158564 5070 158566 5122
rect 158618 5070 158620 5122
rect 158676 6188 158732 6198
rect 158676 5180 158732 6132
rect 158676 5114 158732 5124
rect 158564 5058 158620 5070
rect 158676 5010 158732 5022
rect 158676 4958 158678 5010
rect 158730 4958 158732 5010
rect 158676 4172 158732 4958
rect 158676 4106 158732 4116
rect 158788 4060 158844 9604
rect 158900 9594 158956 9604
rect 158900 8428 158956 8438
rect 159012 8428 159068 10612
rect 159236 10602 159292 10612
rect 159124 10444 159180 10454
rect 159124 9222 159180 10388
rect 159348 9884 159404 12964
rect 159572 12122 159628 13972
rect 159796 13244 159852 14200
rect 159796 13178 159852 13188
rect 160580 12348 160636 14200
rect 161252 14140 161308 14200
rect 161476 14140 161532 14858
rect 162008 14200 162120 15000
rect 162484 14700 162540 14710
rect 162260 14588 162316 14598
rect 161252 14084 161532 14140
rect 161252 13578 161308 13590
rect 161252 13526 161254 13578
rect 161306 13526 161308 13578
rect 160580 12282 160636 12292
rect 161028 13020 161084 13030
rect 159572 12070 159574 12122
rect 159626 12070 159628 12122
rect 159572 12058 159628 12070
rect 159460 11788 159516 11798
rect 159460 11340 159516 11732
rect 159460 11274 159516 11284
rect 160916 11564 160972 11574
rect 159348 9826 159404 9828
rect 159348 9774 159350 9826
rect 159402 9774 159404 9826
rect 160804 9826 160860 9838
rect 159348 9752 159404 9774
rect 159628 9772 159684 9782
rect 159124 9210 159236 9222
rect 159124 9158 159182 9210
rect 159234 9158 159236 9210
rect 159124 9156 159236 9158
rect 159180 9146 159236 9156
rect 159628 9210 159684 9716
rect 160804 9774 160806 9826
rect 160858 9774 160860 9826
rect 160804 9772 160860 9774
rect 160804 9706 160860 9716
rect 159628 9158 159630 9210
rect 159682 9158 159684 9210
rect 159628 9146 159684 9158
rect 160580 9602 160636 9614
rect 160580 9550 160582 9602
rect 160634 9550 160636 9602
rect 158900 8426 159068 8428
rect 158900 8374 158902 8426
rect 158954 8374 159068 8426
rect 158900 8372 159068 8374
rect 158900 8362 158956 8372
rect 160580 8316 160636 9550
rect 160916 9436 160972 11508
rect 160860 9380 160972 9436
rect 160860 9042 160916 9380
rect 160860 8990 160862 9042
rect 160914 8990 160916 9042
rect 160748 8876 160804 8886
rect 159236 8260 159292 8270
rect 159124 8258 159292 8260
rect 159124 8206 159238 8258
rect 159290 8206 159292 8258
rect 160580 8250 160636 8260
rect 160692 8874 160804 8876
rect 160692 8822 160750 8874
rect 160802 8822 160804 8874
rect 160692 8810 160804 8822
rect 159124 8204 159292 8206
rect 159012 6578 159068 6590
rect 159012 6526 159014 6578
rect 159066 6526 159068 6578
rect 159012 5068 159068 6526
rect 159012 5002 159068 5012
rect 158788 4004 159068 4060
rect 158004 3331 158508 3387
rect 158788 3834 158844 3846
rect 158788 3782 158790 3834
rect 158842 3782 158844 3834
rect 158004 800 158060 3331
rect 158788 2828 158844 3782
rect 159012 3387 159068 4004
rect 159124 4058 159180 8204
rect 159236 8194 159292 8204
rect 160692 8204 160748 8810
rect 160860 8540 160916 8990
rect 160692 8138 160748 8148
rect 160804 8484 160916 8540
rect 160804 7980 160860 8484
rect 160468 7924 160860 7980
rect 160916 8258 160972 8270
rect 160916 8206 160918 8258
rect 160970 8206 160972 8258
rect 159460 7644 159516 7654
rect 159460 7474 159516 7588
rect 159460 7422 159462 7474
rect 159514 7422 159516 7474
rect 159460 7196 159516 7422
rect 159460 7130 159516 7140
rect 159348 6690 159404 6702
rect 159348 6638 159350 6690
rect 159402 6638 159404 6690
rect 159348 5292 159404 6638
rect 159460 6076 159516 6086
rect 159460 6018 159516 6020
rect 159460 5966 159462 6018
rect 159514 5966 159516 6018
rect 159460 5954 159516 5966
rect 159348 5068 159404 5236
rect 159348 5002 159404 5012
rect 159460 5180 159516 5190
rect 159124 4006 159126 4058
rect 159178 4006 159180 4058
rect 159124 3994 159180 4006
rect 159236 4172 159292 4182
rect 159012 3331 159180 3387
rect 158676 2772 158844 2828
rect 158676 800 158732 2772
rect 159124 2156 159180 3331
rect 159124 2090 159180 2100
rect 159236 800 159292 4116
rect 159460 3834 159516 5124
rect 159460 3782 159462 3834
rect 159514 3782 159516 3834
rect 159460 3770 159516 3782
rect 159908 4284 159964 4294
rect 159908 800 159964 4228
rect 160468 3276 160524 7924
rect 160916 6636 160972 8206
rect 161028 7306 161084 12964
rect 161252 11116 161308 13526
rect 161252 11050 161308 11060
rect 161476 13356 161532 13366
rect 161476 10220 161532 13300
rect 161924 12908 161980 12918
rect 162036 12908 162092 14200
rect 161980 12852 162092 12908
rect 161924 12842 161980 12852
rect 161476 9894 161532 10164
rect 161420 9882 161532 9894
rect 161420 9830 161422 9882
rect 161474 9830 161532 9882
rect 161420 9828 161532 9830
rect 161420 9818 161476 9828
rect 161588 9772 161644 9782
rect 161308 9436 161364 9446
rect 161308 9210 161364 9380
rect 161308 9158 161310 9210
rect 161362 9158 161364 9210
rect 161308 9146 161364 9158
rect 161476 8258 161532 8270
rect 161476 8206 161478 8258
rect 161530 8206 161532 8258
rect 161028 7254 161030 7306
rect 161082 7254 161084 7306
rect 161028 7242 161084 7254
rect 161364 7644 161420 7654
rect 160916 6570 160972 6580
rect 161140 6690 161196 6702
rect 161140 6638 161142 6690
rect 161194 6638 161196 6690
rect 160636 6524 160692 6534
rect 160636 6076 160692 6468
rect 160580 6074 160692 6076
rect 160580 6022 160638 6074
rect 160690 6022 160692 6074
rect 160580 6010 160692 6022
rect 160580 5740 160636 6010
rect 160580 5674 160636 5684
rect 160748 5740 160804 5750
rect 160748 5404 160804 5684
rect 161140 5628 161196 6638
rect 161364 6524 161420 7588
rect 161476 7532 161532 8206
rect 161476 7466 161532 7476
rect 161364 6458 161420 6468
rect 161588 5908 161644 9716
rect 161756 9100 161812 9110
rect 161756 9006 161812 9044
rect 162260 6074 162316 14532
rect 162372 12010 162428 12022
rect 162372 11958 162374 12010
rect 162426 11958 162428 12010
rect 162372 10556 162428 11958
rect 162372 9826 162428 10500
rect 162372 9774 162374 9826
rect 162426 9774 162428 9826
rect 162372 9762 162428 9774
rect 162484 8764 162540 14644
rect 162680 14200 162792 15000
rect 163268 14700 163324 14710
rect 162708 14028 162764 14200
rect 162708 13962 162764 13972
rect 162820 12458 162876 12470
rect 162820 12406 162822 12458
rect 162874 12406 162876 12458
rect 162708 12124 162764 12134
rect 162708 8876 162764 12068
rect 162820 11900 162876 12406
rect 162820 11834 162876 11844
rect 162932 12236 162988 12246
rect 162932 11116 162988 12180
rect 162932 11050 162988 11060
rect 162820 8876 162876 8886
rect 162708 8874 162876 8876
rect 162708 8822 162822 8874
rect 162874 8822 162876 8874
rect 162708 8820 162876 8822
rect 162820 8810 162876 8820
rect 162484 8708 162764 8764
rect 162260 6022 162262 6074
rect 162314 6022 162316 6074
rect 162260 6010 162316 6022
rect 162372 8146 162428 8158
rect 162372 8094 162374 8146
rect 162426 8094 162428 8146
rect 161140 5562 161196 5572
rect 161476 5852 161644 5908
rect 160748 4954 160804 5348
rect 161476 4966 161532 5852
rect 161084 4956 161140 4966
rect 160748 4902 160750 4954
rect 160802 4902 160804 4954
rect 160748 4890 160804 4902
rect 161028 4954 161140 4956
rect 161028 4902 161086 4954
rect 161138 4902 161140 4954
rect 161028 4890 161140 4902
rect 161476 4954 161588 4966
rect 161476 4902 161534 4954
rect 161586 4902 161588 4954
rect 161476 4900 161588 4902
rect 161532 4890 161588 4900
rect 161028 4058 161084 4890
rect 161028 4006 161030 4058
rect 161082 4006 161084 4058
rect 161028 3994 161084 4006
rect 161700 4620 161756 4630
rect 160468 3210 160524 3220
rect 161140 3276 161196 3286
rect 161028 3162 161084 3174
rect 161028 3110 161030 3162
rect 161082 3110 161084 3162
rect 161028 2380 161084 3110
rect 161028 2314 161084 2324
rect 160468 1596 160524 1606
rect 160468 800 160524 1540
rect 161140 800 161196 3220
rect 161700 800 161756 4564
rect 162260 2044 162316 2054
rect 162260 800 162316 1988
rect 162372 1932 162428 8094
rect 162596 7756 162652 7766
rect 162596 7474 162652 7700
rect 162596 7422 162598 7474
rect 162650 7422 162652 7474
rect 162484 6578 162540 6590
rect 162484 6526 162486 6578
rect 162538 6526 162540 6578
rect 162484 5404 162540 6526
rect 162484 5338 162540 5348
rect 162596 4396 162652 7422
rect 162708 5234 162764 8708
rect 163268 7868 163324 14644
rect 163464 14200 163576 15000
rect 164136 14200 164248 15000
rect 164920 14200 165032 15000
rect 165704 14200 165816 15000
rect 166376 14200 166488 15000
rect 167160 14200 167272 15000
rect 167524 14586 167580 14598
rect 167524 14534 167526 14586
rect 167578 14534 167580 14586
rect 163492 13692 163548 14200
rect 163492 13626 163548 13636
rect 163940 13580 163996 13590
rect 163828 11340 163884 11350
rect 163716 9772 163772 9782
rect 163716 9714 163772 9716
rect 163716 9662 163718 9714
rect 163770 9662 163772 9714
rect 163716 9650 163772 9662
rect 163268 6646 163324 7812
rect 163604 9602 163660 9614
rect 163604 9550 163606 9602
rect 163658 9550 163660 9602
rect 163604 7532 163660 9550
rect 163828 8270 163884 11284
rect 163940 8428 163996 13524
rect 164164 13468 164220 14200
rect 164164 13402 164220 13412
rect 164948 13244 165004 14200
rect 164948 13178 165004 13188
rect 165060 13242 165116 13254
rect 165060 13190 165062 13242
rect 165114 13190 165116 13242
rect 164052 12460 164108 12470
rect 164052 9996 164108 12404
rect 165060 12236 165116 13190
rect 165732 13020 165788 14200
rect 165732 12954 165788 12964
rect 165060 12170 165116 12180
rect 165620 11900 165676 11910
rect 164612 11786 164668 11798
rect 164612 11734 164614 11786
rect 164666 11734 164668 11786
rect 164612 11452 164668 11734
rect 164612 11386 164668 11396
rect 165284 11564 165340 11574
rect 164052 9212 164108 9940
rect 165284 10556 165340 11508
rect 164332 9884 164388 9894
rect 164332 9790 164388 9828
rect 165284 9770 165340 10500
rect 165620 9994 165676 11844
rect 165620 9942 165622 9994
rect 165674 9942 165676 9994
rect 165620 9930 165676 9942
rect 165732 11788 165788 11798
rect 165284 9718 165286 9770
rect 165338 9718 165340 9770
rect 165284 9706 165340 9718
rect 164196 9436 164460 9446
rect 164252 9380 164300 9436
rect 164356 9380 164404 9436
rect 164196 9370 164460 9380
rect 164052 9156 164444 9212
rect 164388 9042 164444 9156
rect 164388 8990 164390 9042
rect 164442 8990 164444 9042
rect 164388 8978 164444 8990
rect 163940 8372 164108 8428
rect 163828 8258 163940 8270
rect 163828 8206 163886 8258
rect 163938 8206 163940 8258
rect 163828 8204 163940 8206
rect 163884 8194 163940 8204
rect 163604 7466 163660 7476
rect 163772 8090 163828 8102
rect 163772 8038 163774 8090
rect 163826 8038 163828 8090
rect 163772 7420 163828 8038
rect 163772 7364 163884 7420
rect 163268 6634 163380 6646
rect 163268 6582 163326 6634
rect 163378 6582 163380 6634
rect 163268 6580 163380 6582
rect 163324 6570 163380 6580
rect 163828 6636 163884 7364
rect 163828 6570 163884 6580
rect 163660 6524 163716 6534
rect 162708 5182 162710 5234
rect 162762 5182 162764 5234
rect 162708 5170 162764 5182
rect 163604 6522 163716 6524
rect 163604 6470 163662 6522
rect 163714 6470 163716 6522
rect 163604 6458 163716 6470
rect 163604 4732 163660 6458
rect 163828 5908 163884 5918
rect 164052 5908 164108 8372
rect 164724 8258 164780 8270
rect 164724 8206 164726 8258
rect 164778 8206 164780 8258
rect 164196 7868 164460 7878
rect 164252 7812 164300 7868
rect 164356 7812 164404 7868
rect 164196 7802 164460 7812
rect 164276 7644 164332 7654
rect 164276 7474 164332 7588
rect 164276 7422 164278 7474
rect 164330 7422 164332 7474
rect 164276 7410 164332 7422
rect 164612 7196 164668 7206
rect 164724 7196 164780 8206
rect 164836 7474 164892 7486
rect 164836 7422 164838 7474
rect 164890 7422 164892 7474
rect 164836 7420 164892 7422
rect 164836 7354 164892 7364
rect 164668 7140 164780 7196
rect 164836 7196 164892 7206
rect 164612 7130 164668 7140
rect 164556 6522 164612 6534
rect 164556 6470 164558 6522
rect 164610 6470 164612 6522
rect 164196 6300 164460 6310
rect 164252 6244 164300 6300
rect 164356 6244 164404 6300
rect 164196 6234 164460 6244
rect 164556 6188 164612 6470
rect 163828 5906 164108 5908
rect 163828 5854 163830 5906
rect 163882 5854 164108 5906
rect 163828 5852 164108 5854
rect 164500 6132 164612 6188
rect 163828 5516 163884 5852
rect 163828 5450 163884 5460
rect 164500 5292 164556 6132
rect 164836 5906 164892 7140
rect 165004 6524 165060 6534
rect 165004 6430 165060 6468
rect 164836 5854 164838 5906
rect 164890 5854 164892 5906
rect 164836 5842 164892 5854
rect 165396 5964 165452 5974
rect 165396 5906 165452 5908
rect 165396 5854 165398 5906
rect 165450 5854 165452 5906
rect 164500 5226 164556 5236
rect 165396 5292 165452 5854
rect 165396 5226 165452 5236
rect 164052 5122 164108 5134
rect 164052 5070 164054 5122
rect 164106 5070 164108 5122
rect 164052 5068 164108 5070
rect 164052 5002 164108 5012
rect 164556 4954 164612 4966
rect 164556 4902 164558 4954
rect 164610 4902 164612 4954
rect 163604 4666 163660 4676
rect 164196 4732 164460 4742
rect 164252 4676 164300 4732
rect 164356 4676 164404 4732
rect 164196 4666 164460 4676
rect 164556 4508 164612 4902
rect 165116 4954 165172 4966
rect 165116 4902 165118 4954
rect 165170 4902 165172 4954
rect 165116 4732 165172 4902
rect 165452 4956 165508 4966
rect 165452 4862 165508 4900
rect 165116 4666 165172 4676
rect 164556 4442 164612 4452
rect 162596 4330 162652 4340
rect 165172 3948 165228 3958
rect 162708 2828 162764 2838
rect 162708 2734 162764 2772
rect 165172 2044 165228 3892
rect 165732 2380 165788 11732
rect 166404 11788 166460 14200
rect 167188 12124 167244 14200
rect 167188 12058 167244 12068
rect 166404 11722 166460 11732
rect 166628 11114 166684 11126
rect 166628 11062 166630 11114
rect 166682 11062 166684 11114
rect 166628 10332 166684 11062
rect 166628 10266 166684 10276
rect 166628 9826 166684 9838
rect 166460 9772 166516 9782
rect 166460 9324 166516 9716
rect 166460 9210 166516 9268
rect 166460 9158 166462 9210
rect 166514 9158 166516 9210
rect 166460 9146 166516 9158
rect 166628 9774 166630 9826
rect 166682 9774 166684 9826
rect 166628 9660 166684 9774
rect 166068 9100 166124 9110
rect 166068 9042 166124 9044
rect 166068 8990 166070 9042
rect 166122 8990 166124 9042
rect 166068 8978 166124 8990
rect 166628 8204 166684 9604
rect 166068 8146 166124 8158
rect 166068 8094 166070 8146
rect 166122 8094 166124 8146
rect 166628 8138 166684 8148
rect 166740 9714 166796 9726
rect 166740 9662 166742 9714
rect 166794 9662 166796 9714
rect 165844 6412 165900 6422
rect 165844 2828 165900 6356
rect 166068 5124 166124 8094
rect 166180 7362 166236 7374
rect 166180 7310 166182 7362
rect 166234 7310 166236 7362
rect 166180 5516 166236 7310
rect 166404 6188 166460 6198
rect 166180 5450 166236 5460
rect 166292 5794 166348 5806
rect 166292 5742 166294 5794
rect 166346 5742 166348 5794
rect 166292 5180 166348 5742
rect 166068 5068 166236 5124
rect 166292 5114 166348 5124
rect 166404 5122 166460 6132
rect 166628 6188 166684 6198
rect 166628 5628 166684 6132
rect 166628 5562 166684 5572
rect 166180 4956 166236 5068
rect 166404 5070 166406 5122
rect 166458 5070 166460 5122
rect 166292 4956 166348 4966
rect 166180 4900 166292 4956
rect 166292 4890 166348 4900
rect 166404 4058 166460 5070
rect 166516 5010 166572 5022
rect 166516 4958 166518 5010
rect 166570 4958 166572 5010
rect 166516 4172 166572 4958
rect 166516 4106 166572 4116
rect 166404 4006 166406 4058
rect 166458 4006 166460 4058
rect 166404 3994 166460 4006
rect 166740 3724 166796 9662
rect 166852 9324 166908 9334
rect 166852 8998 166908 9268
rect 166852 8986 166964 8998
rect 166852 8934 166910 8986
rect 166962 8934 166964 8986
rect 166852 8922 166964 8934
rect 166852 7476 166908 8922
rect 166964 8316 167020 8326
rect 166964 8258 167020 8260
rect 166964 8206 166966 8258
rect 167018 8206 167020 8258
rect 166964 8194 167020 8206
rect 167412 8146 167468 8158
rect 167412 8094 167414 8146
rect 167466 8094 167468 8146
rect 166964 7980 167020 7990
rect 166964 7642 167020 7924
rect 166964 7590 166966 7642
rect 167018 7590 167020 7642
rect 166964 7578 167020 7590
rect 167300 7530 167356 7542
rect 167300 7478 167302 7530
rect 167354 7478 167356 7530
rect 166852 7420 167020 7476
rect 166852 6636 166908 6646
rect 166852 6522 166908 6580
rect 166852 6470 166854 6522
rect 166906 6470 166908 6522
rect 166852 6458 166908 6470
rect 166964 5628 167020 7420
rect 167300 5964 167356 7478
rect 167300 5898 167356 5908
rect 166964 5562 167020 5572
rect 167076 5516 167132 5526
rect 166964 4396 167020 4406
rect 166964 4060 167020 4340
rect 166964 3994 167020 4004
rect 166740 3658 166796 3668
rect 167076 3724 167132 5460
rect 167076 3658 167132 3668
rect 167188 5404 167244 5414
rect 167076 3052 167132 3062
rect 165844 2772 166012 2828
rect 165732 2314 165788 2324
rect 165172 1978 165228 1988
rect 165396 2044 165452 2054
rect 162372 1866 162428 1876
rect 162932 1596 162988 1606
rect 162932 800 162988 1540
rect 164724 1596 164780 1606
rect 163492 1372 163548 1382
rect 163492 800 163548 1316
rect 164164 1260 164220 1270
rect 164164 800 164220 1204
rect 164724 800 164780 1540
rect 165396 800 165452 1988
rect 165956 800 166012 2772
rect 167076 2380 167132 2996
rect 167076 2314 167132 2324
rect 166516 1596 166572 1606
rect 166516 800 166572 1540
rect 167188 800 167244 5348
rect 167412 1596 167468 8094
rect 167524 6074 167580 14534
rect 167832 14200 167944 15000
rect 168616 14200 168728 15000
rect 169092 14252 169148 14262
rect 167860 13132 167916 14200
rect 167860 13066 167916 13076
rect 168644 11900 168700 14200
rect 169288 14200 169400 15000
rect 169764 14476 169820 14486
rect 169092 14140 169148 14196
rect 169316 14140 169372 14200
rect 169092 14084 169372 14140
rect 169764 14140 169820 14420
rect 170072 14200 170184 15000
rect 170744 14200 170856 15000
rect 171332 14364 171388 14374
rect 170100 14140 170156 14200
rect 169764 14084 170156 14140
rect 168644 11834 168700 11844
rect 169428 12460 169484 12470
rect 167636 10556 167692 10566
rect 167636 7476 167692 10500
rect 168868 10332 168924 10342
rect 168700 10220 168756 10230
rect 167860 10108 167916 10118
rect 167860 9660 167916 10052
rect 168700 9882 168756 10164
rect 168700 9830 168702 9882
rect 168754 9830 168756 9882
rect 168700 9818 168756 9830
rect 167860 9604 167972 9660
rect 167916 9154 167972 9604
rect 167916 9102 167918 9154
rect 167970 9102 167972 9154
rect 167916 9090 167972 9102
rect 168868 9042 168924 10276
rect 169148 9660 169204 9670
rect 168868 8990 168870 9042
rect 168922 8990 168924 9042
rect 168868 8978 168924 8990
rect 169092 9658 169204 9660
rect 169092 9606 169150 9658
rect 169202 9606 169204 9658
rect 169092 9594 169204 9606
rect 169316 9660 169372 9670
rect 167804 8876 167860 8886
rect 167748 8874 167860 8876
rect 167748 8822 167806 8874
rect 167858 8822 167860 8874
rect 167748 8810 167860 8822
rect 167748 7644 167804 8810
rect 167748 7578 167804 7588
rect 168756 8540 168812 8550
rect 167860 7532 167916 7542
rect 167636 7420 167916 7476
rect 167804 7418 167860 7420
rect 167804 7366 167806 7418
rect 167858 7366 167860 7418
rect 167804 7354 167860 7366
rect 167524 6022 167526 6074
rect 167578 6022 167580 6074
rect 167524 6010 167580 6022
rect 167636 6690 167692 6702
rect 167636 6638 167638 6690
rect 167690 6638 167692 6690
rect 167636 6636 167692 6638
rect 167636 5180 167692 6580
rect 167860 5962 167916 5974
rect 167860 5910 167862 5962
rect 167914 5910 167916 5962
rect 167860 5516 167916 5910
rect 168756 5906 168812 8484
rect 169092 8316 169148 9594
rect 169204 8988 169260 8998
rect 169204 8874 169260 8932
rect 169204 8822 169206 8874
rect 169258 8822 169260 8874
rect 169204 8810 169260 8822
rect 169316 8540 169372 9604
rect 169092 8250 169148 8260
rect 169204 8484 169372 8540
rect 168868 7308 168924 7318
rect 168868 6300 168924 7252
rect 169204 6709 169260 8484
rect 169204 6657 169206 6709
rect 169258 6657 169260 6709
rect 169204 6645 169260 6657
rect 169316 8146 169372 8158
rect 169316 8094 169318 8146
rect 169370 8094 169372 8146
rect 168868 6234 168924 6244
rect 169316 6076 169372 8094
rect 169428 7642 169484 12404
rect 170660 11898 170716 11910
rect 170660 11846 170662 11898
rect 170714 11846 170716 11898
rect 170212 11564 170268 11574
rect 170100 9772 170156 9782
rect 170100 9042 170156 9716
rect 170100 8990 170102 9042
rect 170154 8990 170156 9042
rect 169428 7590 169430 7642
rect 169482 7590 169484 7642
rect 169428 7578 169484 7590
rect 169540 8316 169596 8326
rect 169540 7084 169596 8260
rect 169540 7018 169596 7028
rect 169316 6010 169372 6020
rect 168756 5854 168758 5906
rect 168810 5854 168812 5906
rect 168756 5842 168812 5854
rect 169204 5964 169260 5974
rect 167860 5450 167916 5460
rect 167636 5114 167692 5124
rect 168644 4954 168700 4966
rect 168644 4902 168646 4954
rect 168698 4902 168700 4954
rect 167972 4732 168028 4742
rect 167748 1932 167804 1942
rect 167972 1932 168028 4676
rect 168644 4060 168700 4902
rect 168644 3994 168700 4004
rect 168868 4956 168924 4966
rect 167804 1876 168028 1932
rect 168420 3724 168476 3734
rect 167748 1866 167804 1876
rect 167412 1530 167468 1540
rect 167748 1484 167804 1494
rect 167748 800 167804 1428
rect 168420 800 168476 3668
rect 168868 3387 168924 4900
rect 168980 4954 169036 4966
rect 168980 4902 168982 4954
rect 169034 4902 169036 4954
rect 168980 4396 169036 4902
rect 168980 4330 169036 4340
rect 169204 4060 169260 5908
rect 169652 5794 169708 5806
rect 169652 5742 169654 5794
rect 169706 5742 169708 5794
rect 169484 5628 169540 5638
rect 169484 5404 169540 5572
rect 169484 4954 169540 5348
rect 169484 4902 169486 4954
rect 169538 4902 169540 4954
rect 169484 4890 169540 4902
rect 169204 3994 169260 4004
rect 168868 3331 169036 3387
rect 168980 800 169036 3331
rect 169652 800 169708 5742
rect 170100 5404 170156 8990
rect 170212 6802 170268 11508
rect 170324 9602 170380 9614
rect 170324 9550 170326 9602
rect 170378 9550 170380 9602
rect 170324 8428 170380 9550
rect 170324 8362 170380 8372
rect 170660 7474 170716 11846
rect 170772 11788 170828 14200
rect 171108 13132 171164 13142
rect 170996 12122 171052 12134
rect 170996 12070 170998 12122
rect 171050 12070 171052 12122
rect 170884 12012 170940 12022
rect 170996 12012 171052 12070
rect 170940 11956 171052 12012
rect 170884 11946 170940 11956
rect 170772 11722 170828 11732
rect 170996 9324 171052 11956
rect 171108 11676 171164 13076
rect 171108 11610 171164 11620
rect 171220 12348 171276 12358
rect 171220 9826 171276 12292
rect 171220 9774 171222 9826
rect 171274 9774 171276 9826
rect 171220 9762 171276 9774
rect 170996 9268 171164 9324
rect 170828 9100 170884 9110
rect 170828 9006 170884 9044
rect 170940 9100 171052 9110
rect 170940 9098 170996 9100
rect 170940 9046 170942 9098
rect 170994 9046 170996 9098
rect 170940 9044 170996 9046
rect 170940 9034 171052 9044
rect 170772 8316 170828 8326
rect 170772 8258 170828 8260
rect 170772 8206 170774 8258
rect 170826 8206 170828 8258
rect 170772 8194 170828 8206
rect 170660 7422 170662 7474
rect 170714 7422 170716 7474
rect 170660 7410 170716 7422
rect 170212 6750 170214 6802
rect 170266 6750 170268 6802
rect 170212 6738 170268 6750
rect 171108 5964 171164 9268
rect 171332 8426 171388 14308
rect 171528 14200 171640 15000
rect 172200 14200 172312 15000
rect 172676 14924 172732 14934
rect 171556 13356 171612 14200
rect 171556 13290 171612 13300
rect 172228 12348 172284 14200
rect 172228 12282 172284 12292
rect 172564 11900 172620 11910
rect 172452 11788 172508 11798
rect 171668 10556 171724 10566
rect 171668 9714 171724 10500
rect 172452 9994 172508 11732
rect 172452 9942 172454 9994
rect 172506 9942 172508 9994
rect 172452 9930 172508 9942
rect 171668 9662 171670 9714
rect 171722 9662 171724 9714
rect 171668 8540 171724 9662
rect 172564 9210 172620 11844
rect 172564 9158 172566 9210
rect 172618 9158 172620 9210
rect 172564 9146 172620 9158
rect 171668 8474 171724 8484
rect 171332 8374 171334 8426
rect 171386 8374 171388 8426
rect 171332 8362 171388 8374
rect 171668 8090 171724 8102
rect 171668 8038 171670 8090
rect 171722 8038 171724 8090
rect 171220 6690 171276 6702
rect 171220 6638 171222 6690
rect 171274 6638 171276 6690
rect 171220 6524 171276 6638
rect 171220 6458 171276 6468
rect 171108 5898 171164 5908
rect 170100 5338 170156 5348
rect 171668 5404 171724 8038
rect 172564 8090 172620 8102
rect 172564 8038 172566 8090
rect 172618 8038 172620 8090
rect 172228 7980 172284 7990
rect 172228 7474 172284 7924
rect 172228 7422 172230 7474
rect 172282 7422 172284 7474
rect 172228 7410 172284 7422
rect 171668 5338 171724 5348
rect 171892 6300 171948 6310
rect 171892 5122 171948 6244
rect 171892 5070 171894 5122
rect 171946 5070 171948 5122
rect 170436 5010 170492 5022
rect 170436 4958 170438 5010
rect 170490 4958 170492 5010
rect 170436 4284 170492 4958
rect 170436 4218 170492 4228
rect 171892 3834 171948 5070
rect 172564 4732 172620 8038
rect 172676 5738 172732 14868
rect 172984 14200 173096 15000
rect 173656 14200 173768 15000
rect 174132 14252 174188 14262
rect 173012 12012 173068 14200
rect 173684 13242 173740 14200
rect 174440 14200 174552 15000
rect 174692 14812 174748 14822
rect 173684 13190 173686 13242
rect 173738 13190 173740 13242
rect 173684 13178 173740 13190
rect 174020 13580 174076 13590
rect 173460 12796 173516 12806
rect 173460 12348 173516 12740
rect 173460 12282 173516 12292
rect 173012 11946 173068 11956
rect 172788 11116 172844 11126
rect 172788 9770 172844 11060
rect 173292 9996 173348 10006
rect 173292 9882 173348 9940
rect 173292 9830 173294 9882
rect 173346 9830 173348 9882
rect 173292 9818 173348 9830
rect 172788 9718 172790 9770
rect 172842 9718 172844 9770
rect 172788 9706 172844 9718
rect 173348 9100 173404 9110
rect 173348 9042 173404 9044
rect 173348 8990 173350 9042
rect 173402 8990 173404 9042
rect 173348 8978 173404 8990
rect 172676 5686 172678 5738
rect 172730 5686 172732 5738
rect 172676 5674 172732 5686
rect 172900 8090 172956 8102
rect 172900 8038 172902 8090
rect 172954 8038 172956 8090
rect 172564 4666 172620 4676
rect 172676 4954 172732 4966
rect 172676 4902 172678 4954
rect 172730 4902 172732 4954
rect 171892 3782 171894 3834
rect 171946 3782 171948 3834
rect 171892 3770 171948 3782
rect 172004 4508 172060 4518
rect 170212 1596 170268 1606
rect 170212 800 170268 1540
rect 170884 1148 170940 1158
rect 170884 800 170940 1092
rect 171444 924 171500 934
rect 171444 800 171500 868
rect 172004 800 172060 4452
rect 172676 3612 172732 4902
rect 172676 3546 172732 3556
rect 172900 2044 172956 8038
rect 173404 8092 173460 8102
rect 173404 7998 173460 8036
rect 173124 7362 173180 7374
rect 173124 7310 173126 7362
rect 173178 7310 173180 7362
rect 173012 5964 173068 5974
rect 173012 5906 173068 5908
rect 173012 5854 173014 5906
rect 173066 5854 173068 5906
rect 173012 5842 173068 5854
rect 173012 4956 173068 4966
rect 173012 4862 173068 4900
rect 173124 3948 173180 7310
rect 174020 6860 174076 13524
rect 174132 13244 174188 14196
rect 174468 13916 174524 14200
rect 174692 14140 174748 14756
rect 175112 14200 175224 15000
rect 175588 14588 175644 14598
rect 174692 14074 174748 14084
rect 174468 13850 174524 13860
rect 174132 13178 174188 13188
rect 174916 13804 174972 13814
rect 174804 9826 174860 9838
rect 174188 9772 174244 9782
rect 174188 9678 174244 9716
rect 174804 9774 174806 9826
rect 174858 9774 174860 9826
rect 174244 9212 174300 9222
rect 174132 6860 174188 6870
rect 174020 6858 174188 6860
rect 174020 6806 174134 6858
rect 174186 6806 174188 6858
rect 174020 6804 174188 6806
rect 174132 6794 174188 6804
rect 173124 3882 173180 3892
rect 174244 5122 174300 9156
rect 174804 7868 174860 9774
rect 174356 7644 174412 7654
rect 174356 7474 174412 7588
rect 174356 7422 174358 7474
rect 174410 7422 174412 7474
rect 174356 7410 174412 7422
rect 174804 6972 174860 7812
rect 174916 7642 174972 13748
rect 175140 12124 175196 14200
rect 175140 12058 175196 12068
rect 175476 14140 175532 14150
rect 175588 14140 175644 14532
rect 175896 14200 176008 15000
rect 176568 14200 176680 15000
rect 176820 14588 176876 14598
rect 175924 14140 175980 14200
rect 175588 14084 175980 14140
rect 176372 14138 176428 14150
rect 176372 14086 176374 14138
rect 176426 14086 176428 14138
rect 175140 9714 175196 9726
rect 175140 9662 175142 9714
rect 175194 9662 175196 9714
rect 175028 9038 175084 9050
rect 175028 8986 175030 9038
rect 175082 8986 175084 9038
rect 175028 8316 175084 8986
rect 175028 8250 175084 8260
rect 175028 8092 175084 8102
rect 175028 7998 175084 8036
rect 174916 7590 174918 7642
rect 174970 7590 174972 7642
rect 174916 7578 174972 7590
rect 174804 6906 174860 6916
rect 174468 6690 174524 6702
rect 174468 6638 174470 6690
rect 174522 6638 174524 6690
rect 174468 6412 174524 6638
rect 175140 6636 175196 9662
rect 175476 9210 175532 14084
rect 175476 9158 175478 9210
rect 175530 9158 175532 9210
rect 175476 9146 175532 9158
rect 175924 12234 175980 12246
rect 175924 12182 175926 12234
rect 175978 12182 175980 12234
rect 175924 11228 175980 12182
rect 175812 9098 175868 9110
rect 175812 9046 175814 9098
rect 175866 9046 175868 9098
rect 175812 7756 175868 9046
rect 175924 8258 175980 11172
rect 176372 9212 176428 14086
rect 176596 14140 176652 14200
rect 176820 14140 176876 14532
rect 177352 14200 177464 15000
rect 178024 14200 178136 15000
rect 178808 14200 178920 15000
rect 179480 14200 179592 15000
rect 180264 14200 180376 15000
rect 180936 14200 181048 15000
rect 181720 14200 181832 15000
rect 181972 14924 182028 14934
rect 181972 14588 182028 14868
rect 181972 14532 182252 14588
rect 176596 14084 176876 14140
rect 177156 13356 177212 13366
rect 176932 12012 176988 12022
rect 176932 9994 176988 11956
rect 176932 9942 176934 9994
rect 176986 9942 176988 9994
rect 176932 9930 176988 9942
rect 176596 9212 176652 9222
rect 176372 9210 176652 9212
rect 176372 9158 176598 9210
rect 176650 9158 176652 9210
rect 176372 9156 176652 9158
rect 176596 9146 176652 9156
rect 176932 9100 176988 9110
rect 176932 9098 177100 9100
rect 176932 9046 176934 9098
rect 176986 9046 177100 9098
rect 176932 9044 177100 9046
rect 176932 9034 176988 9044
rect 175924 8206 175926 8258
rect 175978 8206 175980 8258
rect 175924 8194 175980 8206
rect 175812 7700 175980 7756
rect 175140 6570 175196 6580
rect 175252 7530 175308 7542
rect 175252 7478 175254 7530
rect 175306 7478 175308 7530
rect 174468 6346 174524 6356
rect 175140 6076 175196 6086
rect 175140 5982 175196 6020
rect 174580 5964 174636 5974
rect 174580 5865 174582 5908
rect 174634 5865 174636 5908
rect 174580 5853 174636 5865
rect 174244 5070 174246 5122
rect 174298 5070 174300 5122
rect 174244 3946 174300 5070
rect 174356 5010 174412 5022
rect 174356 4958 174358 5010
rect 174410 4958 174412 5010
rect 174356 4620 174412 4958
rect 174356 4554 174412 4564
rect 174244 3894 174246 3946
rect 174298 3894 174300 3946
rect 174244 3882 174300 3894
rect 175028 4172 175084 4182
rect 172900 1978 172956 1988
rect 173236 3724 173292 3734
rect 172676 1372 172732 1382
rect 172676 800 172732 1316
rect 173236 800 173292 3668
rect 174356 2716 174412 2726
rect 174356 2602 174412 2660
rect 174356 2550 174358 2602
rect 174410 2550 174412 2602
rect 174356 2538 174412 2550
rect 175028 2602 175084 4116
rect 175252 3948 175308 7478
rect 175756 7532 175812 7542
rect 175756 7438 175812 7476
rect 175476 6076 175532 6086
rect 175476 5982 175532 6020
rect 175924 5180 175980 7700
rect 175924 5114 175980 5124
rect 176148 6690 176204 6702
rect 176148 6638 176150 6690
rect 176202 6638 176204 6690
rect 175252 3882 175308 3892
rect 175924 4060 175980 4070
rect 175924 3164 175980 4004
rect 176148 3612 176204 6638
rect 176484 5516 176540 5526
rect 176372 4954 176428 4966
rect 176372 4902 176374 4954
rect 176426 4902 176428 4954
rect 176372 4394 176428 4902
rect 176372 4342 176374 4394
rect 176426 4342 176428 4394
rect 176372 4330 176428 4342
rect 176484 3836 176540 5460
rect 176708 4954 176764 4966
rect 176708 4902 176710 4954
rect 176762 4902 176764 4954
rect 176708 4172 176764 4902
rect 176708 4106 176764 4116
rect 176932 4396 176988 4406
rect 177044 4396 177100 9044
rect 177156 6802 177212 13300
rect 177268 12796 177324 12806
rect 177268 11564 177324 12740
rect 177380 11788 177436 14200
rect 178052 14028 178108 14200
rect 178052 13962 178108 13972
rect 178276 13802 178332 13814
rect 178276 13750 178278 13802
rect 178330 13750 178332 13802
rect 177380 11722 177436 11732
rect 177492 12796 177548 12806
rect 177268 11508 177436 11564
rect 177268 10220 177324 10230
rect 177268 9770 177324 10164
rect 177268 9718 177270 9770
rect 177322 9718 177324 9770
rect 177268 9706 177324 9718
rect 177156 6750 177158 6802
rect 177210 6750 177212 6802
rect 177156 6738 177212 6750
rect 177212 5180 177268 5190
rect 177380 5180 177436 11508
rect 177492 6074 177548 12740
rect 178052 12236 178108 12246
rect 178052 12012 178108 12180
rect 178052 11946 178108 11956
rect 178052 10668 178108 10678
rect 178052 8764 178108 10612
rect 178276 10668 178332 13750
rect 178836 12236 178892 14200
rect 178836 12170 178892 12180
rect 179172 14028 179228 14038
rect 178276 10602 178332 10612
rect 178612 12012 178668 12022
rect 178276 9714 178332 9726
rect 178276 9662 178278 9714
rect 178330 9662 178332 9714
rect 178164 9602 178220 9614
rect 178164 9550 178166 9602
rect 178218 9550 178220 9602
rect 178164 9548 178220 9550
rect 178164 9482 178220 9492
rect 178276 9212 178332 9662
rect 178276 9146 178332 9156
rect 178052 8698 178108 8708
rect 178500 8764 178556 8774
rect 177604 8258 177660 8270
rect 177604 8206 177606 8258
rect 177658 8206 177660 8258
rect 177604 8204 177660 8206
rect 177604 8138 177660 8148
rect 177716 7756 177772 7766
rect 177716 7642 177772 7700
rect 177716 7590 177718 7642
rect 177770 7590 177772 7642
rect 177716 7578 177772 7590
rect 178500 7474 178556 8708
rect 178500 7422 178502 7474
rect 178554 7422 178556 7474
rect 178500 7410 178556 7422
rect 177940 6690 177996 6702
rect 177940 6638 177942 6690
rect 177994 6638 177996 6690
rect 177940 6300 177996 6638
rect 177940 6234 177996 6244
rect 177492 6022 177494 6074
rect 177546 6022 177548 6074
rect 177492 6010 177548 6022
rect 177604 6188 177660 6198
rect 177212 5178 177436 5180
rect 177212 5126 177214 5178
rect 177266 5126 177436 5178
rect 177212 5124 177436 5126
rect 177492 5404 177548 5414
rect 177604 5404 177660 6132
rect 178612 5906 178668 11956
rect 179060 9996 179116 10006
rect 179060 8426 179116 9940
rect 179060 8374 179062 8426
rect 179114 8374 179116 8426
rect 179060 8362 179116 8374
rect 179172 8258 179228 13972
rect 179284 13356 179340 13366
rect 179284 8874 179340 13300
rect 179508 13244 179564 14200
rect 179508 13178 179564 13188
rect 180292 12684 180348 14200
rect 180964 13020 181020 14200
rect 181748 13916 181804 14200
rect 182196 14140 182252 14532
rect 182392 14200 182504 15000
rect 183176 14200 183288 15000
rect 183848 14200 183960 15000
rect 184632 14200 184744 15000
rect 185304 14200 185416 15000
rect 186088 14200 186200 15000
rect 186760 14200 186872 15000
rect 187544 14200 187656 15000
rect 188216 14200 188328 15000
rect 188692 14252 188748 14262
rect 182420 14140 182476 14200
rect 182196 14084 182476 14140
rect 182980 14140 183036 14150
rect 181748 13850 181804 13860
rect 180964 12954 181020 12964
rect 182308 13692 182364 13702
rect 180292 12618 180348 12628
rect 179620 12236 179676 12246
rect 179396 10668 179452 10678
rect 179396 9660 179452 10612
rect 179620 9826 179676 12180
rect 181300 12236 181356 12246
rect 180068 12124 180124 12134
rect 180068 9994 180124 12068
rect 180068 9942 180070 9994
rect 180122 9942 180124 9994
rect 180068 9930 180124 9942
rect 180404 11564 180460 11574
rect 179620 9774 179622 9826
rect 179674 9774 179676 9826
rect 179620 9762 179676 9774
rect 180404 9770 180460 11508
rect 181076 10666 181132 10678
rect 181076 10614 181078 10666
rect 181130 10614 181132 10666
rect 181076 10342 181132 10614
rect 181076 10332 181188 10342
rect 181076 10276 181132 10332
rect 180404 9718 180406 9770
rect 180458 9718 180460 9770
rect 181132 9826 181188 10276
rect 181132 9774 181134 9826
rect 181186 9774 181188 9826
rect 181132 9762 181188 9774
rect 180404 9706 180460 9718
rect 181020 9660 181076 9670
rect 181300 9660 181356 12180
rect 179396 9604 179676 9660
rect 179620 9042 179676 9604
rect 181020 9566 181076 9604
rect 181188 9604 181356 9660
rect 182084 9772 182140 9782
rect 182084 9714 182140 9716
rect 182084 9662 182086 9714
rect 182138 9662 182140 9714
rect 182084 9650 182140 9662
rect 179620 8990 179622 9042
rect 179674 8990 179676 9042
rect 179620 8978 179676 8990
rect 180852 9212 180908 9222
rect 179284 8822 179286 8874
rect 179338 8822 179340 8874
rect 179284 8810 179340 8822
rect 179172 8206 179174 8258
rect 179226 8206 179228 8258
rect 179172 8194 179228 8206
rect 180404 8428 180460 8438
rect 179396 8146 179452 8158
rect 179396 8094 179398 8146
rect 179450 8094 179452 8146
rect 178836 6636 178892 6646
rect 178836 6542 178892 6580
rect 179172 6522 179228 6534
rect 179172 6470 179174 6522
rect 179226 6470 179228 6522
rect 179172 6412 179228 6470
rect 179172 6346 179228 6356
rect 178612 5854 178614 5906
rect 178666 5854 178668 5906
rect 178612 5842 178668 5854
rect 177548 5348 177660 5404
rect 178164 5404 178220 5414
rect 177212 5114 177268 5124
rect 177156 4396 177212 4406
rect 177044 4340 177156 4396
rect 176148 3546 176204 3556
rect 176372 3780 176540 3836
rect 175028 2550 175030 2602
rect 175082 2550 175084 2602
rect 175028 2538 175084 2550
rect 175700 3108 175924 3164
rect 175140 1596 175196 1606
rect 174468 1036 174524 1046
rect 173908 924 173964 934
rect 173908 800 173964 868
rect 174468 800 174524 980
rect 175140 800 175196 1540
rect 175700 800 175756 3108
rect 175924 3098 175980 3108
rect 176372 800 176428 3780
rect 176932 800 176988 4340
rect 177156 4330 177212 4340
rect 177492 800 177548 5348
rect 178164 5122 178220 5348
rect 178164 5070 178166 5122
rect 178218 5070 178220 5122
rect 178164 5058 178220 5070
rect 178276 5010 178332 5022
rect 178276 4958 178278 5010
rect 178330 4958 178332 5010
rect 178276 4284 178332 4958
rect 178276 4218 178332 4228
rect 178724 4620 178780 4630
rect 178724 3948 178780 4564
rect 178052 3276 178108 3286
rect 177716 2156 177772 2166
rect 178052 2156 178108 3220
rect 178388 2828 178444 2838
rect 178388 2492 178444 2772
rect 178388 2426 178444 2436
rect 177772 2100 178108 2156
rect 178164 2268 178220 2278
rect 177716 2090 177772 2100
rect 178164 2044 178220 2212
rect 178164 800 178220 1988
rect 178724 800 178780 3892
rect 178836 3500 178892 3510
rect 178836 2044 178892 3444
rect 178948 3388 179004 3398
rect 178948 3274 179004 3332
rect 178948 3222 178950 3274
rect 179002 3222 179004 3274
rect 178948 3210 179004 3222
rect 179396 3276 179452 8094
rect 180180 7470 180236 7482
rect 180180 7418 180182 7470
rect 180234 7418 180236 7470
rect 180180 7308 180236 7418
rect 180180 7242 180236 7252
rect 180404 6758 180460 8372
rect 180852 7598 180908 9156
rect 181188 8258 181244 9604
rect 181860 9436 181916 9446
rect 181860 9266 181916 9380
rect 181860 9214 181862 9266
rect 181914 9214 181916 9266
rect 181860 9202 181916 9214
rect 181300 9038 181356 9050
rect 181300 8986 181302 9038
rect 181354 8986 181356 9038
rect 181300 8428 181356 8986
rect 181300 8362 181356 8372
rect 181524 8876 181580 8886
rect 181524 8426 181580 8820
rect 181524 8374 181526 8426
rect 181578 8374 181580 8426
rect 181524 8362 181580 8374
rect 181188 8206 181190 8258
rect 181242 8206 181244 8258
rect 181188 8194 181244 8206
rect 180796 7586 180908 7598
rect 180796 7534 180798 7586
rect 180850 7534 180908 7586
rect 180796 7532 180908 7534
rect 180964 8146 181020 8158
rect 180964 8094 180966 8146
rect 181018 8094 181020 8146
rect 180796 7522 180852 7532
rect 180684 7306 180740 7318
rect 180684 7254 180686 7306
rect 180738 7254 180740 7306
rect 180684 7196 180740 7254
rect 180684 7130 180740 7140
rect 180404 6746 180516 6758
rect 180404 6694 180462 6746
rect 180514 6694 180516 6746
rect 180404 6692 180516 6694
rect 180460 6682 180516 6692
rect 179676 6636 179732 6646
rect 179676 6542 179732 6580
rect 179620 6076 179676 6086
rect 179620 3388 179676 6020
rect 180180 6076 180236 6086
rect 180180 5906 180236 6020
rect 180180 5854 180182 5906
rect 180234 5854 180236 5906
rect 180180 5842 180236 5854
rect 180068 4956 180124 4966
rect 179620 3387 179788 3388
rect 179620 3332 180012 3387
rect 179732 3331 180012 3332
rect 179396 3210 179452 3220
rect 179956 3276 180012 3331
rect 178836 1978 178892 1988
rect 179060 2492 179116 2502
rect 179060 2042 179116 2436
rect 179060 1990 179062 2042
rect 179114 1990 179116 2042
rect 179060 1978 179116 1990
rect 179396 1596 179452 1606
rect 179396 800 179452 1540
rect 179956 800 180012 3220
rect 180068 3164 180124 4900
rect 180292 4954 180348 4966
rect 180292 4902 180294 4954
rect 180346 4902 180348 4954
rect 180292 4506 180348 4902
rect 180292 4454 180294 4506
rect 180346 4454 180348 4506
rect 180292 4442 180348 4454
rect 180628 4954 180684 4966
rect 180628 4902 180630 4954
rect 180682 4902 180684 4954
rect 180628 4396 180684 4902
rect 180628 4330 180684 4340
rect 180068 3098 180124 3108
rect 180292 3164 180348 3174
rect 180292 2492 180348 3108
rect 180964 3164 181020 8094
rect 181636 7362 181692 7374
rect 181636 7310 181638 7362
rect 181690 7310 181692 7362
rect 181188 6860 181244 6870
rect 181188 5906 181244 6804
rect 181188 5854 181190 5906
rect 181242 5854 181244 5906
rect 181188 5516 181244 5854
rect 181300 6748 181356 6758
rect 181300 5852 181356 6692
rect 181300 5786 181356 5796
rect 181412 5794 181468 5806
rect 181412 5742 181414 5794
rect 181466 5742 181468 5794
rect 181188 5460 181356 5516
rect 181132 4954 181188 4966
rect 181132 4902 181134 4954
rect 181186 4902 181188 4954
rect 181132 4844 181188 4902
rect 181132 4778 181188 4788
rect 181300 3612 181356 5460
rect 181300 3546 181356 3556
rect 180964 3098 181020 3108
rect 180292 2426 180348 2436
rect 181188 1596 181244 1606
rect 180628 1484 180684 1494
rect 180628 800 180684 1428
rect 181188 800 181244 1540
rect 181412 1260 181468 5742
rect 181636 5180 181692 7310
rect 182308 6188 182364 13636
rect 182868 13692 182924 13702
rect 182532 13578 182588 13590
rect 182532 13526 182534 13578
rect 182586 13526 182588 13578
rect 182532 12908 182588 13526
rect 182420 12852 182532 12908
rect 182420 7868 182476 12852
rect 182532 12842 182588 12852
rect 182532 9994 182588 10006
rect 182532 9942 182534 9994
rect 182586 9942 182588 9994
rect 182532 9100 182588 9942
rect 182756 9884 182812 9894
rect 182756 9826 182812 9828
rect 182756 9774 182758 9826
rect 182810 9774 182812 9826
rect 182756 9762 182812 9774
rect 182532 9034 182588 9044
rect 182756 9436 182812 9446
rect 182756 9154 182812 9380
rect 182756 9102 182758 9154
rect 182810 9102 182812 9154
rect 182756 8540 182812 9102
rect 182756 8474 182812 8484
rect 182868 8258 182924 13636
rect 182980 9042 183036 14084
rect 183204 13804 183260 14200
rect 183204 13738 183260 13748
rect 183876 12124 183932 14200
rect 184660 13580 184716 14200
rect 184660 13514 184716 13524
rect 183876 12058 183932 12068
rect 184548 13466 184604 13478
rect 184548 13414 184550 13466
rect 184602 13414 184604 13466
rect 183988 11788 184044 11798
rect 183876 11340 183932 11350
rect 183876 10780 183932 11284
rect 182980 8990 182982 9042
rect 183034 8990 183036 9042
rect 183652 10108 183708 10118
rect 183652 8998 183708 10052
rect 182980 8978 183036 8990
rect 183428 8988 183484 8998
rect 182868 8206 182870 8258
rect 182922 8206 182924 8258
rect 182868 8194 182924 8206
rect 183652 8988 183764 8998
rect 183652 8932 183708 8988
rect 182980 8146 183036 8158
rect 182980 8094 182982 8146
rect 183034 8094 183036 8146
rect 182420 7812 182812 7868
rect 182532 7644 182588 7654
rect 182308 6122 182364 6132
rect 182420 6412 182476 6422
rect 181636 5114 181692 5124
rect 182196 5010 182252 5022
rect 182196 4958 182198 5010
rect 182250 4958 182252 5010
rect 182196 4844 182252 4958
rect 182196 4778 182252 4788
rect 181412 1194 181468 1204
rect 181860 4172 181916 4182
rect 181860 800 181916 4116
rect 182420 800 182476 6356
rect 182532 5124 182588 7588
rect 182756 6972 182812 7812
rect 182980 7756 183036 8094
rect 182980 7690 183036 7700
rect 182980 7474 183036 7486
rect 182980 7422 182982 7474
rect 183034 7422 183036 7474
rect 182980 7420 183036 7422
rect 182980 7196 183036 7364
rect 182980 7130 183036 7140
rect 182756 6916 183036 6972
rect 182644 6860 182700 6870
rect 182644 6766 182700 6804
rect 182980 6690 183036 6916
rect 182980 6638 182982 6690
rect 183034 6638 183036 6690
rect 182980 6626 183036 6638
rect 182868 6188 182924 6198
rect 182868 6074 182924 6132
rect 183428 6188 183484 8932
rect 183708 8894 183764 8932
rect 183540 8652 183596 8662
rect 183540 8426 183596 8596
rect 183540 8374 183542 8426
rect 183594 8374 183596 8426
rect 183540 8362 183596 8374
rect 183652 8316 183708 8326
rect 183652 7654 183708 8260
rect 183652 7642 183764 7654
rect 183652 7590 183710 7642
rect 183762 7590 183764 7642
rect 183876 7598 183932 10724
rect 183988 9994 184044 11732
rect 183988 9942 183990 9994
rect 184042 9942 184044 9994
rect 183988 9930 184044 9942
rect 184548 10892 184604 13414
rect 185332 13020 185388 14200
rect 185332 12954 185388 12964
rect 185668 13580 185724 13590
rect 184324 9658 184380 9670
rect 184324 9606 184326 9658
rect 184378 9606 184380 9658
rect 184324 9212 184380 9606
rect 184324 9146 184380 9156
rect 184548 9042 184604 10836
rect 184548 8990 184550 9042
rect 184602 8990 184604 9042
rect 184548 8978 184604 8990
rect 184772 9996 184828 10006
rect 184772 7698 184828 9940
rect 185052 9884 185108 9894
rect 185052 9826 185108 9828
rect 185052 9774 185054 9826
rect 185106 9774 185108 9826
rect 185052 9762 185108 9774
rect 184940 9658 184996 9670
rect 184940 9606 184942 9658
rect 184994 9606 184996 9658
rect 184940 9044 184996 9606
rect 185108 9660 185164 9670
rect 185108 9154 185164 9604
rect 185108 9102 185110 9154
rect 185162 9102 185164 9154
rect 185108 9090 185164 9102
rect 185556 9324 185612 9334
rect 184940 8988 185052 9044
rect 184996 7868 185052 8988
rect 185556 8426 185612 9268
rect 185556 8374 185558 8426
rect 185610 8374 185612 8426
rect 185556 8362 185612 8374
rect 184996 7802 185052 7812
rect 185108 8316 185164 8326
rect 184772 7646 184774 7698
rect 184826 7646 184828 7698
rect 184772 7634 184828 7646
rect 183652 7588 183764 7590
rect 183708 7578 183764 7588
rect 183820 7586 183932 7598
rect 183820 7534 183822 7586
rect 183874 7534 183932 7586
rect 183820 7532 183932 7534
rect 183820 7522 183876 7532
rect 184660 7474 184716 7486
rect 184660 7422 184662 7474
rect 184714 7422 184716 7474
rect 184492 6690 184548 6702
rect 184492 6638 184494 6690
rect 184546 6638 184548 6690
rect 184492 6636 184548 6638
rect 183428 6122 183484 6132
rect 184324 6580 184548 6636
rect 182868 6022 182870 6074
rect 182922 6022 182924 6074
rect 182868 6010 182924 6022
rect 183204 5962 183260 5974
rect 183204 5910 183206 5962
rect 183258 5910 183260 5962
rect 183204 5852 183260 5910
rect 183204 5786 183260 5796
rect 183540 5852 183596 5862
rect 182644 5124 182700 5134
rect 182532 5122 182700 5124
rect 182532 5070 182646 5122
rect 182698 5070 182700 5122
rect 182532 5068 182700 5070
rect 182644 3500 182700 5068
rect 182644 3434 182700 3444
rect 182980 4396 183036 4406
rect 182980 800 183036 4340
rect 183540 3387 183596 5796
rect 183708 5850 183764 5862
rect 183708 5798 183710 5850
rect 183762 5798 183764 5850
rect 183708 5292 183764 5798
rect 184324 5404 184380 6580
rect 184660 6076 184716 7422
rect 185108 6802 185164 8260
rect 185108 6750 185110 6802
rect 185162 6750 185164 6802
rect 185108 6738 185164 6750
rect 185220 6860 185276 6870
rect 184324 5338 184380 5348
rect 184436 6020 184716 6076
rect 184772 6188 184828 6198
rect 183708 5226 183764 5236
rect 184212 4954 184268 4966
rect 184212 4902 184214 4954
rect 184266 4902 184268 4954
rect 184212 4282 184268 4902
rect 184212 4230 184214 4282
rect 184266 4230 184268 4282
rect 184212 4218 184268 4230
rect 183540 3331 183708 3387
rect 183092 2492 183148 2502
rect 183092 2378 183148 2436
rect 183092 2326 183094 2378
rect 183146 2326 183148 2378
rect 183092 2314 183148 2326
rect 183652 800 183708 3331
rect 184212 3164 184268 3174
rect 184212 800 184268 3108
rect 184436 3052 184492 6020
rect 184772 5964 184828 6132
rect 184660 5908 184828 5964
rect 184660 5906 184716 5908
rect 184660 5854 184662 5906
rect 184714 5854 184716 5906
rect 184660 5842 184716 5854
rect 184772 5794 184828 5806
rect 184772 5742 184774 5794
rect 184826 5742 184828 5794
rect 184772 5628 184828 5742
rect 184772 5562 184828 5572
rect 185220 5068 185276 6804
rect 185668 6690 185724 13524
rect 185780 13132 185836 13142
rect 185780 7474 185836 13076
rect 185892 13130 185948 13142
rect 185892 13078 185894 13130
rect 185946 13078 185948 13130
rect 185892 10780 185948 13078
rect 186116 11788 186172 14200
rect 186116 11722 186172 11732
rect 186228 13692 186284 13702
rect 185892 9826 185948 10724
rect 185892 9774 185894 9826
rect 185946 9774 185948 9826
rect 185892 9762 185948 9774
rect 186004 9714 186060 9726
rect 186004 9662 186006 9714
rect 186058 9662 186060 9714
rect 186004 9660 186060 9662
rect 186004 9594 186060 9604
rect 186116 8930 186172 8942
rect 186116 8878 186118 8930
rect 186170 8878 186172 8930
rect 186116 8876 186172 8878
rect 186116 8810 186172 8820
rect 186228 8652 186284 13636
rect 186564 13018 186620 13030
rect 186564 12966 186566 13018
rect 186618 12966 186620 13018
rect 186452 11900 186508 11910
rect 186116 8596 186284 8652
rect 186340 11228 186396 11238
rect 186116 8258 186172 8596
rect 186116 8206 186118 8258
rect 186170 8206 186172 8258
rect 186116 8194 186172 8206
rect 185780 7422 185782 7474
rect 185834 7422 185836 7474
rect 185780 7410 185836 7422
rect 185892 8146 185948 8158
rect 186340 8148 186396 11172
rect 186452 8428 186508 11844
rect 186564 10666 186620 12966
rect 186788 12796 186844 14200
rect 186788 12730 186844 12740
rect 187572 14028 187628 14200
rect 186564 10614 186566 10666
rect 186618 10614 186620 10666
rect 186564 9042 186620 10614
rect 187124 12684 187180 12694
rect 186676 9660 186732 9670
rect 186676 9212 186732 9604
rect 186676 9154 186732 9156
rect 186676 9102 186678 9154
rect 186730 9102 186732 9154
rect 186676 9080 186732 9102
rect 186564 8990 186566 9042
rect 186618 8990 186620 9042
rect 186564 8978 186620 8990
rect 186564 8428 186620 8438
rect 186452 8426 186620 8428
rect 186452 8374 186566 8426
rect 186618 8374 186620 8426
rect 186452 8372 186620 8374
rect 186564 8362 186620 8372
rect 185892 8094 185894 8146
rect 185946 8094 185948 8146
rect 185668 6638 185670 6690
rect 185722 6638 185724 6690
rect 185668 6626 185724 6638
rect 185220 4966 185276 5012
rect 184436 2986 184492 2996
rect 184548 4954 184604 4966
rect 184548 4902 184550 4954
rect 184602 4902 184604 4954
rect 184548 2492 184604 4902
rect 185164 4954 185276 4966
rect 185164 4902 185166 4954
rect 185218 4902 185276 4954
rect 185164 4900 185276 4902
rect 185164 4890 185220 4900
rect 185332 4844 185388 4854
rect 185332 4732 185388 4788
rect 185780 4732 185836 4742
rect 185332 4676 185780 4732
rect 185780 4666 185836 4676
rect 185892 2940 185948 8094
rect 186228 8092 186396 8148
rect 186900 8092 186956 8102
rect 186228 5122 186284 8092
rect 186900 8090 187068 8092
rect 186900 8038 186902 8090
rect 186954 8038 187068 8090
rect 186900 8036 187068 8038
rect 186900 8026 186956 8036
rect 186676 7474 186732 7486
rect 186676 7422 186678 7474
rect 186730 7422 186732 7474
rect 186564 7362 186620 7374
rect 186564 7310 186566 7362
rect 186618 7310 186620 7362
rect 186564 7084 186620 7310
rect 186564 7018 186620 7028
rect 186228 5070 186230 5122
rect 186282 5070 186284 5122
rect 186228 5058 186284 5070
rect 186340 6578 186396 6590
rect 186340 6526 186342 6578
rect 186394 6526 186396 6578
rect 186116 5010 186172 5022
rect 186116 4958 186118 5010
rect 186170 4958 186172 5010
rect 186116 4956 186172 4958
rect 186004 4900 186172 4956
rect 186004 4284 186060 4900
rect 186340 4844 186396 6526
rect 186676 5404 186732 7422
rect 187012 6972 187068 8036
rect 186900 6748 186956 6758
rect 186788 5794 186844 5806
rect 186788 5742 186790 5794
rect 186842 5742 186844 5794
rect 186788 5740 186844 5742
rect 186788 5674 186844 5684
rect 186004 4218 186060 4228
rect 186116 4788 186396 4844
rect 186452 5348 186732 5404
rect 184548 2426 184604 2436
rect 185444 2492 185500 2502
rect 184884 2156 184940 2166
rect 184884 800 184940 2100
rect 185444 800 185500 2436
rect 185892 2378 185948 2884
rect 186116 2940 186172 4788
rect 186116 2846 186172 2884
rect 186340 4284 186396 4294
rect 186004 2828 186060 2838
rect 186004 2734 186060 2772
rect 186228 2828 186284 2838
rect 186228 2492 186284 2772
rect 186340 2604 186396 4228
rect 186340 2538 186396 2548
rect 186452 2826 186508 5348
rect 186900 5290 186956 6692
rect 186900 5238 186902 5290
rect 186954 5238 186956 5290
rect 186900 5226 186956 5238
rect 187012 5124 187068 6916
rect 187124 6858 187180 12628
rect 187572 12348 187628 13972
rect 187572 12282 187628 12292
rect 187908 12124 187964 12134
rect 187684 11676 187740 11686
rect 187684 11116 187740 11620
rect 187684 11050 187740 11060
rect 187796 10778 187852 10790
rect 187796 10726 187798 10778
rect 187850 10726 187852 10778
rect 187796 9660 187852 10726
rect 187908 9994 187964 12068
rect 187908 9942 187910 9994
rect 187962 9942 187964 9994
rect 187908 9930 187964 9942
rect 188020 11676 188076 11686
rect 187348 9602 187404 9614
rect 187348 9550 187350 9602
rect 187402 9550 187404 9602
rect 187796 9594 187852 9604
rect 187348 7868 187404 9550
rect 187908 8930 187964 8942
rect 187908 8878 187910 8930
rect 187962 8878 187964 8930
rect 187628 8316 187684 8326
rect 187628 8258 187684 8260
rect 187516 8204 187572 8214
rect 187628 8206 187630 8258
rect 187682 8206 187684 8258
rect 187628 8194 187684 8206
rect 187516 8110 187572 8148
rect 187348 7802 187404 7812
rect 187124 6806 187126 6858
rect 187178 6806 187180 6858
rect 187124 6794 187180 6806
rect 187460 6522 187516 6534
rect 187460 6470 187462 6522
rect 187514 6470 187516 6522
rect 186900 5068 187068 5124
rect 187348 6018 187404 6030
rect 187348 5966 187350 6018
rect 187402 5966 187404 6018
rect 186452 2774 186454 2826
rect 186506 2774 186508 2826
rect 186228 2426 186284 2436
rect 186452 2492 186508 2774
rect 186564 3836 186620 3846
rect 186564 2714 186620 3780
rect 186900 3276 186956 5068
rect 186900 3210 186956 3220
rect 187012 4170 187068 4182
rect 187012 4118 187014 4170
rect 187066 4118 187068 4170
rect 186564 2662 186566 2714
rect 186618 2662 186620 2714
rect 186564 2650 186620 2662
rect 187012 2604 187068 4118
rect 187348 3276 187404 5966
rect 187348 3210 187404 3220
rect 187460 4060 187516 6470
rect 187908 5292 187964 8878
rect 188020 7474 188076 11620
rect 188244 9828 188300 14200
rect 189000 14200 189112 15000
rect 189672 14200 189784 15000
rect 190456 14200 190568 15000
rect 191128 14200 191240 15000
rect 191912 14200 192024 15000
rect 192584 14200 192696 15000
rect 193368 14200 193480 15000
rect 194040 14200 194152 15000
rect 194824 14200 194936 15000
rect 195496 14200 195608 15000
rect 196280 14200 196392 15000
rect 196952 14200 197064 15000
rect 197736 14200 197848 15000
rect 198408 14200 198520 15000
rect 199192 14200 199304 15000
rect 199864 14200 199976 15000
rect 200648 14200 200760 15000
rect 201320 14200 201432 15000
rect 202104 14200 202216 15000
rect 202776 14200 202888 15000
rect 203560 14200 203672 15000
rect 204232 14200 204344 15000
rect 205016 14200 205128 15000
rect 205688 14200 205800 15000
rect 206472 14200 206584 15000
rect 207144 14200 207256 15000
rect 207928 14200 208040 15000
rect 208600 14200 208712 15000
rect 209384 14200 209496 15000
rect 210056 14200 210168 15000
rect 210840 14200 210952 15000
rect 211512 14200 211624 15000
rect 212296 14200 212408 15000
rect 212968 14200 213080 15000
rect 213752 14200 213864 15000
rect 214424 14200 214536 15000
rect 215208 14200 215320 15000
rect 215880 14200 215992 15000
rect 216664 14200 216776 15000
rect 217336 14200 217448 15000
rect 218120 14200 218232 15000
rect 218792 14200 218904 15000
rect 219576 14200 219688 15000
rect 188468 12906 188524 12918
rect 188468 12854 188470 12906
rect 188522 12854 188524 12906
rect 188244 9772 188412 9828
rect 188244 9660 188300 9670
rect 188244 9566 188300 9604
rect 188020 7422 188022 7474
rect 188074 7422 188076 7474
rect 188020 7410 188076 7422
rect 188020 5906 188076 5918
rect 188020 5854 188022 5906
rect 188074 5854 188076 5906
rect 188020 5628 188076 5854
rect 188020 5562 188076 5572
rect 187908 5226 187964 5236
rect 187012 2538 187068 2548
rect 187348 2716 187404 2726
rect 186452 2426 186508 2436
rect 185892 2326 185894 2378
rect 185946 2326 185948 2378
rect 185892 2314 185948 2326
rect 186676 2380 186732 2390
rect 186116 1596 186172 1606
rect 186116 800 186172 1540
rect 186676 800 186732 2324
rect 187348 800 187404 2660
rect 187460 2156 187516 4004
rect 188020 4954 188076 4966
rect 188020 4902 188022 4954
rect 188074 4902 188076 4954
rect 188020 3948 188076 4902
rect 188356 4954 188412 9772
rect 188468 8258 188524 12854
rect 188580 12794 188636 12806
rect 188580 12742 188582 12794
rect 188634 12742 188636 12794
rect 188580 10892 188636 12742
rect 188580 9042 188636 10836
rect 188692 9894 188748 14196
rect 189028 13356 189084 14200
rect 189028 13290 189084 13300
rect 189700 11900 189756 14200
rect 189700 11834 189756 11844
rect 189812 12682 189868 12694
rect 189812 12630 189814 12682
rect 189866 12630 189868 12682
rect 189812 11004 189868 12630
rect 190372 11788 190428 11798
rect 189700 10332 189756 10342
rect 188692 9882 188804 9894
rect 188692 9830 188750 9882
rect 188802 9830 188804 9882
rect 188692 9828 188804 9830
rect 188748 9818 188804 9828
rect 188580 8990 188582 9042
rect 188634 8990 188636 9042
rect 188580 8978 188636 8990
rect 188692 9212 188748 9222
rect 188692 9154 188748 9156
rect 188692 9102 188694 9154
rect 188746 9102 188748 9154
rect 188468 8206 188470 8258
rect 188522 8206 188524 8258
rect 188468 8204 188524 8206
rect 188468 8128 188524 8148
rect 188692 8146 188748 9102
rect 188692 8094 188694 8146
rect 188746 8094 188748 8146
rect 188692 8082 188748 8094
rect 189140 8874 189196 8886
rect 189140 8822 189142 8874
rect 189194 8822 189196 8874
rect 188468 6860 188524 6870
rect 188468 6802 188524 6804
rect 188468 6750 188470 6802
rect 188522 6750 188524 6802
rect 188468 6738 188524 6750
rect 188692 6578 188748 6590
rect 188692 6526 188694 6578
rect 188746 6526 188748 6578
rect 188692 5628 188748 6526
rect 188692 5562 188748 5572
rect 188972 5068 189028 5078
rect 188972 4974 189028 5012
rect 189140 5068 189196 8822
rect 189364 8034 189420 8046
rect 189364 7982 189366 8034
rect 189418 7982 189420 8034
rect 189140 5002 189196 5012
rect 189252 6018 189308 6030
rect 189252 5966 189254 6018
rect 189306 5966 189308 6018
rect 188860 4956 188916 4966
rect 188356 4902 188358 4954
rect 188410 4902 188412 4954
rect 188356 4890 188412 4902
rect 188804 4954 188916 4956
rect 188804 4902 188862 4954
rect 188914 4902 188916 4954
rect 188804 4890 188916 4902
rect 188020 3882 188076 3892
rect 187572 3386 187628 3398
rect 187572 3334 187574 3386
rect 187626 3334 187628 3386
rect 187572 2380 187628 3334
rect 188804 3388 188860 4890
rect 188804 3322 188860 3332
rect 189252 4620 189308 5966
rect 189364 5180 189420 7982
rect 189700 7474 189756 10276
rect 189812 9826 189868 10948
rect 189812 9774 189814 9826
rect 189866 9774 189868 9826
rect 189812 9762 189868 9774
rect 190036 11002 190092 11014
rect 190036 10950 190038 11002
rect 190090 10950 190092 11002
rect 189924 9714 189980 9726
rect 189924 9662 189926 9714
rect 189978 9662 189980 9714
rect 189924 9548 189980 9662
rect 189924 9212 189980 9492
rect 189924 9146 189980 9156
rect 189700 7422 189702 7474
rect 189754 7422 189756 7474
rect 189700 7410 189756 7422
rect 189924 7586 189980 7598
rect 189924 7534 189926 7586
rect 189978 7534 189980 7586
rect 189588 7306 189644 7318
rect 189588 7254 189590 7306
rect 189642 7254 189644 7306
rect 189364 5114 189420 5124
rect 189476 6690 189532 6702
rect 189476 6638 189478 6690
rect 189530 6638 189532 6690
rect 189252 3387 189308 4564
rect 189476 3836 189532 6638
rect 189588 6636 189644 7254
rect 189588 6412 189644 6580
rect 189588 6346 189644 6356
rect 189812 6300 189868 6310
rect 189588 5906 189644 5918
rect 189588 5854 189590 5906
rect 189642 5854 189644 5906
rect 189588 4620 189644 5854
rect 189812 5738 189868 6244
rect 189812 5686 189814 5738
rect 189866 5686 189868 5738
rect 189812 5674 189868 5686
rect 189756 4956 189812 4966
rect 189756 4862 189812 4900
rect 189588 4554 189644 4564
rect 189476 3770 189532 3780
rect 189476 3498 189532 3510
rect 189476 3446 189478 3498
rect 189530 3446 189532 3498
rect 189252 3331 189420 3387
rect 187572 2314 187628 2324
rect 189364 2266 189420 3331
rect 189476 2492 189532 3446
rect 189924 3050 189980 7534
rect 189924 2998 189926 3050
rect 189978 2998 189980 3050
rect 189924 2986 189980 2998
rect 190036 2940 190092 10950
rect 190372 8316 190428 11732
rect 190484 8652 190540 14200
rect 191156 14028 191212 14200
rect 191156 13962 191212 13972
rect 191828 13916 191884 13926
rect 190596 13244 190652 13254
rect 190596 9210 190652 13188
rect 191716 11786 191772 11798
rect 191716 11734 191718 11786
rect 191770 11734 191772 11786
rect 191156 10556 191212 10566
rect 190596 9158 190598 9210
rect 190650 9158 190652 9210
rect 190596 9146 190652 9158
rect 190932 9212 190988 9222
rect 191156 9212 191212 10500
rect 191360 10220 191624 10230
rect 191416 10164 191464 10220
rect 191520 10164 191568 10220
rect 191360 10154 191624 10164
rect 191380 9996 191436 10006
rect 191380 9938 191436 9940
rect 191380 9886 191382 9938
rect 191434 9886 191436 9938
rect 191380 9874 191436 9886
rect 191716 9660 191772 11734
rect 191828 9994 191884 13860
rect 191940 12236 191996 14200
rect 191940 12170 191996 12180
rect 191828 9942 191830 9994
rect 191882 9942 191884 9994
rect 191828 9930 191884 9942
rect 192052 12122 192108 12134
rect 192052 12070 192054 12122
rect 192106 12070 192108 12122
rect 191828 9660 191884 9670
rect 191716 9604 191828 9660
rect 191436 9212 191492 9222
rect 191156 9210 191492 9212
rect 191156 9158 191438 9210
rect 191490 9158 191492 9210
rect 191156 9156 191492 9158
rect 190932 9118 190988 9156
rect 191436 9146 191492 9156
rect 191360 8652 191624 8662
rect 190484 8596 190652 8652
rect 190484 8316 190540 8326
rect 190372 8314 190540 8316
rect 190372 8262 190486 8314
rect 190538 8262 190540 8314
rect 190372 8260 190540 8262
rect 190484 8250 190540 8260
rect 190596 7642 190652 8596
rect 191416 8596 191464 8652
rect 191520 8596 191568 8652
rect 191360 8586 191624 8596
rect 190596 7590 190598 7642
rect 190650 7590 190652 7642
rect 190596 7578 190652 7590
rect 190708 8428 190764 8438
rect 190596 7420 190652 7430
rect 190596 6748 190652 7364
rect 190708 6860 190764 8372
rect 191828 8204 191884 9604
rect 191772 8148 191884 8204
rect 190820 8090 190876 8102
rect 190820 8038 190822 8090
rect 190874 8038 190876 8090
rect 190820 7756 190876 8038
rect 191324 8092 191380 8102
rect 191324 7998 191380 8036
rect 190820 7690 190876 7700
rect 190932 7644 190988 7654
rect 190708 6804 190876 6860
rect 190652 6692 190708 6748
rect 190596 6690 190708 6692
rect 190596 6682 190654 6690
rect 190652 6638 190654 6682
rect 190706 6638 190708 6690
rect 190652 6626 190708 6638
rect 190540 6522 190596 6534
rect 190540 6470 190542 6522
rect 190594 6470 190596 6522
rect 190540 5974 190596 6470
rect 190820 6086 190876 6804
rect 190932 6636 190988 7588
rect 191772 7586 191828 8148
rect 191772 7534 191774 7586
rect 191826 7534 191828 7586
rect 191772 7522 191828 7534
rect 191660 7308 191716 7318
rect 191660 7214 191716 7252
rect 191360 7084 191624 7094
rect 191416 7028 191464 7084
rect 191520 7028 191568 7084
rect 191360 7018 191624 7028
rect 191772 6748 191828 6758
rect 190932 6580 191044 6636
rect 191772 6634 191828 6692
rect 190820 6074 190932 6086
rect 190820 6022 190878 6074
rect 190930 6022 190932 6074
rect 190820 6020 190932 6022
rect 190876 6010 190932 6020
rect 190988 6018 191044 6580
rect 191324 6578 191380 6590
rect 190484 5964 190596 5974
rect 190540 5908 190596 5964
rect 190988 5966 190990 6018
rect 191042 5966 191044 6018
rect 191212 6522 191268 6534
rect 191212 6470 191214 6522
rect 191266 6470 191268 6522
rect 191212 6076 191268 6470
rect 191212 6010 191268 6020
rect 191324 6526 191326 6578
rect 191378 6526 191380 6578
rect 191772 6582 191774 6634
rect 191826 6582 191828 6634
rect 191772 6570 191828 6582
rect 190988 5954 191044 5966
rect 190484 5898 190540 5908
rect 191324 5852 191380 6526
rect 192052 6076 192108 12070
rect 192388 11898 192444 11910
rect 192388 11846 192390 11898
rect 192442 11846 192444 11898
rect 192164 9772 192220 9782
rect 192164 9678 192220 9716
rect 192276 8247 192332 8259
rect 192276 8195 192278 8247
rect 192330 8195 192332 8247
rect 192276 7644 192332 8195
rect 192388 7654 192444 11846
rect 192612 11788 192668 14200
rect 193396 13916 193452 14200
rect 193956 14140 194012 14150
rect 194068 14140 194124 14200
rect 194012 14084 194124 14140
rect 193956 14074 194012 14084
rect 193396 13850 193452 13860
rect 193620 13020 193676 13030
rect 192612 11722 192668 11732
rect 193060 12346 193116 12358
rect 193060 12294 193062 12346
rect 193114 12294 193116 12346
rect 192948 9884 193004 9894
rect 192780 9658 192836 9670
rect 192780 9606 192782 9658
rect 192834 9606 192836 9658
rect 192780 9548 192836 9606
rect 192836 9492 192892 9548
rect 192780 9482 192892 9492
rect 192836 9154 192892 9482
rect 192836 9102 192838 9154
rect 192890 9102 192892 9154
rect 192836 9090 192892 9102
rect 192724 8930 192780 8942
rect 192724 8878 192726 8930
rect 192778 8878 192780 8930
rect 192388 7642 192500 7654
rect 192388 7590 192446 7642
rect 192498 7590 192500 7642
rect 192388 7588 192500 7590
rect 192276 7578 192332 7588
rect 192444 7578 192500 7588
rect 192724 6748 192780 8878
rect 192948 7654 193004 9828
rect 193060 9100 193116 12294
rect 193060 9042 193116 9044
rect 193060 8990 193062 9042
rect 193114 8990 193116 9042
rect 193060 8978 193116 8990
rect 193620 8258 193676 12964
rect 194068 12460 194124 14084
rect 194068 12394 194124 12404
rect 194628 12012 194684 12022
rect 194852 12012 194908 14200
rect 195524 13020 195580 14200
rect 195524 12954 195580 12964
rect 196308 13804 196364 14200
rect 196308 12796 196364 13748
rect 196308 12730 196364 12740
rect 196420 14138 196476 14150
rect 196420 14086 196422 14138
rect 196474 14086 196476 14138
rect 196308 12570 196364 12582
rect 196308 12518 196310 12570
rect 196362 12518 196364 12570
rect 195860 12348 195916 12358
rect 194852 11956 195132 12012
rect 193732 11788 193788 11798
rect 193732 9994 193788 11732
rect 193732 9942 193734 9994
rect 193786 9942 193788 9994
rect 193732 9930 193788 9942
rect 194068 11340 194124 11350
rect 194068 9658 194124 11284
rect 194068 9606 194070 9658
rect 194122 9606 194124 9658
rect 193620 8206 193622 8258
rect 193674 8206 193676 8258
rect 192892 7642 193004 7654
rect 192892 7590 192894 7642
rect 192946 7590 193004 7642
rect 192892 7588 193004 7590
rect 193060 7980 193116 7990
rect 192892 7578 192948 7588
rect 193060 6758 193116 7924
rect 193620 7308 193676 8206
rect 193844 9212 193900 9222
rect 193844 8764 193900 9156
rect 193844 8204 193900 8708
rect 194068 8427 194124 9606
rect 194516 10890 194572 10902
rect 194516 10838 194518 10890
rect 194570 10838 194572 10890
rect 194516 9210 194572 10838
rect 194516 9158 194518 9210
rect 194570 9158 194572 9210
rect 194516 9146 194572 9158
rect 194068 8371 194572 8427
rect 193844 8148 193956 8204
rect 193788 7644 193844 7654
rect 193788 7550 193844 7588
rect 193900 7586 193956 8148
rect 193900 7534 193902 7586
rect 193954 7534 193956 7586
rect 193900 7522 193956 7534
rect 194348 7420 194404 7430
rect 193620 7242 193676 7252
rect 194068 7418 194404 7420
rect 194068 7366 194350 7418
rect 194402 7366 194404 7418
rect 194068 7364 194404 7366
rect 193732 6972 193788 6982
rect 192724 6692 192892 6748
rect 193060 6746 193172 6758
rect 193060 6694 193118 6746
rect 193170 6694 193172 6746
rect 193060 6692 193172 6694
rect 192836 6580 192892 6692
rect 193116 6682 193172 6692
rect 192220 6522 192276 6534
rect 192220 6470 192222 6522
rect 192274 6470 192276 6522
rect 192220 6300 192276 6470
rect 192668 6524 192724 6534
rect 192836 6524 193116 6580
rect 192668 6430 192724 6468
rect 192220 6234 192276 6244
rect 192892 6412 192948 6422
rect 192444 6076 192500 6086
rect 192052 6074 192500 6076
rect 192052 6022 192446 6074
rect 192498 6022 192500 6074
rect 192052 6020 192500 6022
rect 192444 6010 192500 6020
rect 192892 6074 192948 6356
rect 192892 6022 192894 6074
rect 192946 6022 192948 6074
rect 192892 6010 192948 6022
rect 191156 5796 191380 5852
rect 191436 5850 191492 5862
rect 191436 5798 191438 5850
rect 191490 5798 191492 5850
rect 191156 5404 191212 5796
rect 191436 5740 191492 5798
rect 191436 5674 191492 5684
rect 191360 5516 191624 5526
rect 191416 5460 191464 5516
rect 191520 5460 191568 5516
rect 191360 5450 191624 5460
rect 193060 5516 193116 6524
rect 193564 6524 193620 6534
rect 193564 6430 193620 6468
rect 193732 6086 193788 6916
rect 193340 6076 193396 6086
rect 193732 6074 193844 6086
rect 193732 6022 193790 6074
rect 193842 6022 193844 6074
rect 193732 6020 193844 6022
rect 193340 5982 193396 6020
rect 193788 6010 193844 6020
rect 193060 5450 193116 5460
rect 194068 5404 194124 7364
rect 194348 7354 194404 7364
rect 194348 6578 194404 6590
rect 194236 6522 194292 6534
rect 194236 6470 194238 6522
rect 194290 6470 194292 6522
rect 194236 6076 194292 6470
rect 194348 6526 194350 6578
rect 194402 6526 194404 6578
rect 194348 6300 194404 6526
rect 194348 6234 194404 6244
rect 194236 6020 194460 6076
rect 194236 5852 194292 5862
rect 194236 5850 194348 5852
rect 194236 5798 194238 5850
rect 194290 5798 194348 5850
rect 194236 5786 194348 5798
rect 191156 5348 191324 5404
rect 190204 4956 190260 4966
rect 190148 4954 190260 4956
rect 190148 4902 190206 4954
rect 190258 4902 190260 4954
rect 190148 4890 190260 4902
rect 190652 4956 190708 4966
rect 190148 4058 190204 4890
rect 190652 4862 190708 4900
rect 191100 4954 191156 4966
rect 191100 4902 191102 4954
rect 191154 4902 191156 4954
rect 191100 4508 191156 4902
rect 191268 4508 191324 5348
rect 193844 5348 194124 5404
rect 191548 4954 191604 4966
rect 191548 4902 191550 4954
rect 191602 4902 191604 4954
rect 191380 4508 191436 4518
rect 191268 4452 191380 4508
rect 191100 4442 191156 4452
rect 190148 4006 190150 4058
rect 190202 4006 190204 4058
rect 190148 3994 190204 4006
rect 191268 4060 191324 4070
rect 191268 3966 191324 4004
rect 191380 3948 191436 4452
rect 191548 4396 191604 4902
rect 191996 4954 192052 4966
rect 191996 4902 191998 4954
rect 192050 4902 192052 4954
rect 191996 4620 192052 4902
rect 192444 4956 192500 4966
rect 192444 4862 192500 4900
rect 192892 4954 192948 4966
rect 192892 4902 192894 4954
rect 192946 4902 192948 4954
rect 192892 4844 192948 4902
rect 193676 4956 193732 4966
rect 193676 4862 193732 4900
rect 192892 4778 192948 4788
rect 193060 4844 193116 4854
rect 191996 4554 192052 4564
rect 191380 3882 191436 3892
rect 191492 4340 191604 4396
rect 191492 3834 191548 4340
rect 191492 3782 191494 3834
rect 191546 3782 191548 3834
rect 191492 3770 191548 3782
rect 191716 4284 191772 4294
rect 190036 2874 190092 2884
rect 190932 3276 190988 3286
rect 189476 2426 189532 2436
rect 189364 2214 189366 2266
rect 189418 2214 189420 2266
rect 189364 2202 189420 2214
rect 190372 2380 190428 2390
rect 187460 2090 187516 2100
rect 188692 2156 188748 2166
rect 188692 2062 188748 2100
rect 189700 1932 189756 1942
rect 188468 1820 188524 1830
rect 187908 1596 187964 1606
rect 187908 800 187964 1540
rect 188468 800 188524 1764
rect 189140 1596 189196 1606
rect 189140 800 189196 1540
rect 189700 800 189756 1876
rect 190372 800 190428 2324
rect 190596 2380 190652 2390
rect 190596 2286 190652 2324
rect 190932 800 190988 3220
rect 191604 3274 191660 3286
rect 191604 3222 191606 3274
rect 191658 3222 191660 3274
rect 191604 800 191660 3222
rect 191716 3052 191772 4228
rect 193060 4058 193116 4788
rect 193060 4006 193062 4058
rect 193114 4006 193116 4058
rect 193060 3994 193116 4006
rect 191716 2986 191772 2996
rect 192276 3052 192332 3062
rect 192276 2958 192332 2996
rect 193844 2268 193900 5348
rect 194124 4956 194180 4966
rect 194124 4954 194236 4956
rect 194124 4902 194126 4954
rect 194178 4902 194236 4954
rect 194124 4890 194236 4902
rect 194180 3946 194236 4890
rect 194292 4060 194348 5786
rect 194404 5404 194460 6020
rect 194516 5964 194572 8371
rect 194628 8090 194684 11956
rect 194964 10554 195020 10566
rect 194964 10502 194966 10554
rect 195018 10502 195020 10554
rect 194740 9772 194796 9782
rect 194740 9678 194796 9716
rect 194964 9324 195020 10502
rect 195076 9994 195132 11956
rect 195076 9942 195078 9994
rect 195130 9942 195132 9994
rect 195076 9930 195132 9942
rect 195636 9660 195692 9670
rect 195636 9566 195692 9604
rect 194628 8038 194630 8090
rect 194682 8038 194684 8090
rect 194628 8026 194684 8038
rect 194852 9098 194908 9110
rect 194852 9046 194854 9098
rect 194906 9046 194908 9098
rect 194852 6748 194908 9046
rect 194964 8204 195020 9268
rect 195188 9212 195244 9222
rect 195412 9212 195468 9222
rect 195244 9156 195356 9212
rect 195188 9146 195244 9156
rect 195300 8988 195356 9156
rect 195412 9118 195468 9156
rect 195748 9098 195804 9110
rect 195748 9046 195750 9098
rect 195802 9046 195804 9098
rect 195524 8988 195580 8998
rect 195300 8932 195468 8988
rect 194964 8148 195076 8204
rect 195020 7586 195076 8148
rect 195020 7534 195022 7586
rect 195074 7534 195076 7586
rect 195132 7644 195188 7654
rect 195132 7550 195188 7588
rect 195020 7522 195076 7534
rect 194852 6682 194908 6692
rect 194796 6522 194852 6534
rect 194796 6470 194798 6522
rect 194850 6470 194852 6522
rect 194796 6412 194852 6470
rect 195244 6524 195300 6534
rect 195244 6430 195300 6468
rect 194796 6346 194852 6356
rect 195412 6300 195468 8932
rect 195524 7654 195580 8932
rect 195524 7642 195636 7654
rect 195524 7590 195582 7642
rect 195634 7590 195636 7642
rect 195524 7588 195636 7590
rect 195580 7578 195636 7588
rect 195748 6972 195804 9046
rect 195748 6906 195804 6916
rect 195692 6748 195748 6758
rect 195860 6748 195916 12292
rect 196196 11900 196252 11910
rect 195972 11788 196028 11798
rect 195972 9994 196028 11732
rect 195972 9942 195974 9994
rect 196026 9942 196028 9994
rect 195972 9930 196028 9942
rect 195972 9660 196028 9670
rect 195972 8988 196028 9604
rect 195972 8922 196028 8932
rect 196028 7756 196084 7766
rect 196028 7642 196084 7700
rect 196028 7590 196030 7642
rect 196082 7590 196084 7642
rect 196028 7578 196084 7590
rect 196196 7420 196252 11844
rect 196308 9210 196364 12518
rect 196420 9994 196476 14086
rect 196420 9942 196422 9994
rect 196474 9942 196476 9994
rect 196420 9930 196476 9942
rect 196868 12236 196924 12246
rect 196308 9158 196310 9210
rect 196362 9158 196364 9210
rect 196308 9146 196364 9158
rect 196756 9658 196812 9670
rect 196756 9606 196758 9658
rect 196810 9606 196812 9658
rect 196644 9098 196700 9110
rect 196644 9046 196646 9098
rect 196698 9046 196700 9098
rect 196420 8258 196476 8270
rect 196420 8206 196422 8258
rect 196474 8206 196476 8258
rect 196420 7644 196476 8206
rect 196420 7578 196476 7588
rect 196476 7420 196532 7430
rect 196196 7418 196532 7420
rect 196196 7366 196478 7418
rect 196530 7366 196532 7418
rect 196196 7364 196532 7366
rect 196476 7354 196532 7364
rect 195692 6746 195916 6748
rect 195692 6694 195694 6746
rect 195746 6694 195916 6746
rect 195692 6692 195916 6694
rect 196644 6748 196700 9046
rect 196756 8652 196812 9606
rect 196756 8586 196812 8596
rect 196868 8428 196924 12180
rect 196980 11788 197036 14200
rect 196980 11722 197036 11732
rect 197204 14026 197260 14038
rect 197204 13974 197206 14026
rect 197258 13974 197260 14026
rect 197204 9210 197260 13974
rect 197764 12124 197820 14200
rect 197764 12058 197820 12068
rect 198436 13580 198492 14200
rect 198436 11900 198492 13524
rect 198436 11834 198492 11844
rect 198660 12796 198716 12806
rect 198100 11788 198156 11798
rect 198100 9994 198156 11732
rect 198324 11116 198380 11126
rect 198100 9942 198102 9994
rect 198154 9942 198156 9994
rect 198100 9930 198156 9942
rect 198212 10780 198268 10790
rect 197764 9660 197820 9670
rect 197764 9566 197820 9604
rect 197204 9158 197206 9210
rect 197258 9158 197260 9210
rect 197204 9146 197260 9158
rect 198044 9212 198100 9222
rect 198044 9118 198100 9156
rect 197540 9098 197596 9110
rect 197540 9046 197542 9098
rect 197594 9046 197596 9098
rect 197540 8540 197596 9046
rect 197540 8474 197596 8484
rect 197988 8876 198044 8886
rect 196756 8372 196924 8428
rect 196756 6758 196812 8372
rect 197316 8316 197372 8326
rect 197316 7654 197372 8260
rect 197540 8316 197596 8326
rect 197540 8258 197596 8260
rect 197540 8206 197542 8258
rect 197594 8206 197596 8258
rect 196924 7644 196980 7654
rect 197316 7642 197428 7654
rect 197316 7590 197374 7642
rect 197426 7590 197428 7642
rect 197316 7588 197428 7590
rect 196924 7550 196980 7588
rect 197372 7578 197428 7588
rect 197540 7084 197596 8206
rect 197820 7418 197876 7430
rect 197820 7366 197822 7418
rect 197874 7366 197876 7418
rect 197820 7196 197876 7366
rect 197820 7130 197876 7140
rect 197540 7018 197596 7028
rect 196756 6746 196868 6758
rect 196756 6694 196814 6746
rect 196866 6694 196868 6746
rect 196756 6692 196868 6694
rect 195692 6682 195748 6692
rect 196644 6682 196700 6692
rect 196812 6682 196868 6692
rect 196364 6636 196420 6646
rect 196364 6542 196420 6580
rect 197260 6636 197316 6646
rect 197260 6542 197316 6580
rect 195300 6244 195468 6300
rect 197708 6522 197764 6534
rect 197708 6470 197710 6522
rect 197762 6470 197764 6522
rect 195132 6076 195188 6086
rect 195132 5982 195188 6020
rect 194516 5898 194572 5908
rect 194684 5852 194740 5862
rect 194684 5850 194796 5852
rect 194684 5798 194686 5850
rect 194738 5798 194796 5850
rect 194684 5786 194796 5798
rect 194404 5338 194460 5348
rect 194572 4956 194628 4966
rect 194516 4954 194628 4956
rect 194516 4902 194574 4954
rect 194626 4902 194628 4954
rect 194516 4890 194628 4902
rect 194516 4172 194572 4890
rect 194516 4106 194572 4116
rect 194292 3994 194348 4004
rect 194180 3894 194182 3946
rect 194234 3894 194236 3946
rect 194180 3882 194236 3894
rect 194068 3836 194124 3846
rect 194068 3388 194124 3780
rect 194068 3322 194124 3332
rect 193844 2202 193900 2212
rect 193956 3276 194012 3286
rect 192836 1148 192892 1158
rect 191828 868 192220 924
rect 142548 746 142604 756
rect 142744 0 142856 800
rect 143416 0 143528 800
rect 143976 0 144088 800
rect 144648 0 144760 800
rect 145208 0 145320 800
rect 145768 0 145880 800
rect 146440 0 146552 800
rect 147000 0 147112 800
rect 147672 0 147784 800
rect 148232 0 148344 800
rect 148904 0 149016 800
rect 149464 0 149576 800
rect 150136 0 150248 800
rect 150696 0 150808 800
rect 151256 0 151368 800
rect 151928 0 152040 800
rect 152488 0 152600 800
rect 153160 0 153272 800
rect 153720 0 153832 800
rect 154392 0 154504 800
rect 154952 0 155064 800
rect 155624 0 155736 800
rect 156184 0 156296 800
rect 156744 0 156856 800
rect 157416 0 157528 800
rect 157976 0 158088 800
rect 158648 0 158760 800
rect 159208 0 159320 800
rect 159880 0 159992 800
rect 160440 0 160552 800
rect 161112 0 161224 800
rect 161672 0 161784 800
rect 162232 0 162344 800
rect 162904 0 163016 800
rect 163464 0 163576 800
rect 164136 0 164248 800
rect 164696 0 164808 800
rect 165368 0 165480 800
rect 165928 0 166040 800
rect 166488 0 166600 800
rect 167160 0 167272 800
rect 167720 0 167832 800
rect 168392 0 168504 800
rect 168952 0 169064 800
rect 169624 0 169736 800
rect 170184 0 170296 800
rect 170856 0 170968 800
rect 171416 0 171528 800
rect 171976 0 172088 800
rect 172648 0 172760 800
rect 173208 0 173320 800
rect 173880 0 173992 800
rect 174440 0 174552 800
rect 175112 0 175224 800
rect 175672 0 175784 800
rect 176344 0 176456 800
rect 176904 0 177016 800
rect 177464 0 177576 800
rect 178136 0 178248 800
rect 178696 0 178808 800
rect 179368 0 179480 800
rect 179928 0 180040 800
rect 180600 0 180712 800
rect 181160 0 181272 800
rect 181832 0 181944 800
rect 182392 0 182504 800
rect 182952 0 183064 800
rect 183624 0 183736 800
rect 184184 0 184296 800
rect 184856 0 184968 800
rect 185416 0 185528 800
rect 186088 0 186200 800
rect 186648 0 186760 800
rect 187320 0 187432 800
rect 187880 0 187992 800
rect 188440 0 188552 800
rect 189112 0 189224 800
rect 189672 0 189784 800
rect 190344 0 190456 800
rect 190904 0 191016 800
rect 191576 0 191688 800
rect 191828 700 191884 868
rect 192164 800 192220 868
rect 192836 800 192892 1092
rect 193396 1034 193452 1046
rect 193396 982 193398 1034
rect 193450 982 193452 1034
rect 193396 800 193452 982
rect 193956 800 194012 3220
rect 194740 3164 194796 5786
rect 195020 4956 195076 4966
rect 194964 4954 195076 4956
rect 194964 4902 195022 4954
rect 195074 4902 195076 4954
rect 194964 4890 195076 4902
rect 194964 3836 195020 4890
rect 195300 4172 195356 6244
rect 197708 6076 197764 6470
rect 197708 6010 197764 6020
rect 197764 5906 197820 5918
rect 195580 5852 195636 5862
rect 197764 5854 197766 5906
rect 197818 5854 197820 5906
rect 195580 5850 195692 5852
rect 195580 5798 195582 5850
rect 195634 5798 195692 5850
rect 195580 5786 195692 5798
rect 195468 4956 195524 4966
rect 195468 4862 195524 4900
rect 195636 4284 195692 5786
rect 196532 5794 196588 5806
rect 196532 5742 196534 5794
rect 196586 5742 196588 5794
rect 195916 4956 195972 4966
rect 195636 4218 195692 4228
rect 195860 4954 195972 4956
rect 195860 4902 195918 4954
rect 195970 4902 195972 4954
rect 195860 4890 195972 4902
rect 196364 4954 196420 4966
rect 196364 4902 196366 4954
rect 196418 4902 196420 4954
rect 195300 4106 195356 4116
rect 194964 3770 195020 3780
rect 195860 3612 195916 4890
rect 196364 4396 196420 4902
rect 196364 4330 196420 4340
rect 195860 3546 195916 3556
rect 194740 3098 194796 3108
rect 196420 2602 196476 2614
rect 196420 2550 196422 2602
rect 196474 2550 196476 2602
rect 194628 1708 194684 1718
rect 194628 800 194684 1652
rect 196420 1708 196476 2550
rect 196420 1642 196476 1652
rect 196532 1484 196588 5742
rect 196812 4956 196868 4966
rect 196756 4954 196868 4956
rect 196756 4902 196814 4954
rect 196866 4902 196868 4954
rect 196756 4890 196868 4902
rect 196756 3500 196812 4890
rect 197764 4396 197820 5854
rect 197988 5122 198044 8820
rect 198212 7654 198268 10724
rect 198324 9212 198380 11060
rect 198492 9884 198548 9894
rect 198492 9790 198548 9828
rect 198492 9212 198548 9222
rect 198324 9210 198548 9212
rect 198324 9158 198494 9210
rect 198546 9158 198548 9210
rect 198324 9156 198548 9158
rect 198492 9146 198548 9156
rect 198660 7654 198716 12740
rect 199220 11788 199276 14200
rect 199220 11722 199276 11732
rect 199332 12460 199388 12470
rect 199108 9658 199164 9670
rect 199108 9606 199110 9658
rect 199162 9606 199164 9658
rect 199108 9212 199164 9606
rect 199332 9222 199388 12404
rect 199892 12012 199948 14200
rect 200676 13132 200732 14200
rect 200676 12348 200732 13076
rect 199892 11946 199948 11956
rect 200228 12292 200732 12348
rect 199668 11900 199724 11910
rect 199444 11788 199500 11798
rect 199444 9994 199500 11732
rect 199444 9942 199446 9994
rect 199498 9942 199500 9994
rect 199444 9930 199500 9942
rect 199332 9210 199444 9222
rect 199332 9158 199390 9210
rect 199442 9158 199444 9210
rect 199332 9156 199444 9158
rect 198940 8986 198996 8998
rect 198940 8934 198942 8986
rect 198994 8934 198996 8986
rect 198940 8428 198996 8934
rect 199108 8764 199164 9156
rect 199388 9146 199444 9156
rect 199108 8698 199164 8708
rect 198940 8362 198996 8372
rect 199668 8426 199724 11844
rect 199948 9658 200004 9670
rect 199948 9606 199950 9658
rect 200002 9606 200004 9658
rect 199948 9548 200004 9606
rect 199948 9482 200004 9492
rect 199668 8374 199670 8426
rect 199722 8374 199724 8426
rect 199668 8362 199724 8374
rect 198212 7642 198324 7654
rect 198212 7590 198270 7642
rect 198322 7590 198324 7642
rect 198212 7588 198324 7590
rect 198660 7642 198772 7654
rect 198660 7590 198718 7642
rect 198770 7590 198772 7642
rect 198660 7588 198772 7590
rect 198268 7578 198324 7588
rect 198716 7578 198772 7588
rect 199612 7532 199668 7542
rect 199780 7532 199836 7542
rect 199668 7476 199724 7532
rect 199612 7438 199724 7476
rect 199164 7420 199220 7430
rect 199164 7326 199220 7364
rect 198324 6972 198380 6982
rect 198156 6524 198212 6534
rect 197988 5070 197990 5122
rect 198042 5070 198044 5122
rect 197988 5058 198044 5070
rect 198100 6522 198212 6524
rect 198100 6470 198158 6522
rect 198210 6470 198212 6522
rect 198100 6458 198212 6470
rect 197876 5010 197932 5022
rect 197876 4958 197878 5010
rect 197930 4958 197932 5010
rect 197876 4732 197932 4958
rect 197876 4666 197932 4676
rect 197764 4330 197820 4340
rect 196756 3434 196812 3444
rect 198100 2380 198156 6458
rect 198100 2314 198156 2324
rect 196532 1418 196588 1428
rect 197652 1596 197708 1606
rect 195188 1036 195244 1046
rect 195188 800 195244 980
rect 197092 1036 197148 1046
rect 195636 868 195916 924
rect 191828 634 191884 644
rect 192136 0 192248 800
rect 192808 0 192920 800
rect 193368 0 193480 800
rect 193928 0 194040 800
rect 194600 0 194712 800
rect 195160 0 195272 800
rect 195636 700 195692 868
rect 195860 800 195916 868
rect 196196 868 196476 924
rect 196196 810 196252 868
rect 195412 644 195692 700
rect 195412 586 195468 644
rect 195412 534 195414 586
rect 195466 534 195468 586
rect 195412 522 195468 534
rect 195832 0 195944 800
rect 196196 758 196198 810
rect 196250 758 196252 810
rect 196420 800 196476 868
rect 197092 800 197148 980
rect 197652 800 197708 1540
rect 198324 800 198380 6916
rect 198772 6748 198828 6758
rect 198492 5852 198548 5862
rect 198492 5758 198548 5796
rect 198772 1596 198828 6692
rect 199668 6524 199724 7438
rect 199780 6748 199836 7476
rect 199780 6682 199836 6692
rect 199668 6458 199724 6468
rect 199388 6188 199444 6198
rect 199388 6074 199444 6132
rect 199388 6022 199390 6074
rect 199442 6022 199444 6074
rect 199388 6010 199444 6022
rect 200228 6076 200284 12292
rect 200564 12124 200620 12134
rect 200396 9884 200452 9894
rect 200396 9790 200452 9828
rect 200396 9548 200452 9558
rect 200396 9210 200452 9492
rect 200396 9158 200398 9210
rect 200450 9158 200452 9210
rect 200396 8988 200452 9158
rect 200564 9212 200620 12068
rect 201348 11788 201404 14200
rect 201348 11722 201404 11732
rect 201460 13692 201516 13702
rect 200676 10668 200732 10678
rect 200676 9894 200732 10612
rect 200900 10666 200956 10678
rect 200900 10614 200902 10666
rect 200954 10614 200956 10666
rect 200676 9882 200788 9894
rect 200676 9830 200734 9882
rect 200786 9830 200788 9882
rect 200676 9828 200788 9830
rect 200732 9818 200788 9828
rect 200900 9222 200956 10614
rect 200564 9156 200732 9212
rect 200396 8314 200452 8932
rect 200396 8262 200398 8314
rect 200450 8262 200452 8314
rect 200396 8250 200452 8262
rect 200564 7868 200620 7878
rect 200564 7474 200620 7812
rect 200564 7422 200566 7474
rect 200618 7422 200620 7474
rect 200564 7410 200620 7422
rect 200564 6860 200620 6870
rect 200676 6860 200732 9156
rect 200844 9210 200956 9222
rect 200844 9158 200846 9210
rect 200898 9158 200956 9210
rect 200844 9156 200956 9158
rect 201292 9772 201348 9782
rect 201292 9210 201348 9716
rect 201292 9158 201294 9210
rect 201346 9158 201348 9210
rect 200844 9146 200900 9156
rect 201292 8876 201348 9158
rect 201292 8810 201348 8820
rect 201460 8326 201516 13636
rect 201572 12236 201628 12246
rect 201572 11676 201628 12180
rect 202132 11900 202188 14200
rect 202804 13692 202860 14200
rect 202804 13626 202860 13636
rect 203028 12236 203084 12246
rect 202132 11834 202188 11844
rect 202580 12012 202636 12022
rect 201572 11610 201628 11620
rect 202020 11788 202076 11798
rect 202020 9994 202076 11732
rect 202356 11004 202412 11014
rect 202020 9942 202022 9994
rect 202074 9942 202076 9994
rect 202020 9930 202076 9942
rect 202132 10892 202188 10902
rect 201684 9658 201740 9670
rect 201684 9606 201686 9658
rect 201738 9606 201740 9658
rect 201684 9324 201740 9606
rect 201684 9258 201740 9268
rect 202132 9222 202188 10836
rect 202356 9894 202412 10948
rect 202356 9882 202468 9894
rect 202356 9830 202414 9882
rect 202466 9830 202468 9882
rect 202356 9828 202468 9830
rect 202412 9818 202468 9828
rect 202132 9210 202244 9222
rect 202132 9158 202190 9210
rect 202242 9158 202244 9210
rect 202132 9156 202244 9158
rect 202188 9146 202244 9156
rect 201740 8988 201796 8998
rect 201796 8932 202076 8988
rect 201740 8894 201796 8932
rect 201404 8314 201516 8326
rect 201404 8262 201406 8314
rect 201458 8262 201516 8314
rect 201404 8260 201516 8262
rect 201404 8250 201460 8260
rect 200844 8092 200900 8102
rect 200564 6858 200732 6860
rect 200564 6806 200566 6858
rect 200618 6806 200732 6858
rect 200564 6804 200732 6806
rect 200788 8090 200900 8092
rect 200788 8038 200846 8090
rect 200898 8038 200900 8090
rect 200788 8026 200900 8038
rect 201740 8092 201796 8102
rect 202020 8092 202076 8932
rect 202580 8876 202636 11956
rect 202860 9660 202916 9670
rect 202860 9566 202916 9604
rect 202692 9436 202748 9446
rect 202692 9212 202748 9380
rect 203028 9324 203084 12180
rect 203476 11900 203532 11910
rect 203308 9884 203364 9894
rect 203308 9790 203364 9828
rect 202692 9146 202748 9156
rect 202804 9268 203084 9324
rect 202356 8820 202636 8876
rect 202188 8204 202244 8214
rect 202188 8110 202244 8148
rect 201740 8090 201964 8092
rect 201740 8038 201742 8090
rect 201794 8038 201964 8090
rect 201740 8036 201964 8038
rect 201740 8026 201796 8036
rect 200788 6860 200844 8026
rect 200564 6794 200620 6804
rect 200788 6794 200844 6804
rect 201572 7362 201628 7374
rect 201572 7310 201574 7362
rect 201626 7310 201628 7362
rect 200900 6690 200956 6702
rect 200900 6638 200902 6690
rect 200954 6638 200956 6690
rect 200900 6636 200956 6638
rect 200900 6570 200956 6580
rect 200508 6076 200564 6086
rect 200228 6074 200564 6076
rect 200228 6022 200510 6074
rect 200562 6022 200564 6074
rect 200228 6020 200564 6022
rect 200508 6010 200564 6020
rect 198940 5852 198996 5862
rect 198884 5850 198996 5852
rect 198884 5798 198942 5850
rect 198994 5798 198996 5850
rect 198884 5786 198996 5798
rect 200844 5852 200900 5862
rect 200844 5850 200956 5852
rect 200844 5798 200846 5850
rect 200898 5798 200956 5850
rect 200844 5786 200956 5798
rect 198884 2156 198940 5786
rect 199836 4956 199892 4966
rect 199780 4954 199892 4956
rect 199780 4902 199838 4954
rect 199890 4902 199892 4954
rect 199780 4890 199892 4902
rect 200284 4954 200340 4966
rect 200732 4956 200788 4966
rect 200284 4902 200286 4954
rect 200338 4902 200340 4954
rect 199780 2716 199836 4890
rect 200284 4732 200340 4902
rect 200284 4666 200340 4676
rect 200676 4954 200788 4956
rect 200676 4902 200734 4954
rect 200786 4902 200788 4954
rect 200676 4890 200788 4902
rect 200900 4956 200956 5786
rect 200900 4890 200956 4900
rect 200676 3948 200732 4890
rect 200676 3882 200732 3892
rect 201572 3052 201628 7310
rect 201684 5292 201740 5302
rect 201684 5122 201740 5236
rect 201684 5070 201686 5122
rect 201738 5070 201740 5122
rect 201684 4284 201740 5070
rect 201796 5010 201852 5022
rect 201796 4958 201798 5010
rect 201850 4958 201852 5010
rect 201796 4844 201852 4958
rect 201796 4778 201852 4788
rect 201684 4218 201740 4228
rect 201908 4060 201964 8036
rect 202020 8026 202076 8036
rect 202356 6074 202412 8820
rect 202636 8092 202692 8102
rect 202356 6022 202358 6074
rect 202410 6022 202412 6074
rect 202356 6010 202412 6022
rect 202468 8090 202692 8092
rect 202468 8038 202638 8090
rect 202690 8038 202692 8090
rect 202468 8036 202692 8038
rect 202020 5628 202076 5638
rect 202020 4620 202076 5572
rect 202020 4554 202076 4564
rect 201684 4004 201964 4060
rect 201684 3276 201740 4004
rect 201684 3220 201964 3276
rect 201572 2996 201740 3052
rect 199780 2650 199836 2660
rect 200676 2828 200732 2838
rect 198884 2090 198940 2100
rect 199444 1596 199500 1606
rect 198772 1540 198940 1596
rect 198884 800 198940 1540
rect 199444 800 199500 1540
rect 200116 1596 200172 1606
rect 200116 800 200172 1540
rect 200676 800 200732 2772
rect 201572 2714 201628 2726
rect 201572 2662 201574 2714
rect 201626 2662 201628 2714
rect 201348 1036 201404 1046
rect 201348 800 201404 980
rect 201572 1036 201628 2662
rect 201684 1372 201740 2996
rect 201908 1932 201964 3220
rect 202468 3052 202524 8036
rect 202636 8026 202692 8036
rect 202804 7868 202860 9268
rect 203252 9212 203308 9222
rect 203476 9212 203532 11844
rect 203588 11788 203644 14200
rect 204260 12124 204316 14200
rect 204820 12908 204876 12918
rect 204260 12058 204316 12068
rect 204372 12348 204428 12358
rect 203588 11722 203644 11732
rect 204372 11004 204428 12292
rect 204260 10948 204428 11004
rect 204596 11788 204652 11798
rect 204260 10108 204316 10948
rect 204036 9996 204092 10006
rect 203868 9660 203924 9670
rect 203868 9658 203980 9660
rect 203868 9606 203870 9658
rect 203922 9606 203980 9658
rect 203868 9594 203980 9606
rect 203252 9210 203532 9212
rect 203252 9158 203254 9210
rect 203306 9158 203532 9210
rect 203252 9156 203532 9158
rect 203252 9146 203308 9156
rect 202916 9100 202972 9110
rect 202916 9098 203196 9100
rect 202916 9046 202918 9098
rect 202970 9046 203196 9098
rect 202916 9044 203196 9046
rect 202916 9034 202972 9044
rect 203140 8427 203196 9044
rect 203140 8371 203308 8427
rect 203084 8092 203140 8102
rect 203084 7998 203140 8036
rect 202804 7812 203140 7868
rect 203084 7642 203140 7812
rect 203084 7590 203086 7642
rect 203138 7590 203140 7642
rect 203084 7578 203140 7590
rect 202636 7420 202692 7430
rect 202636 7326 202692 7364
rect 203252 7196 203308 8371
rect 203924 8204 203980 9594
rect 204036 9042 204092 9940
rect 204036 8990 204038 9042
rect 204090 8990 204092 9042
rect 204036 8978 204092 8990
rect 203644 8090 203700 8102
rect 203644 8038 203646 8090
rect 203698 8038 203700 8090
rect 203644 7980 203700 8038
rect 203644 7914 203700 7924
rect 203532 7420 203588 7430
rect 203532 7326 203588 7364
rect 203924 7420 203980 8148
rect 203924 7354 203980 7364
rect 204148 8930 204204 8942
rect 204148 8878 204150 8930
rect 204202 8878 204204 8930
rect 203196 7140 203308 7196
rect 202580 6690 202636 6702
rect 202580 6638 202582 6690
rect 202634 6638 202636 6690
rect 202580 6636 202636 6638
rect 202580 6570 202636 6580
rect 203084 6636 203140 6646
rect 203084 6542 203140 6580
rect 203196 6578 203252 7140
rect 203196 6526 203198 6578
rect 203250 6526 203252 6578
rect 203196 5964 203252 6526
rect 203644 6524 203700 6534
rect 203140 5908 203252 5964
rect 203588 6522 203700 6524
rect 203588 6470 203646 6522
rect 203698 6470 203700 6522
rect 203588 6458 203700 6470
rect 203140 5628 203196 5908
rect 203140 5562 203196 5572
rect 202468 2986 202524 2996
rect 203588 2268 203644 6458
rect 203924 6300 203980 6310
rect 203924 5906 203980 6244
rect 203924 5854 203926 5906
rect 203978 5854 203980 5906
rect 203924 5842 203980 5854
rect 203756 4954 203812 4966
rect 203756 4902 203758 4954
rect 203810 4902 203812 4954
rect 203756 4732 203812 4902
rect 203812 4676 203868 4732
rect 203756 4666 203868 4676
rect 203812 4172 203868 4666
rect 203812 4106 203868 4116
rect 203588 2202 203644 2212
rect 201908 1866 201964 1876
rect 201684 1306 201740 1316
rect 201908 1484 201964 1494
rect 201572 970 201628 980
rect 201908 800 201964 1428
rect 202580 1146 202636 1158
rect 202580 1094 202582 1146
rect 202634 1094 202636 1146
rect 202580 800 202636 1094
rect 203028 924 203084 934
rect 203812 924 203868 934
rect 203084 868 203196 924
rect 203028 858 203084 868
rect 203140 800 203196 868
rect 203812 800 203868 868
rect 204148 812 204204 8878
rect 204260 8326 204316 10052
rect 204484 9772 204540 9782
rect 204484 9678 204540 9716
rect 204596 8427 204652 11732
rect 204820 9994 204876 12852
rect 205044 12236 205100 14200
rect 205044 12170 205100 12180
rect 205268 13020 205324 13030
rect 204820 9942 204822 9994
rect 204874 9942 204876 9994
rect 204820 9930 204876 9942
rect 204484 8371 204652 8427
rect 204708 9660 204764 9670
rect 204260 8314 204372 8326
rect 204260 8262 204318 8314
rect 204370 8262 204372 8314
rect 204260 8260 204372 8262
rect 204316 8250 204372 8260
rect 204484 7306 204540 8371
rect 204484 7254 204486 7306
rect 204538 7254 204540 7306
rect 204484 7242 204540 7254
rect 204708 6076 204764 9604
rect 205268 6746 205324 12964
rect 205716 11900 205772 14200
rect 205716 11834 205772 11844
rect 205940 12124 205996 12134
rect 205828 9660 205884 9670
rect 205828 9566 205884 9604
rect 205940 8314 205996 12068
rect 206500 12012 206556 14200
rect 207172 12348 207228 14200
rect 207172 12282 207228 12292
rect 206500 11946 206556 11956
rect 207732 11900 207788 11910
rect 206164 11788 206220 11798
rect 206164 9994 206220 11732
rect 206164 9942 206166 9994
rect 206218 9942 206220 9994
rect 206164 9930 206220 9942
rect 206388 11114 206444 11126
rect 206388 11062 206390 11114
rect 206442 11062 206444 11114
rect 206388 8427 206444 11062
rect 206500 9212 206556 9222
rect 206500 9042 206556 9156
rect 206500 8990 206502 9042
rect 206554 8990 206556 9042
rect 206500 8978 206556 8990
rect 207508 9154 207564 9166
rect 207508 9102 207510 9154
rect 207562 9102 207564 9154
rect 206724 8874 206780 8886
rect 206724 8822 206726 8874
rect 206778 8822 206780 8874
rect 206388 8371 206556 8427
rect 205940 8262 205942 8314
rect 205994 8262 205996 8314
rect 205940 8250 205996 8262
rect 206052 8092 206108 8102
rect 206052 7532 206108 8036
rect 206052 7474 206108 7476
rect 206052 7422 206054 7474
rect 206106 7422 206108 7474
rect 206052 7400 206108 7422
rect 205268 6694 205270 6746
rect 205322 6694 205324 6746
rect 205268 6682 205324 6694
rect 206500 6690 206556 8371
rect 206724 8316 206780 8822
rect 206724 8250 206780 8260
rect 206948 8258 207004 8270
rect 206948 8206 206950 8258
rect 207002 8206 207004 8258
rect 206948 8204 207004 8206
rect 206948 8138 207004 8148
rect 207508 7756 207564 9102
rect 207508 7690 207564 7700
rect 207732 7644 207788 11844
rect 207956 11788 208012 14200
rect 208628 13020 208684 14200
rect 208628 12954 208684 12964
rect 209300 12458 209356 12470
rect 209300 12406 209302 12458
rect 209354 12406 209356 12458
rect 207956 11722 208012 11732
rect 208852 11788 208908 11798
rect 208180 10108 208236 10118
rect 208180 9938 208236 10052
rect 208180 9886 208182 9938
rect 208234 9886 208236 9938
rect 208180 9874 208236 9886
rect 208068 9826 208124 9838
rect 208068 9774 208070 9826
rect 208122 9774 208124 9826
rect 208068 8316 208124 9774
rect 208516 9772 208572 9782
rect 208068 8260 208460 8316
rect 206500 6638 206502 6690
rect 206554 6638 206556 6690
rect 206500 6636 206556 6638
rect 206500 6570 206556 6580
rect 207620 7588 207788 7644
rect 207620 6086 207676 7588
rect 207732 7470 207788 7482
rect 207732 7418 207734 7470
rect 207786 7418 207788 7470
rect 207732 7196 207788 7418
rect 208404 7362 208460 8260
rect 208404 7310 208406 7362
rect 208458 7310 208460 7362
rect 208404 7298 208460 7310
rect 207732 7130 207788 7140
rect 204596 6020 204764 6076
rect 207564 6074 207676 6086
rect 207564 6022 207566 6074
rect 207618 6022 207676 6074
rect 207564 6020 207676 6022
rect 207956 6690 208012 6702
rect 207956 6638 207958 6690
rect 208010 6638 208012 6690
rect 204596 5078 204652 6020
rect 207564 6010 207620 6020
rect 205492 5964 205548 5984
rect 204764 5906 204820 5918
rect 204764 5854 204766 5906
rect 204818 5854 204820 5906
rect 204764 5290 204820 5854
rect 204764 5238 204766 5290
rect 204818 5238 204820 5290
rect 204764 5226 204820 5238
rect 205492 5906 205548 5908
rect 205492 5854 205494 5906
rect 205546 5854 205548 5906
rect 205492 5180 205548 5854
rect 205828 5794 205884 5806
rect 205828 5742 205830 5794
rect 205882 5742 205884 5794
rect 205492 5114 205548 5124
rect 205604 5122 205660 5134
rect 204596 5066 204708 5078
rect 204596 5014 204654 5066
rect 204706 5014 204708 5066
rect 204596 5002 204708 5014
rect 205604 5070 205606 5122
rect 205658 5070 205660 5122
rect 205604 5068 205660 5070
rect 204596 4620 204652 5002
rect 204596 2490 204652 4564
rect 205604 4508 205660 5012
rect 205604 4442 205660 4452
rect 205716 5010 205772 5022
rect 205716 4958 205718 5010
rect 205770 4958 205772 5010
rect 205716 3724 205772 4958
rect 205716 3658 205772 3668
rect 204596 2438 204598 2490
rect 204650 2438 204652 2490
rect 204596 2426 204652 2438
rect 196196 746 196252 758
rect 196392 0 196504 800
rect 197064 0 197176 800
rect 197624 0 197736 800
rect 198296 0 198408 800
rect 198856 0 198968 800
rect 199416 0 199528 800
rect 200088 0 200200 800
rect 200648 0 200760 800
rect 201320 0 201432 800
rect 201880 0 201992 800
rect 202552 0 202664 800
rect 203112 0 203224 800
rect 203784 0 203896 800
rect 204372 1596 204428 1606
rect 204372 800 204428 1540
rect 205828 1372 205884 5742
rect 207956 5180 208012 6638
rect 208516 5180 208572 9716
rect 208628 8258 208684 8270
rect 208628 8206 208630 8258
rect 208682 8206 208684 8258
rect 208628 5292 208684 8206
rect 208740 5740 208796 5750
rect 208852 5740 208908 11732
rect 209300 8427 209356 12406
rect 209412 11900 209468 14200
rect 209412 11834 209468 11844
rect 209860 13692 209916 13702
rect 209524 9602 209580 9614
rect 209524 9550 209526 9602
rect 209578 9550 209580 9602
rect 209524 9042 209580 9550
rect 209860 9154 209916 13636
rect 210084 12908 210140 14200
rect 210084 12842 210140 12852
rect 210420 13690 210476 13702
rect 210420 13638 210422 13690
rect 210474 13638 210476 13690
rect 209860 9102 209862 9154
rect 209914 9102 209916 9154
rect 209860 9090 209916 9102
rect 209524 8990 209526 9042
rect 209578 8990 209580 9042
rect 209524 8978 209580 8990
rect 209300 8371 209468 8427
rect 209188 8316 209244 8326
rect 209188 8258 209244 8260
rect 209188 8206 209190 8258
rect 209242 8206 209244 8258
rect 209188 8194 209244 8206
rect 209412 7532 209468 8371
rect 209860 8370 209916 8382
rect 209860 8318 209862 8370
rect 209914 8318 209916 8370
rect 209860 8316 209916 8318
rect 209860 8250 209916 8260
rect 209860 7644 209916 7654
rect 208740 5738 208908 5740
rect 208740 5686 208742 5738
rect 208794 5686 208908 5738
rect 208740 5684 208908 5686
rect 209300 7476 209468 7532
rect 209636 7586 209692 7598
rect 209636 7534 209638 7586
rect 209690 7534 209692 7586
rect 208740 5674 208796 5684
rect 208628 5236 208796 5292
rect 207956 5124 208236 5180
rect 208516 5124 208628 5180
rect 207788 5068 207844 5078
rect 207732 5012 207788 5068
rect 207732 4936 207844 5012
rect 207900 4956 207956 4966
rect 207732 3162 207788 4936
rect 208180 4956 208236 5124
rect 208572 5066 208628 5124
rect 208572 5014 208574 5066
rect 208626 5014 208628 5066
rect 208460 4956 208516 4966
rect 208180 4954 208516 4956
rect 208180 4902 208462 4954
rect 208514 4902 208516 4954
rect 208180 4900 208516 4902
rect 207900 4862 207956 4900
rect 208460 4890 208516 4900
rect 208572 4732 208628 5014
rect 208740 4956 208796 5236
rect 208740 4890 208796 4900
rect 208572 4666 208628 4676
rect 207732 3110 207734 3162
rect 207786 3110 207788 3162
rect 207732 3098 207788 3110
rect 205828 1306 205884 1316
rect 205604 924 205660 934
rect 206836 924 206892 934
rect 204708 868 204988 924
rect 204148 746 204204 756
rect 204344 0 204456 800
rect 204708 364 204764 868
rect 204932 800 204988 868
rect 205604 800 205660 868
rect 205940 868 206220 924
rect 204708 298 204764 308
rect 204904 0 205016 800
rect 205576 0 205688 800
rect 205940 476 205996 868
rect 206164 800 206220 868
rect 206836 800 206892 868
rect 207172 868 207452 924
rect 205828 420 205996 476
rect 205828 252 205884 420
rect 205828 186 205884 196
rect 206136 0 206248 800
rect 206808 0 206920 800
rect 207172 588 207228 868
rect 207396 800 207452 868
rect 207844 868 208124 924
rect 207060 532 207228 588
rect 207060 362 207116 532
rect 207060 310 207062 362
rect 207114 310 207116 362
rect 207060 298 207116 310
rect 207368 0 207480 800
rect 207844 364 207900 868
rect 208068 800 208124 868
rect 208404 868 208684 924
rect 207620 308 207900 364
rect 207620 140 207676 308
rect 207620 74 207676 84
rect 208040 0 208152 800
rect 208404 364 208460 868
rect 208628 800 208684 868
rect 209300 800 209356 7476
rect 209636 6076 209692 7534
rect 209860 7474 209916 7588
rect 209860 7422 209862 7474
rect 209914 7422 209916 7474
rect 209860 7410 209916 7422
rect 209860 6690 209916 6702
rect 209860 6638 209862 6690
rect 209914 6638 209916 6690
rect 209636 6010 209692 6020
rect 209748 6578 209804 6590
rect 209748 6526 209750 6578
rect 209802 6526 209804 6578
rect 209636 5010 209692 5022
rect 209636 4958 209638 5010
rect 209690 4958 209692 5010
rect 209636 3836 209692 4958
rect 209636 3770 209692 3780
rect 209748 1484 209804 6526
rect 209860 6188 209916 6638
rect 209860 6122 209916 6132
rect 209860 5404 209916 5414
rect 209860 4844 209916 5348
rect 209860 4778 209916 4788
rect 209748 1418 209804 1428
rect 209860 1260 209916 1270
rect 209860 800 209916 1204
rect 210420 800 210476 13638
rect 210868 11788 210924 14200
rect 210868 11722 210924 11732
rect 210980 12348 211036 12358
rect 210980 11340 211036 12292
rect 211540 11788 211596 14200
rect 211652 13356 211708 13366
rect 211652 13262 211708 13300
rect 211540 11722 211596 11732
rect 211764 12460 211820 12470
rect 210868 11284 211036 11340
rect 210756 9772 210812 9782
rect 210756 9714 210812 9716
rect 210756 9662 210758 9714
rect 210810 9662 210812 9714
rect 210756 9650 210812 9662
rect 210868 7642 210924 11284
rect 211428 10442 211484 10454
rect 211428 10390 211430 10442
rect 211482 10390 211484 10442
rect 210980 9884 211036 9894
rect 210980 9826 211036 9828
rect 210980 9774 210982 9826
rect 211034 9774 211036 9826
rect 210980 9762 211036 9774
rect 211092 9154 211148 9166
rect 211092 9102 211094 9154
rect 211146 9102 211148 9154
rect 211092 8427 211148 9102
rect 210868 7590 210870 7642
rect 210922 7590 210924 7642
rect 210868 7578 210924 7590
rect 210980 8371 211148 8427
rect 211204 9100 211260 9110
rect 210980 7868 211036 8371
rect 211204 8326 211260 9044
rect 211428 9100 211484 10390
rect 211764 10220 211820 12404
rect 212324 12012 212380 14200
rect 211428 9042 211484 9044
rect 211428 8990 211430 9042
rect 211482 8990 211484 9042
rect 211428 8978 211484 8990
rect 211540 9658 211596 9670
rect 211540 9606 211542 9658
rect 211594 9606 211596 9658
rect 211204 8314 211316 8326
rect 211204 8262 211262 8314
rect 211314 8262 211316 8314
rect 211204 8260 211316 8262
rect 211260 8250 211316 8260
rect 210532 7530 210588 7542
rect 210532 7478 210534 7530
rect 210586 7478 210588 7530
rect 210532 5068 210588 7478
rect 210980 7420 211036 7812
rect 210980 7354 211036 7364
rect 211260 7420 211316 7430
rect 211260 7326 211316 7364
rect 210700 7196 210756 7206
rect 210700 6858 210756 7140
rect 210700 6806 210702 6858
rect 210754 6806 210756 6858
rect 210700 6794 210756 6806
rect 211540 6692 211596 9606
rect 211764 7654 211820 10164
rect 211876 11956 212380 12012
rect 212772 13914 212828 13926
rect 212772 13862 212774 13914
rect 212826 13862 212828 13914
rect 211876 9994 211932 11956
rect 211876 9942 211878 9994
rect 211930 9942 211932 9994
rect 211876 9930 211932 9942
rect 212268 9660 212324 9670
rect 212268 9566 212324 9604
rect 212660 9436 212716 9446
rect 211988 8930 212044 8942
rect 211988 8878 211990 8930
rect 212042 8878 212044 8930
rect 211708 7642 211820 7654
rect 211708 7590 211710 7642
rect 211762 7590 211820 7642
rect 211708 7588 211820 7590
rect 211876 8092 211932 8102
rect 211708 7578 211764 7588
rect 211372 6636 211596 6692
rect 211876 6748 211932 8036
rect 211876 6682 211932 6692
rect 210812 6578 210868 6590
rect 210812 6526 210814 6578
rect 210866 6526 210868 6578
rect 210812 6300 210868 6526
rect 211372 6578 211428 6636
rect 211372 6526 211374 6578
rect 211426 6526 211428 6578
rect 211372 6524 211428 6526
rect 210532 5002 210588 5012
rect 210756 6244 210868 6300
rect 211316 6468 211428 6524
rect 211484 6524 211540 6534
rect 211484 6522 211820 6524
rect 211484 6470 211486 6522
rect 211538 6470 211820 6522
rect 211484 6468 211820 6470
rect 210756 5516 210812 6244
rect 210980 5906 211036 5918
rect 210980 5854 210982 5906
rect 211034 5854 211036 5906
rect 210980 5852 211036 5854
rect 210980 5786 211036 5796
rect 210756 2044 210812 5460
rect 211316 5404 211372 6468
rect 211484 6458 211540 6468
rect 211764 5964 211820 6468
rect 211988 6188 212044 8878
rect 212212 8652 212268 8662
rect 212212 8316 212268 8596
rect 212660 8316 212716 9380
rect 212772 9212 212828 13862
rect 212996 12124 213052 14200
rect 213780 12460 213836 14200
rect 213780 12394 213836 12404
rect 214452 12348 214508 14200
rect 214452 12282 214508 12292
rect 212996 12058 213052 12068
rect 215236 12124 215292 14200
rect 215236 12058 215292 12068
rect 215684 12348 215740 12358
rect 213668 12010 213724 12022
rect 213668 11958 213670 12010
rect 213722 11958 213724 12010
rect 213108 11900 213164 11910
rect 212772 9080 212828 9156
rect 212884 11788 212940 11798
rect 212156 8260 212268 8316
rect 212604 8260 212716 8316
rect 212156 7642 212212 8260
rect 212268 8092 212324 8102
rect 212268 7998 212324 8036
rect 212156 7590 212158 7642
rect 212210 7590 212212 7642
rect 212156 7578 212212 7590
rect 212604 7642 212660 8260
rect 212716 8092 212772 8102
rect 212716 7868 212772 8036
rect 212716 7802 212772 7812
rect 212604 7590 212606 7642
rect 212658 7590 212660 7642
rect 212604 7578 212660 7590
rect 212324 7420 212380 7430
rect 212324 6692 212380 7364
rect 212324 6636 212436 6692
rect 212268 6524 212324 6534
rect 212268 6430 212324 6468
rect 211988 6122 212044 6132
rect 212380 6074 212436 6636
rect 212716 6524 212772 6534
rect 212884 6524 212940 11732
rect 212996 9324 213052 9334
rect 212996 7654 213052 9268
rect 213108 9210 213164 11844
rect 213444 9660 213500 9670
rect 213108 9158 213110 9210
rect 213162 9158 213164 9210
rect 213108 9146 213164 9158
rect 213332 9658 213500 9660
rect 213332 9606 213446 9658
rect 213498 9606 213500 9658
rect 213332 9604 213500 9606
rect 213164 8090 213220 8102
rect 213164 8038 213166 8090
rect 213218 8038 213220 8090
rect 212996 7642 213108 7654
rect 212996 7590 213054 7642
rect 213106 7590 213108 7642
rect 212996 7588 213108 7590
rect 213052 7578 213108 7588
rect 213164 7420 213220 8038
rect 213108 7364 213220 7420
rect 213108 6860 213164 7364
rect 213108 6794 213164 6804
rect 213164 6524 213220 6534
rect 212380 6022 212382 6074
rect 212434 6022 212436 6074
rect 212380 6010 212436 6022
rect 212660 6522 212940 6524
rect 212660 6470 212718 6522
rect 212770 6470 212940 6522
rect 212660 6468 212940 6470
rect 213108 6522 213220 6524
rect 213108 6470 213166 6522
rect 213218 6470 213220 6522
rect 212660 6458 212772 6468
rect 213108 6458 213220 6470
rect 213332 6524 213388 9604
rect 213444 9594 213500 9604
rect 213500 8986 213556 8998
rect 213500 8934 213502 8986
rect 213554 8934 213556 8986
rect 213500 8652 213556 8934
rect 213500 8586 213556 8596
rect 213668 8427 213724 11958
rect 213780 12012 213836 12022
rect 213780 9994 213836 11956
rect 213780 9942 213782 9994
rect 213834 9942 213836 9994
rect 213780 9930 213836 9942
rect 215012 11788 215068 11798
rect 215012 9828 215068 11732
rect 214900 9772 215068 9828
rect 214172 9660 214228 9670
rect 214116 9658 214228 9660
rect 214116 9606 214174 9658
rect 214226 9606 214228 9658
rect 214116 9594 214228 9606
rect 214620 9658 214676 9670
rect 214620 9606 214622 9658
rect 214674 9606 214676 9658
rect 213948 8988 214004 8998
rect 213948 8894 214004 8932
rect 214116 8876 214172 9594
rect 214620 9548 214676 9606
rect 214620 9482 214676 9492
rect 214900 9436 214956 9772
rect 215068 9660 215124 9670
rect 215068 9658 215292 9660
rect 215068 9606 215070 9658
rect 215122 9606 215292 9658
rect 215068 9604 215292 9606
rect 215068 9594 215124 9604
rect 214900 9380 215180 9436
rect 214788 9324 214844 9334
rect 214788 9222 214844 9268
rect 214788 9210 214900 9222
rect 214788 9158 214846 9210
rect 214898 9158 214900 9210
rect 214788 9156 214900 9158
rect 214844 9146 214900 9156
rect 214116 8810 214172 8820
rect 214396 8986 214452 8998
rect 214396 8934 214398 8986
rect 214450 8934 214452 8986
rect 214396 8540 214452 8934
rect 215124 8764 215180 9380
rect 215236 9324 215292 9604
rect 215516 9658 215572 9670
rect 215516 9606 215518 9658
rect 215570 9606 215572 9658
rect 215516 9436 215572 9606
rect 215516 9370 215572 9380
rect 215236 9258 215292 9268
rect 215292 8988 215348 8998
rect 215572 8988 215628 8998
rect 215292 8986 215404 8988
rect 215292 8934 215294 8986
rect 215346 8934 215404 8986
rect 215292 8922 215404 8934
rect 215124 8708 215292 8764
rect 214396 8474 214452 8484
rect 215124 8540 215180 8550
rect 215124 8427 215180 8484
rect 213668 8371 213836 8427
rect 213612 8090 213668 8102
rect 213612 8038 213614 8090
rect 213666 8038 213668 8090
rect 213612 7980 213668 8038
rect 213612 7914 213668 7924
rect 213500 7420 213556 7430
rect 213332 6458 213388 6468
rect 213444 7418 213556 7420
rect 213444 7366 213502 7418
rect 213554 7366 213556 7418
rect 213444 7354 213556 7366
rect 211764 5908 211876 5964
rect 211820 5906 211876 5908
rect 211820 5854 211822 5906
rect 211874 5854 211876 5906
rect 211820 5842 211876 5854
rect 211316 5338 211372 5348
rect 211092 5122 211148 5134
rect 211092 5070 211094 5122
rect 211146 5070 211148 5122
rect 211092 4844 211148 5070
rect 211596 4956 211652 4966
rect 211596 4862 211652 4900
rect 212044 4956 212100 4966
rect 212044 4862 212100 4900
rect 212492 4954 212548 4966
rect 212492 4902 212494 4954
rect 212546 4902 212548 4954
rect 211092 4778 211148 4788
rect 212492 4396 212548 4902
rect 212492 4330 212548 4340
rect 212660 3388 212716 6458
rect 212828 5850 212884 5862
rect 212828 5798 212830 5850
rect 212882 5798 212884 5850
rect 212828 5740 212884 5798
rect 212828 5674 212884 5684
rect 213108 4172 213164 6458
rect 213276 6300 213332 6310
rect 213276 6074 213332 6244
rect 213276 6022 213278 6074
rect 213330 6022 213332 6074
rect 213276 6010 213332 6022
rect 213444 5628 213500 7354
rect 213612 6522 213668 6534
rect 213612 6470 213614 6522
rect 213666 6470 213668 6522
rect 213612 6300 213668 6470
rect 213612 6234 213668 6244
rect 213780 6076 213836 8371
rect 215068 8371 215180 8427
rect 215068 8314 215124 8371
rect 215068 8262 215070 8314
rect 215122 8262 215124 8314
rect 215068 8250 215124 8262
rect 214508 8204 214564 8214
rect 214508 8110 214564 8148
rect 214060 8092 214116 8102
rect 214060 8090 214172 8092
rect 214060 8038 214062 8090
rect 214114 8038 214172 8090
rect 214060 8026 214172 8038
rect 213948 7532 214004 7542
rect 213948 7438 214004 7476
rect 214116 7084 214172 8026
rect 214396 7756 214452 7766
rect 214396 7420 214452 7700
rect 215236 7654 215292 8708
rect 215348 7868 215404 8922
rect 215572 8427 215628 8932
rect 215684 8540 215740 12292
rect 215908 12236 215964 14200
rect 215908 12170 215964 12180
rect 216580 12124 216636 12134
rect 216580 9884 216636 12068
rect 216692 12012 216748 14200
rect 216692 11946 216748 11956
rect 217364 11900 217420 14200
rect 218148 12348 218204 14200
rect 218148 12282 218204 12292
rect 217364 11834 217420 11844
rect 218820 11788 218876 14200
rect 219604 12124 219660 14200
rect 219604 12058 219660 12068
rect 218820 11722 218876 11732
rect 215964 9660 216020 9670
rect 216412 9660 216468 9670
rect 215964 9658 216188 9660
rect 215964 9606 215966 9658
rect 216018 9606 216188 9658
rect 215964 9604 216188 9606
rect 215964 9594 216020 9604
rect 215684 8474 215740 8484
rect 216020 9324 216076 9334
rect 215516 8371 215628 8427
rect 215516 8314 215572 8371
rect 215516 8262 215518 8314
rect 215570 8262 215572 8314
rect 215516 8250 215572 8262
rect 215852 8092 215908 8102
rect 215796 8090 215908 8092
rect 215796 8038 215854 8090
rect 215906 8038 215908 8090
rect 215796 8026 215908 8038
rect 215348 7812 215516 7868
rect 215236 7644 215348 7654
rect 215236 7588 215292 7644
rect 215292 7550 215348 7588
rect 214844 7420 214900 7430
rect 214396 7326 214452 7364
rect 214788 7418 214900 7420
rect 214788 7366 214846 7418
rect 214898 7366 214900 7418
rect 214788 7354 214900 7366
rect 214116 7018 214172 7028
rect 214508 6636 214564 6646
rect 214508 6542 214564 6580
rect 213444 5562 213500 5572
rect 213556 6020 213836 6076
rect 213892 6524 213948 6534
rect 213276 4956 213332 4966
rect 213220 4954 213332 4956
rect 213220 4902 213278 4954
rect 213330 4902 213332 4954
rect 213220 4890 213332 4902
rect 213220 4284 213276 4890
rect 213220 4218 213276 4228
rect 213108 4106 213164 4116
rect 212660 3322 212716 3332
rect 210756 1978 210812 1988
rect 211652 1596 211708 1606
rect 211092 1372 211148 1382
rect 211092 800 211148 1316
rect 211652 800 211708 1540
rect 212324 1036 212380 1046
rect 212324 800 212380 980
rect 212884 924 212940 934
rect 212884 800 212940 868
rect 213556 800 213612 6020
rect 213724 5850 213780 5862
rect 213724 5798 213726 5850
rect 213778 5798 213780 5850
rect 213724 5628 213780 5798
rect 213724 5562 213780 5572
rect 213892 5516 213948 6468
rect 214060 6522 214116 6534
rect 214060 6470 214062 6522
rect 214114 6470 214116 6522
rect 214060 6412 214116 6470
rect 214060 6346 214116 6356
rect 214172 5964 214228 5974
rect 214172 5870 214228 5908
rect 214620 5852 214676 5862
rect 214620 5758 214676 5796
rect 213892 5450 213948 5460
rect 213724 4954 213780 4966
rect 213724 4902 213726 4954
rect 213778 4902 213780 4954
rect 213724 4620 213780 4902
rect 213724 4554 213780 4564
rect 214172 4954 214228 4966
rect 214172 4902 214174 4954
rect 214226 4902 214228 4954
rect 214172 4508 214228 4902
rect 214620 4956 214676 4966
rect 214788 4956 214844 7354
rect 215460 6692 215516 7812
rect 215236 6636 215516 6692
rect 214956 6524 215012 6534
rect 214676 4900 214844 4956
rect 214900 6522 215012 6524
rect 214900 6470 214958 6522
rect 215010 6470 215012 6522
rect 214900 6458 215012 6470
rect 214900 6076 214956 6458
rect 214620 4862 214676 4900
rect 214172 4442 214228 4452
rect 214900 3836 214956 6020
rect 215068 5850 215124 5862
rect 215068 5798 215070 5850
rect 215122 5798 215124 5850
rect 215068 5404 215124 5798
rect 215068 5338 215124 5348
rect 215068 4956 215124 4966
rect 215068 4732 215124 4900
rect 215068 4666 215124 4676
rect 215236 4620 215292 6636
rect 215404 6524 215460 6534
rect 215404 6430 215460 6468
rect 215796 6524 215852 8026
rect 215796 6458 215852 6468
rect 216020 6300 216076 9268
rect 216020 6234 216076 6244
rect 215516 4954 215572 4966
rect 215516 4902 215518 4954
rect 215570 4902 215572 4954
rect 215516 4844 215572 4902
rect 216132 4956 216188 9604
rect 216412 9658 216524 9660
rect 216412 9606 216414 9658
rect 216466 9606 216524 9658
rect 216412 9594 216524 9606
rect 216300 9100 216356 9110
rect 216300 9006 216356 9044
rect 216300 8092 216356 8102
rect 216300 7998 216356 8036
rect 216468 5404 216524 9594
rect 216580 8988 216636 9828
rect 217308 9772 217364 9782
rect 217364 9716 217420 9772
rect 217308 9678 217420 9716
rect 216748 9212 216804 9222
rect 216748 9118 216804 9156
rect 216580 8922 216636 8932
rect 217364 6300 217420 9678
rect 217364 6234 217420 6244
rect 216468 5338 216524 5348
rect 216132 4890 216188 4900
rect 215516 4778 215572 4788
rect 215236 4554 215292 4564
rect 214900 3770 214956 3780
rect 219044 1484 219100 1494
rect 214116 1148 214172 1158
rect 214116 800 214172 1092
rect 217140 924 217196 934
rect 214564 868 214844 924
rect 208292 308 208460 364
rect 208292 138 208348 308
rect 208292 86 208294 138
rect 208346 86 208348 138
rect 208292 74 208348 86
rect 208600 0 208712 800
rect 209272 0 209384 800
rect 209832 0 209944 800
rect 210392 0 210504 800
rect 211064 0 211176 800
rect 211624 0 211736 800
rect 212296 0 212408 800
rect 212856 0 212968 800
rect 213528 0 213640 800
rect 214088 0 214200 800
rect 214564 700 214620 868
rect 214788 800 214844 868
rect 215124 868 215404 924
rect 214340 644 214620 700
rect 214340 588 214396 644
rect 214340 522 214396 532
rect 214760 0 214872 800
rect 215124 364 215180 868
rect 215348 800 215404 868
rect 215684 868 215964 924
rect 215684 810 215740 868
rect 215012 308 215180 364
rect 215012 250 215068 308
rect 215012 198 215014 250
rect 215066 198 215068 250
rect 215012 186 215068 198
rect 215320 0 215432 800
rect 215684 758 215686 810
rect 215738 758 215740 810
rect 215908 800 215964 868
rect 216356 868 216636 924
rect 215684 746 215740 758
rect 215880 0 215992 800
rect 216356 588 216412 868
rect 216580 800 216636 868
rect 217140 800 217196 868
rect 217588 868 217868 924
rect 216132 532 216412 588
rect 216132 474 216188 532
rect 216132 422 216134 474
rect 216186 422 216188 474
rect 216132 410 216188 422
rect 216552 0 216664 800
rect 217112 0 217224 800
rect 217588 588 217644 868
rect 217812 800 217868 868
rect 218372 922 218428 934
rect 218372 870 218374 922
rect 218426 870 218428 922
rect 218372 800 218428 870
rect 219044 800 219100 1428
rect 219604 1148 219660 1158
rect 219604 800 219660 1092
rect 217364 532 217644 588
rect 217364 476 217420 532
rect 217364 410 217420 420
rect 217784 0 217896 800
rect 218344 0 218456 800
rect 219016 0 219128 800
rect 219576 0 219688 800
<< via2 >>
rect 308 13300 364 13356
rect 980 13188 1036 13244
rect 3892 13076 3948 13132
rect 3220 12964 3276 13020
rect 2436 12292 2492 12348
rect 7700 14084 7756 14140
rect 16660 14420 16716 14476
rect 10500 13524 10556 13580
rect 10612 13300 10668 13356
rect 6132 12852 6188 12908
rect 9828 12964 9884 13020
rect 6692 12404 6748 12460
rect 84 7924 140 7980
rect 9716 12292 9772 12348
rect 6692 9716 6748 9772
rect 8316 9770 8372 9772
rect 8316 9718 8318 9770
rect 8318 9718 8370 9770
rect 8370 9718 8372 9770
rect 8316 9716 8372 9718
rect 8876 9658 8932 9660
rect 8876 9606 8878 9658
rect 8878 9606 8930 9658
rect 8930 9606 8932 9658
rect 8876 9604 8932 9606
rect 10164 9658 10220 9660
rect 10164 9606 10166 9658
rect 10166 9606 10218 9658
rect 10218 9606 10220 9658
rect 10164 9604 10220 9606
rect 10724 13188 10780 13244
rect 11620 13076 11676 13132
rect 10836 10948 10892 11004
rect 8988 9098 9044 9100
rect 8988 9046 8990 9098
rect 8990 9046 9042 9098
rect 9042 9046 9044 9098
rect 8988 9044 9044 9046
rect 10052 9098 10108 9100
rect 10052 9046 10054 9098
rect 10054 9046 10106 9098
rect 10106 9046 10108 9098
rect 10052 9044 10108 9046
rect 9716 8372 9772 8428
rect 8932 7588 8988 7644
rect 9548 7642 9604 7644
rect 9548 7590 9550 7642
rect 9550 7590 9602 7642
rect 9602 7590 9604 7642
rect 9548 7588 9604 7590
rect 7924 7252 7980 7308
rect 8764 7252 8820 7308
rect 10276 8314 10332 8316
rect 10276 8262 10278 8314
rect 10278 8262 10330 8314
rect 10330 8262 10332 8314
rect 10276 8260 10332 8262
rect 4452 6356 4508 6412
rect 3780 4788 3836 4844
rect 756 868 812 924
rect 1316 868 1372 924
rect 1988 868 2044 924
rect 2548 868 2604 924
rect 3220 868 3276 924
rect 10332 7418 10388 7420
rect 10332 7366 10334 7418
rect 10334 7366 10386 7418
rect 10386 7366 10388 7418
rect 10332 7364 10388 7366
rect 8820 6020 8876 6076
rect 5012 4676 5068 4732
rect 8708 4900 8764 4956
rect 8260 1540 8316 1596
rect 8708 3332 8764 3388
rect 8148 1428 8204 1484
rect 8036 1316 8092 1372
rect 532 196 588 252
rect 6580 532 6636 588
rect 7812 308 7868 364
rect 9548 6074 9604 6076
rect 9548 6022 9550 6074
rect 9550 6022 9602 6074
rect 9602 6022 9604 6074
rect 9548 6020 9604 6022
rect 9548 4954 9604 4956
rect 9548 4902 9550 4954
rect 9550 4902 9602 4954
rect 9602 4902 9604 4954
rect 9548 4900 9604 4902
rect 12628 13748 12684 13804
rect 11956 12628 12012 12684
rect 14868 13972 14924 14028
rect 14084 13860 14140 13916
rect 23380 14756 23436 14812
rect 17108 14084 17164 14140
rect 17780 13972 17836 14028
rect 19236 13300 19292 13356
rect 18452 13188 18508 13244
rect 15540 13076 15596 13132
rect 13412 12404 13468 12460
rect 18116 11732 18172 11788
rect 14420 11060 14476 11116
rect 13076 10836 13132 10892
rect 11060 9770 11116 9772
rect 11060 9718 11062 9770
rect 11062 9718 11114 9770
rect 11114 9718 11116 9770
rect 11060 9716 11116 9718
rect 11956 9380 12012 9436
rect 12572 9380 12628 9436
rect 13748 9828 13804 9884
rect 13636 8820 13692 8876
rect 12852 8262 12908 8316
rect 12852 8260 12854 8262
rect 12854 8260 12906 8262
rect 12906 8260 12908 8262
rect 13580 8314 13636 8316
rect 13580 8262 13582 8314
rect 13582 8262 13634 8314
rect 13634 8262 13636 8314
rect 13580 8260 13636 8262
rect 11620 8036 11676 8092
rect 10948 7364 11004 7420
rect 12740 7476 12796 7532
rect 14084 8932 14140 8988
rect 13916 8090 13972 8092
rect 13916 8038 13918 8090
rect 13918 8038 13970 8090
rect 13970 8038 13972 8090
rect 13916 8036 13972 8038
rect 13748 7476 13804 7532
rect 10668 6074 10724 6076
rect 10668 6022 10670 6074
rect 10670 6022 10722 6074
rect 10722 6022 10724 6074
rect 10668 6020 10724 6022
rect 10556 4954 10612 4956
rect 10556 4902 10558 4954
rect 10558 4902 10610 4954
rect 10610 4902 10612 4954
rect 10556 4900 10612 4902
rect 11172 3332 11228 3388
rect 10276 2548 10332 2604
rect 9940 1540 9996 1596
rect 9268 1204 9324 1260
rect 11060 1540 11116 1596
rect 10500 1428 10556 1484
rect 10164 1146 10220 1148
rect 10164 1094 10166 1146
rect 10166 1094 10218 1146
rect 10218 1094 10220 1146
rect 10164 1092 10220 1094
rect 12852 6468 12908 6524
rect 14028 6522 14084 6524
rect 14028 6470 14030 6522
rect 14030 6470 14082 6522
rect 14082 6470 14084 6522
rect 14028 6468 14084 6470
rect 12740 6020 12796 6076
rect 11620 4900 11676 4956
rect 11508 4564 11564 4620
rect 11396 1204 11452 1260
rect 11732 1428 11788 1484
rect 14868 10612 14924 10668
rect 16212 10052 16268 10108
rect 15596 9716 15652 9772
rect 15092 9156 15148 9212
rect 15596 9210 15652 9212
rect 15596 9158 15598 9210
rect 15598 9158 15650 9210
rect 15650 9158 15652 9210
rect 15596 9156 15652 9158
rect 16044 8986 16100 8988
rect 16044 8934 16046 8986
rect 16046 8934 16098 8986
rect 16098 8934 16100 8986
rect 16044 8932 16100 8934
rect 15876 7364 15932 7420
rect 17780 9210 17836 9212
rect 17780 9158 17782 9210
rect 17782 9158 17834 9210
rect 17834 9158 17836 9210
rect 17780 9156 17836 9158
rect 21476 14084 21532 14140
rect 19908 11732 19964 11788
rect 20244 11732 20300 11788
rect 19908 9268 19964 9324
rect 18508 9210 18564 9212
rect 18508 9158 18510 9210
rect 18510 9158 18562 9210
rect 18562 9158 18564 9210
rect 18508 9156 18564 9158
rect 23604 13188 23660 13244
rect 22148 11732 22204 11788
rect 22260 11844 22316 11900
rect 20636 9268 20692 9324
rect 16660 8036 16716 8092
rect 16884 7252 16940 7308
rect 18060 7418 18116 7420
rect 18060 7366 18062 7418
rect 18062 7366 18114 7418
rect 18114 7366 18116 7418
rect 18060 7364 18116 7366
rect 18620 7418 18676 7420
rect 18620 7366 18622 7418
rect 18622 7366 18674 7418
rect 18674 7366 18676 7418
rect 18620 7364 18676 7366
rect 17612 7252 17668 7308
rect 16660 6580 16716 6636
rect 15876 5684 15932 5740
rect 14084 5236 14140 5292
rect 13300 4564 13356 4620
rect 11956 1316 12012 1372
rect 12964 4452 13020 4508
rect 12292 1092 12348 1148
rect 13300 4004 13356 4060
rect 14196 2996 14252 3052
rect 15764 4900 15820 4956
rect 14420 1540 14476 1596
rect 14756 2660 14812 2716
rect 15428 2548 15484 2604
rect 15988 868 16044 924
rect 16884 5850 16886 5852
rect 16886 5850 16938 5852
rect 16938 5850 16940 5852
rect 16884 5796 16940 5850
rect 17500 5850 17556 5852
rect 17500 5798 17502 5850
rect 17502 5798 17554 5850
rect 17554 5798 17556 5850
rect 17500 5796 17556 5798
rect 18060 5684 18116 5740
rect 19180 8090 19236 8092
rect 19180 8038 19182 8090
rect 19182 8038 19234 8090
rect 19234 8038 19236 8090
rect 19180 8036 19236 8038
rect 21476 7700 21532 7756
rect 19236 6580 19292 6636
rect 25060 13860 25116 13916
rect 25732 13412 25788 13468
rect 24276 11844 24332 11900
rect 25732 10388 25788 10444
rect 22372 9940 22428 9996
rect 21924 8708 21980 8764
rect 23380 9492 23436 9548
rect 25228 9492 25284 9548
rect 22484 8708 22540 8764
rect 25620 8932 25676 8988
rect 20020 6692 20076 6748
rect 18788 5572 18844 5628
rect 16380 4954 16436 4956
rect 16380 4902 16382 4954
rect 16382 4902 16434 4954
rect 16434 4902 16436 4954
rect 16380 4900 16436 4902
rect 16548 2436 16604 2492
rect 17780 1540 17836 1596
rect 18452 980 18508 1036
rect 19236 5124 19292 5180
rect 20692 6468 20748 6524
rect 21476 6692 21532 6748
rect 20468 5124 20524 5180
rect 19348 1428 19404 1484
rect 21140 5012 21196 5068
rect 21700 6804 21756 6860
rect 21532 6522 21588 6524
rect 21532 6470 21534 6522
rect 21534 6470 21586 6522
rect 21586 6470 21588 6522
rect 21532 6468 21588 6470
rect 18900 868 18956 924
rect 19684 868 19740 924
rect 19236 84 19292 140
rect 21700 5124 21756 5180
rect 19908 196 19964 252
rect 20692 196 20748 252
rect 22708 1540 22764 1596
rect 25060 8036 25116 8092
rect 25452 8090 25508 8092
rect 25452 8038 25454 8090
rect 25454 8038 25506 8090
rect 25506 8038 25508 8090
rect 25452 8036 25508 8038
rect 23380 7924 23436 7980
rect 23044 7140 23100 7196
rect 25564 7140 25620 7196
rect 24612 6468 24668 6524
rect 24388 6244 24444 6300
rect 25004 6244 25060 6300
rect 24724 5908 24780 5964
rect 25452 5908 25508 5964
rect 23044 5124 23100 5180
rect 25452 5348 25508 5404
rect 23380 5012 23436 5068
rect 24388 5012 24444 5068
rect 25228 5012 25284 5068
rect 23044 4788 23100 4844
rect 25284 3556 25340 3612
rect 24500 3108 24556 3164
rect 22932 644 22988 700
rect 25172 1428 25228 1484
rect 42308 14868 42364 14924
rect 27972 12964 28028 13020
rect 27188 12740 27244 12796
rect 26964 11732 27020 11788
rect 26740 10052 26796 10108
rect 26348 8986 26404 8988
rect 26348 8934 26350 8986
rect 26350 8934 26402 8986
rect 26402 8934 26404 8986
rect 26348 8932 26404 8934
rect 26628 8202 26684 8204
rect 26628 8150 26630 8202
rect 26630 8150 26682 8202
rect 26682 8150 26684 8202
rect 26628 8148 26684 8150
rect 25900 7924 25956 7980
rect 30100 12516 30156 12572
rect 28644 11732 28700 11788
rect 29876 11732 29932 11788
rect 28376 10218 28432 10220
rect 28376 10166 28378 10218
rect 28378 10166 28430 10218
rect 28430 10166 28432 10218
rect 28376 10164 28432 10166
rect 28480 10218 28536 10220
rect 28480 10166 28482 10218
rect 28482 10166 28534 10218
rect 28534 10166 28536 10218
rect 28480 10164 28536 10166
rect 28584 10218 28640 10220
rect 28584 10166 28586 10218
rect 28586 10166 28638 10218
rect 28638 10166 28640 10218
rect 28584 10164 28640 10166
rect 28376 8650 28432 8652
rect 28376 8598 28378 8650
rect 28378 8598 28430 8650
rect 28430 8598 28432 8650
rect 28376 8596 28432 8598
rect 28480 8650 28536 8652
rect 28480 8598 28482 8650
rect 28482 8598 28534 8650
rect 28534 8598 28536 8650
rect 28480 8596 28536 8598
rect 28584 8650 28640 8652
rect 28584 8598 28586 8650
rect 28586 8598 28638 8650
rect 28638 8598 28640 8650
rect 28584 8596 28640 8598
rect 32340 13636 32396 13692
rect 31556 12516 31612 12572
rect 30884 11732 30940 11788
rect 34468 12964 34524 13020
rect 34356 11732 34412 11788
rect 32676 10164 32732 10220
rect 27468 8148 27524 8204
rect 29540 8202 29596 8204
rect 29540 8150 29542 8202
rect 29542 8150 29594 8202
rect 29594 8150 29596 8202
rect 29540 8148 29596 8150
rect 30324 8148 30380 8204
rect 31556 8202 31612 8204
rect 31556 8150 31558 8202
rect 31558 8150 31610 8202
rect 31610 8150 31612 8202
rect 31556 8148 31612 8150
rect 32340 8148 32396 8204
rect 26404 6356 26460 6412
rect 26404 1652 26460 1708
rect 26964 4676 27020 4732
rect 28196 7140 28252 7196
rect 28376 7082 28432 7084
rect 28376 7030 28378 7082
rect 28378 7030 28430 7082
rect 28430 7030 28432 7082
rect 28376 7028 28432 7030
rect 28480 7082 28536 7084
rect 28480 7030 28482 7082
rect 28482 7030 28534 7082
rect 28534 7030 28536 7082
rect 28480 7028 28536 7030
rect 28584 7082 28640 7084
rect 28584 7030 28586 7082
rect 28586 7030 28638 7082
rect 28638 7030 28640 7082
rect 28584 7028 28640 7030
rect 28700 6634 28756 6636
rect 28700 6582 28702 6634
rect 28702 6582 28754 6634
rect 28754 6582 28756 6634
rect 28700 6580 28756 6582
rect 27748 6132 27804 6188
rect 28364 6132 28420 6188
rect 30100 6020 30156 6076
rect 28376 5514 28432 5516
rect 28376 5462 28378 5514
rect 28378 5462 28430 5514
rect 28430 5462 28432 5514
rect 28376 5460 28432 5462
rect 28480 5514 28536 5516
rect 28480 5462 28482 5514
rect 28482 5462 28534 5514
rect 28534 5462 28536 5514
rect 28480 5460 28536 5462
rect 28584 5514 28640 5516
rect 28584 5462 28586 5514
rect 28586 5462 28638 5514
rect 28638 5462 28640 5514
rect 28584 5460 28640 5462
rect 28308 4900 28364 4956
rect 28196 2884 28252 2940
rect 26852 1092 26908 1148
rect 26964 2772 27020 2828
rect 28756 1540 28812 1596
rect 29148 4954 29204 4956
rect 29148 4902 29150 4954
rect 29150 4902 29202 4954
rect 29202 4902 29204 4954
rect 29148 4900 29204 4902
rect 30604 7140 30660 7196
rect 30604 6916 30660 6972
rect 30884 4564 30940 4620
rect 30324 4228 30380 4284
rect 29204 3892 29260 3948
rect 31220 3444 31276 3500
rect 30660 3332 30716 3388
rect 29988 1540 30044 1596
rect 29652 644 29708 700
rect 31780 5460 31836 5516
rect 35252 11732 35308 11788
rect 36708 12740 36764 12796
rect 36708 11732 36764 11788
rect 37380 11732 37436 11788
rect 38836 13524 38892 13580
rect 36820 10052 36876 10108
rect 34916 8202 34972 8204
rect 34916 8150 34918 8202
rect 34918 8150 34970 8202
rect 34970 8150 34972 8202
rect 34916 8148 34972 8150
rect 35756 8148 35812 8204
rect 36372 8148 36428 8204
rect 34020 7140 34076 7196
rect 34524 7140 34580 7196
rect 34692 6356 34748 6412
rect 35084 6356 35140 6412
rect 33460 6020 33516 6076
rect 35532 6020 35588 6076
rect 32676 5684 32732 5740
rect 33460 5684 33516 5740
rect 33852 5684 33908 5740
rect 33460 4676 33516 4732
rect 32452 3220 32508 3276
rect 33684 1204 33740 1260
rect 31444 532 31500 588
rect 35028 4900 35084 4956
rect 35644 4954 35700 4956
rect 35644 4902 35646 4954
rect 35646 4902 35698 4954
rect 35698 4902 35700 4954
rect 35644 4900 35700 4902
rect 34244 1540 34300 1596
rect 35476 1540 35532 1596
rect 35924 4452 35980 4508
rect 36932 8148 36988 8204
rect 38724 7028 38780 7084
rect 37828 6580 37884 6636
rect 39004 6580 39060 6636
rect 38500 5572 38556 5628
rect 37604 2324 37660 2380
rect 39228 5572 39284 5628
rect 39060 1428 39116 1484
rect 39172 980 39228 1036
rect 40740 7924 40796 7980
rect 39788 7028 39844 7084
rect 40068 6132 40124 6188
rect 40068 5572 40124 5628
rect 41972 10052 42028 10108
rect 42980 14644 43036 14700
rect 45668 14532 45724 14588
rect 43652 12628 43708 12684
rect 42980 11732 43036 11788
rect 42644 11284 42700 11340
rect 42644 10052 42700 10108
rect 42532 9268 42588 9324
rect 40180 4228 40236 4284
rect 42868 9098 42924 9100
rect 42868 9046 42870 9098
rect 42870 9046 42922 9098
rect 42922 9046 42924 9098
rect 42868 9044 42924 9046
rect 42196 7642 42252 7644
rect 42196 7590 42198 7642
rect 42198 7590 42250 7642
rect 42250 7590 42252 7642
rect 42196 7588 42252 7590
rect 41972 5796 42028 5852
rect 42364 5850 42420 5852
rect 42364 5798 42366 5850
rect 42366 5798 42418 5850
rect 42418 5798 42420 5850
rect 42364 5796 42420 5798
rect 41860 4676 41916 4732
rect 41748 2996 41804 3052
rect 42196 4004 42252 4060
rect 41636 2212 41692 2268
rect 35812 308 35868 364
rect 39396 756 39452 812
rect 39732 868 39788 924
rect 40404 868 40460 924
rect 40964 868 41020 924
rect 43988 11732 44044 11788
rect 44884 12068 44940 12124
rect 44660 11732 44716 11788
rect 43204 9604 43260 9660
rect 43484 9044 43540 9100
rect 43204 8260 43260 8316
rect 43932 9268 43988 9324
rect 44100 9268 44156 9324
rect 44548 9268 44604 9324
rect 45444 11396 45500 11452
rect 45220 9658 45276 9660
rect 45220 9606 45222 9658
rect 45222 9606 45274 9658
rect 45274 9606 45276 9658
rect 45220 9604 45276 9606
rect 46116 11732 46172 11788
rect 46452 12964 46508 13020
rect 47684 12292 47740 12348
rect 46900 11844 46956 11900
rect 46060 9658 46116 9660
rect 46060 9606 46062 9658
rect 46062 9606 46114 9658
rect 46114 9606 46116 9658
rect 46060 9604 46116 9606
rect 46676 9604 46732 9660
rect 43428 6692 43484 6748
rect 43316 6627 43318 6636
rect 43318 6627 43370 6636
rect 43370 6627 43372 6636
rect 43316 6580 43372 6627
rect 43204 6132 43260 6188
rect 42756 5796 42812 5852
rect 43260 5850 43316 5852
rect 43260 5798 43262 5850
rect 43262 5798 43314 5850
rect 43314 5798 43316 5850
rect 43260 5796 43316 5798
rect 43092 4788 43148 4844
rect 43932 6746 43988 6748
rect 43932 6694 43934 6746
rect 43934 6694 43986 6746
rect 43986 6694 43988 6746
rect 43932 6692 43988 6694
rect 43652 6468 43708 6524
rect 43820 6580 43876 6636
rect 43876 5124 43932 5180
rect 43708 4788 43764 4844
rect 43316 1988 43372 2044
rect 43988 1316 44044 1372
rect 41188 420 41244 476
rect 44604 7140 44660 7196
rect 44380 6522 44436 6524
rect 44380 6470 44382 6522
rect 44382 6470 44434 6522
rect 44434 6470 44436 6522
rect 44380 6468 44436 6470
rect 44324 4676 44380 4732
rect 45108 4788 45164 4844
rect 45108 2996 45164 3052
rect 45220 2660 45276 2716
rect 45892 1428 45948 1484
rect 45220 1316 45276 1372
rect 44660 1092 44716 1148
rect 47348 10276 47404 10332
rect 47068 9658 47124 9660
rect 47068 9606 47070 9658
rect 47070 9606 47122 9658
rect 47122 9606 47124 9658
rect 47068 9604 47124 9606
rect 46844 9098 46900 9100
rect 46844 9046 46846 9098
rect 46846 9046 46898 9098
rect 46898 9046 46900 9098
rect 46844 9044 46900 9046
rect 48580 12180 48636 12236
rect 48356 11844 48412 11900
rect 48468 11956 48524 12012
rect 47796 11732 47852 11788
rect 48020 11172 48076 11228
rect 48020 10276 48076 10332
rect 48244 8932 48300 8988
rect 48244 8596 48300 8652
rect 50260 11844 50316 11900
rect 49028 11732 49084 11788
rect 49812 11732 49868 11788
rect 48860 10276 48916 10332
rect 48804 8596 48860 8652
rect 46228 7642 46284 7644
rect 46228 7590 46230 7642
rect 46230 7590 46282 7642
rect 46282 7590 46284 7642
rect 46228 7588 46284 7590
rect 46564 5796 46620 5852
rect 46564 2548 46620 2604
rect 46452 1540 46508 1596
rect 44212 308 44268 364
rect 47348 8090 47404 8092
rect 47348 8038 47350 8090
rect 47350 8038 47402 8090
rect 47402 8038 47404 8090
rect 47348 8036 47404 8038
rect 47124 7588 47180 7644
rect 47404 6746 47460 6748
rect 47404 6694 47406 6746
rect 47406 6694 47458 6746
rect 47458 6694 47460 6746
rect 47404 6692 47460 6694
rect 47068 5796 47124 5852
rect 48356 6858 48412 6860
rect 48356 6806 48358 6858
rect 48358 6806 48410 6858
rect 48410 6806 48412 6858
rect 48356 6804 48412 6806
rect 46900 4564 46956 4620
rect 49308 8986 49364 8988
rect 49308 8934 49310 8986
rect 49310 8934 49362 8986
rect 49362 8934 49364 8986
rect 49308 8932 49364 8934
rect 49924 9268 49980 9324
rect 52948 14644 53004 14700
rect 51044 13188 51100 13244
rect 53620 14644 53676 14700
rect 53060 13188 53116 13244
rect 52724 12068 52780 12124
rect 51268 11956 51324 12012
rect 52500 11956 52556 12012
rect 50372 11732 50428 11788
rect 51156 11620 51212 11676
rect 50820 10276 50876 10332
rect 50540 9268 50596 9324
rect 50708 9492 50764 9548
rect 49028 6692 49084 6748
rect 51828 10388 51884 10444
rect 51604 10276 51660 10332
rect 52164 10052 52220 10108
rect 54404 14868 54460 14924
rect 53844 13466 53900 13468
rect 53844 13414 53846 13466
rect 53846 13414 53898 13466
rect 53898 13414 53900 13466
rect 53844 13412 53900 13414
rect 58324 14308 58380 14364
rect 54404 13300 54460 13356
rect 55748 13300 55804 13356
rect 55972 12852 56028 12908
rect 57092 13748 57148 13804
rect 55636 12292 55692 12348
rect 53620 11956 53676 12012
rect 54404 11956 54460 12012
rect 53284 10500 53340 10556
rect 52780 10052 52836 10108
rect 52500 8932 52556 8988
rect 51828 8148 51884 8204
rect 52164 8484 52220 8540
rect 51604 6804 51660 6860
rect 48636 6132 48692 6188
rect 48356 4788 48412 4844
rect 48748 4564 48804 4620
rect 51772 6746 51828 6748
rect 51772 6694 51774 6746
rect 51774 6694 51826 6746
rect 51826 6694 51828 6746
rect 51772 6692 51828 6694
rect 52164 6692 52220 6748
rect 50372 5796 50428 5852
rect 51044 5796 51100 5852
rect 51548 5850 51604 5852
rect 51548 5798 51550 5850
rect 51550 5798 51602 5850
rect 51602 5798 51604 5850
rect 51548 5796 51604 5798
rect 52052 5572 52108 5628
rect 49812 5012 49868 5068
rect 49644 4788 49700 4844
rect 49700 3668 49756 3724
rect 49588 2884 49644 2940
rect 52052 4676 52108 4732
rect 52276 4788 52332 4844
rect 54180 10276 54236 10332
rect 53564 9770 53620 9772
rect 53564 9718 53566 9770
rect 53566 9718 53618 9770
rect 53618 9718 53620 9770
rect 53564 9716 53620 9718
rect 54068 7924 54124 7980
rect 52668 7028 52724 7084
rect 52556 6804 52612 6860
rect 52556 6522 52612 6524
rect 52556 6470 52558 6522
rect 52558 6470 52610 6522
rect 52610 6470 52612 6522
rect 52556 6468 52612 6470
rect 53844 6580 53900 6636
rect 52388 3892 52444 3948
rect 52724 4676 52780 4732
rect 52724 3892 52780 3948
rect 50484 2436 50540 2492
rect 50708 2548 50764 2604
rect 48356 1876 48412 1932
rect 47684 1540 47740 1596
rect 49476 1428 49532 1484
rect 48916 1316 48972 1372
rect 50148 1092 50204 1148
rect 52500 3108 52556 3164
rect 52164 1540 52220 1596
rect 53172 1652 53228 1708
rect 46676 532 46732 588
rect 49924 474 49980 476
rect 49924 422 49926 474
rect 49926 422 49978 474
rect 49978 422 49980 474
rect 49924 420 49980 422
rect 54516 9994 54572 9996
rect 54516 9942 54518 9994
rect 54518 9942 54570 9994
rect 54570 9942 54572 9994
rect 54516 9940 54572 9942
rect 57092 12068 57148 12124
rect 56308 10388 56364 10444
rect 55188 9716 55244 9772
rect 55412 9716 55468 9772
rect 55540 9434 55596 9436
rect 55540 9382 55542 9434
rect 55542 9382 55594 9434
rect 55594 9382 55596 9434
rect 55540 9380 55596 9382
rect 55644 9434 55700 9436
rect 55644 9382 55646 9434
rect 55646 9382 55698 9434
rect 55698 9382 55700 9434
rect 55644 9380 55700 9382
rect 55748 9434 55804 9436
rect 55748 9382 55750 9434
rect 55750 9382 55802 9434
rect 55802 9382 55804 9434
rect 55748 9380 55804 9382
rect 54852 9156 54908 9212
rect 56588 9770 56644 9772
rect 56588 9718 56590 9770
rect 56590 9718 56642 9770
rect 56642 9718 56644 9770
rect 56588 9716 56644 9718
rect 56420 9492 56476 9548
rect 57036 9492 57092 9548
rect 57316 9156 57372 9212
rect 57428 8932 57484 8988
rect 56644 7924 56700 7980
rect 55540 7866 55596 7868
rect 55540 7814 55542 7866
rect 55542 7814 55594 7866
rect 55594 7814 55596 7866
rect 55540 7812 55596 7814
rect 55644 7866 55700 7868
rect 55644 7814 55646 7866
rect 55646 7814 55698 7866
rect 55698 7814 55700 7866
rect 55644 7812 55700 7814
rect 55748 7866 55804 7868
rect 55748 7814 55750 7866
rect 55750 7814 55802 7866
rect 55802 7814 55804 7866
rect 55748 7812 55804 7814
rect 54964 6580 55020 6636
rect 54516 4788 54572 4844
rect 54628 4676 54684 4732
rect 54628 1652 54684 1708
rect 52164 532 52220 588
rect 55540 6298 55596 6300
rect 55540 6246 55542 6298
rect 55542 6246 55594 6298
rect 55594 6246 55596 6298
rect 55540 6244 55596 6246
rect 55644 6298 55700 6300
rect 55644 6246 55646 6298
rect 55646 6246 55698 6298
rect 55698 6246 55700 6298
rect 55644 6244 55700 6246
rect 55748 6298 55804 6300
rect 55748 6246 55750 6298
rect 55750 6246 55802 6298
rect 55802 6246 55804 6298
rect 55748 6244 55804 6246
rect 55748 5124 55804 5180
rect 55188 4676 55244 4732
rect 55540 4730 55596 4732
rect 55540 4678 55542 4730
rect 55542 4678 55594 4730
rect 55594 4678 55596 4730
rect 55540 4676 55596 4678
rect 55644 4730 55700 4732
rect 55644 4678 55646 4730
rect 55646 4678 55698 4730
rect 55698 4678 55700 4730
rect 55644 4676 55700 4678
rect 55748 4730 55804 4732
rect 55748 4678 55750 4730
rect 55750 4678 55802 4730
rect 55802 4678 55804 4730
rect 55748 4676 55804 4678
rect 55188 4228 55244 4284
rect 55076 3834 55132 3836
rect 55076 3782 55078 3834
rect 55078 3782 55130 3834
rect 55130 3782 55132 3834
rect 55076 3780 55132 3782
rect 55636 1764 55692 1820
rect 55076 1540 55132 1596
rect 56756 6804 56812 6860
rect 56868 7700 56924 7756
rect 56588 6580 56644 6636
rect 56420 6468 56476 6524
rect 56196 5572 56252 5628
rect 56196 5124 56252 5180
rect 56196 4004 56252 4060
rect 56196 3274 56252 3276
rect 56196 3222 56198 3274
rect 56198 3222 56250 3274
rect 56250 3222 56252 3274
rect 56196 3220 56252 3222
rect 56196 1876 56252 1932
rect 55972 1540 56028 1596
rect 57764 13188 57820 13244
rect 57540 7700 57596 7756
rect 57652 10724 57708 10780
rect 56868 6580 56924 6636
rect 56980 6692 57036 6748
rect 58772 14532 58828 14588
rect 58324 14084 58380 14140
rect 58212 13076 58268 13132
rect 63140 14868 63196 14924
rect 60004 12964 60060 13020
rect 60452 13412 60508 13468
rect 59220 12628 59276 12684
rect 57876 11732 57932 11788
rect 58100 11732 58156 11788
rect 58100 11284 58156 11340
rect 58324 11284 58380 11340
rect 58828 9098 58884 9100
rect 58828 9046 58830 9098
rect 58830 9046 58882 9098
rect 58882 9046 58884 9098
rect 58828 9044 58884 9046
rect 57988 8932 58044 8988
rect 58268 8874 58324 8876
rect 58268 8822 58270 8874
rect 58270 8822 58322 8874
rect 58322 8822 58324 8874
rect 58268 8820 58324 8822
rect 58996 8372 59052 8428
rect 60788 12964 60844 13020
rect 61236 13636 61292 13692
rect 61460 12180 61516 12236
rect 60452 11844 60508 11900
rect 60788 10612 60844 10668
rect 60788 10052 60844 10108
rect 60564 9716 60620 9772
rect 60452 9044 60508 9100
rect 59388 8986 59444 8988
rect 59388 8934 59390 8986
rect 59390 8934 59442 8986
rect 59442 8934 59444 8986
rect 59388 8932 59444 8934
rect 60564 8596 60620 8652
rect 61012 9156 61068 9212
rect 61236 9210 61292 9212
rect 61236 9158 61238 9210
rect 61238 9158 61290 9210
rect 61290 9158 61292 9210
rect 61236 9156 61292 9158
rect 61796 13636 61852 13692
rect 64148 14308 64204 14364
rect 65380 14532 65436 14588
rect 63700 13412 63756 13468
rect 64260 13524 64316 13580
rect 62244 12852 62300 12908
rect 63700 12122 63756 12124
rect 63700 12070 63702 12122
rect 63702 12070 63754 12122
rect 63754 12070 63756 12122
rect 63700 12068 63756 12070
rect 63364 11844 63420 11900
rect 62356 11732 62412 11788
rect 62356 11508 62412 11564
rect 61964 9210 62020 9212
rect 61964 9158 61966 9210
rect 61966 9158 62018 9210
rect 62018 9158 62020 9210
rect 61964 9156 62020 9158
rect 60788 8596 60844 8652
rect 60452 8484 60508 8540
rect 59444 8372 59500 8428
rect 58436 7812 58492 7868
rect 58324 7700 58380 7756
rect 58044 7252 58100 7308
rect 58660 7700 58716 7756
rect 59332 7700 59388 7756
rect 58324 7252 58380 7308
rect 58604 6804 58660 6860
rect 57372 6244 57428 6300
rect 63924 11508 63980 11564
rect 60508 8148 60564 8204
rect 63252 8148 63308 8204
rect 59780 7364 59836 7420
rect 62916 7700 62972 7756
rect 63420 7700 63476 7756
rect 58996 6468 59052 6524
rect 59948 6522 60004 6524
rect 59948 6470 59950 6522
rect 59950 6470 60002 6522
rect 60002 6470 60004 6522
rect 59948 6468 60004 6470
rect 58380 6244 58436 6300
rect 60676 6580 60732 6636
rect 57204 5460 57260 5516
rect 57092 5348 57148 5404
rect 58660 5348 58716 5404
rect 56588 4954 56644 4956
rect 56588 4902 56590 4954
rect 56590 4902 56642 4954
rect 56642 4902 56644 4954
rect 56588 4900 56644 4902
rect 57988 4900 58044 4956
rect 57092 4058 57148 4060
rect 57092 4006 57094 4058
rect 57094 4006 57146 4058
rect 57146 4006 57148 4058
rect 57092 4004 57148 4006
rect 57316 4004 57372 4060
rect 57316 3556 57372 3612
rect 56980 2660 57036 2716
rect 56420 1652 56476 1708
rect 56868 2212 56924 2268
rect 58772 4228 58828 4284
rect 58884 4116 58940 4172
rect 59444 4116 59500 4172
rect 60508 5348 60564 5404
rect 60676 5124 60732 5180
rect 60228 4676 60284 4732
rect 60676 4004 60732 4060
rect 60340 3780 60396 3836
rect 63028 7364 63084 7420
rect 60340 3220 60396 3276
rect 60900 7252 60956 7308
rect 60228 3108 60284 3164
rect 60116 2996 60172 3052
rect 59892 2660 59948 2716
rect 59668 2548 59724 2604
rect 60116 2436 60172 2492
rect 57988 2100 58044 2156
rect 58660 2212 58716 2268
rect 57876 1988 57932 2044
rect 57428 1652 57484 1708
rect 59220 1204 59276 1260
rect 56532 420 56588 476
rect 60116 1876 60172 1932
rect 62356 7252 62412 7308
rect 62244 6804 62300 6860
rect 61740 6244 61796 6300
rect 62692 6692 62748 6748
rect 62692 6244 62748 6300
rect 62468 6132 62524 6188
rect 60900 2996 60956 3052
rect 60676 1764 60732 1820
rect 60452 1652 60508 1708
rect 61908 2436 61964 2492
rect 61796 2324 61852 2380
rect 62020 2378 62076 2380
rect 62020 2326 62022 2378
rect 62022 2326 62074 2378
rect 62074 2326 62076 2378
rect 62020 2324 62076 2326
rect 62132 2100 62188 2156
rect 61796 1988 61852 2044
rect 63476 4788 63532 4844
rect 62804 4116 62860 4172
rect 62804 3332 62860 3388
rect 63868 7364 63924 7420
rect 67900 14868 67956 14924
rect 65940 13636 65996 13692
rect 66500 13076 66556 13132
rect 65716 12292 65772 12348
rect 65268 12068 65324 12124
rect 64372 11732 64428 11788
rect 66724 13636 66780 13692
rect 68068 13524 68124 13580
rect 66724 12292 66780 12348
rect 66948 12292 67004 12348
rect 66612 11956 66668 12012
rect 68292 13188 68348 13244
rect 67844 12180 67900 12236
rect 67396 11956 67452 12012
rect 66276 11172 66332 11228
rect 66500 11172 66556 11228
rect 64260 8260 64316 8316
rect 64932 8932 64988 8988
rect 65324 8986 65380 8988
rect 65324 8934 65326 8986
rect 65326 8934 65378 8986
rect 65378 8934 65380 8986
rect 65324 8932 65380 8934
rect 64148 6692 64204 6748
rect 63812 5124 63868 5180
rect 64428 4788 64484 4844
rect 65268 4676 65324 4732
rect 64820 4564 64876 4620
rect 67060 10612 67116 10668
rect 66500 10276 66556 10332
rect 67172 9940 67228 9996
rect 67284 10612 67340 10668
rect 66388 9268 66444 9324
rect 65604 8372 65660 8428
rect 65716 8260 65772 8316
rect 66052 8202 66108 8204
rect 66052 8150 66054 8202
rect 66054 8150 66106 8202
rect 66106 8150 66108 8202
rect 66052 8148 66108 8150
rect 66556 8314 66612 8316
rect 66556 8262 66558 8314
rect 66558 8262 66610 8314
rect 66610 8262 66612 8314
rect 66556 8260 66612 8262
rect 66724 7700 66780 7756
rect 66836 8372 66892 8428
rect 66276 6804 66332 6860
rect 66724 6804 66780 6860
rect 65828 6694 65884 6748
rect 65828 6692 65830 6694
rect 65830 6692 65882 6694
rect 65882 6692 65884 6694
rect 65604 5796 65660 5852
rect 66724 6132 66780 6188
rect 63700 3556 63756 3612
rect 62580 2884 62636 2940
rect 62468 2548 62524 2604
rect 62580 2212 62636 2268
rect 62468 1876 62524 1932
rect 62804 1930 62860 1932
rect 62804 1878 62806 1930
rect 62806 1878 62858 1930
rect 62858 1878 62860 1930
rect 62804 1876 62860 1878
rect 62244 1540 62300 1596
rect 62468 1540 62524 1596
rect 62244 1316 62300 1372
rect 62580 1204 62636 1260
rect 65156 1988 65212 2044
rect 64148 980 64204 1036
rect 69860 14308 69916 14364
rect 68628 12628 68684 12684
rect 69076 12068 69132 12124
rect 70420 14756 70476 14812
rect 71876 14756 71932 14812
rect 68180 11172 68236 11228
rect 69188 11284 69244 11340
rect 67620 10388 67676 10444
rect 67844 10388 67900 10444
rect 67508 9268 67564 9324
rect 68964 10388 69020 10444
rect 68964 10164 69020 10220
rect 69300 10164 69356 10220
rect 69188 9828 69244 9884
rect 69300 9604 69356 9660
rect 67956 8372 68012 8428
rect 67060 7700 67116 7756
rect 67172 6804 67228 6860
rect 67452 5850 67508 5852
rect 67452 5798 67454 5850
rect 67454 5798 67506 5850
rect 67506 5798 67508 5850
rect 67452 5796 67508 5798
rect 67060 4900 67116 4956
rect 66612 4228 66668 4284
rect 66500 4004 66556 4060
rect 66052 3108 66108 3164
rect 66164 3332 66220 3388
rect 65492 2324 65548 2380
rect 65268 1876 65324 1932
rect 66724 3780 66780 3836
rect 66276 1540 66332 1596
rect 59668 308 59724 364
rect 66164 756 66220 812
rect 67060 3834 67116 3836
rect 67060 3782 67062 3834
rect 67062 3782 67114 3834
rect 67114 3782 67116 3834
rect 67060 3780 67116 3782
rect 67900 7700 67956 7756
rect 68348 7476 68404 7532
rect 68964 7700 69020 7756
rect 68124 7418 68180 7420
rect 68124 7366 68126 7418
rect 68126 7366 68178 7418
rect 68178 7366 68180 7418
rect 68124 7364 68180 7366
rect 67900 6804 67956 6860
rect 68348 6244 68404 6300
rect 68180 5236 68236 5292
rect 68796 6132 68852 6188
rect 67620 4788 67676 4844
rect 67284 3444 67340 3500
rect 67396 4004 67452 4060
rect 67844 2212 67900 2268
rect 68404 4900 68460 4956
rect 68404 3610 68460 3612
rect 68404 3558 68406 3610
rect 68406 3558 68458 3610
rect 68458 3558 68460 3610
rect 68404 3556 68460 3558
rect 68292 2100 68348 2156
rect 68404 2772 68460 2828
rect 68628 2548 68684 2604
rect 68740 2324 68796 2380
rect 68516 1204 68572 1260
rect 68740 532 68796 588
rect 68964 4900 69020 4956
rect 69412 8148 69468 8204
rect 69524 7700 69580 7756
rect 69524 7252 69580 7308
rect 69412 5796 69468 5852
rect 69244 5738 69300 5740
rect 69244 5686 69246 5738
rect 69246 5686 69298 5738
rect 69298 5686 69300 5738
rect 69244 5684 69300 5686
rect 69076 4452 69132 4508
rect 69188 3556 69244 3612
rect 69860 12234 69916 12236
rect 69860 12182 69862 12234
rect 69862 12182 69914 12234
rect 69914 12182 69916 12234
rect 69860 12180 69916 12182
rect 71764 14084 71820 14140
rect 71876 13860 71932 13916
rect 71764 12068 71820 12124
rect 70980 11844 71036 11900
rect 71204 11844 71260 11900
rect 70980 10612 71036 10668
rect 69972 9268 70028 9324
rect 70196 9268 70252 9324
rect 70588 8820 70644 8876
rect 70196 8596 70252 8652
rect 69748 8372 69804 8428
rect 71204 9268 71260 9324
rect 70644 8148 70700 8204
rect 74004 13412 74060 13468
rect 74004 13188 74060 13244
rect 74228 13412 74284 13468
rect 74228 13076 74284 13132
rect 74452 13076 74508 13132
rect 73556 12852 73612 12908
rect 73556 12628 73612 12684
rect 73108 11956 73164 12012
rect 74116 12068 74172 12124
rect 72100 9940 72156 9996
rect 72660 11172 72716 11228
rect 72660 9828 72716 9884
rect 72772 9716 72828 9772
rect 71204 8148 71260 8204
rect 71428 8202 71484 8204
rect 71428 8150 71430 8202
rect 71430 8150 71482 8202
rect 71482 8150 71484 8202
rect 71428 8148 71484 8150
rect 74340 12068 74396 12124
rect 73444 11172 73500 11228
rect 73220 9604 73276 9660
rect 72772 8484 72828 8540
rect 71988 8148 72044 8204
rect 72100 8372 72156 8428
rect 71764 7588 71820 7644
rect 70868 7364 70924 7420
rect 71428 7364 71484 7420
rect 69860 7140 69916 7196
rect 70532 6916 70588 6972
rect 70140 6804 70196 6860
rect 70588 6356 70644 6412
rect 69916 5962 69972 5964
rect 69916 5910 69918 5962
rect 69918 5910 69970 5962
rect 69970 5910 69972 5962
rect 70700 6244 70756 6300
rect 69916 5908 69972 5910
rect 69636 5796 69692 5852
rect 70308 5796 70364 5852
rect 71428 6132 71484 6188
rect 69524 4788 69580 4844
rect 69636 3892 69692 3948
rect 70196 3220 70252 3276
rect 69076 2548 69132 2604
rect 69076 1764 69132 1820
rect 69636 2100 69692 2156
rect 68964 980 69020 1036
rect 70308 2660 70364 2716
rect 72212 7924 72268 7980
rect 72324 7140 72380 7196
rect 72100 6356 72156 6412
rect 71932 6074 71988 6076
rect 71932 6022 71934 6074
rect 71934 6022 71986 6074
rect 71986 6022 71988 6074
rect 71932 6020 71988 6022
rect 71764 5236 71820 5292
rect 71204 5012 71260 5068
rect 70868 4900 70924 4956
rect 70756 4004 70812 4060
rect 72100 4228 72156 4284
rect 70532 3108 70588 3164
rect 70756 3108 70812 3164
rect 71876 3332 71932 3388
rect 70868 1764 70924 1820
rect 70532 1428 70588 1484
rect 71988 1428 72044 1484
rect 72324 2884 72380 2940
rect 73332 6020 73388 6076
rect 73276 5572 73332 5628
rect 72548 5236 72604 5292
rect 72436 2324 72492 2380
rect 72548 4788 72604 4844
rect 73332 4004 73388 4060
rect 73220 3668 73276 3724
rect 72772 3556 72828 3612
rect 72884 3444 72940 3500
rect 72772 3332 72828 3388
rect 72884 3220 72940 3276
rect 73108 2436 73164 2492
rect 72548 1316 72604 1372
rect 72660 2324 72716 2380
rect 73892 11172 73948 11228
rect 73668 9156 73724 9212
rect 74116 9210 74172 9212
rect 74116 9158 74118 9210
rect 74118 9158 74170 9210
rect 74170 9158 74172 9210
rect 74116 9156 74172 9158
rect 73892 7476 73948 7532
rect 74116 7588 74172 7644
rect 74676 13860 74732 13916
rect 77700 14532 77756 14588
rect 74900 13860 74956 13916
rect 75012 12852 75068 12908
rect 74788 11956 74844 12012
rect 74564 11844 74620 11900
rect 74452 11732 74508 11788
rect 77252 14084 77308 14140
rect 78036 14138 78092 14140
rect 78036 14086 78038 14138
rect 78038 14086 78090 14138
rect 78090 14086 78092 14138
rect 78036 14084 78092 14086
rect 76916 13748 76972 13804
rect 77140 13748 77196 13804
rect 76916 13412 76972 13468
rect 76580 11732 76636 11788
rect 75236 10052 75292 10108
rect 77140 13412 77196 13468
rect 77252 13188 77308 13244
rect 77140 13076 77196 13132
rect 77028 12852 77084 12908
rect 77364 12964 77420 13020
rect 78036 12740 78092 12796
rect 77924 12458 77980 12460
rect 77924 12406 77926 12458
rect 77926 12406 77978 12458
rect 77978 12406 77980 12458
rect 77924 12404 77980 12406
rect 78260 12346 78316 12348
rect 78260 12294 78262 12346
rect 78262 12294 78314 12346
rect 78314 12294 78316 12346
rect 78260 12292 78316 12294
rect 77252 10724 77308 10780
rect 79156 14644 79212 14700
rect 78484 13972 78540 14028
rect 78484 13076 78540 13132
rect 78708 13972 78764 14028
rect 79156 13972 79212 14028
rect 78708 12404 78764 12460
rect 79268 12964 79324 13020
rect 78820 12292 78876 12348
rect 78932 12404 78988 12460
rect 78036 10948 78092 11004
rect 78148 11060 78204 11116
rect 76804 10052 76860 10108
rect 76020 9604 76076 9660
rect 74844 9156 74900 9212
rect 74676 8372 74732 8428
rect 74900 8260 74956 8316
rect 74676 7364 74732 7420
rect 74564 7252 74620 7308
rect 75012 7364 75068 7420
rect 74788 7140 74844 7196
rect 75068 6804 75124 6860
rect 75628 7252 75684 7308
rect 75628 6916 75684 6972
rect 76076 7418 76132 7420
rect 76076 7366 76078 7418
rect 76078 7366 76130 7418
rect 76130 7366 76132 7418
rect 76076 7364 76132 7366
rect 75180 6634 75236 6636
rect 75180 6582 75182 6634
rect 75182 6582 75234 6634
rect 75234 6582 75236 6634
rect 75180 6580 75236 6582
rect 76020 6804 76076 6860
rect 76300 7140 76356 7196
rect 75740 6522 75796 6524
rect 75740 6470 75742 6522
rect 75742 6470 75794 6522
rect 75794 6470 75796 6522
rect 75740 6468 75796 6470
rect 76020 6356 76076 6412
rect 75572 6244 75628 6300
rect 75572 5572 75628 5628
rect 75180 5460 75236 5516
rect 73892 5012 73948 5068
rect 75180 5012 75236 5068
rect 73668 4900 73724 4956
rect 73556 4004 73612 4060
rect 74004 4788 74060 4844
rect 74116 4564 74172 4620
rect 74452 4228 74508 4284
rect 74004 4004 74060 4060
rect 74676 3780 74732 3836
rect 73444 2884 73500 2940
rect 73668 3332 73724 3388
rect 75348 3780 75404 3836
rect 75012 3556 75068 3612
rect 73556 2660 73612 2716
rect 73444 2100 73500 2156
rect 71876 196 71932 252
rect 73668 2436 73724 2492
rect 74564 1876 74620 1932
rect 75012 2996 75068 3052
rect 75348 3220 75404 3276
rect 75908 4228 75964 4284
rect 75796 3220 75852 3276
rect 75684 2772 75740 2828
rect 75908 2548 75964 2604
rect 75236 2212 75292 2268
rect 75012 2100 75068 2156
rect 74900 1204 74956 1260
rect 74788 644 74844 700
rect 75460 1876 75516 1932
rect 75348 1316 75404 1372
rect 75348 756 75404 812
rect 76804 8260 76860 8316
rect 76468 6020 76524 6076
rect 76692 4564 76748 4620
rect 76468 4340 76524 4396
rect 76692 2996 76748 3052
rect 76468 1988 76524 2044
rect 76692 1988 76748 2044
rect 76020 980 76076 1036
rect 76468 1428 76524 1484
rect 76244 868 76300 924
rect 76916 6468 76972 6524
rect 77140 9716 77196 9772
rect 77140 8260 77196 8316
rect 77588 9994 77644 9996
rect 77588 9942 77590 9994
rect 77590 9942 77642 9994
rect 77642 9942 77644 9994
rect 77588 9940 77644 9942
rect 78596 11620 78652 11676
rect 78820 11620 78876 11676
rect 78372 10276 78428 10332
rect 79156 12516 79212 12572
rect 78260 9940 78316 9996
rect 78372 10052 78428 10108
rect 78820 11060 78876 11116
rect 79380 12516 79436 12572
rect 80948 13972 81004 14028
rect 79604 12740 79660 12796
rect 79716 12180 79772 12236
rect 79380 11284 79436 11340
rect 79604 11284 79660 11340
rect 78596 10052 78652 10108
rect 78652 9268 78708 9324
rect 79044 10164 79100 10220
rect 78932 10052 78988 10108
rect 77588 8708 77644 8764
rect 78204 8986 78260 8988
rect 78204 8934 78206 8986
rect 78206 8934 78258 8986
rect 78258 8934 78260 8986
rect 78204 8932 78260 8934
rect 77476 8036 77532 8092
rect 77980 8596 78036 8652
rect 77924 8036 77980 8092
rect 77588 7924 77644 7980
rect 77812 7924 77868 7980
rect 77924 7306 77980 7308
rect 77924 7254 77926 7306
rect 77926 7254 77978 7306
rect 77978 7254 77980 7306
rect 77924 7252 77980 7254
rect 77812 5908 77868 5964
rect 78876 8090 78932 8092
rect 78876 8038 78878 8090
rect 78878 8038 78930 8090
rect 78930 8038 78932 8090
rect 78876 8036 78932 8038
rect 79268 10052 79324 10108
rect 79156 9156 79212 9212
rect 79268 8932 79324 8988
rect 79604 10164 79660 10220
rect 79492 8932 79548 8988
rect 79268 8260 79324 8316
rect 79436 8596 79492 8652
rect 80164 12516 80220 12572
rect 80052 12404 80108 12460
rect 82068 13860 82124 13916
rect 82852 14756 82908 14812
rect 82852 14420 82908 14476
rect 83524 14868 83580 14924
rect 82292 13412 82348 13468
rect 83076 13860 83132 13916
rect 82404 13300 82460 13356
rect 82516 13412 82572 13468
rect 82740 13354 82796 13356
rect 82740 13302 82742 13354
rect 82742 13302 82794 13354
rect 82794 13302 82796 13354
rect 82740 13300 82796 13302
rect 80948 12516 81004 12572
rect 81732 12068 81788 12124
rect 81508 11844 81564 11900
rect 83076 12570 83132 12572
rect 83076 12518 83078 12570
rect 83078 12518 83130 12570
rect 83130 12518 83132 12570
rect 83076 12516 83132 12518
rect 83188 12292 83244 12348
rect 82852 12068 82908 12124
rect 83076 12068 83132 12124
rect 82740 11844 82796 11900
rect 83412 12740 83468 12796
rect 83412 12516 83468 12572
rect 83412 11956 83468 12012
rect 81732 10724 81788 10780
rect 83188 11396 83244 11452
rect 82964 11172 83020 11228
rect 83748 14868 83804 14924
rect 83748 13524 83804 13580
rect 83636 13300 83692 13356
rect 83636 12404 83692 12460
rect 83860 13300 83916 13356
rect 83860 12740 83916 12796
rect 84980 13524 85036 13580
rect 84868 13076 84924 13132
rect 84756 12516 84812 12572
rect 84980 12516 85036 12572
rect 83972 11732 84028 11788
rect 83860 11396 83916 11452
rect 84196 11284 84252 11340
rect 84420 11284 84476 11340
rect 82292 10276 82348 10332
rect 79828 9604 79884 9660
rect 80612 9156 80668 9212
rect 79716 8596 79772 8652
rect 79940 8708 79996 8764
rect 78708 7252 78764 7308
rect 78876 7252 78932 7308
rect 79436 7642 79492 7644
rect 79436 7590 79438 7642
rect 79438 7590 79490 7642
rect 79490 7590 79492 7642
rect 79436 7588 79492 7590
rect 78092 6468 78148 6524
rect 77364 5012 77420 5068
rect 77700 4564 77756 4620
rect 77028 3892 77084 3948
rect 77364 3946 77420 3948
rect 77364 3894 77366 3946
rect 77366 3894 77418 3946
rect 77418 3894 77420 3946
rect 77364 3892 77420 3894
rect 77812 3444 77868 3500
rect 76916 2996 76972 3052
rect 76692 1316 76748 1372
rect 76692 980 76748 1036
rect 76580 868 76636 924
rect 76692 810 76748 812
rect 76692 758 76694 810
rect 76694 758 76746 810
rect 76746 758 76748 810
rect 76692 756 76748 758
rect 77252 756 77308 812
rect 77140 532 77196 588
rect 78036 3444 78092 3500
rect 78260 4564 78316 4620
rect 78260 4340 78316 4396
rect 78260 4116 78316 4172
rect 78484 6356 78540 6412
rect 78596 6804 78652 6860
rect 79268 7028 79324 7084
rect 79268 6692 79324 6748
rect 78820 6580 78876 6636
rect 79828 7028 79884 7084
rect 79828 6804 79884 6860
rect 78484 4900 78540 4956
rect 79268 4900 79324 4956
rect 79044 4340 79100 4396
rect 79492 4452 79548 4508
rect 78596 4004 78652 4060
rect 79380 4004 79436 4060
rect 78260 3556 78316 3612
rect 78596 3444 78652 3500
rect 79380 3556 79436 3612
rect 79156 3444 79212 3500
rect 78484 3220 78540 3276
rect 79716 4452 79772 4508
rect 80724 8932 80780 8988
rect 80052 8090 80108 8092
rect 80052 8038 80054 8090
rect 80054 8038 80106 8090
rect 80106 8038 80108 8090
rect 80052 8036 80108 8038
rect 80388 8090 80444 8092
rect 80388 8038 80390 8090
rect 80390 8038 80442 8090
rect 80442 8038 80444 8090
rect 80388 8036 80444 8038
rect 80052 6916 80108 6972
rect 80164 7252 80220 7308
rect 80276 7364 80332 7420
rect 80500 7306 80556 7308
rect 80500 7254 80502 7306
rect 80502 7254 80554 7306
rect 80554 7254 80556 7306
rect 80500 7252 80556 7254
rect 80276 6356 80332 6412
rect 80500 6356 80556 6412
rect 80052 5124 80108 5180
rect 80500 5572 80556 5628
rect 80108 4954 80164 4956
rect 80108 4902 80110 4954
rect 80110 4902 80162 4954
rect 80162 4902 80164 4954
rect 80108 4900 80164 4902
rect 80052 4116 80108 4172
rect 79940 3556 79996 3612
rect 79940 2996 79996 3052
rect 79828 2324 79884 2380
rect 78708 1316 78764 1372
rect 79492 1428 79548 1484
rect 79044 1316 79100 1372
rect 78596 644 78652 700
rect 80276 3780 80332 3836
rect 80388 3444 80444 3500
rect 80164 1316 80220 1372
rect 80164 868 80220 924
rect 81060 9604 81116 9660
rect 81284 9940 81340 9996
rect 82180 10164 82236 10220
rect 82704 10218 82760 10220
rect 82704 10166 82706 10218
rect 82706 10166 82758 10218
rect 82758 10166 82760 10218
rect 82704 10164 82760 10166
rect 82808 10218 82864 10220
rect 82808 10166 82810 10218
rect 82810 10166 82862 10218
rect 82862 10166 82864 10218
rect 82808 10164 82864 10166
rect 82912 10218 82968 10220
rect 82912 10166 82914 10218
rect 82914 10166 82966 10218
rect 82966 10166 82968 10218
rect 82912 10164 82968 10166
rect 83188 10164 83244 10220
rect 83748 10276 83804 10332
rect 84308 9940 84364 9996
rect 81396 9604 81452 9660
rect 81620 9604 81676 9660
rect 83916 9658 83972 9660
rect 83916 9606 83918 9658
rect 83918 9606 83970 9658
rect 83970 9606 83972 9658
rect 83916 9604 83972 9606
rect 84084 9604 84140 9660
rect 84644 10724 84700 10780
rect 84644 9380 84700 9436
rect 82292 9156 82348 9212
rect 82516 9210 82572 9212
rect 82516 9158 82518 9210
rect 82518 9158 82570 9210
rect 82570 9158 82572 9210
rect 82516 9156 82572 9158
rect 81060 8932 81116 8988
rect 85092 10836 85148 10892
rect 82180 8932 82236 8988
rect 81508 8820 81564 8876
rect 82516 8596 82572 8652
rect 82704 8650 82760 8652
rect 82704 8598 82706 8650
rect 82706 8598 82758 8650
rect 82758 8598 82760 8650
rect 82704 8596 82760 8598
rect 82808 8650 82864 8652
rect 82808 8598 82810 8650
rect 82810 8598 82862 8650
rect 82862 8598 82864 8650
rect 82808 8596 82864 8598
rect 82912 8650 82968 8652
rect 82912 8598 82914 8650
rect 82914 8598 82966 8650
rect 82966 8598 82968 8650
rect 82912 8596 82968 8598
rect 83076 8596 83132 8652
rect 81284 8148 81340 8204
rect 81172 7252 81228 7308
rect 80836 4900 80892 4956
rect 80724 3780 80780 3836
rect 80948 3668 81004 3724
rect 80836 2324 80892 2380
rect 80948 1876 81004 1932
rect 81844 8260 81900 8316
rect 81732 8148 81788 8204
rect 81284 4900 81340 4956
rect 81284 3220 81340 3276
rect 81396 3444 81452 3500
rect 81620 5460 81676 5516
rect 82068 8260 82124 8316
rect 84252 8986 84308 8988
rect 84252 8934 84254 8986
rect 84254 8934 84306 8986
rect 84306 8934 84308 8986
rect 84252 8932 84308 8934
rect 84700 8708 84756 8764
rect 84868 8708 84924 8764
rect 83748 8596 83804 8652
rect 85988 10836 86044 10892
rect 86660 13076 86716 13132
rect 86212 10836 86268 10892
rect 86996 11508 87052 11564
rect 87220 11508 87276 11564
rect 86436 10836 86492 10892
rect 86548 10724 86604 10780
rect 86100 10052 86156 10108
rect 85540 9156 85596 9212
rect 85932 9658 85988 9660
rect 85932 9606 85934 9658
rect 85934 9606 85986 9658
rect 85986 9606 85988 9658
rect 85932 9604 85988 9606
rect 86436 9658 86492 9660
rect 86436 9606 86438 9658
rect 86438 9606 86490 9658
rect 86490 9606 86492 9658
rect 86436 9604 86492 9606
rect 86772 10052 86828 10108
rect 88676 13076 88732 13132
rect 87668 9940 87724 9996
rect 87780 12516 87836 12572
rect 87332 9604 87388 9660
rect 87220 9156 87276 9212
rect 85652 8932 85708 8988
rect 85652 8596 85708 8652
rect 86212 8708 86268 8764
rect 85932 8372 85988 8428
rect 86100 8372 86156 8428
rect 82180 8036 82236 8092
rect 84084 7924 84140 7980
rect 83300 7588 83356 7644
rect 85316 8260 85372 8316
rect 84420 8036 84476 8092
rect 85260 7924 85316 7980
rect 81844 6468 81900 6524
rect 82292 7140 82348 7196
rect 83636 7140 83692 7196
rect 82704 7082 82760 7084
rect 82704 7030 82706 7082
rect 82706 7030 82758 7082
rect 82758 7030 82760 7082
rect 82704 7028 82760 7030
rect 82808 7082 82864 7084
rect 82808 7030 82810 7082
rect 82810 7030 82862 7082
rect 82862 7030 82864 7082
rect 82808 7028 82864 7030
rect 82912 7082 82968 7084
rect 82912 7030 82914 7082
rect 82914 7030 82966 7082
rect 82966 7030 82968 7082
rect 82912 7028 82968 7030
rect 83412 6916 83468 6972
rect 84420 7588 84476 7644
rect 85820 7924 85876 7980
rect 85708 7700 85764 7756
rect 84420 7306 84476 7308
rect 84420 7254 84422 7306
rect 84422 7254 84474 7306
rect 84474 7254 84476 7306
rect 84420 7252 84476 7254
rect 84308 6916 84364 6972
rect 82628 6804 82684 6860
rect 84196 6804 84252 6860
rect 82516 6580 82572 6636
rect 82740 6692 82796 6748
rect 82292 6468 82348 6524
rect 82180 6356 82236 6412
rect 82180 5684 82236 5740
rect 83188 6020 83244 6076
rect 83748 6692 83804 6748
rect 82740 5684 82796 5740
rect 82516 5460 82572 5516
rect 82704 5514 82760 5516
rect 82704 5462 82706 5514
rect 82706 5462 82758 5514
rect 82758 5462 82760 5514
rect 82704 5460 82760 5462
rect 82808 5514 82864 5516
rect 82808 5462 82810 5514
rect 82810 5462 82862 5514
rect 82862 5462 82864 5514
rect 82808 5460 82864 5462
rect 82912 5514 82968 5516
rect 82912 5462 82914 5514
rect 82914 5462 82966 5514
rect 82966 5462 82968 5514
rect 82912 5460 82968 5462
rect 82292 5124 82348 5180
rect 83188 5124 83244 5180
rect 81956 4900 82012 4956
rect 82068 4788 82124 4844
rect 82292 4676 82348 4732
rect 82180 4228 82236 4284
rect 82516 3668 82572 3724
rect 81172 2324 81228 2380
rect 81620 2324 81676 2380
rect 81172 1652 81228 1708
rect 80724 980 80780 1036
rect 81732 1988 81788 2044
rect 81172 868 81228 924
rect 81396 868 81452 924
rect 81508 810 81564 812
rect 79044 420 79100 476
rect 81508 758 81510 810
rect 81510 758 81562 810
rect 81562 758 81564 810
rect 81508 756 81564 758
rect 81732 868 81788 924
rect 82068 2212 82124 2268
rect 81956 1876 82012 1932
rect 82628 3444 82684 3500
rect 82740 3220 82796 3276
rect 82404 2772 82460 2828
rect 82628 2772 82684 2828
rect 82292 1876 82348 1932
rect 82516 2100 82572 2156
rect 82628 1316 82684 1372
rect 83076 4676 83132 4732
rect 83300 4676 83356 4732
rect 83748 5796 83804 5852
rect 84084 6468 84140 6524
rect 84308 6580 84364 6636
rect 83972 6132 84028 6188
rect 83524 4228 83580 4284
rect 83636 4900 83692 4956
rect 83188 3668 83244 3724
rect 83916 5460 83972 5516
rect 84196 4004 84252 4060
rect 84476 5684 84532 5740
rect 84476 5460 84532 5516
rect 84420 4004 84476 4060
rect 83972 2772 84028 2828
rect 83860 2266 83916 2268
rect 83860 2214 83862 2266
rect 83862 2214 83914 2266
rect 83914 2214 83916 2266
rect 83860 2212 83916 2214
rect 83972 1764 84028 1820
rect 84644 4340 84700 4396
rect 84420 1876 84476 1932
rect 86100 7588 86156 7644
rect 84868 7252 84924 7308
rect 85372 7252 85428 7308
rect 84980 7028 85036 7084
rect 85764 7028 85820 7084
rect 84868 6132 84924 6188
rect 84868 5908 84924 5964
rect 84924 5124 84980 5180
rect 84924 4954 84980 4956
rect 84924 4902 84926 4954
rect 84926 4902 84978 4954
rect 84978 4902 84980 4954
rect 84924 4900 84980 4902
rect 86212 6580 86268 6636
rect 86212 6356 86268 6412
rect 85540 5908 85596 5964
rect 85428 5796 85484 5852
rect 85204 5348 85260 5404
rect 85428 5348 85484 5404
rect 85820 5850 85876 5852
rect 85820 5798 85822 5850
rect 85822 5798 85874 5850
rect 85874 5798 85876 5850
rect 85820 5796 85876 5798
rect 84868 2548 84924 2604
rect 84868 2100 84924 2156
rect 85428 4676 85484 4732
rect 85652 4564 85708 4620
rect 85652 3780 85708 3836
rect 85652 2996 85708 3052
rect 85988 4900 86044 4956
rect 86436 8484 86492 8540
rect 86436 7588 86492 7644
rect 86548 7924 86604 7980
rect 86212 4564 86268 4620
rect 85988 4340 86044 4396
rect 85876 4058 85932 4060
rect 85876 4006 85878 4058
rect 85878 4006 85930 4058
rect 85930 4006 85932 4058
rect 85876 4004 85932 4006
rect 85764 2660 85820 2716
rect 86660 5012 86716 5068
rect 86548 4564 86604 4620
rect 86436 4004 86492 4060
rect 86548 4340 86604 4396
rect 86548 3780 86604 3836
rect 85988 2660 86044 2716
rect 85988 2212 86044 2268
rect 86100 2100 86156 2156
rect 84420 980 84476 1036
rect 85428 1652 85484 1708
rect 85652 1652 85708 1708
rect 85652 1316 85708 1372
rect 85540 980 85596 1036
rect 86996 6132 87052 6188
rect 86996 5796 87052 5852
rect 87556 9492 87612 9548
rect 87444 9156 87500 9212
rect 89460 12964 89516 13020
rect 89124 12292 89180 12348
rect 88788 12180 88844 12236
rect 88788 11396 88844 11452
rect 89908 12068 89964 12124
rect 89012 11956 89068 12012
rect 89348 11284 89404 11340
rect 90356 13412 90412 13468
rect 98084 14756 98140 14812
rect 91028 13748 91084 13804
rect 88676 9604 88732 9660
rect 88900 9940 88956 9996
rect 88900 9604 88956 9660
rect 87892 9492 87948 9548
rect 87724 9210 87780 9212
rect 87724 9158 87726 9210
rect 87726 9158 87778 9210
rect 87778 9158 87780 9210
rect 87724 9156 87780 9158
rect 90692 9828 90748 9884
rect 88116 8820 88172 8876
rect 88900 8596 88956 8652
rect 88452 8484 88508 8540
rect 88508 8260 88564 8316
rect 87556 8148 87612 8204
rect 87556 7924 87612 7980
rect 87332 6132 87388 6188
rect 87668 8036 87724 8092
rect 88396 7812 88452 7868
rect 88004 7700 88060 7756
rect 89068 7924 89124 7980
rect 89236 8036 89292 8092
rect 88676 7588 88732 7644
rect 88116 7476 88172 7532
rect 87668 6916 87724 6972
rect 87780 7028 87836 7084
rect 87780 6692 87836 6748
rect 87668 6580 87724 6636
rect 88004 6580 88060 6636
rect 87220 5796 87276 5852
rect 87108 5012 87164 5068
rect 86884 4004 86940 4060
rect 86996 4564 87052 4620
rect 86884 3780 86940 3836
rect 86884 1652 86940 1708
rect 87108 2660 87164 2716
rect 87108 2436 87164 2492
rect 87948 5850 88004 5852
rect 87948 5798 87950 5850
rect 87950 5798 88002 5850
rect 88002 5798 88004 5850
rect 87948 5796 88004 5798
rect 87780 5684 87836 5740
rect 87948 5012 88004 5068
rect 88340 6916 88396 6972
rect 89124 6916 89180 6972
rect 88564 5796 88620 5852
rect 88564 5348 88620 5404
rect 88788 5796 88844 5852
rect 88228 5012 88284 5068
rect 87892 2884 87948 2940
rect 87444 1146 87500 1148
rect 87444 1094 87446 1146
rect 87446 1094 87498 1146
rect 87498 1094 87500 1146
rect 87444 1092 87500 1094
rect 88340 4004 88396 4060
rect 89572 7924 89628 7980
rect 89460 5796 89516 5852
rect 89572 4900 89628 4956
rect 88452 1764 88508 1820
rect 88564 3780 88620 3836
rect 88340 1652 88396 1708
rect 88676 2772 88732 2828
rect 88788 2212 88844 2268
rect 88900 1428 88956 1484
rect 89236 2212 89292 2268
rect 89012 1316 89068 1372
rect 90412 8708 90468 8764
rect 89908 8314 89964 8316
rect 89908 8262 89910 8314
rect 89910 8262 89962 8314
rect 89962 8262 89964 8314
rect 89908 8260 89964 8262
rect 90356 8148 90412 8204
rect 90356 7700 90412 7756
rect 91476 12964 91532 13020
rect 91476 12740 91532 12796
rect 91924 12516 91980 12572
rect 92708 13860 92764 13916
rect 92036 11396 92092 11452
rect 91476 11284 91532 11340
rect 91140 10612 91196 10668
rect 91364 10836 91420 10892
rect 91364 10612 91420 10668
rect 92932 12516 92988 12572
rect 93492 12292 93548 12348
rect 94164 12292 94220 12348
rect 93828 11844 93884 11900
rect 92820 11060 92876 11116
rect 93044 11060 93100 11116
rect 91812 10724 91868 10780
rect 91476 10164 91532 10220
rect 91252 9716 91308 9772
rect 91252 9492 91308 9548
rect 91700 9492 91756 9548
rect 91196 8484 91252 8540
rect 91084 8090 91140 8092
rect 91084 8038 91086 8090
rect 91086 8038 91138 8090
rect 91138 8038 91140 8090
rect 91084 8036 91140 8038
rect 90804 7924 90860 7980
rect 91532 7700 91588 7756
rect 90468 7252 90524 7308
rect 90468 6468 90524 6524
rect 90244 6356 90300 6412
rect 91252 7476 91308 7532
rect 90580 6356 90636 6412
rect 90748 6916 90804 6972
rect 90860 6634 90916 6636
rect 90860 6582 90862 6634
rect 90862 6582 90914 6634
rect 90914 6582 90916 6634
rect 90860 6580 90916 6582
rect 89908 5124 89964 5180
rect 90580 5124 90636 5180
rect 89908 4900 89964 4956
rect 89796 3220 89852 3276
rect 91252 7140 91308 7196
rect 91476 7140 91532 7196
rect 91252 6916 91308 6972
rect 91476 6916 91532 6972
rect 91364 6692 91420 6748
rect 91420 6356 91476 6412
rect 91196 5684 91252 5740
rect 91196 5178 91252 5180
rect 91196 5126 91198 5178
rect 91198 5126 91250 5178
rect 91250 5126 91252 5178
rect 91196 5124 91252 5126
rect 91364 5124 91420 5180
rect 91028 4676 91084 4732
rect 90020 4340 90076 4396
rect 90020 4116 90076 4172
rect 90580 2996 90636 3052
rect 90132 2324 90188 2380
rect 89796 1316 89852 1372
rect 90580 1370 90636 1372
rect 90580 1318 90582 1370
rect 90582 1318 90634 1370
rect 90634 1318 90636 1370
rect 90580 1316 90636 1318
rect 89908 1204 89964 1260
rect 91252 4452 91308 4508
rect 91756 7140 91812 7196
rect 91924 4900 91980 4956
rect 91700 4340 91756 4396
rect 92820 6468 92876 6524
rect 92372 6132 92428 6188
rect 92148 4228 92204 4284
rect 91364 3444 91420 3500
rect 91588 3780 91644 3836
rect 91476 3162 91532 3164
rect 91476 3110 91478 3162
rect 91478 3110 91530 3162
rect 91530 3110 91532 3162
rect 91476 3108 91532 3110
rect 92036 3332 92092 3388
rect 91924 3050 91980 3052
rect 91924 2998 91926 3050
rect 91926 2998 91978 3050
rect 91978 2998 91980 3050
rect 91924 2996 91980 2998
rect 93268 8484 93324 8540
rect 94276 10052 94332 10108
rect 93940 8820 93996 8876
rect 93268 8036 93324 8092
rect 92148 2100 92204 2156
rect 92372 1092 92428 1148
rect 93828 6132 93884 6188
rect 93940 5348 93996 5404
rect 93380 4564 93436 4620
rect 94836 10276 94892 10332
rect 94724 8148 94780 8204
rect 95340 8986 95396 8988
rect 95340 8934 95342 8986
rect 95342 8934 95394 8986
rect 95394 8934 95396 8986
rect 95340 8932 95396 8934
rect 95172 5572 95228 5628
rect 94780 5348 94836 5404
rect 95956 8932 96012 8988
rect 95396 7924 95452 7980
rect 95732 8036 95788 8092
rect 95620 7642 95676 7644
rect 95620 7590 95622 7642
rect 95622 7590 95674 7642
rect 95674 7590 95676 7642
rect 95620 7588 95676 7590
rect 95284 5236 95340 5292
rect 95172 4004 95228 4060
rect 95284 4228 95340 4284
rect 94164 2996 94220 3052
rect 94388 2996 94444 3052
rect 94164 2378 94220 2380
rect 94164 2326 94166 2378
rect 94166 2326 94218 2378
rect 94218 2326 94220 2378
rect 94164 2324 94220 2326
rect 94612 2100 94668 2156
rect 93380 1764 93436 1820
rect 95732 2266 95788 2268
rect 95732 2214 95734 2266
rect 95734 2214 95786 2266
rect 95786 2214 95788 2266
rect 95732 2212 95788 2214
rect 96292 8484 96348 8540
rect 96068 7924 96124 7980
rect 97076 12516 97132 12572
rect 97524 13972 97580 14028
rect 100436 14756 100492 14812
rect 97412 12404 97468 12460
rect 96740 10948 96796 11004
rect 96852 11396 96908 11452
rect 96628 10724 96684 10780
rect 96852 10724 96908 10780
rect 97300 11396 97356 11452
rect 97300 10052 97356 10108
rect 97412 9604 97468 9660
rect 98084 11956 98140 12012
rect 98308 11732 98364 11788
rect 98196 11060 98252 11116
rect 96404 8036 96460 8092
rect 97636 7924 97692 7980
rect 97524 7364 97580 7420
rect 97692 7418 97748 7420
rect 97692 7366 97694 7418
rect 97694 7366 97746 7418
rect 97746 7366 97748 7418
rect 97692 7364 97748 7366
rect 96068 6468 96124 6524
rect 96852 7140 96908 7196
rect 96068 5124 96124 5180
rect 96180 4676 96236 4732
rect 96068 2436 96124 2492
rect 96404 4676 96460 4732
rect 96404 4228 96460 4284
rect 96292 3220 96348 3276
rect 96740 4004 96796 4060
rect 95956 2212 96012 2268
rect 95956 1652 96012 1708
rect 96292 980 96348 1036
rect 96516 2100 96572 2156
rect 96628 1764 96684 1820
rect 97412 6132 97468 6188
rect 97412 5124 97468 5180
rect 96964 5012 97020 5068
rect 96964 3780 97020 3836
rect 97076 4900 97132 4956
rect 97972 5460 98028 5516
rect 98028 5178 98084 5180
rect 98028 5126 98030 5178
rect 98030 5126 98082 5178
rect 98082 5126 98084 5178
rect 98028 5124 98084 5126
rect 98420 10948 98476 11004
rect 98644 12180 98700 12236
rect 98980 13524 99036 13580
rect 98532 10052 98588 10108
rect 98532 8932 98588 8988
rect 98364 6356 98420 6412
rect 98364 6132 98420 6188
rect 97860 3220 97916 3276
rect 97972 3668 98028 3724
rect 97636 2100 97692 2156
rect 97412 1764 97468 1820
rect 97636 1764 97692 1820
rect 97412 980 97468 1036
rect 85764 308 85820 364
rect 97300 308 97356 364
rect 99204 13524 99260 13580
rect 99204 12068 99260 12124
rect 99652 13860 99708 13916
rect 101332 14756 101388 14812
rect 101108 14532 101164 14588
rect 99316 11620 99372 11676
rect 100436 12404 100492 12460
rect 100324 12068 100380 12124
rect 100212 11732 100268 11788
rect 99540 11620 99596 11676
rect 99204 10948 99260 11004
rect 98924 10052 98980 10108
rect 99092 9380 99148 9436
rect 99204 7812 99260 7868
rect 99092 7364 99148 7420
rect 101780 12740 101836 12796
rect 102676 14868 102732 14924
rect 102564 14532 102620 14588
rect 104020 14196 104076 14252
rect 102004 12740 102060 12796
rect 101556 12404 101612 12460
rect 100548 12068 100604 12124
rect 101892 11732 101948 11788
rect 100212 11172 100268 11228
rect 100436 11172 100492 11228
rect 100548 11060 100604 11116
rect 100772 10836 100828 10892
rect 100212 10724 100268 10780
rect 101444 10724 101500 10780
rect 99652 10612 99708 10668
rect 100436 10612 100492 10668
rect 99876 10164 99932 10220
rect 99708 9380 99764 9436
rect 99540 8260 99596 8316
rect 100884 9492 100940 9548
rect 101220 9380 101276 9436
rect 99316 6916 99372 6972
rect 98644 6468 98700 6524
rect 99204 5012 99260 5068
rect 99428 4452 99484 4508
rect 99204 3668 99260 3724
rect 101668 9044 101724 9100
rect 99876 8596 99932 8652
rect 100100 8260 100156 8316
rect 100436 8596 100492 8652
rect 99876 7812 99932 7868
rect 100100 7476 100156 7532
rect 100100 6916 100156 6972
rect 100212 6468 100268 6524
rect 100100 4900 100156 4956
rect 100436 5796 100492 5852
rect 100548 8260 100604 8316
rect 100324 4900 100380 4956
rect 100436 5572 100492 5628
rect 100212 4340 100268 4396
rect 99540 4058 99596 4060
rect 99540 4006 99542 4058
rect 99542 4006 99594 4058
rect 99594 4006 99596 4058
rect 99540 4004 99596 4006
rect 99988 4004 100044 4060
rect 99092 3556 99148 3612
rect 99876 3556 99932 3612
rect 98644 2548 98700 2604
rect 99316 2548 99372 2604
rect 99764 2548 99820 2604
rect 99540 2212 99596 2268
rect 98868 1988 98924 2044
rect 99428 1316 99484 1372
rect 99876 1764 99932 1820
rect 99988 1204 100044 1260
rect 100100 1652 100156 1708
rect 100772 8260 100828 8316
rect 101892 9044 101948 9100
rect 101220 8260 101276 8316
rect 101444 8260 101500 8316
rect 101444 7924 101500 7980
rect 101780 8036 101836 8092
rect 100772 7140 100828 7196
rect 101052 6522 101108 6524
rect 101052 6470 101054 6522
rect 101054 6470 101106 6522
rect 101106 6470 101108 6522
rect 101052 6468 101108 6470
rect 101612 6522 101668 6524
rect 101612 6470 101614 6522
rect 101614 6470 101666 6522
rect 101666 6470 101668 6522
rect 101612 6468 101668 6470
rect 100660 6132 100716 6188
rect 100660 5796 100716 5852
rect 100996 5236 101052 5292
rect 100772 3780 100828 3836
rect 101724 5850 101780 5852
rect 101724 5798 101726 5850
rect 101726 5798 101778 5850
rect 101778 5798 101780 5850
rect 101724 5796 101780 5798
rect 101556 5012 101612 5068
rect 101780 5012 101836 5068
rect 103012 13300 103068 13356
rect 103348 13076 103404 13132
rect 104244 12852 104300 12908
rect 104356 12964 104412 13020
rect 103124 12292 103180 12348
rect 102900 11284 102956 11340
rect 103460 12068 103516 12124
rect 104132 12292 104188 12348
rect 104244 12516 104300 12572
rect 104132 12068 104188 12124
rect 104020 11898 104076 11900
rect 104020 11846 104022 11898
rect 104022 11846 104074 11898
rect 104074 11846 104076 11898
rect 104020 11844 104076 11846
rect 103796 10052 103852 10108
rect 103460 9940 103516 9996
rect 102956 9770 103012 9772
rect 102956 9718 102958 9770
rect 102958 9718 103010 9770
rect 103010 9718 103012 9770
rect 102956 9716 103012 9718
rect 102228 9492 102284 9548
rect 102452 8484 102508 8540
rect 102116 6580 102172 6636
rect 102564 8036 102620 8092
rect 101332 4900 101388 4956
rect 101780 4676 101836 4732
rect 101444 4340 101500 4396
rect 101108 3892 101164 3948
rect 101220 4004 101276 4060
rect 100884 3444 100940 3500
rect 100996 3332 101052 3388
rect 100660 1540 100716 1596
rect 101108 3108 101164 3164
rect 101220 1652 101276 1708
rect 101332 3892 101388 3948
rect 100996 1316 101052 1372
rect 100212 1204 100268 1260
rect 101556 3108 101612 3164
rect 102004 4676 102060 4732
rect 101892 4564 101948 4620
rect 102900 8932 102956 8988
rect 103684 9770 103740 9772
rect 103684 9718 103686 9770
rect 103686 9718 103738 9770
rect 103738 9718 103740 9770
rect 103684 9716 103740 9718
rect 103460 8932 103516 8988
rect 102676 7364 102732 7420
rect 103348 7812 103404 7868
rect 104020 10052 104076 10108
rect 104692 12852 104748 12908
rect 113652 14756 113708 14812
rect 104468 10948 104524 11004
rect 105364 12852 105420 12908
rect 105140 9716 105196 9772
rect 105252 12516 105308 12572
rect 104356 9380 104412 9436
rect 103908 8260 103964 8316
rect 104076 8090 104132 8092
rect 104076 8038 104078 8090
rect 104078 8038 104130 8090
rect 104130 8038 104132 8090
rect 104076 8036 104132 8038
rect 103348 7252 103404 7308
rect 102788 6916 102844 6972
rect 103012 7140 103068 7196
rect 103012 6916 103068 6972
rect 103796 6804 103852 6860
rect 103124 6468 103180 6524
rect 103684 5796 103740 5852
rect 102676 5460 102732 5516
rect 102004 3220 102060 3276
rect 101780 2212 101836 2268
rect 101556 1988 101612 2044
rect 102452 2436 102508 2492
rect 102004 1988 102060 2044
rect 102340 2324 102396 2380
rect 102676 3332 102732 3388
rect 102900 3332 102956 3388
rect 102676 2772 102732 2828
rect 103684 2548 103740 2604
rect 103684 2324 103740 2380
rect 102900 2212 102956 2268
rect 103012 1764 103068 1820
rect 103124 1652 103180 1708
rect 104132 7476 104188 7532
rect 104972 7476 105028 7532
rect 104020 7028 104076 7084
rect 104132 7140 104188 7196
rect 104020 6692 104076 6748
rect 104132 5796 104188 5852
rect 104020 5124 104076 5180
rect 104356 5796 104412 5852
rect 103908 2324 103964 2380
rect 104916 5796 104972 5852
rect 105028 6468 105084 6524
rect 105588 10948 105644 11004
rect 105364 6468 105420 6524
rect 105364 5684 105420 5740
rect 105924 11732 105980 11788
rect 106372 12068 106428 12124
rect 105812 10388 105868 10444
rect 105700 8372 105756 8428
rect 105700 6858 105756 6860
rect 105700 6806 105702 6858
rect 105702 6806 105754 6858
rect 105754 6806 105756 6858
rect 105700 6804 105756 6806
rect 105700 6356 105756 6412
rect 105700 5684 105756 5740
rect 107380 12740 107436 12796
rect 107940 12740 107996 12796
rect 106596 11956 106652 12012
rect 106484 11284 106540 11340
rect 106484 10276 106540 10332
rect 106708 5124 106764 5180
rect 109172 12906 109228 12908
rect 109172 12854 109174 12906
rect 109174 12854 109226 12906
rect 109226 12854 109228 12906
rect 109172 12852 109228 12854
rect 108948 11956 109004 12012
rect 109620 12404 109676 12460
rect 109844 12404 109900 12460
rect 109620 12180 109676 12236
rect 109508 11508 109564 11564
rect 108836 10724 108892 10780
rect 109396 10612 109452 10668
rect 108164 9658 108220 9660
rect 108164 9606 108166 9658
rect 108166 9606 108218 9658
rect 108218 9606 108220 9658
rect 108164 9604 108220 9606
rect 108836 9828 108892 9884
rect 109060 9882 109116 9884
rect 109060 9830 109062 9882
rect 109062 9830 109114 9882
rect 109114 9830 109116 9882
rect 109060 9828 109116 9830
rect 109284 9380 109340 9436
rect 110964 11508 111020 11564
rect 110852 11284 110908 11340
rect 111636 10388 111692 10444
rect 110180 9940 110236 9996
rect 107268 8260 107324 8316
rect 107884 8314 107940 8316
rect 107884 8262 107886 8314
rect 107886 8262 107938 8314
rect 107938 8262 107940 8314
rect 107884 8260 107940 8262
rect 107828 6916 107884 6972
rect 107548 5124 107604 5180
rect 106932 3892 106988 3948
rect 105812 1204 105868 1260
rect 105924 980 105980 1036
rect 106148 1034 106204 1036
rect 106148 982 106150 1034
rect 106150 982 106202 1034
rect 106202 982 106204 1034
rect 106148 980 106204 982
rect 106820 2436 106876 2492
rect 106372 1034 106428 1036
rect 106372 982 106374 1034
rect 106374 982 106426 1034
rect 106426 982 106428 1034
rect 106372 980 106428 982
rect 107604 3220 107660 3276
rect 107492 2660 107548 2716
rect 108500 6580 108556 6636
rect 108500 5908 108556 5964
rect 107716 2660 107772 2716
rect 109172 8260 109228 8316
rect 109868 9434 109924 9436
rect 109868 9382 109870 9434
rect 109870 9382 109922 9434
rect 109922 9382 109924 9434
rect 109868 9380 109924 9382
rect 109972 9434 110028 9436
rect 109972 9382 109974 9434
rect 109974 9382 110026 9434
rect 110026 9382 110028 9434
rect 109972 9380 110028 9382
rect 110076 9434 110132 9436
rect 110076 9382 110078 9434
rect 110078 9382 110130 9434
rect 110130 9382 110132 9434
rect 110076 9380 110132 9382
rect 110628 9044 110684 9100
rect 109620 8260 109676 8316
rect 110460 8260 110516 8316
rect 109868 7866 109924 7868
rect 109868 7814 109870 7866
rect 109870 7814 109922 7866
rect 109922 7814 109924 7866
rect 109868 7812 109924 7814
rect 109972 7866 110028 7868
rect 109972 7814 109974 7866
rect 109974 7814 110026 7866
rect 110026 7814 110028 7866
rect 109972 7812 110028 7814
rect 110076 7866 110132 7868
rect 110076 7814 110078 7866
rect 110078 7814 110130 7866
rect 110130 7814 110132 7866
rect 110076 7812 110132 7814
rect 110964 9492 111020 9548
rect 110964 9156 111020 9212
rect 111188 9044 111244 9100
rect 110740 8036 110796 8092
rect 110908 8090 110964 8092
rect 110908 8038 110910 8090
rect 110910 8038 110962 8090
rect 110962 8038 110964 8090
rect 110908 8036 110964 8038
rect 109508 7700 109564 7756
rect 111076 7700 111132 7756
rect 111860 11508 111916 11564
rect 111748 7924 111804 7980
rect 109172 6916 109228 6972
rect 110180 6804 110236 6860
rect 110068 6580 110124 6636
rect 109868 6298 109924 6300
rect 109868 6246 109870 6298
rect 109870 6246 109922 6298
rect 109922 6246 109924 6298
rect 109868 6244 109924 6246
rect 109972 6298 110028 6300
rect 109972 6246 109974 6298
rect 109974 6246 110026 6298
rect 110026 6246 110028 6298
rect 109972 6244 110028 6246
rect 110076 6298 110132 6300
rect 110076 6246 110078 6298
rect 110078 6246 110130 6298
rect 110130 6246 110132 6298
rect 110076 6244 110132 6246
rect 109732 6132 109788 6188
rect 110516 6132 110572 6188
rect 109732 5908 109788 5964
rect 110068 5908 110124 5964
rect 109732 5572 109788 5628
rect 109396 4676 109452 4732
rect 110068 5012 110124 5068
rect 110292 5012 110348 5068
rect 111300 6468 111356 6524
rect 111636 7028 111692 7084
rect 110516 4900 110572 4956
rect 110964 4900 111020 4956
rect 111468 5012 111524 5068
rect 113652 13748 113708 13804
rect 113764 14532 113820 14588
rect 113876 13748 113932 13804
rect 112084 12516 112140 12572
rect 115220 14868 115276 14924
rect 114884 14474 114940 14476
rect 114884 14422 114886 14474
rect 114886 14422 114938 14474
rect 114938 14422 114940 14474
rect 114884 14420 114940 14422
rect 115220 14420 115276 14476
rect 115444 13972 115500 14028
rect 114212 12516 114268 12572
rect 112308 11060 112364 11116
rect 112420 12180 112476 12236
rect 111972 6132 112028 6188
rect 114212 12180 114268 12236
rect 113092 11732 113148 11788
rect 112756 11508 112812 11564
rect 112756 11172 112812 11228
rect 112532 10052 112588 10108
rect 112532 8036 112588 8092
rect 113092 8036 113148 8092
rect 113428 11284 113484 11340
rect 113204 7588 113260 7644
rect 113316 11060 113372 11116
rect 113428 10948 113484 11004
rect 114324 11620 114380 11676
rect 113652 8148 113708 8204
rect 113652 7812 113708 7868
rect 113764 7588 113820 7644
rect 112308 6132 112364 6188
rect 112644 5012 112700 5068
rect 109868 4730 109924 4732
rect 109868 4678 109870 4730
rect 109870 4678 109922 4730
rect 109922 4678 109924 4730
rect 109868 4676 109924 4678
rect 109972 4730 110028 4732
rect 109972 4678 109974 4730
rect 109974 4678 110026 4730
rect 110026 4678 110028 4730
rect 109972 4676 110028 4678
rect 110076 4730 110132 4732
rect 110076 4678 110078 4730
rect 110078 4678 110130 4730
rect 110130 4678 110132 4730
rect 110076 4676 110132 4678
rect 110516 4676 110572 4732
rect 110516 4340 110572 4396
rect 110628 4564 110684 4620
rect 112532 4900 112588 4956
rect 112420 4788 112476 4844
rect 109060 3220 109116 3276
rect 109172 3108 109228 3164
rect 109060 2884 109116 2940
rect 109060 2548 109116 2604
rect 108948 2324 109004 2380
rect 108388 1988 108444 2044
rect 108612 1988 108668 2044
rect 108388 1652 108444 1708
rect 108276 1316 108332 1372
rect 98140 420 98196 476
rect 108276 756 108332 812
rect 109172 1764 109228 1820
rect 109284 1316 109340 1372
rect 110292 2772 110348 2828
rect 109956 1988 110012 2044
rect 110628 2996 110684 3052
rect 111412 1370 111468 1372
rect 111412 1318 111414 1370
rect 111414 1318 111466 1370
rect 111466 1318 111468 1370
rect 111412 1316 111468 1318
rect 111636 1316 111692 1372
rect 110740 1092 110796 1148
rect 112420 3556 112476 3612
rect 112308 3332 112364 3388
rect 112084 756 112140 812
rect 112644 4676 112700 4732
rect 113204 6132 113260 6188
rect 112868 4676 112924 4732
rect 112644 3610 112700 3612
rect 112644 3558 112646 3610
rect 112646 3558 112698 3610
rect 112698 3558 112700 3610
rect 112644 3556 112700 3558
rect 113428 5236 113484 5292
rect 113708 6132 113764 6188
rect 113540 4228 113596 4284
rect 113988 10164 114044 10220
rect 114436 11172 114492 11228
rect 115556 13076 115612 13132
rect 115892 13748 115948 13804
rect 116340 13748 116396 13804
rect 116564 13748 116620 13804
rect 115892 13076 115948 13132
rect 114996 11786 115052 11788
rect 114996 11734 114998 11786
rect 114998 11734 115050 11786
rect 115050 11734 115052 11786
rect 114996 11732 115052 11734
rect 115668 12122 115724 12124
rect 115668 12070 115670 12122
rect 115670 12070 115722 12122
rect 115722 12070 115724 12122
rect 115668 12068 115724 12070
rect 115892 11844 115948 11900
rect 115332 11396 115388 11452
rect 116228 12516 116284 12572
rect 116004 11284 116060 11340
rect 118020 14868 118076 14924
rect 117796 14420 117852 14476
rect 117124 12516 117180 12572
rect 117012 12292 117068 12348
rect 116228 11956 116284 12012
rect 116564 11620 116620 11676
rect 115556 10052 115612 10108
rect 115780 10052 115836 10108
rect 116676 10388 116732 10444
rect 116004 9940 116060 9996
rect 114772 9492 114828 9548
rect 115332 9492 115388 9548
rect 115220 9380 115276 9436
rect 117684 13860 117740 13916
rect 118020 14420 118076 14476
rect 118132 14196 118188 14252
rect 118580 14868 118636 14924
rect 117908 13860 117964 13916
rect 118580 13860 118636 13916
rect 118020 13412 118076 13468
rect 116900 9940 116956 9996
rect 118020 11956 118076 12012
rect 118244 11956 118300 12012
rect 116676 9268 116732 9324
rect 116228 9156 116284 9212
rect 115220 8596 115276 8652
rect 114324 7700 114380 7756
rect 115444 8596 115500 8652
rect 114156 5236 114212 5292
rect 114100 4228 114156 4284
rect 112644 3220 112700 3276
rect 112532 3108 112588 3164
rect 112420 2996 112476 3052
rect 113540 3332 113596 3388
rect 113428 3108 113484 3164
rect 113652 2212 113708 2268
rect 113540 2100 113596 2156
rect 114324 4340 114380 4396
rect 114772 7700 114828 7756
rect 117684 11338 117740 11340
rect 117684 11286 117686 11338
rect 117686 11286 117738 11338
rect 117738 11286 117740 11338
rect 117684 11284 117740 11286
rect 117348 10948 117404 11004
rect 117124 10724 117180 10780
rect 115780 8596 115836 8652
rect 115108 6804 115164 6860
rect 115556 7588 115612 7644
rect 116004 8372 116060 8428
rect 116228 8372 116284 8428
rect 115948 7642 116004 7644
rect 115948 7590 115950 7642
rect 115950 7590 116002 7642
rect 116002 7590 116004 7642
rect 115948 7588 116004 7590
rect 115780 6580 115836 6636
rect 117012 8372 117068 8428
rect 116452 8260 116508 8316
rect 115892 5012 115948 5068
rect 116228 6244 116284 6300
rect 116116 4564 116172 4620
rect 115668 4116 115724 4172
rect 115556 3892 115612 3948
rect 115220 3780 115276 3836
rect 114884 3220 114940 3276
rect 115220 3498 115276 3500
rect 115220 3446 115222 3498
rect 115222 3446 115274 3498
rect 115274 3446 115276 3498
rect 115220 3444 115276 3446
rect 114548 2884 114604 2940
rect 114324 2212 114380 2268
rect 113316 1988 113372 2044
rect 113652 1988 113708 2044
rect 114324 1876 114380 1932
rect 115108 2884 115164 2940
rect 114772 2548 114828 2604
rect 115444 3332 115500 3388
rect 116116 3780 116172 3836
rect 115668 1764 115724 1820
rect 115556 1540 115612 1596
rect 115892 1764 115948 1820
rect 116340 6132 116396 6188
rect 116340 4564 116396 4620
rect 116564 6244 116620 6300
rect 116900 7812 116956 7868
rect 116676 4900 116732 4956
rect 116564 4564 116620 4620
rect 116452 1034 116508 1036
rect 116452 982 116454 1034
rect 116454 982 116506 1034
rect 116506 982 116508 1034
rect 116452 980 116508 982
rect 117684 10666 117740 10668
rect 117684 10614 117686 10666
rect 117686 10614 117738 10666
rect 117738 10614 117740 10666
rect 117684 10612 117740 10614
rect 117572 10388 117628 10444
rect 117460 9828 117516 9884
rect 120148 14868 120204 14924
rect 118804 13188 118860 13244
rect 118580 12292 118636 12348
rect 118468 12068 118524 12124
rect 119252 13524 119308 13580
rect 119364 12964 119420 13020
rect 119700 13076 119756 13132
rect 119140 12180 119196 12236
rect 119364 12180 119420 12236
rect 118468 11898 118524 11900
rect 118468 11846 118470 11898
rect 118470 11846 118522 11898
rect 118522 11846 118524 11898
rect 118468 11844 118524 11846
rect 118804 11732 118860 11788
rect 119028 11732 119084 11788
rect 119252 11284 119308 11340
rect 118580 10052 118636 10108
rect 118580 9716 118636 9772
rect 118804 9716 118860 9772
rect 118356 9380 118412 9436
rect 117572 8484 117628 8540
rect 117460 8260 117516 8316
rect 117908 8148 117964 8204
rect 118132 8148 118188 8204
rect 118468 8036 118524 8092
rect 118580 7924 118636 7980
rect 119252 8932 119308 8988
rect 117460 7140 117516 7196
rect 118020 7476 118076 7532
rect 117012 6692 117068 6748
rect 117124 6804 117180 6860
rect 117796 6692 117852 6748
rect 117684 6580 117740 6636
rect 117684 5908 117740 5964
rect 117348 5236 117404 5292
rect 116900 2826 116956 2828
rect 116900 2774 116902 2826
rect 116902 2774 116954 2826
rect 116954 2774 116956 2826
rect 116900 2772 116956 2774
rect 117124 3108 117180 3164
rect 117236 3220 117292 3276
rect 118916 7364 118972 7420
rect 119028 7588 119084 7644
rect 118132 6692 118188 6748
rect 118412 6692 118468 6748
rect 117460 4452 117516 4508
rect 117908 4452 117964 4508
rect 118468 4004 118524 4060
rect 118244 3668 118300 3724
rect 118020 3444 118076 3500
rect 117572 3220 117628 3276
rect 117236 2772 117292 2828
rect 117236 2154 117292 2156
rect 117236 2102 117238 2154
rect 117238 2102 117290 2154
rect 117290 2102 117292 2154
rect 117236 2100 117292 2102
rect 117684 2548 117740 2604
rect 117908 2548 117964 2604
rect 117460 2324 117516 2380
rect 117796 1540 117852 1596
rect 116788 1204 116844 1260
rect 117012 1204 117068 1260
rect 118132 2548 118188 2604
rect 118356 3444 118412 3500
rect 118692 3780 118748 3836
rect 119028 5908 119084 5964
rect 118468 2996 118524 3052
rect 118356 2324 118412 2380
rect 118356 1876 118412 1932
rect 119476 11284 119532 11340
rect 119588 9268 119644 9324
rect 119364 8036 119420 8092
rect 119812 12740 119868 12796
rect 120148 13860 120204 13916
rect 120708 14532 120764 14588
rect 121044 14420 121100 14476
rect 121492 14420 121548 14476
rect 120036 12740 120092 12796
rect 120708 12740 120764 12796
rect 120484 12516 120540 12572
rect 121268 12404 121324 12460
rect 120820 12292 120876 12348
rect 120372 12180 120428 12236
rect 119812 12068 119868 12124
rect 119812 10164 119868 10220
rect 119812 9156 119868 9212
rect 119924 7812 119980 7868
rect 120148 11956 120204 12012
rect 120372 11956 120428 12012
rect 120372 11786 120428 11788
rect 120372 11734 120374 11786
rect 120374 11734 120426 11786
rect 120426 11734 120428 11786
rect 120372 11732 120428 11734
rect 120708 10836 120764 10892
rect 120260 10612 120316 10668
rect 120260 9492 120316 9548
rect 120540 9770 120596 9772
rect 120540 9718 120542 9770
rect 120542 9718 120594 9770
rect 120594 9718 120596 9770
rect 120540 9716 120596 9718
rect 120372 8596 120428 8652
rect 122948 14420 123004 14476
rect 121940 12180 121996 12236
rect 122164 12180 122220 12236
rect 121380 11732 121436 11788
rect 120932 10948 120988 11004
rect 121044 10836 121100 10892
rect 120932 10612 120988 10668
rect 121044 9770 121100 9772
rect 121044 9718 121046 9770
rect 121046 9718 121098 9770
rect 121098 9718 121100 9770
rect 121044 9716 121100 9718
rect 124404 14420 124460 14476
rect 122724 12292 122780 12348
rect 122948 12964 123004 13020
rect 121268 9716 121324 9772
rect 120708 8596 120764 8652
rect 120932 9268 120988 9324
rect 120260 7700 120316 7756
rect 119700 7588 119756 7644
rect 119364 6244 119420 6300
rect 119252 5908 119308 5964
rect 119364 4004 119420 4060
rect 118916 2548 118972 2604
rect 119028 2772 119084 2828
rect 118916 1652 118972 1708
rect 118468 1540 118524 1596
rect 119140 2212 119196 2268
rect 119364 2212 119420 2268
rect 119700 7364 119756 7420
rect 121156 8484 121212 8540
rect 119924 7364 119980 7420
rect 121044 7252 121100 7308
rect 120372 6916 120428 6972
rect 119700 6244 119756 6300
rect 120708 6020 120764 6076
rect 119756 5962 119812 5964
rect 119756 5910 119758 5962
rect 119758 5910 119810 5962
rect 119810 5910 119812 5962
rect 119756 5908 119812 5910
rect 120372 5796 120428 5852
rect 119812 4340 119868 4396
rect 119476 980 119532 1036
rect 119924 4004 119980 4060
rect 120148 4340 120204 4396
rect 120148 4116 120204 4172
rect 121324 7418 121380 7420
rect 121324 7366 121326 7418
rect 121326 7366 121378 7418
rect 121378 7366 121380 7418
rect 121324 7364 121380 7366
rect 121324 7028 121380 7084
rect 121380 4900 121436 4956
rect 120260 4004 120316 4060
rect 121156 4058 121212 4060
rect 121156 4006 121158 4058
rect 121158 4006 121210 4058
rect 121210 4006 121212 4058
rect 121156 4004 121212 4006
rect 121380 4004 121436 4060
rect 119924 2548 119980 2604
rect 121716 8260 121772 8316
rect 121716 7364 121772 7420
rect 122164 8596 122220 8652
rect 122052 8036 122108 8092
rect 122388 8596 122444 8652
rect 121604 5908 121660 5964
rect 121940 7252 121996 7308
rect 121828 5684 121884 5740
rect 121716 5236 121772 5292
rect 121604 4900 121660 4956
rect 121828 4900 121884 4956
rect 122276 7252 122332 7308
rect 122276 6692 122332 6748
rect 122164 6468 122220 6524
rect 122164 6244 122220 6300
rect 122500 8484 122556 8540
rect 122836 7364 122892 7420
rect 124516 13748 124572 13804
rect 124516 12852 124572 12908
rect 124964 12964 125020 13020
rect 124180 11060 124236 11116
rect 124292 10836 124348 10892
rect 123396 9044 123452 9100
rect 123732 9268 123788 9324
rect 123732 8596 123788 8652
rect 123956 9268 124012 9324
rect 123340 8148 123396 8204
rect 123228 8090 123284 8092
rect 123228 8038 123230 8090
rect 123230 8038 123282 8090
rect 123282 8038 123284 8090
rect 123228 8036 123284 8038
rect 122948 7028 123004 7084
rect 123284 7028 123340 7084
rect 122500 6692 122556 6748
rect 122500 6468 122556 6524
rect 122948 6020 123004 6076
rect 122612 5908 122668 5964
rect 122612 5236 122668 5292
rect 122836 5908 122892 5964
rect 120260 3220 120316 3276
rect 121268 2884 121324 2940
rect 121492 2660 121548 2716
rect 120372 2324 120428 2380
rect 119700 980 119756 1036
rect 120820 2324 120876 2380
rect 121604 2324 121660 2380
rect 120932 2212 120988 2268
rect 121156 2212 121212 2268
rect 120932 1988 120988 2044
rect 121156 1988 121212 2044
rect 121044 1764 121100 1820
rect 120708 1540 120764 1596
rect 120820 1428 120876 1484
rect 120708 1370 120764 1372
rect 120708 1318 120710 1370
rect 120710 1318 120762 1370
rect 120762 1318 120764 1370
rect 120708 1316 120764 1318
rect 117012 644 117068 700
rect 121268 308 121324 364
rect 122612 3444 122668 3500
rect 122164 2772 122220 2828
rect 122164 2548 122220 2604
rect 123564 6522 123620 6524
rect 123564 6470 123566 6522
rect 123566 6470 123618 6522
rect 123618 6470 123620 6522
rect 123564 6468 123620 6470
rect 123284 5796 123340 5852
rect 123172 5460 123228 5516
rect 123284 4900 123340 4956
rect 123060 3668 123116 3724
rect 123284 3220 123340 3276
rect 121716 644 121772 700
rect 123844 6468 123900 6524
rect 123732 5572 123788 5628
rect 124068 8484 124124 8540
rect 126756 13860 126812 13916
rect 126756 13412 126812 13468
rect 126980 13188 127036 13244
rect 126980 12516 127036 12572
rect 127092 11844 127148 11900
rect 127316 12740 127372 12796
rect 125636 9828 125692 9884
rect 126532 10388 126588 10444
rect 125860 10276 125916 10332
rect 125748 9492 125804 9548
rect 127988 11844 128044 11900
rect 127316 10164 127372 10220
rect 124740 8260 124796 8316
rect 124852 8708 124908 8764
rect 127092 8708 127148 8764
rect 126532 8484 126588 8540
rect 125076 8372 125132 8428
rect 125972 8260 126028 8316
rect 126644 8260 126700 8316
rect 126420 8148 126476 8204
rect 125412 7476 125468 7532
rect 125412 7252 125468 7308
rect 127652 8260 127708 8316
rect 127540 8090 127596 8092
rect 127540 8038 127542 8090
rect 127542 8038 127594 8090
rect 127594 8038 127596 8090
rect 127540 8036 127596 8038
rect 124740 6580 124796 6636
rect 124404 6132 124460 6188
rect 126532 4900 126588 4956
rect 125636 4340 125692 4396
rect 123956 4116 124012 4172
rect 124180 4116 124236 4172
rect 126756 4900 126812 4956
rect 126756 4676 126812 4732
rect 127204 4004 127260 4060
rect 125636 3780 125692 3836
rect 128548 11844 128604 11900
rect 129556 11620 129612 11676
rect 129108 11172 129164 11228
rect 129220 10388 129276 10444
rect 129108 10052 129164 10108
rect 130452 10612 130508 10668
rect 129556 10388 129612 10444
rect 130004 10500 130060 10556
rect 128380 9380 128436 9436
rect 127876 7364 127932 7420
rect 127988 8372 128044 8428
rect 128436 7812 128492 7868
rect 128268 7418 128324 7420
rect 128268 7366 128270 7418
rect 128270 7366 128322 7418
rect 128322 7366 128324 7418
rect 128268 7364 128324 7366
rect 128268 6580 128324 6636
rect 129052 7812 129108 7868
rect 130004 9156 130060 9212
rect 129444 7700 129500 7756
rect 128548 6580 128604 6636
rect 129220 6132 129276 6188
rect 129444 6132 129500 6188
rect 128772 5236 128828 5292
rect 129444 5236 129500 5292
rect 130340 9156 130396 9212
rect 131012 12292 131068 12348
rect 130900 10666 130956 10668
rect 130900 10614 130902 10666
rect 130902 10614 130954 10666
rect 130954 10614 130956 10666
rect 130900 10612 130956 10614
rect 134148 14308 134204 14364
rect 130900 10164 130956 10220
rect 131236 11844 131292 11900
rect 131348 10724 131404 10780
rect 131348 10276 131404 10332
rect 131236 9380 131292 9436
rect 131460 10052 131516 10108
rect 131124 9268 131180 9324
rect 130676 8596 130732 8652
rect 130396 7700 130452 7756
rect 130228 7364 130284 7420
rect 130452 7364 130508 7420
rect 130452 6916 130508 6972
rect 130900 6580 130956 6636
rect 130788 6468 130844 6524
rect 131572 10724 131628 10780
rect 131684 10612 131740 10668
rect 131796 9716 131852 9772
rect 132132 10276 132188 10332
rect 132356 13076 132412 13132
rect 132020 10052 132076 10108
rect 132916 11732 132972 11788
rect 132692 11620 132748 11676
rect 132468 11396 132524 11452
rect 132916 10164 132972 10220
rect 132356 8148 132412 8204
rect 132468 7924 132524 7980
rect 132916 9940 132972 9996
rect 132916 8372 132972 8428
rect 132580 6916 132636 6972
rect 132804 7700 132860 7756
rect 131404 6634 131460 6636
rect 131404 6582 131406 6634
rect 131406 6582 131458 6634
rect 131458 6582 131460 6634
rect 131404 6580 131460 6582
rect 131852 6522 131908 6524
rect 131852 6470 131854 6522
rect 131854 6470 131906 6522
rect 131906 6470 131908 6522
rect 131852 6468 131908 6470
rect 130900 6020 130956 6076
rect 130564 5908 130620 5964
rect 130004 4788 130060 4844
rect 128100 4116 128156 4172
rect 129556 3780 129612 3836
rect 125860 2996 125916 3052
rect 125860 2660 125916 2716
rect 126084 2660 126140 2716
rect 125412 2436 125468 2492
rect 123844 1876 123900 1932
rect 124516 1764 124572 1820
rect 123508 644 123564 700
rect 124740 420 124796 476
rect 125860 1876 125916 1932
rect 129332 2884 129388 2940
rect 127652 2660 127708 2716
rect 128772 2772 128828 2828
rect 127764 2436 127820 2492
rect 126084 1316 126140 1372
rect 127652 2154 127708 2156
rect 127652 2102 127654 2154
rect 127654 2102 127706 2154
rect 127706 2102 127708 2154
rect 127652 2100 127708 2102
rect 127876 2100 127932 2156
rect 126308 1316 126364 1372
rect 128212 1764 128268 1820
rect 125748 1204 125804 1260
rect 127540 1204 127596 1260
rect 126980 1092 127036 1148
rect 131068 5908 131124 5964
rect 129556 2324 129612 2380
rect 130900 2772 130956 2828
rect 130564 1092 130620 1148
rect 131684 3108 131740 3164
rect 132020 3780 132076 3836
rect 131908 2884 131964 2940
rect 131796 1652 131852 1708
rect 125300 532 125356 588
rect 132524 5572 132580 5628
rect 132356 5236 132412 5292
rect 132580 4788 132636 4844
rect 132692 3444 132748 3500
rect 132244 3220 132300 3276
rect 132691 2996 132747 3052
rect 134708 14308 134764 14364
rect 134148 12068 134204 12124
rect 133588 11620 133644 11676
rect 133588 11114 133644 11116
rect 133588 11062 133590 11114
rect 133590 11062 133642 11114
rect 133642 11062 133644 11114
rect 133588 11060 133644 11062
rect 133924 10554 133980 10556
rect 133924 10502 133926 10554
rect 133926 10502 133978 10554
rect 133978 10502 133980 10554
rect 133924 10500 133980 10502
rect 133140 10388 133196 10444
rect 133140 9940 133196 9996
rect 133588 10388 133644 10444
rect 133476 9044 133532 9100
rect 134484 12964 134540 13020
rect 134372 12068 134428 12124
rect 134932 11956 134988 12012
rect 134260 11844 134316 11900
rect 134260 11172 134316 11228
rect 134148 10500 134204 10556
rect 134036 10388 134092 10444
rect 134260 10442 134316 10444
rect 134260 10390 134262 10442
rect 134262 10390 134314 10442
rect 134314 10390 134316 10442
rect 134260 10388 134316 10390
rect 134484 10388 134540 10444
rect 134372 10276 134428 10332
rect 133924 9044 133980 9100
rect 133364 8596 133420 8652
rect 133252 8202 133308 8204
rect 133252 8150 133254 8202
rect 133254 8150 133306 8202
rect 133306 8150 133308 8202
rect 133252 8148 133308 8150
rect 133140 8036 133196 8092
rect 133140 5684 133196 5740
rect 133028 5460 133084 5516
rect 133700 8708 133756 8764
rect 134092 9044 134148 9100
rect 134260 8932 134316 8988
rect 133812 7476 133868 7532
rect 135380 12068 135436 12124
rect 135044 11060 135100 11116
rect 135268 11060 135324 11116
rect 135492 10948 135548 11004
rect 135604 13524 135660 13580
rect 135380 10836 135436 10892
rect 135828 12964 135884 13020
rect 135604 10836 135660 10892
rect 135940 11396 135996 11452
rect 135828 10724 135884 10780
rect 134932 9828 134988 9884
rect 135492 9716 135548 9772
rect 134820 8260 134876 8316
rect 134484 7924 134540 7980
rect 134932 9380 134988 9436
rect 134596 7588 134652 7644
rect 134820 6804 134876 6860
rect 134148 6244 134204 6300
rect 134260 5572 134316 5628
rect 134260 5348 134316 5404
rect 134148 5236 134204 5292
rect 133420 4788 133476 4844
rect 132132 2660 132188 2716
rect 132692 2772 132748 2828
rect 132916 2660 132972 2716
rect 132804 1764 132860 1820
rect 132916 1540 132972 1596
rect 133364 2324 133420 2380
rect 133364 1988 133420 2044
rect 133700 4452 133756 4508
rect 133700 3220 133756 3276
rect 134148 4058 134204 4060
rect 134148 4006 134150 4058
rect 134150 4006 134202 4058
rect 134202 4006 134204 4058
rect 134148 4004 134204 4006
rect 134820 4004 134876 4060
rect 134036 3444 134092 3500
rect 134260 3444 134316 3500
rect 134148 3220 134204 3276
rect 134036 2772 134092 2828
rect 134148 2884 134204 2940
rect 133924 1652 133980 1708
rect 133924 868 133980 924
rect 134260 2378 134316 2380
rect 134260 2326 134262 2378
rect 134262 2326 134314 2378
rect 134314 2326 134316 2378
rect 134260 2324 134316 2326
rect 135268 9044 135324 9100
rect 135156 8596 135212 8652
rect 135380 8372 135436 8428
rect 135772 8986 135828 8988
rect 135772 8934 135774 8986
rect 135774 8934 135826 8986
rect 135826 8934 135828 8986
rect 135772 8932 135828 8934
rect 135940 8932 135996 8988
rect 135100 5908 135156 5964
rect 135268 5012 135324 5068
rect 135548 5962 135604 5964
rect 135548 5910 135550 5962
rect 135550 5910 135602 5962
rect 135602 5910 135604 5962
rect 135548 5908 135604 5910
rect 135604 5684 135660 5740
rect 134372 1540 134428 1596
rect 134484 3332 134540 3388
rect 132020 532 132076 588
rect 134820 3220 134876 3276
rect 135380 3220 135436 3276
rect 134596 3108 134652 3164
rect 134596 2884 134652 2940
rect 135604 4900 135660 4956
rect 136276 8708 136332 8764
rect 135996 7642 136052 7644
rect 135996 7590 135998 7642
rect 135998 7590 136050 7642
rect 136050 7590 136052 7642
rect 135996 7588 136052 7590
rect 136108 6916 136164 6972
rect 135940 5908 135996 5964
rect 136276 6580 136332 6636
rect 135716 3332 135772 3388
rect 136164 3780 136220 3836
rect 135492 2884 135548 2940
rect 134820 1652 134876 1708
rect 135044 1370 135100 1372
rect 135044 1318 135046 1370
rect 135046 1318 135098 1370
rect 135098 1318 135100 1370
rect 135044 1316 135100 1318
rect 136052 3220 136108 3276
rect 136276 2212 136332 2268
rect 136500 10164 136556 10220
rect 136500 6916 136556 6972
rect 137396 12852 137452 12908
rect 137844 12740 137900 12796
rect 137620 11956 137676 12012
rect 136724 9940 136780 9996
rect 137032 10218 137088 10220
rect 137032 10166 137034 10218
rect 137034 10166 137086 10218
rect 137086 10166 137088 10218
rect 137032 10164 137088 10166
rect 137136 10218 137192 10220
rect 137136 10166 137138 10218
rect 137138 10166 137190 10218
rect 137190 10166 137192 10218
rect 137136 10164 137192 10166
rect 137240 10218 137296 10220
rect 137240 10166 137242 10218
rect 137242 10166 137294 10218
rect 137294 10166 137296 10218
rect 137240 10164 137296 10166
rect 137956 11844 138012 11900
rect 138292 13860 138348 13916
rect 137732 11620 137788 11676
rect 138740 13860 138796 13916
rect 138852 11732 138908 11788
rect 138292 11674 138348 11676
rect 138292 11622 138294 11674
rect 138294 11622 138346 11674
rect 138346 11622 138348 11674
rect 138292 11620 138348 11622
rect 137620 10164 137676 10220
rect 137060 9940 137116 9996
rect 137396 9994 137452 9996
rect 137396 9942 137398 9994
rect 137398 9942 137450 9994
rect 137450 9942 137452 9994
rect 137396 9940 137452 9942
rect 137396 9156 137452 9212
rect 137788 9882 137844 9884
rect 137788 9830 137790 9882
rect 137790 9830 137842 9882
rect 137842 9830 137844 9882
rect 137788 9828 137844 9830
rect 137956 9380 138012 9436
rect 137032 8650 137088 8652
rect 137032 8598 137034 8650
rect 137034 8598 137086 8650
rect 137086 8598 137088 8650
rect 137032 8596 137088 8598
rect 137136 8650 137192 8652
rect 137136 8598 137138 8650
rect 137138 8598 137190 8650
rect 137190 8598 137192 8650
rect 137136 8596 137192 8598
rect 137240 8650 137296 8652
rect 137240 8598 137242 8650
rect 137242 8598 137294 8650
rect 137294 8598 137296 8650
rect 137240 8596 137296 8598
rect 137620 8260 137676 8316
rect 136948 8036 137004 8092
rect 137032 7082 137088 7084
rect 137032 7030 137034 7082
rect 137034 7030 137086 7082
rect 137086 7030 137088 7082
rect 137032 7028 137088 7030
rect 137136 7082 137192 7084
rect 137136 7030 137138 7082
rect 137138 7030 137190 7082
rect 137190 7030 137192 7082
rect 137136 7028 137192 7030
rect 137240 7082 137296 7084
rect 137240 7030 137242 7082
rect 137242 7030 137294 7082
rect 137294 7030 137296 7082
rect 137240 7028 137296 7030
rect 136612 5908 136668 5964
rect 137508 7028 137564 7084
rect 137732 6020 137788 6076
rect 136612 5124 136668 5180
rect 136500 4676 136556 4732
rect 136724 3668 136780 3724
rect 136500 3220 136556 3276
rect 136724 3220 136780 3276
rect 137508 5572 137564 5628
rect 137032 5514 137088 5516
rect 137032 5462 137034 5514
rect 137034 5462 137086 5514
rect 137086 5462 137088 5514
rect 137032 5460 137088 5462
rect 137136 5514 137192 5516
rect 137136 5462 137138 5514
rect 137138 5462 137190 5514
rect 137190 5462 137192 5514
rect 137136 5460 137192 5462
rect 137240 5514 137296 5516
rect 137240 5462 137242 5514
rect 137242 5462 137294 5514
rect 137294 5462 137296 5514
rect 137240 5460 137296 5462
rect 137620 5460 137676 5516
rect 137116 4676 137172 4732
rect 137284 4676 137340 4732
rect 136724 2212 136780 2268
rect 136388 1876 136444 1932
rect 136164 1652 136220 1708
rect 137172 1316 137228 1372
rect 137172 980 137228 1036
rect 137844 5796 137900 5852
rect 138292 8932 138348 8988
rect 138852 8484 138908 8540
rect 138068 5684 138124 5740
rect 138292 6356 138348 6412
rect 137956 4788 138012 4844
rect 138628 6356 138684 6412
rect 138740 5796 138796 5852
rect 138628 5236 138684 5292
rect 138964 4676 139020 4732
rect 139300 12068 139356 12124
rect 139524 13860 139580 13916
rect 140084 13748 140140 13804
rect 139748 11844 139804 11900
rect 139524 11620 139580 11676
rect 139412 10612 139468 10668
rect 139748 8932 139804 8988
rect 139524 8820 139580 8876
rect 139636 8596 139692 8652
rect 139412 6804 139468 6860
rect 138516 3332 138572 3388
rect 138180 2548 138236 2604
rect 138180 1764 138236 1820
rect 139412 6020 139468 6076
rect 139300 5908 139356 5964
rect 139412 4788 139468 4844
rect 139412 4564 139468 4620
rect 139076 2884 139132 2940
rect 139860 7140 139916 7196
rect 139860 6804 139916 6860
rect 139860 4452 139916 4508
rect 139524 3668 139580 3724
rect 139636 4116 139692 4172
rect 139636 3444 139692 3500
rect 139748 3668 139804 3724
rect 139412 2884 139468 2940
rect 139636 3108 139692 3164
rect 139636 2660 139692 2716
rect 140756 14084 140812 14140
rect 140196 13076 140252 13132
rect 140308 8932 140364 8988
rect 140196 8708 140252 8764
rect 140420 7364 140476 7420
rect 141092 11620 141148 11676
rect 141204 10276 141260 10332
rect 142660 13636 142716 13692
rect 140756 10052 140812 10108
rect 140980 9380 141036 9436
rect 140756 9156 140812 9212
rect 142660 12852 142716 12908
rect 142996 13188 143052 13244
rect 142324 10836 142380 10892
rect 141540 10164 141596 10220
rect 141708 9940 141764 9996
rect 140756 8932 140812 8988
rect 142772 11732 142828 11788
rect 142436 10164 142492 10220
rect 140980 8708 141036 8764
rect 141092 8484 141148 8540
rect 141092 8148 141148 8204
rect 141876 7924 141932 7980
rect 142884 9770 142940 9772
rect 142884 9718 142886 9770
rect 142886 9718 142938 9770
rect 142938 9718 142940 9770
rect 142884 9716 142940 9718
rect 143108 12628 143164 12684
rect 143220 12180 143276 12236
rect 143332 11844 143388 11900
rect 143332 11396 143388 11452
rect 143668 11060 143724 11116
rect 142996 8484 143052 8540
rect 143108 9716 143164 9772
rect 141876 7306 141932 7308
rect 141876 7254 141878 7306
rect 141878 7254 141930 7306
rect 141930 7254 141932 7306
rect 141876 7252 141932 7254
rect 142660 6916 142716 6972
rect 141764 6858 141820 6860
rect 141764 6806 141766 6858
rect 141766 6806 141818 6858
rect 141818 6806 141820 6858
rect 141764 6804 141820 6806
rect 140644 6692 140700 6748
rect 142996 6916 143052 6972
rect 140868 5908 140924 5964
rect 140644 5012 140700 5068
rect 140532 4900 140588 4956
rect 140308 3444 140364 3500
rect 139860 3108 139916 3164
rect 139860 2212 139916 2268
rect 141148 4676 141204 4732
rect 140980 4452 141036 4508
rect 140980 4228 141036 4284
rect 140756 3444 140812 3500
rect 140868 4116 140924 4172
rect 140644 3332 140700 3388
rect 140532 3108 140588 3164
rect 140756 3108 140812 3164
rect 140756 2660 140812 2716
rect 141204 4228 141260 4284
rect 142156 5460 142212 5516
rect 142156 5124 142212 5180
rect 141596 4954 141652 4956
rect 141596 4902 141598 4954
rect 141598 4902 141650 4954
rect 141650 4902 141652 4954
rect 141596 4900 141652 4902
rect 141764 4900 141820 4956
rect 141540 3946 141596 3948
rect 141540 3894 141542 3946
rect 141542 3894 141594 3946
rect 141594 3894 141596 3946
rect 141540 3892 141596 3894
rect 141428 3668 141484 3724
rect 141316 3444 141372 3500
rect 141764 3444 141820 3500
rect 140980 2324 141036 2380
rect 141540 3332 141596 3388
rect 141764 3220 141820 3276
rect 141540 2324 141596 2380
rect 141540 2100 141596 2156
rect 134484 532 134540 588
rect 142828 4788 142884 4844
rect 142660 4676 142716 4732
rect 142996 4452 143052 4508
rect 142772 4340 142828 4396
rect 142548 3556 142604 3612
rect 142212 1428 142268 1484
rect 142772 3444 142828 3500
rect 144116 13860 144172 13916
rect 144228 12852 144284 12908
rect 144452 11844 144508 11900
rect 144564 11732 144620 11788
rect 143780 9156 143836 9212
rect 143892 8932 143948 8988
rect 143668 8372 143724 8428
rect 143724 7642 143780 7644
rect 143724 7590 143726 7642
rect 143726 7590 143778 7642
rect 143778 7590 143780 7642
rect 143724 7588 143780 7590
rect 143556 6804 143612 6860
rect 141988 420 142044 476
rect 142548 756 142604 812
rect 142772 2772 142828 2828
rect 143780 5348 143836 5404
rect 143612 4564 143668 4620
rect 143780 4564 143836 4620
rect 144956 9770 145012 9772
rect 144956 9718 144958 9770
rect 144958 9718 145010 9770
rect 145010 9718 145012 9770
rect 144956 9716 145012 9718
rect 144676 9156 144732 9212
rect 144452 8820 144508 8876
rect 144452 8260 144508 8316
rect 144676 8820 144732 8876
rect 144228 7588 144284 7644
rect 144564 8036 144620 8092
rect 145012 9156 145068 9212
rect 144788 8148 144844 8204
rect 144788 7588 144844 7644
rect 144676 7028 144732 7084
rect 144564 6804 144620 6860
rect 144228 5796 144284 5852
rect 144452 5796 144508 5852
rect 144452 5236 144508 5292
rect 145236 11956 145292 12012
rect 145348 12852 145404 12908
rect 145236 8260 145292 8316
rect 145124 8148 145180 8204
rect 146692 12964 146748 13020
rect 147140 13188 147196 13244
rect 147028 12852 147084 12908
rect 146132 11284 146188 11340
rect 146020 8820 146076 8876
rect 145684 8426 145740 8428
rect 145684 8374 145686 8426
rect 145686 8374 145738 8426
rect 145738 8374 145740 8426
rect 145684 8372 145740 8374
rect 145572 7364 145628 7420
rect 145796 6858 145852 6860
rect 145796 6806 145798 6858
rect 145798 6806 145850 6858
rect 145850 6806 145852 6858
rect 145796 6804 145852 6806
rect 145012 6468 145068 6524
rect 145236 6580 145292 6636
rect 144788 6020 144844 6076
rect 145124 6020 145180 6076
rect 144676 5908 144732 5964
rect 145236 5908 145292 5964
rect 145012 5572 145068 5628
rect 144452 4788 144508 4844
rect 144900 4788 144956 4844
rect 144004 3722 144060 3724
rect 144004 3670 144006 3722
rect 144006 3670 144058 3722
rect 144058 3670 144060 3722
rect 144004 3668 144060 3670
rect 145572 4564 145628 4620
rect 145348 4228 145404 4284
rect 145908 5236 145964 5292
rect 146020 4788 146076 4844
rect 145572 4228 145628 4284
rect 146916 10836 146972 10892
rect 146804 10724 146860 10780
rect 146580 10388 146636 10444
rect 146580 10164 146636 10220
rect 146804 10164 146860 10220
rect 147924 13636 147980 13692
rect 148372 13748 148428 13804
rect 148372 13466 148428 13468
rect 148372 13414 148374 13466
rect 148374 13414 148426 13466
rect 148426 13414 148428 13466
rect 148372 13412 148428 13414
rect 149156 14420 149212 14476
rect 148708 13972 148764 14028
rect 149268 14250 149324 14252
rect 149268 14198 149270 14250
rect 149270 14198 149322 14250
rect 149322 14198 149324 14250
rect 149268 14196 149324 14198
rect 149268 13524 149324 13580
rect 148932 13076 148988 13132
rect 149492 13524 149548 13580
rect 149380 13354 149436 13356
rect 149380 13302 149382 13354
rect 149382 13302 149434 13354
rect 149434 13302 149436 13354
rect 149380 13300 149436 13302
rect 149156 12964 149212 13020
rect 148708 12570 148764 12572
rect 148708 12518 148710 12570
rect 148710 12518 148762 12570
rect 148762 12518 148764 12570
rect 148708 12516 148764 12518
rect 149044 12516 149100 12572
rect 148708 12292 148764 12348
rect 147812 11844 147868 11900
rect 147700 11732 147756 11788
rect 147700 10948 147756 11004
rect 147812 10500 147868 10556
rect 147924 11060 147980 11116
rect 147252 10388 147308 10444
rect 146580 8820 146636 8876
rect 146356 8148 146412 8204
rect 146244 7476 146300 7532
rect 146244 6244 146300 6300
rect 146468 4116 146524 4172
rect 144900 2100 144956 2156
rect 143444 1876 143500 1932
rect 145796 1764 145852 1820
rect 143444 1540 143500 1596
rect 144004 1540 144060 1596
rect 145236 1540 145292 1596
rect 147532 10052 147588 10108
rect 148148 9828 148204 9884
rect 147420 8820 147476 8876
rect 147532 8314 147588 8316
rect 147532 8262 147534 8314
rect 147534 8262 147586 8314
rect 147586 8262 147588 8314
rect 147532 8260 147588 8262
rect 147588 7476 147644 7532
rect 147812 6916 147868 6972
rect 147924 7476 147980 7532
rect 147644 6804 147700 6860
rect 146916 6132 146972 6188
rect 146580 3892 146636 3948
rect 147084 4954 147140 4956
rect 147084 4902 147086 4954
rect 147086 4902 147138 4954
rect 147138 4902 147140 4954
rect 147084 4900 147140 4902
rect 146916 4676 146972 4732
rect 147644 6522 147700 6524
rect 147644 6470 147646 6522
rect 147646 6470 147698 6522
rect 147698 6470 147700 6522
rect 147644 6468 147700 6470
rect 147252 4340 147308 4396
rect 147644 4954 147700 4956
rect 147644 4902 147646 4954
rect 147646 4902 147698 4954
rect 147698 4902 147700 4954
rect 147644 4900 147700 4902
rect 147700 4452 147756 4508
rect 147476 4340 147532 4396
rect 146916 3780 146972 3836
rect 147476 4004 147532 4060
rect 147364 1652 147420 1708
rect 148428 10164 148484 10220
rect 149492 12292 149548 12348
rect 148932 11898 148988 11900
rect 148932 11846 148934 11898
rect 148934 11846 148986 11898
rect 148986 11846 148988 11898
rect 148932 11844 148988 11846
rect 148708 11060 148764 11116
rect 149380 9940 149436 9996
rect 148876 9658 148932 9660
rect 148876 9606 148878 9658
rect 148878 9606 148930 9658
rect 148930 9606 148932 9658
rect 148876 9604 148932 9606
rect 149828 14196 149884 14252
rect 150724 14308 150780 14364
rect 150164 13412 150220 13468
rect 149716 13076 149772 13132
rect 150052 11284 150108 11340
rect 149716 10388 149772 10444
rect 149772 9882 149828 9884
rect 149772 9830 149774 9882
rect 149774 9830 149826 9882
rect 149826 9830 149828 9882
rect 149772 9828 149828 9830
rect 149604 9044 149660 9100
rect 148820 8820 148876 8876
rect 148708 8484 148764 8540
rect 149268 8708 149324 8764
rect 149604 8372 149660 8428
rect 150052 8372 150108 8428
rect 151396 14868 151452 14924
rect 151284 14532 151340 14588
rect 150500 13972 150556 14028
rect 150388 11284 150444 11340
rect 150276 11002 150332 11004
rect 150276 10950 150278 11002
rect 150278 10950 150330 11002
rect 150330 10950 150332 11002
rect 150276 10948 150332 10950
rect 150164 8148 150220 8204
rect 148708 7812 148764 7868
rect 149996 7530 150052 7532
rect 149996 7478 149998 7530
rect 149998 7478 150050 7530
rect 150050 7478 150052 7530
rect 149996 7476 150052 7478
rect 150164 7476 150220 7532
rect 150276 9828 150332 9884
rect 148820 6916 148876 6972
rect 148596 6244 148652 6300
rect 150388 9716 150444 9772
rect 150388 9044 150444 9100
rect 150724 10052 150780 10108
rect 151060 12628 151116 12684
rect 151172 12740 151228 12796
rect 151060 11620 151116 11676
rect 151172 11060 151228 11116
rect 151060 9994 151116 9996
rect 151060 9942 151062 9994
rect 151062 9942 151114 9994
rect 151114 9942 151116 9994
rect 151060 9940 151116 9942
rect 150948 9828 151004 9884
rect 151172 9828 151228 9884
rect 150500 8372 150556 8428
rect 150668 8202 150724 8204
rect 150668 8150 150670 8202
rect 150670 8150 150722 8202
rect 150722 8150 150724 8202
rect 150668 8148 150724 8150
rect 150948 8372 151004 8428
rect 151116 8484 151172 8540
rect 151508 14420 151564 14476
rect 151844 13636 151900 13692
rect 152068 13636 152124 13692
rect 152068 13412 152124 13468
rect 152516 12852 152572 12908
rect 152852 14196 152908 14252
rect 155204 14420 155260 14476
rect 152964 13748 153020 13804
rect 151508 11898 151564 11900
rect 151508 11846 151510 11898
rect 151510 11846 151562 11898
rect 151562 11846 151564 11898
rect 151508 11844 151564 11846
rect 151732 11508 151788 11564
rect 151732 10724 151788 10780
rect 152068 10836 152124 10892
rect 151452 10052 151508 10108
rect 151396 8484 151452 8540
rect 151844 8484 151900 8540
rect 151396 8148 151452 8204
rect 149604 6580 149660 6636
rect 150724 7476 150780 7532
rect 149268 6468 149324 6524
rect 150500 6692 150556 6748
rect 151900 8148 151956 8204
rect 148540 5066 148596 5068
rect 148540 5014 148542 5066
rect 148542 5014 148594 5066
rect 148594 5014 148596 5066
rect 148540 5012 148596 5014
rect 148876 4788 148932 4844
rect 148708 3668 148764 3724
rect 147812 3220 147868 3276
rect 149716 5348 149772 5404
rect 149436 5012 149492 5068
rect 149940 4788 149996 4844
rect 149772 4676 149828 4732
rect 150052 4676 150108 4732
rect 150164 3332 150220 3388
rect 149268 2772 149324 2828
rect 149492 3220 149548 3276
rect 148932 2100 148988 2156
rect 148260 1876 148316 1932
rect 147700 980 147756 1036
rect 150052 2884 150108 2940
rect 151116 6522 151172 6524
rect 151116 6470 151118 6522
rect 151118 6470 151170 6522
rect 151170 6470 151172 6522
rect 151116 6468 151172 6470
rect 150948 5796 151004 5852
rect 152404 10388 152460 10444
rect 152292 8484 152348 8540
rect 151508 6580 151564 6636
rect 151732 6580 151788 6636
rect 151788 5850 151844 5852
rect 151788 5798 151790 5850
rect 151790 5798 151842 5850
rect 151842 5798 151844 5850
rect 151788 5796 151844 5798
rect 151788 5236 151844 5292
rect 151284 4564 151340 4620
rect 151508 4564 151564 4620
rect 151060 3610 151116 3612
rect 151060 3558 151062 3610
rect 151062 3558 151114 3610
rect 151114 3558 151116 3610
rect 151060 3556 151116 3558
rect 152180 6916 152236 6972
rect 153188 13802 153244 13804
rect 153188 13750 153190 13802
rect 153190 13750 153242 13802
rect 153242 13750 153244 13802
rect 153188 13748 153244 13750
rect 153860 14084 153916 14140
rect 154756 13412 154812 13468
rect 154980 13412 155036 13468
rect 154644 13076 154700 13132
rect 153300 12068 153356 12124
rect 153524 12068 153580 12124
rect 154532 11956 154588 12012
rect 154532 11172 154588 11228
rect 154756 12516 154812 12572
rect 154868 11732 154924 11788
rect 154756 11620 154812 11676
rect 154644 10836 154700 10892
rect 153412 10388 153468 10444
rect 152516 9604 152572 9660
rect 153076 8484 153132 8540
rect 152964 8372 153020 8428
rect 152628 8148 152684 8204
rect 152852 6020 152908 6076
rect 152628 5348 152684 5404
rect 151956 4340 152012 4396
rect 152852 4900 152908 4956
rect 152852 4452 152908 4508
rect 152180 3892 152236 3948
rect 152292 4340 152348 4396
rect 150164 2660 150220 2716
rect 150276 2772 150332 2828
rect 150052 2212 150108 2268
rect 150276 1706 150332 1708
rect 150276 1654 150278 1706
rect 150278 1654 150330 1706
rect 150330 1654 150332 1706
rect 150276 1652 150332 1654
rect 150164 1316 150220 1372
rect 153300 7588 153356 7644
rect 154644 9940 154700 9996
rect 155092 13300 155148 13356
rect 155092 11956 155148 12012
rect 157108 14644 157164 14700
rect 157108 14308 157164 14364
rect 155316 13300 155372 13356
rect 156212 13972 156268 14028
rect 155428 12180 155484 12236
rect 155540 13748 155596 13804
rect 155372 9940 155428 9996
rect 153972 8426 154028 8428
rect 153972 8374 153974 8426
rect 153974 8374 154026 8426
rect 154026 8374 154028 8426
rect 153972 8372 154028 8374
rect 153076 6692 153132 6748
rect 153132 4788 153188 4844
rect 153300 4452 153356 4508
rect 153076 4116 153132 4172
rect 152516 3892 152572 3948
rect 151060 1930 151116 1932
rect 151060 1878 151062 1930
rect 151062 1878 151114 1930
rect 151114 1878 151116 1930
rect 151060 1876 151116 1878
rect 153076 3892 153132 3948
rect 152628 2996 152684 3052
rect 152628 2490 152684 2492
rect 152628 2438 152630 2490
rect 152630 2438 152682 2490
rect 152682 2438 152684 2490
rect 152628 2436 152684 2438
rect 152404 1764 152460 1820
rect 152516 2324 152572 2380
rect 151956 868 152012 924
rect 153188 3668 153244 3724
rect 153748 7140 153804 7196
rect 154420 7364 154476 7420
rect 153692 6634 153748 6636
rect 153692 6582 153694 6634
rect 153694 6582 153746 6634
rect 153746 6582 153748 6634
rect 153692 6580 153748 6582
rect 153580 4676 153636 4732
rect 153188 3444 153244 3500
rect 152852 2212 152908 2268
rect 153188 2548 153244 2604
rect 154980 6580 155036 6636
rect 154308 6468 154364 6524
rect 154532 6356 154588 6412
rect 154700 6356 154756 6412
rect 154980 6356 155036 6412
rect 155428 7252 155484 7308
rect 157668 13860 157724 13916
rect 158340 13860 158396 13916
rect 158900 14196 158956 14252
rect 161532 14868 161588 14924
rect 156884 12404 156940 12460
rect 157220 13524 157276 13580
rect 156436 11620 156492 11676
rect 157108 11620 157164 11676
rect 156212 10388 156268 10444
rect 156436 10388 156492 10444
rect 155988 8148 156044 8204
rect 156324 9380 156380 9436
rect 155316 6692 155372 6748
rect 155540 6580 155596 6636
rect 155988 7588 156044 7644
rect 156100 6356 156156 6412
rect 154476 4954 154532 4956
rect 154476 4902 154478 4954
rect 154478 4902 154530 4954
rect 154530 4902 154532 4954
rect 154476 4900 154532 4902
rect 155652 5572 155708 5628
rect 154644 4676 154700 4732
rect 154420 4116 154476 4172
rect 155652 4452 155708 4508
rect 155988 4676 156044 4732
rect 155316 4004 155372 4060
rect 154644 3332 154700 3388
rect 154532 3108 154588 3164
rect 154532 2490 154588 2492
rect 154532 2438 154534 2490
rect 154534 2438 154586 2490
rect 154586 2438 154588 2490
rect 154532 2436 154588 2438
rect 154756 2436 154812 2492
rect 153860 2266 153916 2268
rect 153860 2214 153862 2266
rect 153862 2214 153914 2266
rect 153914 2214 153916 2266
rect 153860 2212 153916 2214
rect 153748 980 153804 1036
rect 154868 1428 154924 1484
rect 156100 4452 156156 4508
rect 156100 4282 156156 4284
rect 156100 4230 156102 4282
rect 156102 4230 156154 4282
rect 156154 4230 156156 4282
rect 156100 4228 156156 4230
rect 155988 2660 156044 2716
rect 155988 1652 156044 1708
rect 158788 10836 158844 10892
rect 159572 13972 159628 14028
rect 159124 13300 159180 13356
rect 159012 11844 159068 11900
rect 159236 11508 159292 11564
rect 159348 12964 159404 13020
rect 159012 10836 159068 10892
rect 159236 11060 159292 11116
rect 157780 10164 157836 10220
rect 158676 9716 158732 9772
rect 157220 9380 157276 9436
rect 158564 9044 158620 9100
rect 157780 8484 157836 8540
rect 158564 8372 158620 8428
rect 156548 6468 156604 6524
rect 156436 4900 156492 4956
rect 157332 6858 157388 6860
rect 157332 6806 157334 6858
rect 157334 6806 157386 6858
rect 157386 6806 157388 6858
rect 157332 6804 157388 6806
rect 157556 6580 157612 6636
rect 158564 8036 158620 8092
rect 158564 7588 158620 7644
rect 158228 6468 158284 6524
rect 156772 6356 156828 6412
rect 157556 6356 157612 6412
rect 158116 6132 158172 6188
rect 156996 5738 157052 5740
rect 156996 5686 156998 5738
rect 156998 5686 157050 5738
rect 157050 5686 157052 5738
rect 156996 5684 157052 5686
rect 157444 5012 157500 5068
rect 156660 4004 156716 4060
rect 156772 4116 156828 4172
rect 156436 1652 156492 1708
rect 158676 6132 158732 6188
rect 158676 5124 158732 5180
rect 158676 4116 158732 4172
rect 159236 10612 159292 10668
rect 159124 10388 159180 10444
rect 159796 13188 159852 13244
rect 162484 14644 162540 14700
rect 162260 14532 162316 14588
rect 160580 12292 160636 12348
rect 161028 12964 161084 13020
rect 159460 11732 159516 11788
rect 159460 11284 159516 11340
rect 160916 11508 160972 11564
rect 159348 9828 159404 9884
rect 159628 9716 159684 9772
rect 160804 9716 160860 9772
rect 160580 8260 160636 8316
rect 159012 5012 159068 5068
rect 160692 8148 160748 8204
rect 159460 7588 159516 7644
rect 159460 7140 159516 7196
rect 159460 6020 159516 6076
rect 159348 5236 159404 5292
rect 159348 5012 159404 5068
rect 159460 5124 159516 5180
rect 159236 4116 159292 4172
rect 159124 2100 159180 2156
rect 159908 4228 159964 4284
rect 161252 11060 161308 11116
rect 161476 13300 161532 13356
rect 161924 12852 161980 12908
rect 161476 10164 161532 10220
rect 161588 9716 161644 9772
rect 161308 9380 161364 9436
rect 161364 7588 161420 7644
rect 160916 6580 160972 6636
rect 160636 6468 160692 6524
rect 160580 5684 160636 5740
rect 160748 5684 160804 5740
rect 161476 7476 161532 7532
rect 161364 6468 161420 6524
rect 161756 9098 161812 9100
rect 161756 9046 161758 9098
rect 161758 9046 161810 9098
rect 161810 9046 161812 9098
rect 161756 9044 161812 9046
rect 162372 10500 162428 10556
rect 163268 14644 163324 14700
rect 162708 13972 162764 14028
rect 162708 12068 162764 12124
rect 162820 11844 162876 11900
rect 162932 12180 162988 12236
rect 162932 11060 162988 11116
rect 161140 5572 161196 5628
rect 160748 5348 160804 5404
rect 161700 4564 161756 4620
rect 160468 3220 160524 3276
rect 161140 3220 161196 3276
rect 161028 2324 161084 2380
rect 160468 1540 160524 1596
rect 162260 1988 162316 2044
rect 162596 7700 162652 7756
rect 162484 5348 162540 5404
rect 163492 13636 163548 13692
rect 163940 13524 163996 13580
rect 163828 11284 163884 11340
rect 163716 9716 163772 9772
rect 163268 7812 163324 7868
rect 164164 13412 164220 13468
rect 164948 13188 165004 13244
rect 164052 12404 164108 12460
rect 165732 12964 165788 13020
rect 165060 12180 165116 12236
rect 165620 11844 165676 11900
rect 164612 11396 164668 11452
rect 165284 11508 165340 11564
rect 164052 9940 164108 9996
rect 165284 10500 165340 10556
rect 164332 9882 164388 9884
rect 164332 9830 164334 9882
rect 164334 9830 164386 9882
rect 164386 9830 164388 9882
rect 164332 9828 164388 9830
rect 165732 11732 165788 11788
rect 164196 9434 164252 9436
rect 164196 9382 164198 9434
rect 164198 9382 164250 9434
rect 164250 9382 164252 9434
rect 164196 9380 164252 9382
rect 164300 9434 164356 9436
rect 164300 9382 164302 9434
rect 164302 9382 164354 9434
rect 164354 9382 164356 9434
rect 164300 9380 164356 9382
rect 164404 9434 164460 9436
rect 164404 9382 164406 9434
rect 164406 9382 164458 9434
rect 164458 9382 164460 9434
rect 164404 9380 164460 9382
rect 163604 7476 163660 7532
rect 163828 6580 163884 6636
rect 164196 7866 164252 7868
rect 164196 7814 164198 7866
rect 164198 7814 164250 7866
rect 164250 7814 164252 7866
rect 164196 7812 164252 7814
rect 164300 7866 164356 7868
rect 164300 7814 164302 7866
rect 164302 7814 164354 7866
rect 164354 7814 164356 7866
rect 164300 7812 164356 7814
rect 164404 7866 164460 7868
rect 164404 7814 164406 7866
rect 164406 7814 164458 7866
rect 164458 7814 164460 7866
rect 164404 7812 164460 7814
rect 164276 7588 164332 7644
rect 164836 7364 164892 7420
rect 164612 7140 164668 7196
rect 164836 7140 164892 7196
rect 164196 6298 164252 6300
rect 164196 6246 164198 6298
rect 164198 6246 164250 6298
rect 164250 6246 164252 6298
rect 164196 6244 164252 6246
rect 164300 6298 164356 6300
rect 164300 6246 164302 6298
rect 164302 6246 164354 6298
rect 164354 6246 164356 6298
rect 164300 6244 164356 6246
rect 164404 6298 164460 6300
rect 164404 6246 164406 6298
rect 164406 6246 164458 6298
rect 164458 6246 164460 6298
rect 164404 6244 164460 6246
rect 163828 5460 163884 5516
rect 165004 6522 165060 6524
rect 165004 6470 165006 6522
rect 165006 6470 165058 6522
rect 165058 6470 165060 6522
rect 165004 6468 165060 6470
rect 165396 5908 165452 5964
rect 164500 5236 164556 5292
rect 165396 5236 165452 5292
rect 164052 5012 164108 5068
rect 163604 4676 163660 4732
rect 164196 4730 164252 4732
rect 164196 4678 164198 4730
rect 164198 4678 164250 4730
rect 164250 4678 164252 4730
rect 164196 4676 164252 4678
rect 164300 4730 164356 4732
rect 164300 4678 164302 4730
rect 164302 4678 164354 4730
rect 164354 4678 164356 4730
rect 164300 4676 164356 4678
rect 164404 4730 164460 4732
rect 164404 4678 164406 4730
rect 164406 4678 164458 4730
rect 164458 4678 164460 4730
rect 164404 4676 164460 4678
rect 165452 4954 165508 4956
rect 165452 4902 165454 4954
rect 165454 4902 165506 4954
rect 165506 4902 165508 4954
rect 165452 4900 165508 4902
rect 165116 4676 165172 4732
rect 164556 4452 164612 4508
rect 162596 4340 162652 4396
rect 165172 3892 165228 3948
rect 162708 2826 162764 2828
rect 162708 2774 162710 2826
rect 162710 2774 162762 2826
rect 162762 2774 162764 2826
rect 162708 2772 162764 2774
rect 167188 12068 167244 12124
rect 166404 11732 166460 11788
rect 166628 10276 166684 10332
rect 166460 9716 166516 9772
rect 166460 9268 166516 9324
rect 166628 9604 166684 9660
rect 166068 9044 166124 9100
rect 166628 8148 166684 8204
rect 165844 6356 165900 6412
rect 166404 6132 166460 6188
rect 166180 5460 166236 5516
rect 166292 5124 166348 5180
rect 166628 6132 166684 6188
rect 166628 5572 166684 5628
rect 166292 4900 166348 4956
rect 166516 4116 166572 4172
rect 166852 9268 166908 9324
rect 166964 8260 167020 8316
rect 166964 7924 167020 7980
rect 166852 6580 166908 6636
rect 167300 5908 167356 5964
rect 166964 5572 167020 5628
rect 167076 5460 167132 5516
rect 166964 4340 167020 4396
rect 166964 4004 167020 4060
rect 166740 3668 166796 3724
rect 167076 3668 167132 3724
rect 167188 5348 167244 5404
rect 167076 2996 167132 3052
rect 165732 2324 165788 2380
rect 165172 1988 165228 2044
rect 165396 1988 165452 2044
rect 162372 1876 162428 1932
rect 162932 1540 162988 1596
rect 164724 1540 164780 1596
rect 163492 1316 163548 1372
rect 164164 1204 164220 1260
rect 167076 2324 167132 2380
rect 166516 1540 166572 1596
rect 167860 13076 167916 13132
rect 169092 14196 169148 14252
rect 169764 14420 169820 14476
rect 171332 14308 171388 14364
rect 168644 11844 168700 11900
rect 169428 12404 169484 12460
rect 167636 10500 167692 10556
rect 168868 10276 168924 10332
rect 168700 10164 168756 10220
rect 167860 10052 167916 10108
rect 169316 9604 169372 9660
rect 167748 7588 167804 7644
rect 168756 8484 168812 8540
rect 167860 7476 167916 7532
rect 167636 6580 167692 6636
rect 169204 8932 169260 8988
rect 169092 8260 169148 8316
rect 168868 7252 168924 7308
rect 168868 6244 168924 6300
rect 170212 11508 170268 11564
rect 170100 9716 170156 9772
rect 169540 8260 169596 8316
rect 169540 7028 169596 7084
rect 169316 6020 169372 6076
rect 169204 5908 169260 5964
rect 167860 5460 167916 5516
rect 167636 5124 167692 5180
rect 167972 4676 168028 4732
rect 168644 4004 168700 4060
rect 168868 4900 168924 4956
rect 167748 1876 167804 1932
rect 168420 3668 168476 3724
rect 167412 1540 167468 1596
rect 167748 1428 167804 1484
rect 168980 4340 169036 4396
rect 169484 5572 169540 5628
rect 169484 5348 169540 5404
rect 169204 4004 169260 4060
rect 170324 8372 170380 8428
rect 171108 13076 171164 13132
rect 170884 11956 170940 12012
rect 170772 11732 170828 11788
rect 171108 11620 171164 11676
rect 171220 12292 171276 12348
rect 170828 9098 170884 9100
rect 170828 9046 170830 9098
rect 170830 9046 170882 9098
rect 170882 9046 170884 9098
rect 170828 9044 170884 9046
rect 170996 9044 171052 9100
rect 170772 8260 170828 8316
rect 172676 14868 172732 14924
rect 171556 13300 171612 13356
rect 172228 12292 172284 12348
rect 172564 11844 172620 11900
rect 172452 11732 172508 11788
rect 171668 10500 171724 10556
rect 171668 8484 171724 8540
rect 171220 6468 171276 6524
rect 171108 5908 171164 5964
rect 170100 5348 170156 5404
rect 172228 7924 172284 7980
rect 171668 5348 171724 5404
rect 171892 6244 171948 6300
rect 170436 4228 170492 4284
rect 174132 14196 174188 14252
rect 174692 14756 174748 14812
rect 174020 13524 174076 13580
rect 173460 12740 173516 12796
rect 173460 12292 173516 12348
rect 173012 11956 173068 12012
rect 172788 11060 172844 11116
rect 173292 9940 173348 9996
rect 173348 9044 173404 9100
rect 172564 4676 172620 4732
rect 172004 4452 172060 4508
rect 170212 1540 170268 1596
rect 170884 1092 170940 1148
rect 171444 868 171500 924
rect 172676 3556 172732 3612
rect 173404 8090 173460 8092
rect 173404 8038 173406 8090
rect 173406 8038 173458 8090
rect 173458 8038 173460 8090
rect 173404 8036 173460 8038
rect 173012 5908 173068 5964
rect 173012 4954 173068 4956
rect 173012 4902 173014 4954
rect 173014 4902 173066 4954
rect 173066 4902 173068 4954
rect 173012 4900 173068 4902
rect 175588 14532 175644 14588
rect 174692 14084 174748 14140
rect 174468 13860 174524 13916
rect 174132 13188 174188 13244
rect 174916 13748 174972 13804
rect 174188 9770 174244 9772
rect 174188 9718 174190 9770
rect 174190 9718 174242 9770
rect 174242 9718 174244 9770
rect 174188 9716 174244 9718
rect 174244 9156 174300 9212
rect 173124 3892 173180 3948
rect 174804 7812 174860 7868
rect 174356 7588 174412 7644
rect 175140 12068 175196 12124
rect 175476 14084 175532 14140
rect 176820 14532 176876 14588
rect 175028 8260 175084 8316
rect 175028 8090 175084 8092
rect 175028 8038 175030 8090
rect 175030 8038 175082 8090
rect 175082 8038 175084 8090
rect 175028 8036 175084 8038
rect 174804 6916 174860 6972
rect 175924 11172 175980 11228
rect 181972 14868 182028 14924
rect 177156 13300 177212 13356
rect 176932 11956 176988 12012
rect 175140 6580 175196 6636
rect 174468 6356 174524 6412
rect 175140 6074 175196 6076
rect 175140 6022 175142 6074
rect 175142 6022 175194 6074
rect 175194 6022 175196 6074
rect 175140 6020 175196 6022
rect 174580 5917 174636 5964
rect 174580 5908 174582 5917
rect 174582 5908 174634 5917
rect 174634 5908 174636 5917
rect 174356 4564 174412 4620
rect 175028 4116 175084 4172
rect 172900 1988 172956 2044
rect 173236 3668 173292 3724
rect 172676 1316 172732 1372
rect 174356 2660 174412 2716
rect 175756 7530 175812 7532
rect 175756 7478 175758 7530
rect 175758 7478 175810 7530
rect 175810 7478 175812 7530
rect 175756 7476 175812 7478
rect 175476 6074 175532 6076
rect 175476 6022 175478 6074
rect 175478 6022 175530 6074
rect 175530 6022 175532 6074
rect 175476 6020 175532 6022
rect 175924 5124 175980 5180
rect 175252 3892 175308 3948
rect 175924 4004 175980 4060
rect 176484 5460 176540 5516
rect 176708 4116 176764 4172
rect 176932 4340 176988 4396
rect 177268 12740 177324 12796
rect 178052 13972 178108 14028
rect 177380 11732 177436 11788
rect 177492 12740 177548 12796
rect 177268 10164 177324 10220
rect 178052 12180 178108 12236
rect 178052 11956 178108 12012
rect 178052 10612 178108 10668
rect 178836 12180 178892 12236
rect 179172 13972 179228 14028
rect 178276 10612 178332 10668
rect 178612 11956 178668 12012
rect 178164 9492 178220 9548
rect 178276 9156 178332 9212
rect 178052 8708 178108 8764
rect 178500 8708 178556 8764
rect 177604 8148 177660 8204
rect 177716 7700 177772 7756
rect 177940 6244 177996 6300
rect 177604 6132 177660 6188
rect 179060 9940 179116 9996
rect 179284 13300 179340 13356
rect 179508 13188 179564 13244
rect 182980 14084 183036 14140
rect 181748 13860 181804 13916
rect 180964 12964 181020 13020
rect 182308 13636 182364 13692
rect 180292 12628 180348 12684
rect 179620 12180 179676 12236
rect 179396 10612 179452 10668
rect 181300 12180 181356 12236
rect 180068 12068 180124 12124
rect 180404 11508 180460 11564
rect 181132 10276 181188 10332
rect 181020 9658 181076 9660
rect 181020 9606 181022 9658
rect 181022 9606 181074 9658
rect 181074 9606 181076 9658
rect 181020 9604 181076 9606
rect 182084 9716 182140 9772
rect 180852 9156 180908 9212
rect 180404 8372 180460 8428
rect 178836 6634 178892 6636
rect 178836 6582 178838 6634
rect 178838 6582 178890 6634
rect 178890 6582 178892 6634
rect 178836 6580 178892 6582
rect 179172 6356 179228 6412
rect 177492 5348 177548 5404
rect 178164 5348 178220 5404
rect 177156 4340 177212 4396
rect 176148 3556 176204 3612
rect 175924 3108 175980 3164
rect 175140 1540 175196 1596
rect 174468 980 174524 1036
rect 173908 868 173964 924
rect 178276 4228 178332 4284
rect 178724 4564 178780 4620
rect 178724 3892 178780 3948
rect 178052 3220 178108 3276
rect 178388 2772 178444 2828
rect 178388 2436 178444 2492
rect 177716 2100 177772 2156
rect 178164 2212 178220 2268
rect 178164 1988 178220 2044
rect 178836 3444 178892 3500
rect 178948 3332 179004 3388
rect 180180 7252 180236 7308
rect 181860 9380 181916 9436
rect 181300 8372 181356 8428
rect 181524 8820 181580 8876
rect 180684 7140 180740 7196
rect 179676 6634 179732 6636
rect 179676 6582 179678 6634
rect 179678 6582 179730 6634
rect 179730 6582 179732 6634
rect 179676 6580 179732 6582
rect 179620 6020 179676 6076
rect 180180 6020 180236 6076
rect 180068 4900 180124 4956
rect 179396 3220 179452 3276
rect 179956 3220 180012 3276
rect 178836 1988 178892 2044
rect 179060 2436 179116 2492
rect 179396 1540 179452 1596
rect 180628 4340 180684 4396
rect 180068 3108 180124 3164
rect 180292 3108 180348 3164
rect 181188 6804 181244 6860
rect 181300 6692 181356 6748
rect 181300 5796 181356 5852
rect 181132 4788 181188 4844
rect 181300 3556 181356 3612
rect 180964 3108 181020 3164
rect 180292 2436 180348 2492
rect 181188 1540 181244 1596
rect 180628 1428 180684 1484
rect 182868 13636 182924 13692
rect 182532 12852 182588 12908
rect 182756 9828 182812 9884
rect 182532 9044 182588 9100
rect 182756 9380 182812 9436
rect 182756 8484 182812 8540
rect 183204 13748 183260 13804
rect 184660 13524 184716 13580
rect 183876 12068 183932 12124
rect 183988 11732 184044 11788
rect 183876 11284 183932 11340
rect 183876 10724 183932 10780
rect 183652 10052 183708 10108
rect 183428 8932 183484 8988
rect 183708 8986 183764 8988
rect 183708 8934 183710 8986
rect 183710 8934 183762 8986
rect 183762 8934 183764 8986
rect 183708 8932 183764 8934
rect 182532 7588 182588 7644
rect 182308 6132 182364 6188
rect 182420 6356 182476 6412
rect 181636 5124 181692 5180
rect 182196 4788 182252 4844
rect 181412 1204 181468 1260
rect 181860 4116 181916 4172
rect 182980 7700 183036 7756
rect 182980 7364 183036 7420
rect 182980 7140 183036 7196
rect 182644 6858 182700 6860
rect 182644 6806 182646 6858
rect 182646 6806 182698 6858
rect 182698 6806 182700 6858
rect 182644 6804 182700 6806
rect 182868 6132 182924 6188
rect 183540 8596 183596 8652
rect 183652 8260 183708 8316
rect 185332 12964 185388 13020
rect 185668 13524 185724 13580
rect 184548 10836 184604 10892
rect 184324 9156 184380 9212
rect 184772 9940 184828 9996
rect 185052 9828 185108 9884
rect 185108 9604 185164 9660
rect 185556 9268 185612 9324
rect 184996 7812 185052 7868
rect 185108 8260 185164 8316
rect 183428 6132 183484 6188
rect 183204 5796 183260 5852
rect 183540 5796 183596 5852
rect 182644 3444 182700 3500
rect 182980 4340 183036 4396
rect 185220 6804 185276 6860
rect 184324 5348 184380 5404
rect 184772 6132 184828 6188
rect 183708 5236 183764 5292
rect 183092 2436 183148 2492
rect 184212 3108 184268 3164
rect 184772 5572 184828 5628
rect 185780 13076 185836 13132
rect 186116 11732 186172 11788
rect 186228 13636 186284 13692
rect 185892 10724 185948 10780
rect 186004 9604 186060 9660
rect 186116 8820 186172 8876
rect 186452 11844 186508 11900
rect 186340 11172 186396 11228
rect 186788 12740 186844 12796
rect 187572 13972 187628 14028
rect 187124 12628 187180 12684
rect 186676 9604 186732 9660
rect 186676 9156 186732 9212
rect 185220 5012 185276 5068
rect 184436 2996 184492 3052
rect 185332 4788 185388 4844
rect 185780 4676 185836 4732
rect 186564 7028 186620 7084
rect 187012 6916 187068 6972
rect 186900 6692 186956 6748
rect 186788 5684 186844 5740
rect 186004 4228 186060 4284
rect 185892 2884 185948 2940
rect 184548 2436 184604 2492
rect 185444 2436 185500 2492
rect 184884 2100 184940 2156
rect 186116 2938 186172 2940
rect 186116 2886 186118 2938
rect 186118 2886 186170 2938
rect 186170 2886 186172 2938
rect 186116 2884 186172 2886
rect 186340 4228 186396 4284
rect 186004 2826 186060 2828
rect 186004 2774 186006 2826
rect 186006 2774 186058 2826
rect 186058 2774 186060 2826
rect 186004 2772 186060 2774
rect 186228 2772 186284 2828
rect 186340 2548 186396 2604
rect 187572 12292 187628 12348
rect 187908 12068 187964 12124
rect 187684 11620 187740 11676
rect 187684 11060 187740 11116
rect 188020 11620 188076 11676
rect 187796 9604 187852 9660
rect 187628 8260 187684 8316
rect 187516 8202 187572 8204
rect 187516 8150 187518 8202
rect 187518 8150 187570 8202
rect 187570 8150 187572 8202
rect 187516 8148 187572 8150
rect 187348 7812 187404 7868
rect 186228 2436 186284 2492
rect 186564 3780 186620 3836
rect 186900 3220 186956 3276
rect 187348 3220 187404 3276
rect 188692 14196 188748 14252
rect 188244 9658 188300 9660
rect 188244 9606 188246 9658
rect 188246 9606 188298 9658
rect 188298 9606 188300 9658
rect 188244 9604 188300 9606
rect 188020 5572 188076 5628
rect 187908 5236 187964 5292
rect 187460 4004 187516 4060
rect 187012 2548 187068 2604
rect 187348 2660 187404 2716
rect 186452 2436 186508 2492
rect 186676 2324 186732 2380
rect 186116 1540 186172 1596
rect 188580 10836 188636 10892
rect 189028 13300 189084 13356
rect 189700 11844 189756 11900
rect 190372 11732 190428 11788
rect 189812 10948 189868 11004
rect 189700 10276 189756 10332
rect 188692 9156 188748 9212
rect 188468 8148 188524 8204
rect 188468 6804 188524 6860
rect 188692 5572 188748 5628
rect 188972 5066 189028 5068
rect 188972 5014 188974 5066
rect 188974 5014 189026 5066
rect 189026 5014 189028 5066
rect 188972 5012 189028 5014
rect 189140 5012 189196 5068
rect 188020 3892 188076 3948
rect 188804 3332 188860 3388
rect 189924 9492 189980 9548
rect 189924 9156 189980 9212
rect 189364 5124 189420 5180
rect 189252 4564 189308 4620
rect 189588 6580 189644 6636
rect 189588 6356 189644 6412
rect 189812 6244 189868 6300
rect 189756 4954 189812 4956
rect 189756 4902 189758 4954
rect 189758 4902 189810 4954
rect 189810 4902 189812 4954
rect 189756 4900 189812 4902
rect 189588 4564 189644 4620
rect 189476 3780 189532 3836
rect 187572 2324 187628 2380
rect 191156 13972 191212 14028
rect 191828 13860 191884 13916
rect 190596 13188 190652 13244
rect 191156 10500 191212 10556
rect 190932 9210 190988 9212
rect 190932 9158 190934 9210
rect 190934 9158 190986 9210
rect 190986 9158 190988 9210
rect 190932 9156 190988 9158
rect 191360 10218 191416 10220
rect 191360 10166 191362 10218
rect 191362 10166 191414 10218
rect 191414 10166 191416 10218
rect 191360 10164 191416 10166
rect 191464 10218 191520 10220
rect 191464 10166 191466 10218
rect 191466 10166 191518 10218
rect 191518 10166 191520 10218
rect 191464 10164 191520 10166
rect 191568 10218 191624 10220
rect 191568 10166 191570 10218
rect 191570 10166 191622 10218
rect 191622 10166 191624 10218
rect 191568 10164 191624 10166
rect 191380 9940 191436 9996
rect 191940 12180 191996 12236
rect 191828 9604 191884 9660
rect 191360 8650 191416 8652
rect 191360 8598 191362 8650
rect 191362 8598 191414 8650
rect 191414 8598 191416 8650
rect 191360 8596 191416 8598
rect 191464 8650 191520 8652
rect 191464 8598 191466 8650
rect 191466 8598 191518 8650
rect 191518 8598 191520 8650
rect 191464 8596 191520 8598
rect 191568 8650 191624 8652
rect 191568 8598 191570 8650
rect 191570 8598 191622 8650
rect 191622 8598 191624 8650
rect 191568 8596 191624 8598
rect 190708 8372 190764 8428
rect 190596 7364 190652 7420
rect 191324 8090 191380 8092
rect 191324 8038 191326 8090
rect 191326 8038 191378 8090
rect 191378 8038 191380 8090
rect 191324 8036 191380 8038
rect 190820 7700 190876 7756
rect 190932 7642 190988 7644
rect 190932 7590 190934 7642
rect 190934 7590 190986 7642
rect 190986 7590 190988 7642
rect 190932 7588 190988 7590
rect 190596 6692 190652 6748
rect 191660 7306 191716 7308
rect 191660 7254 191662 7306
rect 191662 7254 191714 7306
rect 191714 7254 191716 7306
rect 191660 7252 191716 7254
rect 191360 7082 191416 7084
rect 191360 7030 191362 7082
rect 191362 7030 191414 7082
rect 191414 7030 191416 7082
rect 191360 7028 191416 7030
rect 191464 7082 191520 7084
rect 191464 7030 191466 7082
rect 191466 7030 191518 7082
rect 191518 7030 191520 7082
rect 191464 7028 191520 7030
rect 191568 7082 191624 7084
rect 191568 7030 191570 7082
rect 191570 7030 191622 7082
rect 191622 7030 191624 7082
rect 191568 7028 191624 7030
rect 191772 6692 191828 6748
rect 190484 5908 190540 5964
rect 191212 6020 191268 6076
rect 192164 9770 192220 9772
rect 192164 9718 192166 9770
rect 192166 9718 192218 9770
rect 192218 9718 192220 9770
rect 192164 9716 192220 9718
rect 192276 7588 192332 7644
rect 193956 14084 194012 14140
rect 193396 13860 193452 13916
rect 193620 12964 193676 13020
rect 192612 11732 192668 11788
rect 192948 9828 193004 9884
rect 192780 9492 192836 9548
rect 193060 9044 193116 9100
rect 194068 12404 194124 12460
rect 194628 11956 194684 12012
rect 195524 12964 195580 13020
rect 196308 13748 196364 13804
rect 196308 12740 196364 12796
rect 195860 12292 195916 12348
rect 193732 11732 193788 11788
rect 194068 11284 194124 11340
rect 193060 7924 193116 7980
rect 193844 9156 193900 9212
rect 193844 8708 193900 8764
rect 193788 7642 193844 7644
rect 193788 7590 193790 7642
rect 193790 7590 193842 7642
rect 193842 7590 193844 7642
rect 193788 7588 193844 7590
rect 193620 7252 193676 7308
rect 193732 6916 193788 6972
rect 192668 6522 192724 6524
rect 192668 6470 192670 6522
rect 192670 6470 192722 6522
rect 192722 6470 192724 6522
rect 192668 6468 192724 6470
rect 192220 6244 192276 6300
rect 192892 6356 192948 6412
rect 191436 5684 191492 5740
rect 191360 5514 191416 5516
rect 191360 5462 191362 5514
rect 191362 5462 191414 5514
rect 191414 5462 191416 5514
rect 191360 5460 191416 5462
rect 191464 5514 191520 5516
rect 191464 5462 191466 5514
rect 191466 5462 191518 5514
rect 191518 5462 191520 5514
rect 191464 5460 191520 5462
rect 191568 5514 191624 5516
rect 191568 5462 191570 5514
rect 191570 5462 191622 5514
rect 191622 5462 191624 5514
rect 191568 5460 191624 5462
rect 193564 6522 193620 6524
rect 193564 6470 193566 6522
rect 193566 6470 193618 6522
rect 193618 6470 193620 6522
rect 193564 6468 193620 6470
rect 193340 6074 193396 6076
rect 193340 6022 193342 6074
rect 193342 6022 193394 6074
rect 193394 6022 193396 6074
rect 193340 6020 193396 6022
rect 193060 5460 193116 5516
rect 194348 6244 194404 6300
rect 190652 4954 190708 4956
rect 190652 4902 190654 4954
rect 190654 4902 190706 4954
rect 190706 4902 190708 4954
rect 190652 4900 190708 4902
rect 191100 4452 191156 4508
rect 191380 4452 191436 4508
rect 191268 4058 191324 4060
rect 191268 4006 191270 4058
rect 191270 4006 191322 4058
rect 191322 4006 191324 4058
rect 191268 4004 191324 4006
rect 192444 4954 192500 4956
rect 192444 4902 192446 4954
rect 192446 4902 192498 4954
rect 192498 4902 192500 4954
rect 192444 4900 192500 4902
rect 193676 4954 193732 4956
rect 193676 4902 193678 4954
rect 193678 4902 193730 4954
rect 193730 4902 193732 4954
rect 193676 4900 193732 4902
rect 192892 4788 192948 4844
rect 193060 4788 193116 4844
rect 191996 4564 192052 4620
rect 191380 3892 191436 3948
rect 191716 4228 191772 4284
rect 190036 2884 190092 2940
rect 190932 3220 190988 3276
rect 189476 2436 189532 2492
rect 190372 2324 190428 2380
rect 187460 2100 187516 2156
rect 188692 2154 188748 2156
rect 188692 2102 188694 2154
rect 188694 2102 188746 2154
rect 188746 2102 188748 2154
rect 188692 2100 188748 2102
rect 189700 1876 189756 1932
rect 188468 1764 188524 1820
rect 187908 1540 187964 1596
rect 189140 1540 189196 1596
rect 190596 2378 190652 2380
rect 190596 2326 190598 2378
rect 190598 2326 190650 2378
rect 190650 2326 190652 2378
rect 190596 2324 190652 2326
rect 191716 2996 191772 3052
rect 192276 3050 192332 3052
rect 192276 2998 192278 3050
rect 192278 2998 192330 3050
rect 192330 2998 192332 3050
rect 192276 2996 192332 2998
rect 194740 9770 194796 9772
rect 194740 9718 194742 9770
rect 194742 9718 194794 9770
rect 194794 9718 194796 9770
rect 194740 9716 194796 9718
rect 195636 9658 195692 9660
rect 195636 9606 195638 9658
rect 195638 9606 195690 9658
rect 195690 9606 195692 9658
rect 195636 9604 195692 9606
rect 194964 9268 195020 9324
rect 195188 9156 195244 9212
rect 195412 9210 195468 9212
rect 195412 9158 195414 9210
rect 195414 9158 195466 9210
rect 195466 9158 195468 9210
rect 195412 9156 195468 9158
rect 195132 7642 195188 7644
rect 195132 7590 195134 7642
rect 195134 7590 195186 7642
rect 195186 7590 195188 7642
rect 195132 7588 195188 7590
rect 194852 6692 194908 6748
rect 195244 6522 195300 6524
rect 195244 6470 195246 6522
rect 195246 6470 195298 6522
rect 195298 6470 195300 6522
rect 195244 6468 195300 6470
rect 194796 6356 194852 6412
rect 195524 8932 195580 8988
rect 195748 6916 195804 6972
rect 196196 11844 196252 11900
rect 195972 11732 196028 11788
rect 195972 9604 196028 9660
rect 195972 8932 196028 8988
rect 196028 7700 196084 7756
rect 196868 12180 196924 12236
rect 196420 7588 196476 7644
rect 196756 8596 196812 8652
rect 196980 11732 197036 11788
rect 197764 12068 197820 12124
rect 198436 13524 198492 13580
rect 198436 11844 198492 11900
rect 198660 12740 198716 12796
rect 198100 11732 198156 11788
rect 198324 11060 198380 11116
rect 198212 10724 198268 10780
rect 197764 9658 197820 9660
rect 197764 9606 197766 9658
rect 197766 9606 197818 9658
rect 197818 9606 197820 9658
rect 197764 9604 197820 9606
rect 198044 9210 198100 9212
rect 198044 9158 198046 9210
rect 198046 9158 198098 9210
rect 198098 9158 198100 9210
rect 198044 9156 198100 9158
rect 197540 8484 197596 8540
rect 197988 8820 198044 8876
rect 196644 6692 196700 6748
rect 197316 8260 197372 8316
rect 197540 8260 197596 8316
rect 196924 7642 196980 7644
rect 196924 7590 196926 7642
rect 196926 7590 196978 7642
rect 196978 7590 196980 7642
rect 196924 7588 196980 7590
rect 197820 7140 197876 7196
rect 197540 7028 197596 7084
rect 196364 6634 196420 6636
rect 196364 6582 196366 6634
rect 196366 6582 196418 6634
rect 196418 6582 196420 6634
rect 196364 6580 196420 6582
rect 197260 6634 197316 6636
rect 197260 6582 197262 6634
rect 197262 6582 197314 6634
rect 197314 6582 197316 6634
rect 197260 6580 197316 6582
rect 195132 6074 195188 6076
rect 195132 6022 195134 6074
rect 195134 6022 195186 6074
rect 195186 6022 195188 6074
rect 195132 6020 195188 6022
rect 194516 5908 194572 5964
rect 194404 5348 194460 5404
rect 194516 4116 194572 4172
rect 194292 4004 194348 4060
rect 194068 3780 194124 3836
rect 194068 3332 194124 3388
rect 193844 2212 193900 2268
rect 193956 3220 194012 3276
rect 192836 1092 192892 1148
rect 197708 6020 197764 6076
rect 195468 4954 195524 4956
rect 195468 4902 195470 4954
rect 195470 4902 195522 4954
rect 195522 4902 195524 4954
rect 195468 4900 195524 4902
rect 195636 4228 195692 4284
rect 195300 4116 195356 4172
rect 194964 3780 195020 3836
rect 196364 4340 196420 4396
rect 195860 3556 195916 3612
rect 194740 3108 194796 3164
rect 194628 1652 194684 1708
rect 196420 1652 196476 1708
rect 198492 9882 198548 9884
rect 198492 9830 198494 9882
rect 198494 9830 198546 9882
rect 198546 9830 198548 9882
rect 198492 9828 198548 9830
rect 199220 11732 199276 11788
rect 199332 12404 199388 12460
rect 199108 9156 199164 9212
rect 200676 13076 200732 13132
rect 199892 11956 199948 12012
rect 199668 11844 199724 11900
rect 199444 11732 199500 11788
rect 199108 8708 199164 8764
rect 198940 8372 198996 8428
rect 199948 9492 200004 9548
rect 199612 7530 199668 7532
rect 199612 7478 199614 7530
rect 199614 7478 199666 7530
rect 199666 7478 199668 7530
rect 199612 7476 199668 7478
rect 199164 7418 199220 7420
rect 199164 7366 199166 7418
rect 199166 7366 199218 7418
rect 199218 7366 199220 7418
rect 199164 7364 199220 7366
rect 198324 6916 198380 6972
rect 197876 4676 197932 4732
rect 197764 4340 197820 4396
rect 196756 3444 196812 3500
rect 198100 2324 198156 2380
rect 196532 1428 196588 1484
rect 197652 1540 197708 1596
rect 195188 980 195244 1036
rect 197092 980 197148 1036
rect 191828 644 191884 700
rect 198772 6692 198828 6748
rect 198492 5850 198548 5852
rect 198492 5798 198494 5850
rect 198494 5798 198546 5850
rect 198546 5798 198548 5850
rect 198492 5796 198548 5798
rect 199780 7476 199836 7532
rect 199780 6692 199836 6748
rect 199668 6468 199724 6524
rect 199388 6132 199444 6188
rect 200564 12068 200620 12124
rect 200396 9882 200452 9884
rect 200396 9830 200398 9882
rect 200398 9830 200450 9882
rect 200450 9830 200452 9882
rect 200396 9828 200452 9830
rect 200396 9492 200452 9548
rect 201348 11732 201404 11788
rect 201460 13636 201516 13692
rect 200676 10612 200732 10668
rect 200396 8932 200452 8988
rect 200564 7812 200620 7868
rect 201292 9716 201348 9772
rect 201292 8820 201348 8876
rect 201572 12180 201628 12236
rect 202804 13636 202860 13692
rect 203028 12180 203084 12236
rect 202132 11844 202188 11900
rect 202580 11956 202636 12012
rect 201572 11620 201628 11676
rect 202020 11732 202076 11788
rect 202356 10948 202412 11004
rect 202132 10836 202188 10892
rect 201684 9268 201740 9324
rect 201740 8986 201796 8988
rect 201740 8934 201742 8986
rect 201742 8934 201794 8986
rect 201794 8934 201796 8986
rect 201740 8932 201796 8934
rect 202860 9658 202916 9660
rect 202860 9606 202862 9658
rect 202862 9606 202914 9658
rect 202914 9606 202916 9658
rect 202860 9604 202916 9606
rect 202692 9380 202748 9436
rect 203476 11844 203532 11900
rect 203308 9882 203364 9884
rect 203308 9830 203310 9882
rect 203310 9830 203362 9882
rect 203362 9830 203364 9882
rect 203308 9828 203364 9830
rect 202692 9156 202748 9212
rect 202188 8202 202244 8204
rect 202188 8150 202190 8202
rect 202190 8150 202242 8202
rect 202242 8150 202244 8202
rect 202188 8148 202244 8150
rect 200788 6804 200844 6860
rect 200900 6580 200956 6636
rect 200284 4676 200340 4732
rect 200900 4900 200956 4956
rect 200676 3892 200732 3948
rect 201684 5236 201740 5292
rect 201796 4788 201852 4844
rect 201684 4228 201740 4284
rect 202020 8036 202076 8092
rect 202020 5572 202076 5628
rect 202020 4564 202076 4620
rect 199780 2660 199836 2716
rect 200676 2772 200732 2828
rect 198884 2100 198940 2156
rect 199444 1540 199500 1596
rect 200116 1540 200172 1596
rect 201348 980 201404 1036
rect 204820 12852 204876 12908
rect 204260 12068 204316 12124
rect 204372 12292 204428 12348
rect 203588 11732 203644 11788
rect 204596 11732 204652 11788
rect 204260 10052 204316 10108
rect 204036 9940 204092 9996
rect 203084 8090 203140 8092
rect 203084 8038 203086 8090
rect 203086 8038 203138 8090
rect 203138 8038 203140 8090
rect 203084 8036 203140 8038
rect 202636 7418 202692 7420
rect 202636 7366 202638 7418
rect 202638 7366 202690 7418
rect 202690 7366 202692 7418
rect 202636 7364 202692 7366
rect 203924 8148 203980 8204
rect 203644 7924 203700 7980
rect 203532 7418 203588 7420
rect 203532 7366 203534 7418
rect 203534 7366 203586 7418
rect 203586 7366 203588 7418
rect 203532 7364 203588 7366
rect 203924 7364 203980 7420
rect 202580 6580 202636 6636
rect 203084 6634 203140 6636
rect 203084 6582 203086 6634
rect 203086 6582 203138 6634
rect 203138 6582 203140 6634
rect 203084 6580 203140 6582
rect 203140 5572 203196 5628
rect 202468 2996 202524 3052
rect 203924 6244 203980 6300
rect 203756 4676 203812 4732
rect 203812 4116 203868 4172
rect 203588 2212 203644 2268
rect 201908 1876 201964 1932
rect 201684 1316 201740 1372
rect 201908 1428 201964 1484
rect 201572 980 201628 1036
rect 203028 868 203084 924
rect 203812 868 203868 924
rect 204484 9770 204540 9772
rect 204484 9718 204486 9770
rect 204486 9718 204538 9770
rect 204538 9718 204540 9770
rect 204484 9716 204540 9718
rect 205044 12180 205100 12236
rect 205268 12964 205324 13020
rect 204708 9604 204764 9660
rect 205716 11844 205772 11900
rect 205940 12068 205996 12124
rect 205828 9658 205884 9660
rect 205828 9606 205830 9658
rect 205830 9606 205882 9658
rect 205882 9606 205884 9658
rect 205828 9604 205884 9606
rect 207172 12292 207228 12348
rect 206500 11956 206556 12012
rect 207732 11844 207788 11900
rect 206164 11732 206220 11788
rect 206500 9156 206556 9212
rect 206052 8036 206108 8092
rect 206052 7476 206108 7532
rect 206724 8260 206780 8316
rect 206948 8148 207004 8204
rect 207508 7700 207564 7756
rect 208628 12964 208684 13020
rect 207956 11732 208012 11788
rect 208852 11732 208908 11788
rect 208180 10052 208236 10108
rect 208516 9716 208572 9772
rect 206500 6580 206556 6636
rect 207732 7140 207788 7196
rect 205492 5908 205548 5964
rect 205492 5124 205548 5180
rect 205604 5012 205660 5068
rect 204596 4564 204652 4620
rect 205604 4452 205660 4508
rect 205716 3668 205772 3724
rect 204148 756 204204 812
rect 204372 1540 204428 1596
rect 209412 11844 209468 11900
rect 209860 13636 209916 13692
rect 210084 12852 210140 12908
rect 209188 8260 209244 8316
rect 209860 8260 209916 8316
rect 207788 5066 207844 5068
rect 207788 5014 207790 5066
rect 207790 5014 207842 5066
rect 207842 5014 207844 5066
rect 207788 5012 207844 5014
rect 207900 4954 207956 4956
rect 207900 4902 207902 4954
rect 207902 4902 207954 4954
rect 207954 4902 207956 4954
rect 207900 4900 207956 4902
rect 208740 4900 208796 4956
rect 208572 4676 208628 4732
rect 205828 1316 205884 1372
rect 205604 868 205660 924
rect 204708 308 204764 364
rect 206836 868 206892 924
rect 205828 196 205884 252
rect 207620 84 207676 140
rect 209860 7588 209916 7644
rect 209636 6020 209692 6076
rect 209636 3780 209692 3836
rect 209860 6132 209916 6188
rect 209860 5348 209916 5404
rect 209860 4788 209916 4844
rect 209748 1428 209804 1484
rect 209860 1204 209916 1260
rect 210868 11732 210924 11788
rect 210980 12292 211036 12348
rect 211652 13354 211708 13356
rect 211652 13302 211654 13354
rect 211654 13302 211706 13354
rect 211706 13302 211708 13354
rect 211652 13300 211708 13302
rect 211540 11732 211596 11788
rect 211764 12404 211820 12460
rect 210756 9716 210812 9772
rect 210980 9828 211036 9884
rect 211204 9044 211260 9100
rect 211764 10164 211820 10220
rect 211428 9044 211484 9100
rect 210980 7812 211036 7868
rect 210980 7364 211036 7420
rect 211260 7418 211316 7420
rect 211260 7366 211262 7418
rect 211262 7366 211314 7418
rect 211314 7366 211316 7418
rect 211260 7364 211316 7366
rect 210700 7140 210756 7196
rect 212268 9658 212324 9660
rect 212268 9606 212270 9658
rect 212270 9606 212322 9658
rect 212322 9606 212324 9658
rect 212268 9604 212324 9606
rect 212660 9380 212716 9436
rect 211876 8036 211932 8092
rect 211876 6692 211932 6748
rect 210532 5012 210588 5068
rect 210980 5796 211036 5852
rect 210756 5460 210812 5516
rect 212212 8596 212268 8652
rect 213780 12404 213836 12460
rect 214452 12292 214508 12348
rect 212996 12068 213052 12124
rect 215236 12068 215292 12124
rect 215684 12292 215740 12348
rect 213108 11844 213164 11900
rect 212772 9210 212828 9212
rect 212772 9158 212774 9210
rect 212774 9158 212826 9210
rect 212826 9158 212828 9210
rect 212772 9156 212828 9158
rect 212884 11732 212940 11788
rect 212268 8090 212324 8092
rect 212268 8038 212270 8090
rect 212270 8038 212322 8090
rect 212322 8038 212324 8090
rect 212268 8036 212324 8038
rect 212716 8090 212772 8092
rect 212716 8038 212718 8090
rect 212718 8038 212770 8090
rect 212770 8038 212772 8090
rect 212716 8036 212772 8038
rect 212716 7812 212772 7868
rect 212324 7364 212380 7420
rect 212268 6522 212324 6524
rect 212268 6470 212270 6522
rect 212270 6470 212322 6522
rect 212322 6470 212324 6522
rect 212268 6468 212324 6470
rect 211988 6132 212044 6188
rect 212996 9268 213052 9324
rect 213108 6804 213164 6860
rect 213500 8596 213556 8652
rect 213780 11956 213836 12012
rect 215012 11732 215068 11788
rect 213948 8986 214004 8988
rect 213948 8934 213950 8986
rect 213950 8934 214002 8986
rect 214002 8934 214004 8986
rect 213948 8932 214004 8934
rect 214620 9492 214676 9548
rect 214788 9268 214844 9324
rect 214116 8820 214172 8876
rect 215516 9380 215572 9436
rect 215236 9268 215292 9324
rect 214396 8484 214452 8540
rect 215124 8484 215180 8540
rect 213612 7924 213668 7980
rect 213332 6468 213388 6524
rect 211316 5348 211372 5404
rect 211596 4954 211652 4956
rect 211596 4902 211598 4954
rect 211598 4902 211650 4954
rect 211650 4902 211652 4954
rect 211596 4900 211652 4902
rect 212044 4954 212100 4956
rect 212044 4902 212046 4954
rect 212046 4902 212098 4954
rect 212098 4902 212100 4954
rect 212044 4900 212100 4902
rect 211092 4788 211148 4844
rect 212492 4340 212548 4396
rect 212828 5684 212884 5740
rect 213276 6244 213332 6300
rect 213612 6244 213668 6300
rect 214508 8202 214564 8204
rect 214508 8150 214510 8202
rect 214510 8150 214562 8202
rect 214562 8150 214564 8202
rect 214508 8148 214564 8150
rect 213948 7530 214004 7532
rect 213948 7478 213950 7530
rect 213950 7478 214002 7530
rect 214002 7478 214004 7530
rect 213948 7476 214004 7478
rect 214396 7700 214452 7756
rect 215572 8932 215628 8988
rect 215908 12180 215964 12236
rect 216580 12068 216636 12124
rect 216692 11956 216748 12012
rect 218148 12292 218204 12348
rect 217364 11844 217420 11900
rect 219604 12068 219660 12124
rect 218820 11732 218876 11788
rect 216580 9828 216636 9884
rect 215684 8484 215740 8540
rect 216020 9268 216076 9324
rect 215292 7642 215348 7644
rect 215292 7590 215294 7642
rect 215294 7590 215346 7642
rect 215346 7590 215348 7642
rect 215292 7588 215348 7590
rect 214396 7418 214452 7420
rect 214396 7366 214398 7418
rect 214398 7366 214450 7418
rect 214450 7366 214452 7418
rect 214396 7364 214452 7366
rect 214116 7028 214172 7084
rect 214508 6634 214564 6636
rect 214508 6582 214510 6634
rect 214510 6582 214562 6634
rect 214562 6582 214564 6634
rect 214508 6580 214564 6582
rect 213444 5572 213500 5628
rect 213892 6468 213948 6524
rect 213220 4228 213276 4284
rect 213108 4116 213164 4172
rect 212660 3332 212716 3388
rect 210756 1988 210812 2044
rect 211652 1540 211708 1596
rect 211092 1316 211148 1372
rect 212324 980 212380 1036
rect 212884 868 212940 924
rect 213724 5572 213780 5628
rect 214060 6356 214116 6412
rect 214172 5962 214228 5964
rect 214172 5910 214174 5962
rect 214174 5910 214226 5962
rect 214226 5910 214228 5962
rect 214172 5908 214228 5910
rect 214620 5850 214676 5852
rect 214620 5798 214622 5850
rect 214622 5798 214674 5850
rect 214674 5798 214676 5850
rect 214620 5796 214676 5798
rect 213892 5460 213948 5516
rect 213724 4564 213780 4620
rect 214620 4954 214676 4956
rect 214620 4902 214622 4954
rect 214622 4902 214674 4954
rect 214674 4902 214676 4954
rect 214620 4900 214676 4902
rect 214900 6020 214956 6076
rect 214172 4452 214228 4508
rect 215068 5348 215124 5404
rect 215068 4954 215124 4956
rect 215068 4902 215070 4954
rect 215070 4902 215122 4954
rect 215122 4902 215124 4954
rect 215068 4900 215124 4902
rect 215068 4676 215124 4732
rect 215404 6522 215460 6524
rect 215404 6470 215406 6522
rect 215406 6470 215458 6522
rect 215458 6470 215460 6522
rect 215404 6468 215460 6470
rect 215796 6468 215852 6524
rect 216020 6244 216076 6300
rect 216300 9098 216356 9100
rect 216300 9046 216302 9098
rect 216302 9046 216354 9098
rect 216354 9046 216356 9098
rect 216300 9044 216356 9046
rect 216300 8090 216356 8092
rect 216300 8038 216302 8090
rect 216302 8038 216354 8090
rect 216354 8038 216356 8090
rect 216300 8036 216356 8038
rect 217308 9770 217364 9772
rect 217308 9718 217310 9770
rect 217310 9718 217362 9770
rect 217362 9718 217364 9770
rect 217308 9716 217364 9718
rect 216748 9210 216804 9212
rect 216748 9158 216750 9210
rect 216750 9158 216802 9210
rect 216802 9158 216804 9210
rect 216748 9156 216804 9158
rect 216580 8932 216636 8988
rect 217364 6244 217420 6300
rect 216468 5348 216524 5404
rect 216132 4900 216188 4956
rect 215516 4788 215572 4844
rect 215236 4564 215292 4620
rect 214900 3780 214956 3836
rect 219044 1428 219100 1484
rect 214116 1092 214172 1148
rect 214340 532 214396 588
rect 217140 868 217196 924
rect 219604 1092 219660 1148
rect 217364 420 217420 476
<< metal3 >>
rect 42298 14868 42308 14924
rect 42364 14868 54404 14924
rect 54460 14868 54470 14924
rect 63130 14868 63140 14924
rect 63196 14868 67004 14924
rect 67890 14868 67900 14924
rect 67956 14868 83524 14924
rect 83580 14868 83590 14924
rect 83738 14868 83748 14924
rect 83804 14868 102452 14924
rect 102508 14868 102518 14924
rect 102666 14868 102676 14924
rect 102732 14868 103012 14924
rect 103068 14868 103078 14924
rect 103236 14868 115220 14924
rect 115276 14868 115286 14924
rect 115434 14868 115444 14924
rect 115500 14868 118020 14924
rect 118076 14868 118086 14924
rect 118570 14868 118580 14924
rect 118636 14868 120148 14924
rect 120204 14868 120214 14924
rect 120922 14868 120932 14924
rect 120988 14868 151396 14924
rect 151452 14868 151462 14924
rect 151610 14868 151620 14924
rect 151676 14868 161532 14924
rect 161588 14868 161598 14924
rect 172666 14868 172676 14924
rect 172732 14868 181972 14924
rect 182028 14868 182038 14924
rect 66948 14812 67004 14868
rect 103236 14812 103292 14868
rect 23370 14756 23380 14812
rect 23436 14756 66892 14812
rect 66948 14756 70196 14812
rect 70252 14756 70262 14812
rect 70410 14756 70420 14812
rect 70476 14756 71652 14812
rect 71708 14756 71718 14812
rect 71866 14756 71876 14812
rect 71932 14756 77588 14812
rect 77644 14756 77654 14812
rect 77812 14756 80836 14812
rect 80892 14756 80902 14812
rect 81060 14756 82180 14812
rect 82236 14756 82246 14812
rect 82842 14756 82852 14812
rect 82908 14756 98084 14812
rect 98140 14756 98150 14812
rect 98298 14756 98308 14812
rect 98364 14756 100436 14812
rect 100492 14756 100502 14812
rect 101322 14756 101332 14812
rect 101388 14756 103292 14812
rect 103348 14756 111412 14812
rect 111468 14756 111478 14812
rect 113642 14756 113652 14812
rect 113708 14756 174692 14812
rect 174748 14756 174758 14812
rect 66836 14700 66892 14756
rect 77812 14700 77868 14756
rect 81060 14700 81116 14756
rect 103348 14700 103404 14756
rect 42970 14644 42980 14700
rect 43036 14644 52948 14700
rect 53004 14644 53014 14700
rect 53610 14644 53620 14700
rect 53676 14644 63980 14700
rect 66836 14644 77868 14700
rect 77924 14644 79156 14700
rect 79212 14644 79222 14700
rect 79380 14644 81116 14700
rect 81274 14644 81284 14700
rect 81340 14644 100660 14700
rect 100716 14644 100726 14700
rect 100884 14644 103404 14700
rect 103898 14644 103908 14700
rect 103964 14644 121044 14700
rect 121100 14644 121110 14700
rect 121258 14644 121268 14700
rect 121324 14644 124628 14700
rect 124684 14644 124694 14700
rect 126756 14644 149660 14700
rect 151050 14644 151060 14700
rect 151116 14644 153076 14700
rect 153132 14644 153142 14700
rect 153514 14644 153524 14700
rect 153580 14644 155596 14700
rect 156090 14644 156100 14700
rect 156156 14644 157108 14700
rect 157164 14644 157174 14700
rect 159460 14644 162484 14700
rect 162540 14644 162550 14700
rect 163258 14644 163268 14700
rect 163324 14644 176427 14700
rect 63924 14588 63980 14644
rect 77924 14588 77980 14644
rect 79380 14588 79436 14644
rect 100884 14588 100940 14644
rect 126756 14588 126812 14644
rect 45658 14532 45668 14588
rect 45724 14532 58772 14588
rect 58828 14532 58838 14588
rect 63924 14532 65380 14588
rect 65436 14532 65446 14588
rect 65594 14532 65604 14588
rect 65660 14532 77700 14588
rect 77756 14532 77766 14588
rect 77914 14532 77924 14588
rect 77980 14532 77990 14588
rect 78138 14532 78148 14588
rect 78204 14532 79436 14588
rect 79594 14532 79604 14588
rect 79660 14532 80388 14588
rect 80444 14532 80454 14588
rect 80602 14532 80612 14588
rect 80668 14532 92596 14588
rect 92652 14532 92662 14588
rect 92810 14532 92820 14588
rect 92876 14532 98308 14588
rect 98364 14532 98374 14588
rect 98522 14532 98532 14588
rect 98588 14532 100940 14588
rect 101098 14532 101108 14588
rect 101164 14532 102564 14588
rect 102620 14532 102630 14588
rect 102778 14532 102788 14588
rect 102844 14532 113764 14588
rect 113820 14532 113830 14588
rect 113978 14532 113988 14588
rect 114044 14532 120372 14588
rect 120428 14532 120438 14588
rect 120698 14532 120708 14588
rect 120764 14532 126812 14588
rect 126868 14532 149380 14588
rect 149436 14532 149446 14588
rect 126868 14476 126924 14532
rect 149604 14476 149660 14644
rect 155540 14588 155596 14644
rect 159460 14588 159516 14644
rect 176371 14588 176427 14644
rect 151274 14532 151284 14588
rect 151340 14532 155484 14588
rect 155540 14532 159516 14588
rect 162250 14532 162260 14588
rect 162316 14532 175588 14588
rect 175644 14532 175654 14588
rect 176371 14532 176820 14588
rect 176876 14532 176886 14588
rect 155428 14476 155484 14532
rect 16650 14420 16660 14476
rect 16716 14420 82068 14476
rect 82124 14420 82134 14476
rect 82282 14420 82292 14476
rect 82348 14420 82628 14476
rect 82684 14420 82694 14476
rect 82842 14420 82852 14476
rect 82908 14420 114492 14476
rect 114874 14420 114884 14476
rect 114940 14420 114996 14476
rect 115052 14420 115062 14476
rect 115210 14420 115220 14476
rect 115276 14420 117796 14476
rect 117852 14420 117862 14476
rect 118010 14420 118020 14476
rect 118076 14420 118804 14476
rect 118860 14420 118870 14476
rect 119354 14420 119364 14476
rect 119420 14420 119924 14476
rect 119980 14420 119990 14476
rect 120474 14420 120484 14476
rect 120540 14420 121044 14476
rect 121100 14420 121110 14476
rect 121482 14420 121492 14476
rect 121548 14420 122948 14476
rect 123004 14420 123014 14476
rect 124366 14420 124404 14476
rect 124460 14420 124470 14476
rect 124618 14420 124628 14476
rect 124684 14420 126924 14476
rect 132691 14420 149156 14476
rect 149212 14420 149222 14476
rect 149604 14420 151004 14476
rect 151498 14420 151508 14476
rect 151564 14420 155204 14476
rect 155260 14420 155270 14476
rect 155428 14420 156212 14476
rect 156268 14420 156278 14476
rect 156426 14420 156436 14476
rect 156492 14420 169764 14476
rect 169820 14420 169830 14476
rect 114436 14364 114492 14420
rect 132691 14364 132747 14420
rect 150948 14364 151004 14420
rect 8371 14308 58324 14364
rect 58380 14308 58390 14364
rect 64138 14308 64148 14364
rect 64204 14308 69860 14364
rect 69916 14308 69926 14364
rect 70074 14308 70084 14364
rect 70140 14308 77476 14364
rect 77532 14308 77542 14364
rect 77812 14308 114212 14364
rect 114268 14308 114278 14364
rect 114436 14308 120708 14364
rect 120764 14308 120774 14364
rect 121034 14308 121044 14364
rect 121100 14308 132747 14364
rect 134138 14308 134148 14364
rect 134204 14308 134708 14364
rect 134764 14308 134774 14364
rect 139402 14308 139412 14364
rect 139468 14308 150724 14364
rect 150780 14308 150790 14364
rect 150948 14308 156772 14364
rect 156828 14308 156838 14364
rect 157098 14308 157108 14364
rect 157164 14308 171332 14364
rect 171388 14308 171398 14364
rect 173572 14308 182756 14364
rect 182812 14308 182822 14364
rect 8371 14140 8427 14308
rect 20131 14196 77588 14252
rect 77644 14196 77654 14252
rect 20131 14140 20187 14196
rect 77812 14140 77868 14308
rect 78138 14196 78148 14252
rect 78204 14196 79492 14252
rect 79548 14196 79558 14252
rect 79706 14196 79716 14252
rect 79772 14196 103348 14252
rect 103404 14196 103414 14252
rect 104010 14196 104020 14252
rect 104076 14196 116340 14252
rect 116396 14196 116406 14252
rect 116554 14196 116564 14252
rect 116620 14196 117236 14252
rect 117292 14196 117302 14252
rect 117786 14196 117796 14252
rect 117852 14196 118132 14252
rect 118188 14196 118198 14252
rect 118346 14196 118356 14252
rect 118412 14196 142660 14252
rect 142716 14196 142726 14252
rect 149230 14196 149268 14252
rect 149324 14196 149334 14252
rect 149818 14196 149828 14252
rect 149884 14196 151284 14252
rect 151340 14196 151350 14252
rect 152730 14196 152740 14252
rect 152796 14196 152852 14252
rect 152908 14196 152918 14252
rect 153066 14196 153076 14252
rect 153132 14196 158676 14252
rect 158732 14196 158742 14252
rect 158890 14196 158900 14252
rect 158956 14196 169092 14252
rect 169148 14196 169158 14252
rect 173572 14140 173628 14308
rect 174122 14196 174132 14252
rect 174188 14196 188692 14252
rect 188748 14196 188758 14252
rect 7690 14084 7700 14140
rect 7756 14084 8427 14140
rect 17098 14084 17108 14140
rect 17164 14084 20187 14140
rect 21438 14084 21476 14140
rect 21532 14084 21542 14140
rect 58314 14084 58324 14140
rect 58380 14084 69636 14140
rect 69692 14084 69702 14140
rect 71754 14084 71764 14140
rect 71820 14084 77252 14140
rect 77308 14084 77318 14140
rect 77476 14084 77868 14140
rect 78026 14084 78036 14140
rect 78092 14084 79044 14140
rect 79100 14084 79110 14140
rect 79594 14084 79604 14140
rect 79660 14084 80612 14140
rect 80668 14084 80678 14140
rect 80826 14084 80836 14140
rect 80892 14084 124516 14140
rect 124572 14084 124582 14140
rect 124730 14084 124740 14140
rect 124796 14084 140756 14140
rect 140812 14084 140822 14140
rect 144451 14084 153860 14140
rect 153916 14084 153926 14140
rect 154074 14084 154084 14140
rect 154140 14084 173628 14140
rect 174682 14084 174692 14140
rect 174748 14084 175476 14140
rect 175532 14084 175542 14140
rect 182970 14084 182980 14140
rect 183036 14084 193956 14140
rect 194012 14084 194022 14140
rect 77476 14028 77532 14084
rect 144451 14028 144507 14084
rect 14830 13972 14868 14028
rect 14924 13972 14934 14028
rect 17742 13972 17780 14028
rect 17836 13972 17846 14028
rect 20131 13972 77532 14028
rect 77690 13972 77700 14028
rect 77756 13972 78484 14028
rect 78540 13972 78550 14028
rect 78698 13972 78708 14028
rect 78764 13972 78802 14028
rect 79146 13972 79156 14028
rect 79212 13972 80948 14028
rect 81004 13972 81014 14028
rect 81274 13972 81284 14028
rect 81340 13972 92372 14028
rect 92428 13972 92438 14028
rect 92586 13972 92596 14028
rect 92652 13972 97300 14028
rect 97356 13972 97366 14028
rect 97514 13972 97524 14028
rect 97580 13972 115052 14028
rect 115406 13972 115444 14028
rect 115500 13972 115510 14028
rect 115994 13972 116004 14028
rect 116060 13972 134036 14028
rect 134092 13972 134102 14028
rect 134250 13972 134260 14028
rect 134316 13972 144507 14028
rect 148698 13972 148708 14028
rect 148764 13972 150500 14028
rect 150556 13972 150566 14028
rect 151162 13972 151172 14028
rect 151228 13972 156212 14028
rect 156268 13972 156278 14028
rect 156426 13972 156436 14028
rect 156492 13972 159180 14028
rect 159450 13972 159460 14028
rect 159516 13972 159572 14028
rect 159628 13972 159638 14028
rect 162670 13972 162708 14028
rect 162764 13972 162774 14028
rect 166842 13972 166852 14028
rect 166908 13972 178052 14028
rect 178108 13972 178118 14028
rect 179162 13972 179172 14028
rect 179228 13972 187572 14028
rect 187628 13972 187638 14028
rect 191118 13972 191156 14028
rect 191212 13972 191222 14028
rect 20131 13916 20187 13972
rect 114996 13916 115052 13972
rect 159124 13916 159180 13972
rect 14074 13860 14084 13916
rect 14140 13860 20187 13916
rect 25022 13860 25060 13916
rect 25116 13860 25126 13916
rect 31891 13860 59612 13916
rect 61450 13860 61460 13916
rect 61516 13860 71876 13916
rect 71932 13860 71942 13916
rect 73098 13860 73108 13916
rect 73164 13860 74508 13916
rect 74638 13860 74676 13916
rect 74732 13860 74742 13916
rect 74890 13860 74900 13916
rect 74956 13860 77140 13916
rect 77196 13860 77206 13916
rect 77354 13860 77364 13916
rect 77420 13860 81732 13916
rect 81788 13860 81798 13916
rect 82058 13860 82068 13916
rect 82124 13860 82292 13916
rect 82348 13860 82358 13916
rect 83066 13860 83076 13916
rect 83132 13860 92484 13916
rect 92540 13860 92550 13916
rect 92698 13860 92708 13916
rect 92764 13860 99652 13916
rect 99708 13860 99718 13916
rect 99866 13860 99876 13916
rect 99932 13860 114772 13916
rect 114828 13860 114838 13916
rect 114996 13860 117684 13916
rect 117740 13860 117750 13916
rect 117898 13860 117908 13916
rect 117964 13860 118002 13916
rect 118122 13860 118132 13916
rect 118188 13860 118580 13916
rect 118636 13860 118646 13916
rect 118794 13860 118804 13916
rect 118860 13860 119700 13916
rect 119756 13860 119766 13916
rect 120138 13860 120148 13916
rect 120204 13860 126756 13916
rect 126812 13860 126822 13916
rect 126970 13860 126980 13916
rect 127036 13860 138068 13916
rect 138124 13860 138134 13916
rect 138282 13860 138292 13916
rect 138348 13860 138740 13916
rect 138796 13860 138806 13916
rect 139486 13860 139524 13916
rect 139580 13860 139590 13916
rect 144106 13860 144116 13916
rect 144172 13860 157668 13916
rect 157724 13860 157734 13916
rect 158302 13860 158340 13916
rect 158396 13860 158406 13916
rect 159124 13860 172452 13916
rect 172508 13860 172518 13916
rect 174430 13860 174468 13916
rect 174524 13860 174534 13916
rect 181738 13860 181748 13916
rect 181804 13860 191828 13916
rect 191884 13860 191894 13916
rect 193358 13860 193396 13916
rect 193452 13860 193462 13916
rect 31891 13804 31947 13860
rect 59556 13804 59612 13860
rect 74452 13804 74508 13860
rect 12618 13748 12628 13804
rect 12684 13748 31947 13804
rect 57054 13748 57092 13804
rect 57148 13748 57158 13804
rect 59556 13748 74228 13804
rect 74284 13748 74294 13804
rect 74452 13748 76916 13804
rect 76972 13748 76982 13804
rect 77130 13748 77140 13804
rect 77196 13748 82852 13804
rect 82908 13748 82918 13804
rect 83066 13748 83076 13804
rect 83132 13748 91028 13804
rect 91084 13748 91094 13804
rect 91196 13748 113652 13804
rect 113708 13748 113718 13804
rect 113866 13748 113876 13804
rect 113932 13748 115892 13804
rect 115948 13748 115958 13804
rect 116228 13748 116340 13804
rect 116396 13748 116406 13804
rect 116554 13748 116564 13804
rect 116620 13748 120596 13804
rect 120652 13748 120662 13804
rect 120810 13748 120820 13804
rect 120876 13748 124292 13804
rect 124348 13748 124358 13804
rect 124506 13748 124516 13804
rect 124572 13748 140084 13804
rect 140140 13748 140150 13804
rect 148362 13748 148372 13804
rect 148428 13748 152964 13804
rect 153020 13748 153030 13804
rect 153178 13748 153188 13804
rect 153244 13748 155540 13804
rect 155596 13748 155606 13804
rect 155866 13748 155876 13804
rect 155932 13748 174916 13804
rect 174972 13748 174982 13804
rect 183166 13748 183204 13804
rect 183260 13748 183270 13804
rect 183428 13748 196308 13804
rect 196364 13748 196374 13804
rect 91196 13692 91252 13748
rect 116228 13692 116284 13748
rect 183428 13692 183484 13748
rect 219200 13692 220000 13720
rect 32330 13636 32340 13692
rect 32396 13636 61236 13692
rect 61292 13636 61302 13692
rect 61786 13636 61796 13692
rect 61852 13636 65604 13692
rect 65660 13636 65670 13692
rect 65902 13636 65940 13692
rect 65996 13636 66006 13692
rect 66714 13636 66724 13692
rect 66780 13636 67732 13692
rect 67788 13636 67798 13692
rect 67900 13636 81844 13692
rect 81900 13636 81910 13692
rect 82058 13636 82068 13692
rect 82124 13636 91252 13692
rect 92474 13636 92484 13692
rect 92540 13636 102788 13692
rect 102844 13636 102854 13692
rect 102956 13636 116284 13692
rect 116442 13636 116452 13692
rect 116508 13636 138572 13692
rect 142650 13636 142660 13692
rect 142716 13636 146020 13692
rect 146076 13636 146086 13692
rect 147886 13636 147924 13692
rect 147980 13636 147990 13692
rect 148138 13636 148148 13692
rect 148204 13636 151844 13692
rect 151900 13636 151910 13692
rect 152058 13636 152068 13692
rect 152124 13636 163492 13692
rect 163548 13636 163558 13692
rect 163716 13636 173852 13692
rect 174010 13636 174020 13692
rect 174076 13636 182308 13692
rect 182364 13636 182374 13692
rect 182858 13636 182868 13692
rect 182924 13636 183484 13692
rect 186218 13636 186228 13692
rect 186284 13636 201460 13692
rect 201516 13636 202804 13692
rect 202860 13636 202870 13692
rect 209850 13636 209860 13692
rect 209916 13636 220000 13692
rect 67900 13580 67956 13636
rect 102956 13580 103012 13636
rect 138516 13580 138572 13636
rect 163716 13580 163772 13636
rect 10462 13524 10500 13580
rect 10556 13524 10566 13580
rect 38826 13524 38836 13580
rect 38892 13524 64036 13580
rect 64092 13524 64102 13580
rect 64250 13524 64260 13580
rect 64316 13524 67956 13580
rect 68058 13524 68068 13580
rect 68124 13524 68162 13580
rect 68282 13524 68292 13580
rect 68348 13524 83188 13580
rect 83244 13524 83254 13580
rect 83402 13524 83412 13580
rect 83468 13524 83748 13580
rect 83804 13524 83814 13580
rect 83962 13524 83972 13580
rect 84028 13524 84980 13580
rect 85036 13524 85046 13580
rect 85194 13524 85204 13580
rect 85260 13524 90636 13580
rect 91242 13524 91252 13580
rect 91308 13524 97076 13580
rect 97132 13524 97142 13580
rect 97290 13524 97300 13580
rect 97356 13524 98980 13580
rect 99036 13524 99046 13580
rect 99194 13524 99204 13580
rect 99260 13524 103012 13580
rect 103786 13524 103796 13580
rect 103852 13524 119252 13580
rect 119308 13524 119318 13580
rect 119466 13524 119476 13580
rect 119532 13524 120372 13580
rect 120428 13524 120438 13580
rect 120586 13524 120596 13580
rect 120652 13524 135604 13580
rect 135660 13524 135670 13580
rect 138516 13524 149268 13580
rect 149324 13524 149334 13580
rect 149482 13524 149492 13580
rect 149548 13524 157220 13580
rect 157276 13524 157286 13580
rect 162250 13524 162260 13580
rect 162316 13524 163772 13580
rect 163930 13524 163940 13580
rect 163996 13524 173572 13580
rect 173628 13524 173638 13580
rect 90580 13468 90636 13524
rect 173796 13468 173852 13636
rect 219200 13608 220000 13636
rect 174010 13524 174020 13580
rect 174076 13524 184660 13580
rect 184716 13524 184726 13580
rect 185658 13524 185668 13580
rect 185724 13524 198436 13580
rect 198492 13524 198502 13580
rect 25694 13412 25732 13468
rect 25788 13412 25798 13468
rect 53806 13412 53844 13468
rect 53900 13412 53910 13468
rect 60442 13412 60452 13468
rect 60508 13412 63700 13468
rect 63756 13412 63766 13468
rect 63914 13412 63924 13468
rect 63980 13412 74004 13468
rect 74060 13412 74070 13468
rect 74218 13412 74228 13468
rect 74284 13412 76916 13468
rect 76972 13412 76982 13468
rect 77130 13412 77140 13468
rect 77196 13412 77588 13468
rect 77644 13412 77654 13468
rect 77802 13412 77812 13468
rect 77868 13412 82292 13468
rect 82348 13412 82358 13468
rect 82506 13412 82516 13468
rect 82572 13412 90356 13468
rect 90412 13412 90422 13468
rect 90580 13412 117796 13468
rect 117852 13412 117862 13468
rect 118010 13412 118020 13468
rect 118076 13412 124740 13468
rect 124796 13412 124806 13468
rect 126746 13412 126756 13468
rect 126812 13412 136500 13468
rect 136556 13412 136566 13468
rect 137946 13412 137956 13468
rect 138012 13412 148148 13468
rect 148204 13412 148214 13468
rect 148334 13412 148372 13468
rect 148428 13412 148438 13468
rect 150154 13412 150164 13468
rect 150220 13412 152068 13468
rect 152124 13412 152134 13468
rect 152282 13412 152292 13468
rect 152348 13412 154756 13468
rect 154812 13412 154822 13468
rect 154970 13412 154980 13468
rect 155036 13412 164164 13468
rect 164220 13412 164230 13468
rect 167962 13412 167972 13468
rect 168028 13412 171836 13468
rect 173796 13412 187572 13468
rect 187628 13412 187638 13468
rect 298 13300 308 13356
rect 364 13300 10612 13356
rect 10668 13300 10678 13356
rect 19226 13300 19236 13356
rect 19292 13300 54404 13356
rect 54460 13300 54470 13356
rect 55738 13300 55748 13356
rect 55804 13300 82404 13356
rect 82460 13300 82470 13356
rect 82730 13300 82740 13356
rect 82796 13300 82834 13356
rect 83290 13300 83300 13356
rect 83356 13300 83636 13356
rect 83692 13300 83702 13356
rect 83850 13300 83860 13356
rect 83916 13300 103012 13356
rect 103068 13300 103078 13356
rect 103226 13300 103236 13356
rect 103292 13300 149380 13356
rect 149436 13300 149446 13356
rect 149818 13300 149828 13356
rect 149884 13300 155092 13356
rect 155148 13300 155158 13356
rect 155306 13300 155316 13356
rect 155372 13300 159124 13356
rect 159180 13300 159190 13356
rect 161466 13300 161476 13356
rect 161532 13300 165228 13356
rect 165386 13300 165396 13356
rect 165452 13300 171556 13356
rect 171612 13300 171622 13356
rect 165172 13244 165228 13300
rect 171780 13244 171836 13412
rect 172442 13300 172452 13356
rect 172508 13300 177156 13356
rect 177212 13300 177222 13356
rect 179274 13300 179284 13356
rect 179340 13300 189028 13356
rect 189084 13300 189094 13356
rect 211614 13300 211652 13356
rect 211708 13300 211718 13356
rect 970 13188 980 13244
rect 1036 13188 10724 13244
rect 10780 13188 10790 13244
rect 18414 13188 18452 13244
rect 18508 13188 18518 13244
rect 23594 13188 23604 13244
rect 23660 13188 51044 13244
rect 51100 13188 51110 13244
rect 53022 13188 53060 13244
rect 53116 13188 53126 13244
rect 57754 13188 57764 13244
rect 57820 13188 68068 13244
rect 68124 13188 68134 13244
rect 68282 13188 68292 13244
rect 68348 13188 73780 13244
rect 73836 13188 73846 13244
rect 73994 13188 74004 13244
rect 74060 13188 77252 13244
rect 77308 13188 77318 13244
rect 77466 13188 77476 13244
rect 77532 13188 118804 13244
rect 118860 13188 118870 13244
rect 119028 13188 126980 13244
rect 127036 13188 127046 13244
rect 133466 13188 133476 13244
rect 133532 13188 134260 13244
rect 134316 13188 134326 13244
rect 135594 13188 135604 13244
rect 135660 13188 140476 13244
rect 142986 13188 142996 13244
rect 143052 13188 146916 13244
rect 146972 13188 146982 13244
rect 147130 13188 147140 13244
rect 147196 13188 159796 13244
rect 159852 13188 159862 13244
rect 161018 13188 161028 13244
rect 161084 13188 162596 13244
rect 162652 13188 162662 13244
rect 164910 13188 164948 13244
rect 165004 13188 165014 13244
rect 165172 13188 170940 13244
rect 171780 13188 174132 13244
rect 174188 13188 174198 13244
rect 179498 13188 179508 13244
rect 179564 13188 190596 13244
rect 190652 13188 190662 13244
rect 119028 13132 119084 13188
rect 140420 13132 140476 13188
rect 3882 13076 3892 13132
rect 3948 13076 11620 13132
rect 11676 13076 11686 13132
rect 15530 13076 15540 13132
rect 15596 13076 58212 13132
rect 58268 13076 58278 13132
rect 66490 13076 66500 13132
rect 66556 13076 73220 13132
rect 73276 13076 73286 13132
rect 73434 13076 73444 13132
rect 73500 13076 74228 13132
rect 74284 13076 74294 13132
rect 74442 13076 74452 13132
rect 74508 13076 77140 13132
rect 77196 13076 77206 13132
rect 77578 13076 77588 13132
rect 77644 13076 78148 13132
rect 78474 13076 78484 13132
rect 78540 13076 80724 13132
rect 80780 13076 80790 13132
rect 81050 13076 81060 13132
rect 81116 13076 83524 13132
rect 83580 13076 83590 13132
rect 83738 13076 83748 13132
rect 83804 13076 84644 13132
rect 84700 13076 84710 13132
rect 84858 13076 84868 13132
rect 84924 13076 84962 13132
rect 85194 13076 85204 13132
rect 85260 13076 86660 13132
rect 86716 13076 86726 13132
rect 86986 13076 86996 13132
rect 87052 13076 88676 13132
rect 88732 13076 88742 13132
rect 88900 13076 103012 13132
rect 103068 13076 103078 13132
rect 103338 13076 103348 13132
rect 103404 13076 115556 13132
rect 115612 13076 115622 13132
rect 115882 13076 115892 13132
rect 115948 13076 119084 13132
rect 119140 13076 119700 13132
rect 119756 13076 119766 13132
rect 119914 13076 119924 13132
rect 119980 13076 132356 13132
rect 132412 13076 132422 13132
rect 132682 13076 132692 13132
rect 132748 13076 140196 13132
rect 140252 13076 140262 13132
rect 140420 13076 148932 13132
rect 148988 13076 148998 13132
rect 149146 13076 149156 13132
rect 149212 13076 149492 13132
rect 149548 13076 149558 13132
rect 149706 13076 149716 13132
rect 149772 13076 154308 13132
rect 154364 13076 154374 13132
rect 154634 13076 154644 13132
rect 154700 13076 167860 13132
rect 167916 13076 167926 13132
rect 78092 13020 78148 13076
rect 88900 13020 88956 13076
rect 119140 13020 119196 13076
rect 170884 13020 170940 13188
rect 171098 13076 171108 13132
rect 171164 13076 185612 13132
rect 185770 13076 185780 13132
rect 185836 13076 200676 13132
rect 200732 13076 200742 13132
rect 185556 13020 185612 13076
rect 3210 12964 3220 13020
rect 3276 12964 9828 13020
rect 9884 12964 9894 13020
rect 27934 12964 27972 13020
rect 28028 12964 28038 13020
rect 34430 12964 34468 13020
rect 34524 12964 34534 13020
rect 46442 12964 46452 13020
rect 46508 12964 60004 13020
rect 60060 12964 60070 13020
rect 60778 12964 60788 13020
rect 60844 12964 63924 13020
rect 64026 12964 64036 13020
rect 64092 12964 77140 13020
rect 77196 12964 77206 13020
rect 77354 12964 77364 13020
rect 77420 12964 77924 13020
rect 77980 12964 77990 13020
rect 78092 12964 78932 13020
rect 78988 12964 78998 13020
rect 79258 12964 79268 13020
rect 79324 12964 88956 13020
rect 89450 12964 89460 13020
rect 89516 12964 91252 13020
rect 91308 12964 91318 13020
rect 91466 12964 91476 13020
rect 91532 12964 103236 13020
rect 103292 12964 103302 13020
rect 103562 12964 103572 13020
rect 103628 12964 104132 13020
rect 104188 12964 104198 13020
rect 104346 12964 104356 13020
rect 104412 12964 109452 13020
rect 109610 12964 109620 13020
rect 109676 12964 119196 13020
rect 119354 12964 119364 13020
rect 119420 12964 122724 13020
rect 122780 12964 122790 13020
rect 122938 12964 122948 13020
rect 123004 12964 124796 13020
rect 124954 12964 124964 13020
rect 125020 12964 134484 13020
rect 134540 12964 134550 13020
rect 135818 12964 135828 13020
rect 135884 12964 146692 13020
rect 146748 12964 146758 13020
rect 146906 12964 146916 13020
rect 146972 12964 148932 13020
rect 148988 12964 148998 13020
rect 149146 12964 149156 13020
rect 149212 12964 159348 13020
rect 159404 12964 159414 13020
rect 161018 12964 161028 13020
rect 161084 12964 165396 13020
rect 165452 12964 165462 13020
rect 165694 12964 165732 13020
rect 165788 12964 165798 13020
rect 170884 12964 180964 13020
rect 181020 12964 181030 13020
rect 185294 12964 185332 13020
rect 185388 12964 185398 13020
rect 185556 12964 193620 13020
rect 193676 12964 193686 13020
rect 195486 12964 195524 13020
rect 195580 12964 195590 13020
rect 205258 12964 205268 13020
rect 205324 12964 208628 13020
rect 208684 12964 208694 13020
rect 63868 12908 63924 12964
rect 109396 12908 109452 12964
rect 124740 12908 124796 12964
rect 6122 12852 6132 12908
rect 6188 12852 55972 12908
rect 56028 12852 56038 12908
rect 56186 12852 56196 12908
rect 56252 12852 62244 12908
rect 62300 12852 62310 12908
rect 63868 12852 73556 12908
rect 73612 12852 73622 12908
rect 73770 12852 73780 12908
rect 73836 12852 75012 12908
rect 75068 12852 75078 12908
rect 75226 12852 75236 12908
rect 75292 12852 77028 12908
rect 77084 12852 77094 12908
rect 77364 12852 103684 12908
rect 103740 12852 103750 12908
rect 103898 12852 103908 12908
rect 103964 12852 104244 12908
rect 104300 12852 104310 12908
rect 104654 12852 104692 12908
rect 104748 12852 104758 12908
rect 105354 12852 105364 12908
rect 105420 12852 109172 12908
rect 109228 12852 109238 12908
rect 109396 12852 114324 12908
rect 114380 12852 114390 12908
rect 114538 12852 114548 12908
rect 114604 12852 119140 12908
rect 119196 12852 119206 12908
rect 119354 12852 119364 12908
rect 119420 12852 124516 12908
rect 124572 12852 124582 12908
rect 124740 12852 137396 12908
rect 137452 12852 137462 12908
rect 137610 12852 137620 12908
rect 137676 12852 142436 12908
rect 142492 12852 142502 12908
rect 142650 12852 142660 12908
rect 142716 12852 142772 12908
rect 142828 12852 142838 12908
rect 144218 12852 144228 12908
rect 144284 12852 145348 12908
rect 145404 12852 145414 12908
rect 147018 12852 147028 12908
rect 147084 12852 152516 12908
rect 152572 12852 152582 12908
rect 152842 12852 152852 12908
rect 152908 12852 161924 12908
rect 161980 12852 161990 12908
rect 162138 12852 162148 12908
rect 162204 12852 173796 12908
rect 173852 12852 173862 12908
rect 182522 12852 182532 12908
rect 182588 12852 196532 12908
rect 196588 12852 196598 12908
rect 204810 12852 204820 12908
rect 204876 12852 210084 12908
rect 210140 12852 210150 12908
rect 77364 12796 77420 12852
rect 27150 12740 27188 12796
rect 27244 12740 27254 12796
rect 36698 12740 36708 12796
rect 36764 12740 77420 12796
rect 77756 12684 77812 12796
rect 77868 12740 77878 12796
rect 78026 12740 78036 12796
rect 78092 12740 78820 12796
rect 78876 12740 78886 12796
rect 79594 12740 79604 12796
rect 79660 12740 80500 12796
rect 80556 12740 80566 12796
rect 80826 12740 80836 12796
rect 80892 12740 83412 12796
rect 83468 12740 83478 12796
rect 83850 12740 83860 12796
rect 83916 12740 91476 12796
rect 91532 12740 91542 12796
rect 91690 12740 91700 12796
rect 91756 12740 101780 12796
rect 101836 12740 101846 12796
rect 101994 12740 102004 12796
rect 102060 12740 102564 12796
rect 102620 12740 102630 12796
rect 102778 12740 102788 12796
rect 102844 12740 107380 12796
rect 107436 12740 107446 12796
rect 107930 12740 107940 12796
rect 107996 12740 119812 12796
rect 119868 12740 119878 12796
rect 120026 12740 120036 12796
rect 120092 12740 120708 12796
rect 120764 12740 120774 12796
rect 120922 12740 120932 12796
rect 120988 12740 127316 12796
rect 127372 12740 127382 12796
rect 137834 12740 137844 12796
rect 137900 12740 149156 12796
rect 149212 12740 149222 12796
rect 149482 12740 149492 12796
rect 149548 12740 150948 12796
rect 151004 12740 151014 12796
rect 151162 12740 151172 12796
rect 151228 12740 173460 12796
rect 173516 12740 173526 12796
rect 173674 12740 173684 12796
rect 173740 12740 177268 12796
rect 177324 12740 177334 12796
rect 177482 12740 177492 12796
rect 177548 12740 186788 12796
rect 186844 12740 186854 12796
rect 196298 12740 196308 12796
rect 196364 12740 198660 12796
rect 198716 12740 198726 12796
rect 11946 12628 11956 12684
rect 12012 12628 43652 12684
rect 43708 12628 43718 12684
rect 59210 12628 59220 12684
rect 59276 12628 68628 12684
rect 68684 12628 68694 12684
rect 69514 12628 69524 12684
rect 69580 12628 73108 12684
rect 73164 12628 73174 12684
rect 73546 12628 73556 12684
rect 73612 12628 77812 12684
rect 77914 12628 77924 12684
rect 77980 12628 94948 12684
rect 95004 12628 95014 12684
rect 96058 12628 96068 12684
rect 96124 12628 102004 12684
rect 102060 12628 102070 12684
rect 102330 12628 102340 12684
rect 102396 12628 114772 12684
rect 114828 12628 114838 12684
rect 114986 12628 114996 12684
rect 115052 12628 137620 12684
rect 137676 12628 137686 12684
rect 137834 12628 137844 12684
rect 137900 12628 143108 12684
rect 143164 12628 143174 12684
rect 144451 12628 149268 12684
rect 149324 12628 149334 12684
rect 149930 12628 149940 12684
rect 149996 12628 151060 12684
rect 151116 12628 151126 12684
rect 151274 12628 151284 12684
rect 151340 12628 174020 12684
rect 174076 12628 174086 12684
rect 174234 12628 174244 12684
rect 174300 12628 180292 12684
rect 180348 12628 180358 12684
rect 180842 12628 180852 12684
rect 180908 12628 187124 12684
rect 187180 12628 187190 12684
rect 193834 12628 193844 12684
rect 193900 12628 200900 12684
rect 200956 12628 200966 12684
rect 144451 12572 144507 12628
rect 30062 12516 30100 12572
rect 30156 12516 30166 12572
rect 31546 12516 31556 12572
rect 31612 12516 68852 12572
rect 68908 12516 68918 12572
rect 69066 12516 69076 12572
rect 69132 12516 78148 12572
rect 78204 12516 78214 12572
rect 78362 12516 78372 12572
rect 78428 12516 78932 12572
rect 78988 12516 78998 12572
rect 79146 12516 79156 12572
rect 79212 12516 79380 12572
rect 79436 12516 79446 12572
rect 80042 12516 80052 12572
rect 80108 12516 80164 12572
rect 80220 12516 80230 12572
rect 80378 12516 80388 12572
rect 80444 12516 80948 12572
rect 81004 12516 81014 12572
rect 81274 12516 81284 12572
rect 81340 12516 81350 12572
rect 81722 12516 81732 12572
rect 81788 12516 83076 12572
rect 83132 12516 83142 12572
rect 83402 12516 83412 12572
rect 83468 12516 84308 12572
rect 84364 12516 84374 12572
rect 84718 12516 84756 12572
rect 84812 12516 84822 12572
rect 84970 12516 84980 12572
rect 85036 12516 86548 12572
rect 86604 12516 86614 12572
rect 87770 12516 87780 12572
rect 87836 12516 91700 12572
rect 91756 12516 91766 12572
rect 91914 12516 91924 12572
rect 91980 12516 92932 12572
rect 92988 12516 92998 12572
rect 97066 12516 97076 12572
rect 97132 12516 104244 12572
rect 104300 12516 104310 12572
rect 105242 12516 105252 12572
rect 105308 12516 111748 12572
rect 111804 12516 111814 12572
rect 112074 12516 112084 12572
rect 112140 12516 114212 12572
rect 114268 12516 114278 12572
rect 114426 12516 114436 12572
rect 114492 12516 116228 12572
rect 116284 12516 116294 12572
rect 117114 12516 117124 12572
rect 117180 12516 120484 12572
rect 120540 12516 120550 12572
rect 120698 12516 120708 12572
rect 120764 12516 126812 12572
rect 126970 12516 126980 12572
rect 127036 12516 144507 12572
rect 148670 12516 148708 12572
rect 148764 12516 148774 12572
rect 149034 12516 149044 12572
rect 149100 12516 154756 12572
rect 154812 12516 154822 12572
rect 154980 12516 156492 12572
rect 0 12460 800 12488
rect 81284 12460 81340 12516
rect 126756 12460 126812 12516
rect 154980 12460 155036 12516
rect 156436 12460 156492 12516
rect 158452 12516 195412 12572
rect 195468 12516 195478 12572
rect 0 12404 6692 12460
rect 6748 12404 6758 12460
rect 13402 12404 13412 12460
rect 13468 12404 62972 12460
rect 63242 12404 63252 12460
rect 63308 12404 69748 12460
rect 69804 12404 69814 12460
rect 69962 12404 69972 12460
rect 70028 12404 73556 12460
rect 73612 12404 73622 12460
rect 73994 12404 74004 12460
rect 74060 12404 77364 12460
rect 77420 12404 77430 12460
rect 77914 12404 77924 12460
rect 77980 12404 78708 12460
rect 78764 12404 78774 12460
rect 78922 12404 78932 12460
rect 78988 12404 80052 12460
rect 80108 12404 80118 12460
rect 80266 12404 80276 12460
rect 80332 12404 81340 12460
rect 81498 12404 81508 12460
rect 81564 12404 83300 12460
rect 83356 12404 83366 12460
rect 83626 12404 83636 12460
rect 83692 12404 97412 12460
rect 97468 12404 97478 12460
rect 97626 12404 97636 12460
rect 97692 12404 99876 12460
rect 99932 12404 99942 12460
rect 100426 12404 100436 12460
rect 100492 12404 101556 12460
rect 101612 12404 101622 12460
rect 102106 12404 102116 12460
rect 102172 12404 109620 12460
rect 109676 12404 109686 12460
rect 109834 12404 109844 12460
rect 109900 12404 114548 12460
rect 114604 12404 114614 12460
rect 114762 12404 114772 12460
rect 114828 12404 119028 12460
rect 119084 12404 119094 12460
rect 119354 12404 119364 12460
rect 119420 12404 121268 12460
rect 121324 12404 121334 12460
rect 122714 12404 122724 12460
rect 122780 12404 123004 12460
rect 125514 12404 125524 12460
rect 125580 12404 126532 12460
rect 126588 12404 126598 12460
rect 126756 12404 154084 12460
rect 154140 12404 154150 12460
rect 154298 12404 154308 12460
rect 154364 12404 155036 12460
rect 155754 12404 155764 12460
rect 155820 12404 156212 12460
rect 156268 12404 156278 12460
rect 156436 12404 156884 12460
rect 156940 12404 156950 12460
rect 0 12376 800 12404
rect 2426 12292 2436 12348
rect 2492 12292 9716 12348
rect 9772 12292 9782 12348
rect 47674 12292 47684 12348
rect 47740 12292 55412 12348
rect 55468 12292 55478 12348
rect 55598 12292 55636 12348
rect 55692 12292 55702 12348
rect 62916 12236 62972 12404
rect 122948 12348 123004 12404
rect 158452 12348 158508 12516
rect 158666 12404 158676 12460
rect 158732 12404 164052 12460
rect 164108 12404 164118 12460
rect 164266 12404 164276 12460
rect 164332 12404 166516 12460
rect 166572 12404 166582 12460
rect 169418 12404 169428 12460
rect 169484 12404 174244 12460
rect 174300 12404 174310 12460
rect 174458 12404 174468 12460
rect 174524 12404 193844 12460
rect 193900 12404 193910 12460
rect 194058 12404 194068 12460
rect 194124 12404 199332 12460
rect 199388 12404 199398 12460
rect 211754 12404 211764 12460
rect 211820 12404 213780 12460
rect 213836 12404 213846 12460
rect 65706 12292 65716 12348
rect 65772 12292 66724 12348
rect 66780 12292 66790 12348
rect 66938 12292 66948 12348
rect 67004 12292 70084 12348
rect 70140 12292 70150 12348
rect 70298 12292 70308 12348
rect 70364 12292 78260 12348
rect 78316 12292 78326 12348
rect 78474 12292 78484 12348
rect 78540 12292 78820 12348
rect 78876 12292 78886 12348
rect 79818 12292 79828 12348
rect 79884 12292 83188 12348
rect 83244 12292 83254 12348
rect 83402 12292 83412 12348
rect 83468 12292 83748 12348
rect 83804 12292 83814 12348
rect 83962 12292 83972 12348
rect 84028 12292 84644 12348
rect 84700 12292 84710 12348
rect 84858 12292 84868 12348
rect 84924 12292 89124 12348
rect 89180 12292 89190 12348
rect 89450 12292 89460 12348
rect 89516 12292 93492 12348
rect 93548 12292 93558 12348
rect 94154 12292 94164 12348
rect 94220 12292 103124 12348
rect 103180 12292 103190 12348
rect 103898 12292 103908 12348
rect 103964 12292 104132 12348
rect 104188 12292 104198 12348
rect 104458 12292 104468 12348
rect 104524 12292 113652 12348
rect 113708 12292 113718 12348
rect 114202 12292 114212 12348
rect 114268 12292 116788 12348
rect 116844 12292 116854 12348
rect 117002 12292 117012 12348
rect 117068 12292 117908 12348
rect 117964 12292 117974 12348
rect 118570 12292 118580 12348
rect 118636 12292 120820 12348
rect 120876 12292 120886 12348
rect 121034 12292 121044 12348
rect 121100 12292 122724 12348
rect 122780 12292 122790 12348
rect 122948 12292 130788 12348
rect 130844 12292 130854 12348
rect 131002 12292 131012 12348
rect 131068 12292 138292 12348
rect 138348 12292 138358 12348
rect 138516 12292 148708 12348
rect 148764 12292 148774 12348
rect 149482 12292 149492 12348
rect 149548 12292 158508 12348
rect 160542 12292 160580 12348
rect 160636 12292 160646 12348
rect 162698 12292 162708 12348
rect 162764 12292 167692 12348
rect 171182 12292 171220 12348
rect 171276 12292 171286 12348
rect 172190 12292 172228 12348
rect 172284 12292 172294 12348
rect 173450 12292 173460 12348
rect 173516 12292 180852 12348
rect 180908 12292 180918 12348
rect 181076 12292 187012 12348
rect 187068 12292 187078 12348
rect 187562 12292 187572 12348
rect 187628 12292 195860 12348
rect 195916 12292 195926 12348
rect 204362 12292 204372 12348
rect 204428 12292 207172 12348
rect 207228 12292 207238 12348
rect 210970 12292 210980 12348
rect 211036 12292 214452 12348
rect 214508 12292 214518 12348
rect 215674 12292 215684 12348
rect 215740 12292 218148 12348
rect 218204 12292 218214 12348
rect 138516 12236 138572 12292
rect 48570 12180 48580 12236
rect 48636 12180 56196 12236
rect 56252 12180 56262 12236
rect 56420 12180 61460 12236
rect 61516 12180 61526 12236
rect 62916 12180 67508 12236
rect 67564 12180 67574 12236
rect 67834 12180 67844 12236
rect 67900 12180 69860 12236
rect 69916 12180 69926 12236
rect 70084 12180 71988 12236
rect 72044 12180 72054 12236
rect 73546 12180 73556 12236
rect 73612 12180 79716 12236
rect 79772 12180 79782 12236
rect 79930 12180 79940 12236
rect 79996 12180 80388 12236
rect 80444 12180 80454 12236
rect 80612 12180 88788 12236
rect 88844 12180 88854 12236
rect 89002 12180 89012 12236
rect 89068 12180 90188 12236
rect 90346 12180 90356 12236
rect 90412 12180 97636 12236
rect 97692 12180 97702 12236
rect 98074 12180 98084 12236
rect 98140 12180 98644 12236
rect 98700 12180 98710 12236
rect 99082 12180 99092 12236
rect 99148 12180 102564 12236
rect 102620 12180 102630 12236
rect 103002 12180 103012 12236
rect 103068 12180 109396 12236
rect 109452 12180 109462 12236
rect 109610 12180 109620 12236
rect 109676 12180 112420 12236
rect 112476 12180 112486 12236
rect 114202 12180 114212 12236
rect 114268 12180 119140 12236
rect 119196 12180 119206 12236
rect 119354 12180 119364 12236
rect 119420 12180 120092 12236
rect 120250 12180 120260 12236
rect 120316 12180 120372 12236
rect 120428 12180 120438 12236
rect 120586 12180 120596 12236
rect 120652 12180 121940 12236
rect 121996 12180 122006 12236
rect 122154 12180 122164 12236
rect 122220 12180 125524 12236
rect 125580 12180 125590 12236
rect 125738 12180 125748 12236
rect 125804 12180 131460 12236
rect 131516 12180 131526 12236
rect 132458 12180 132468 12236
rect 132524 12180 138572 12236
rect 138628 12180 141204 12236
rect 141260 12180 141270 12236
rect 143210 12180 143220 12236
rect 143276 12180 155428 12236
rect 155484 12180 155494 12236
rect 156202 12180 156212 12236
rect 156268 12180 162932 12236
rect 162988 12180 162998 12236
rect 163156 12180 165060 12236
rect 165116 12180 165126 12236
rect 56420 12124 56476 12180
rect 70084 12124 70140 12180
rect 80612 12124 80668 12180
rect 90132 12124 90188 12180
rect 120036 12124 120092 12180
rect 138628 12124 138684 12180
rect 163156 12124 163212 12180
rect 167636 12124 167692 12292
rect 181076 12236 181132 12292
rect 171108 12180 178052 12236
rect 178108 12180 178118 12236
rect 178798 12180 178836 12236
rect 178892 12180 178902 12236
rect 179610 12180 179620 12236
rect 179676 12180 181132 12236
rect 181290 12180 181300 12236
rect 181356 12180 191940 12236
rect 191996 12180 196868 12236
rect 196924 12180 196934 12236
rect 201562 12180 201572 12236
rect 201628 12180 203028 12236
rect 203084 12180 205044 12236
rect 205100 12180 205110 12236
rect 212986 12180 212996 12236
rect 213052 12180 215908 12236
rect 215964 12180 215974 12236
rect 171108 12124 171164 12180
rect 44874 12068 44884 12124
rect 44940 12068 52724 12124
rect 52780 12068 52790 12124
rect 55402 12068 55412 12124
rect 55468 12068 56476 12124
rect 57082 12068 57092 12124
rect 57148 12068 63476 12124
rect 63532 12068 63542 12124
rect 63690 12068 63700 12124
rect 63756 12068 63794 12124
rect 65258 12068 65268 12124
rect 65324 12068 68852 12124
rect 68908 12068 68918 12124
rect 69066 12068 69076 12124
rect 69132 12068 70140 12124
rect 71754 12068 71764 12124
rect 71820 12068 73388 12124
rect 74078 12068 74116 12124
rect 74172 12068 74182 12124
rect 74330 12068 74340 12124
rect 74396 12068 80668 12124
rect 80826 12068 80836 12124
rect 80892 12068 81172 12124
rect 81228 12068 81238 12124
rect 81722 12068 81732 12124
rect 81788 12068 82852 12124
rect 82908 12068 82918 12124
rect 83066 12068 83076 12124
rect 83132 12068 89908 12124
rect 89964 12068 89974 12124
rect 90132 12068 98980 12124
rect 99036 12068 99046 12124
rect 99194 12068 99204 12124
rect 99260 12068 100324 12124
rect 100380 12068 100390 12124
rect 100538 12068 100548 12124
rect 100604 12068 103460 12124
rect 103516 12068 103526 12124
rect 104122 12068 104132 12124
rect 104188 12068 106148 12124
rect 106204 12068 106214 12124
rect 106362 12068 106372 12124
rect 106428 12068 114100 12124
rect 114156 12068 114166 12124
rect 114314 12068 114324 12124
rect 114380 12068 115500 12124
rect 115630 12068 115668 12124
rect 115724 12068 115734 12124
rect 115882 12068 115892 12124
rect 115948 12068 117180 12124
rect 117338 12068 117348 12124
rect 117404 12068 118244 12124
rect 118300 12068 118310 12124
rect 118458 12068 118468 12124
rect 118524 12068 119812 12124
rect 119868 12068 119878 12124
rect 120036 12068 134148 12124
rect 134204 12068 134214 12124
rect 134362 12068 134372 12124
rect 134428 12068 135212 12124
rect 135370 12068 135380 12124
rect 135436 12068 138684 12124
rect 139290 12068 139300 12124
rect 139356 12068 153300 12124
rect 153356 12068 153366 12124
rect 153514 12068 153524 12124
rect 153580 12068 162036 12124
rect 162092 12068 162102 12124
rect 162698 12068 162708 12124
rect 162764 12068 163212 12124
rect 163268 12068 164276 12124
rect 164332 12068 164342 12124
rect 164490 12068 164500 12124
rect 164556 12068 167188 12124
rect 167244 12068 167254 12124
rect 167636 12068 171164 12124
rect 175130 12068 175140 12124
rect 175196 12068 180068 12124
rect 180124 12068 180134 12124
rect 183866 12068 183876 12124
rect 183932 12068 187908 12124
rect 187964 12068 187974 12124
rect 191491 12068 194852 12124
rect 194908 12068 194918 12124
rect 197726 12068 197764 12124
rect 197820 12068 197830 12124
rect 200554 12068 200564 12124
rect 200620 12068 204260 12124
rect 204316 12068 204326 12124
rect 205930 12068 205940 12124
rect 205996 12068 212996 12124
rect 213052 12068 213062 12124
rect 213220 12068 215236 12124
rect 215292 12068 215302 12124
rect 216570 12068 216580 12124
rect 216636 12068 219604 12124
rect 219660 12068 219670 12124
rect 73332 12012 73388 12068
rect 115444 12012 115500 12068
rect 117124 12012 117180 12068
rect 135156 12012 135212 12068
rect 163268 12012 163324 12068
rect 191491 12012 191547 12068
rect 213220 12012 213276 12068
rect 48458 11956 48468 12012
rect 48524 11956 51268 12012
rect 51324 11956 51334 12012
rect 52490 11956 52500 12012
rect 52556 11956 53620 12012
rect 53676 11956 53686 12012
rect 54394 11956 54404 12012
rect 54460 11956 66612 12012
rect 66668 11956 66678 12012
rect 67386 11956 67396 12012
rect 67452 11956 73108 12012
rect 73164 11956 73174 12012
rect 73332 11956 74788 12012
rect 74844 11956 74854 12012
rect 75002 11956 75012 12012
rect 75068 11956 80276 12012
rect 80332 11956 80342 12012
rect 80490 11956 80500 12012
rect 80556 11956 82292 12012
rect 82348 11956 82358 12012
rect 82506 11956 82516 12012
rect 82572 11956 83020 12012
rect 83402 11956 83412 12012
rect 83468 11956 89012 12012
rect 89068 11956 89078 12012
rect 89226 11956 89236 12012
rect 89292 11956 97748 12012
rect 97804 11956 97814 12012
rect 98074 11956 98084 12012
rect 98140 11956 106596 12012
rect 106652 11956 106662 12012
rect 106820 11956 108724 12012
rect 108780 11956 108790 12012
rect 108938 11956 108948 12012
rect 109004 11956 109042 12012
rect 109274 11956 109284 12012
rect 109340 11956 115220 12012
rect 115276 11956 115286 12012
rect 115444 11956 116228 12012
rect 116284 11956 116294 12012
rect 117124 11956 118020 12012
rect 118076 11956 118086 12012
rect 118234 11956 118244 12012
rect 118300 11956 120148 12012
rect 120204 11956 120214 12012
rect 120362 11956 120372 12012
rect 120428 11956 134932 12012
rect 134988 11956 134998 12012
rect 135156 11956 137620 12012
rect 137676 11956 137686 12012
rect 138170 11956 138180 12012
rect 138236 11956 145236 12012
rect 145292 11956 145302 12012
rect 147466 11956 147476 12012
rect 147532 11956 149044 12012
rect 149100 11956 149110 12012
rect 149370 11956 149380 12012
rect 149436 11956 154532 12012
rect 154588 11956 154598 12012
rect 155082 11956 155092 12012
rect 155148 11956 162148 12012
rect 162204 11956 162214 12012
rect 162474 11956 162484 12012
rect 162540 11956 163324 12012
rect 163706 11956 163716 12012
rect 163772 11956 166292 12012
rect 166348 11956 166358 12012
rect 166506 11956 166516 12012
rect 166572 11956 170884 12012
rect 170940 11956 170950 12012
rect 171108 11956 172844 12012
rect 173002 11956 173012 12012
rect 173068 11956 176932 12012
rect 176988 11956 176998 12012
rect 178042 11956 178052 12012
rect 178108 11956 178612 12012
rect 178668 11956 191547 12012
rect 194618 11956 194628 12012
rect 194684 11956 199892 12012
rect 199948 11956 199958 12012
rect 202570 11956 202580 12012
rect 202636 11956 206500 12012
rect 206556 11956 206566 12012
rect 206724 11956 213276 12012
rect 213770 11956 213780 12012
rect 213836 11956 216692 12012
rect 216748 11956 216758 12012
rect 82964 11900 83020 11956
rect 106820 11900 106876 11956
rect 171108 11900 171164 11956
rect 22250 11844 22260 11900
rect 22316 11844 24276 11900
rect 24332 11844 24342 11900
rect 46890 11844 46900 11900
rect 46956 11844 48356 11900
rect 48412 11844 48422 11900
rect 50250 11844 50260 11900
rect 50316 11844 60452 11900
rect 60508 11844 60518 11900
rect 63354 11844 63364 11900
rect 63420 11844 70980 11900
rect 71036 11844 71046 11900
rect 71194 11844 71204 11900
rect 71260 11844 74564 11900
rect 74620 11844 74630 11900
rect 75114 11844 75124 11900
rect 75180 11844 78708 11900
rect 78764 11844 78774 11900
rect 79034 11844 79044 11900
rect 79100 11844 81508 11900
rect 81564 11844 81574 11900
rect 82058 11844 82068 11900
rect 82124 11844 82740 11900
rect 82796 11844 82806 11900
rect 82964 11844 84252 11900
rect 84522 11844 84532 11900
rect 84588 11844 93828 11900
rect 93884 11844 93894 11900
rect 95274 11844 95284 11900
rect 95340 11844 98588 11900
rect 98858 11844 98868 11900
rect 98924 11844 104020 11900
rect 104076 11844 104086 11900
rect 104234 11844 104244 11900
rect 104300 11844 106876 11900
rect 107482 11844 107492 11900
rect 107548 11844 115892 11900
rect 115948 11844 115958 11900
rect 116330 11844 116340 11900
rect 116396 11844 118468 11900
rect 118524 11844 118534 11900
rect 119242 11844 119252 11900
rect 119308 11844 121380 11900
rect 121436 11844 121446 11900
rect 126298 11844 126308 11900
rect 126364 11844 127092 11900
rect 127148 11844 127158 11900
rect 127978 11844 127988 11900
rect 128044 11844 128548 11900
rect 128604 11844 128614 11900
rect 130788 11844 131236 11900
rect 131292 11844 131302 11900
rect 131450 11844 131460 11900
rect 131516 11844 134260 11900
rect 134316 11844 134326 11900
rect 135482 11844 135492 11900
rect 135548 11844 137956 11900
rect 138012 11844 138022 11900
rect 139738 11844 139748 11900
rect 139804 11844 141316 11900
rect 141372 11844 141382 11900
rect 141530 11844 141540 11900
rect 141596 11844 143052 11900
rect 143322 11844 143332 11900
rect 143388 11844 144452 11900
rect 144508 11844 144518 11900
rect 146122 11844 146132 11900
rect 146188 11844 147812 11900
rect 147868 11844 147878 11900
rect 148026 11844 148036 11900
rect 148092 11844 148932 11900
rect 148988 11844 148998 11900
rect 149146 11844 149156 11900
rect 149212 11844 151172 11900
rect 151228 11844 151238 11900
rect 151498 11844 151508 11900
rect 151564 11844 153524 11900
rect 153580 11844 153590 11900
rect 154532 11844 159012 11900
rect 159068 11844 159078 11900
rect 159236 11844 162820 11900
rect 162876 11844 162886 11900
rect 165610 11844 165620 11900
rect 165676 11844 168644 11900
rect 168700 11844 168710 11900
rect 168858 11844 168868 11900
rect 168924 11844 171164 11900
rect 172526 11844 172564 11900
rect 172620 11844 172630 11900
rect 84196 11788 84252 11844
rect 98532 11788 98588 11844
rect 130788 11788 130844 11844
rect 142996 11788 143052 11844
rect 18106 11732 18116 11788
rect 18172 11732 19908 11788
rect 19964 11732 19974 11788
rect 20234 11732 20244 11788
rect 20300 11732 22148 11788
rect 22204 11732 22214 11788
rect 26954 11732 26964 11788
rect 27020 11732 28644 11788
rect 28700 11732 28710 11788
rect 29866 11732 29876 11788
rect 29932 11732 30884 11788
rect 30940 11732 30950 11788
rect 34346 11732 34356 11788
rect 34412 11732 35252 11788
rect 35308 11732 35318 11788
rect 36698 11732 36708 11788
rect 36764 11732 37380 11788
rect 37436 11732 37446 11788
rect 42970 11732 42980 11788
rect 43036 11732 43988 11788
rect 44044 11732 44054 11788
rect 44650 11732 44660 11788
rect 44716 11732 46116 11788
rect 46172 11732 46182 11788
rect 47786 11732 47796 11788
rect 47852 11732 49028 11788
rect 49084 11732 49094 11788
rect 49802 11732 49812 11788
rect 49868 11732 50372 11788
rect 50428 11732 50438 11788
rect 52052 11732 57092 11788
rect 57148 11732 57158 11788
rect 57754 11732 57764 11788
rect 57820 11732 57876 11788
rect 57932 11732 57942 11788
rect 58090 11732 58100 11788
rect 58156 11732 62132 11788
rect 62188 11732 62198 11788
rect 62346 11732 62356 11788
rect 62412 11732 64372 11788
rect 64428 11732 64438 11788
rect 65370 11732 65380 11788
rect 65436 11732 67172 11788
rect 67228 11732 67238 11788
rect 67498 11732 67508 11788
rect 67564 11732 74116 11788
rect 74172 11732 74182 11788
rect 74442 11732 74452 11788
rect 74508 11732 76580 11788
rect 76636 11732 76646 11788
rect 76804 11732 77700 11788
rect 77756 11732 77766 11788
rect 77914 11732 77924 11788
rect 77980 11732 83972 11788
rect 84028 11732 84038 11788
rect 84196 11732 96068 11788
rect 96124 11732 96134 11788
rect 97066 11732 97076 11788
rect 97132 11732 98308 11788
rect 98364 11732 98374 11788
rect 98532 11732 100212 11788
rect 100268 11732 100278 11788
rect 100426 11732 100436 11788
rect 100492 11732 101892 11788
rect 101948 11732 101958 11788
rect 102116 11732 105924 11788
rect 105980 11732 105990 11788
rect 106138 11732 106148 11788
rect 106204 11732 113092 11788
rect 113148 11732 113158 11788
rect 113306 11732 113316 11788
rect 113372 11732 113820 11788
rect 114986 11732 114996 11788
rect 115052 11732 117124 11788
rect 117180 11732 117190 11788
rect 117348 11732 118804 11788
rect 118860 11732 118870 11788
rect 119018 11732 119028 11788
rect 119084 11732 119364 11788
rect 119420 11732 119430 11788
rect 120362 11732 120372 11788
rect 120428 11732 120932 11788
rect 120988 11732 120998 11788
rect 121370 11732 121380 11788
rect 121436 11732 122276 11788
rect 122332 11732 122342 11788
rect 122490 11732 122500 11788
rect 122556 11732 130844 11788
rect 130900 11732 132692 11788
rect 132748 11732 132758 11788
rect 132906 11732 132916 11788
rect 132972 11732 137732 11788
rect 137788 11732 137798 11788
rect 138842 11732 138852 11788
rect 138908 11732 142772 11788
rect 142828 11732 142838 11788
rect 142996 11732 144564 11788
rect 144620 11732 144630 11788
rect 147690 11732 147700 11788
rect 147756 11732 151340 11788
rect 52052 11676 52108 11732
rect 76804 11676 76860 11732
rect 102116 11676 102172 11732
rect 113764 11676 113820 11732
rect 117348 11676 117404 11732
rect 130900 11676 130956 11732
rect 151284 11676 151340 11732
rect 154532 11676 154588 11844
rect 159236 11788 159292 11844
rect 172788 11788 172844 11956
rect 206724 11900 206780 11956
rect 173786 11844 173796 11900
rect 173852 11844 186452 11900
rect 186508 11844 186518 11900
rect 187002 11844 187012 11900
rect 187068 11844 189700 11900
rect 189756 11844 196196 11900
rect 196252 11844 196262 11900
rect 198398 11844 198436 11900
rect 198492 11844 198502 11900
rect 199658 11844 199668 11900
rect 199724 11844 202132 11900
rect 202188 11844 202198 11900
rect 203466 11844 203476 11900
rect 203532 11844 205716 11900
rect 205772 11844 205782 11900
rect 205940 11844 206780 11900
rect 206938 11844 206948 11900
rect 207004 11844 207732 11900
rect 207788 11844 209412 11900
rect 209468 11844 209478 11900
rect 213098 11844 213108 11900
rect 213164 11844 217364 11900
rect 217420 11844 217430 11900
rect 205940 11788 205996 11844
rect 154830 11732 154868 11788
rect 154924 11732 154934 11788
rect 155082 11732 155092 11788
rect 155148 11732 159292 11788
rect 159450 11732 159460 11788
rect 159516 11732 162988 11788
rect 165722 11732 165732 11788
rect 165788 11732 166404 11788
rect 166460 11732 166470 11788
rect 170762 11732 170772 11788
rect 170828 11732 172452 11788
rect 172508 11732 172518 11788
rect 172788 11732 174468 11788
rect 174524 11732 174534 11788
rect 177370 11732 177380 11788
rect 177436 11732 183988 11788
rect 184044 11732 184054 11788
rect 186106 11732 186116 11788
rect 186172 11732 190372 11788
rect 190428 11732 190438 11788
rect 192602 11732 192612 11788
rect 192668 11732 193732 11788
rect 193788 11732 193798 11788
rect 195962 11732 195972 11788
rect 196028 11732 196980 11788
rect 197036 11732 197046 11788
rect 198090 11732 198100 11788
rect 198156 11732 199220 11788
rect 199276 11732 199286 11788
rect 199434 11732 199444 11788
rect 199500 11732 201348 11788
rect 201404 11732 201414 11788
rect 202010 11732 202020 11788
rect 202076 11732 203588 11788
rect 203644 11732 203654 11788
rect 204586 11732 204596 11788
rect 204652 11732 205996 11788
rect 206154 11732 206164 11788
rect 206220 11732 207956 11788
rect 208012 11732 208022 11788
rect 208842 11732 208852 11788
rect 208908 11732 210868 11788
rect 210924 11732 210934 11788
rect 211530 11732 211540 11788
rect 211596 11732 212884 11788
rect 212940 11732 212950 11788
rect 215002 11732 215012 11788
rect 215068 11732 218820 11788
rect 218876 11732 218886 11788
rect 162932 11676 162988 11732
rect 51146 11620 51156 11676
rect 51212 11620 52108 11676
rect 55738 11620 55748 11676
rect 55804 11620 66612 11676
rect 66668 11620 66678 11676
rect 66826 11620 66836 11676
rect 66892 11620 67396 11676
rect 67452 11620 67462 11676
rect 68170 11620 68180 11676
rect 68236 11620 69524 11676
rect 69580 11620 69590 11676
rect 69738 11620 69748 11676
rect 69804 11620 76860 11676
rect 77242 11620 77252 11676
rect 77308 11620 78596 11676
rect 78652 11620 78662 11676
rect 78810 11620 78820 11676
rect 78876 11620 99316 11676
rect 99372 11620 99382 11676
rect 99530 11620 99540 11676
rect 99596 11620 102172 11676
rect 102330 11620 102340 11676
rect 102396 11620 103012 11676
rect 103068 11620 103078 11676
rect 103236 11620 112756 11676
rect 112812 11620 112822 11676
rect 113764 11620 114212 11676
rect 114314 11620 114324 11676
rect 114380 11620 116004 11676
rect 116060 11620 116070 11676
rect 116218 11620 116228 11676
rect 116284 11620 116564 11676
rect 116620 11620 116630 11676
rect 116778 11620 116788 11676
rect 116844 11620 117404 11676
rect 117460 11620 119924 11676
rect 119980 11620 119990 11676
rect 120138 11620 120148 11676
rect 120204 11620 126812 11676
rect 129546 11620 129556 11676
rect 129612 11620 130956 11676
rect 132682 11620 132692 11676
rect 132748 11620 133588 11676
rect 133644 11620 133654 11676
rect 134250 11620 134260 11676
rect 134316 11620 137732 11676
rect 137788 11620 137798 11676
rect 138282 11620 138292 11676
rect 138348 11620 139524 11676
rect 139580 11620 139590 11676
rect 141082 11620 141092 11676
rect 141148 11620 151060 11676
rect 151116 11620 151126 11676
rect 151284 11620 154588 11676
rect 154746 11620 154756 11676
rect 154812 11620 156212 11676
rect 156268 11620 156278 11676
rect 156426 11620 156436 11676
rect 156492 11620 157108 11676
rect 157164 11620 158564 11676
rect 158620 11620 158630 11676
rect 158778 11620 158788 11676
rect 158844 11620 162260 11676
rect 162316 11620 162326 11676
rect 162932 11620 171108 11676
rect 171164 11620 171174 11676
rect 182970 11620 182980 11676
rect 183036 11620 187684 11676
rect 187740 11620 187750 11676
rect 188010 11620 188020 11676
rect 188076 11620 201572 11676
rect 201628 11620 201638 11676
rect 103236 11564 103292 11620
rect 51706 11508 51716 11564
rect 51772 11508 56196 11564
rect 56252 11508 56262 11564
rect 57082 11508 57092 11564
rect 57148 11508 62356 11564
rect 62412 11508 62422 11564
rect 63914 11508 63924 11564
rect 63980 11508 86996 11564
rect 87052 11508 87062 11564
rect 87210 11508 87220 11564
rect 87276 11508 103292 11564
rect 103450 11508 103460 11564
rect 103516 11508 107940 11564
rect 107996 11508 108006 11564
rect 109050 11508 109060 11564
rect 109116 11508 109508 11564
rect 109564 11508 109574 11564
rect 110926 11508 110964 11564
rect 111020 11508 111030 11564
rect 111850 11508 111860 11564
rect 111916 11508 112532 11564
rect 112588 11508 112598 11564
rect 112746 11508 112756 11564
rect 112812 11508 113988 11564
rect 114044 11508 114054 11564
rect 114156 11452 114212 11620
rect 117460 11564 117516 11620
rect 126756 11564 126812 11620
rect 114314 11508 114324 11564
rect 114380 11508 115612 11564
rect 115770 11508 115780 11564
rect 115836 11508 116340 11564
rect 116396 11508 116406 11564
rect 116554 11508 116564 11564
rect 116620 11508 117516 11564
rect 117674 11508 117684 11564
rect 117740 11508 126532 11564
rect 126588 11508 126598 11564
rect 126756 11508 140756 11564
rect 140812 11508 140822 11564
rect 140980 11508 151732 11564
rect 151788 11508 151798 11564
rect 152730 11508 152740 11564
rect 152796 11508 159236 11564
rect 159292 11508 159302 11564
rect 160906 11508 160916 11564
rect 160972 11508 165284 11564
rect 165340 11508 165350 11564
rect 168522 11508 168532 11564
rect 168588 11508 170212 11564
rect 170268 11508 170278 11564
rect 170986 11508 170996 11564
rect 171052 11508 180404 11564
rect 180460 11508 191716 11564
rect 191772 11508 191782 11564
rect 115556 11452 115612 11508
rect 140980 11452 141036 11508
rect 45434 11396 45444 11452
rect 45500 11396 63924 11452
rect 63980 11396 63990 11452
rect 64148 11396 66836 11452
rect 66892 11396 66902 11452
rect 67162 11396 67172 11452
rect 67228 11396 82068 11452
rect 82124 11396 82134 11452
rect 82291 11396 82964 11452
rect 83020 11396 83030 11452
rect 83178 11396 83188 11452
rect 83244 11396 83300 11452
rect 83356 11396 83366 11452
rect 83514 11396 83524 11452
rect 83580 11396 83860 11452
rect 83916 11396 83926 11452
rect 84074 11396 84084 11452
rect 84140 11396 88564 11452
rect 88620 11396 88630 11452
rect 88778 11396 88788 11452
rect 88844 11396 88882 11452
rect 89011 11396 92036 11452
rect 92092 11396 92102 11452
rect 92698 11396 92708 11452
rect 92764 11396 96852 11452
rect 96908 11396 96918 11452
rect 97290 11396 97300 11452
rect 97356 11396 99092 11452
rect 99148 11396 99158 11452
rect 99306 11396 99316 11452
rect 99372 11396 113540 11452
rect 113596 11396 113606 11452
rect 114156 11396 115332 11452
rect 115388 11396 115398 11452
rect 115556 11396 118580 11452
rect 118636 11396 118646 11452
rect 119130 11396 119140 11452
rect 119196 11396 132468 11452
rect 132524 11396 132534 11452
rect 132691 11396 135940 11452
rect 135996 11396 136006 11452
rect 138618 11396 138628 11452
rect 138684 11396 141036 11452
rect 141306 11396 141316 11452
rect 141372 11396 143332 11452
rect 143388 11396 143398 11452
rect 146010 11396 146020 11452
rect 146076 11396 164612 11452
rect 164668 11396 164678 11452
rect 164826 11396 164836 11452
rect 164892 11396 183428 11452
rect 183484 11396 183494 11452
rect 183652 11396 189812 11452
rect 189868 11396 189878 11452
rect 64148 11340 64204 11396
rect 42634 11284 42644 11340
rect 42700 11284 51716 11340
rect 51772 11284 51782 11340
rect 51930 11284 51940 11340
rect 51996 11284 55300 11340
rect 55356 11284 55366 11340
rect 56186 11284 56196 11340
rect 56252 11284 58100 11340
rect 58156 11284 58166 11340
rect 58314 11284 58324 11340
rect 58380 11284 64204 11340
rect 65034 11284 65044 11340
rect 65100 11284 69188 11340
rect 69244 11284 69254 11340
rect 69402 11284 69412 11340
rect 69468 11284 79380 11340
rect 79436 11284 79446 11340
rect 79594 11284 79604 11340
rect 79660 11284 79828 11340
rect 79884 11284 79894 11340
rect 80378 11284 80388 11340
rect 80444 11284 81956 11340
rect 82012 11284 82022 11340
rect 82291 11228 82347 11396
rect 89011 11340 89067 11396
rect 132691 11340 132747 11396
rect 183652 11340 183708 11396
rect 82506 11284 82516 11340
rect 82572 11284 84196 11340
rect 84252 11284 84262 11340
rect 84410 11284 84420 11340
rect 84476 11284 89067 11340
rect 89338 11284 89348 11340
rect 89404 11284 91140 11340
rect 91196 11284 91206 11340
rect 91466 11284 91476 11340
rect 91532 11284 102676 11340
rect 102732 11284 102742 11340
rect 102890 11284 102900 11340
rect 102956 11284 103572 11340
rect 103628 11284 103638 11340
rect 103796 11284 104804 11340
rect 104860 11284 104870 11340
rect 105018 11284 105028 11340
rect 105084 11284 106484 11340
rect 106540 11284 106550 11340
rect 109498 11284 109508 11340
rect 109564 11284 110852 11340
rect 110908 11284 110918 11340
rect 111066 11284 111076 11340
rect 111132 11284 113036 11340
rect 113418 11284 113428 11340
rect 113484 11284 116004 11340
rect 116060 11284 116070 11340
rect 116218 11284 116228 11340
rect 116284 11284 117684 11340
rect 117740 11284 117750 11340
rect 118794 11284 118804 11340
rect 118860 11284 119252 11340
rect 119308 11284 119318 11340
rect 119466 11284 119476 11340
rect 119532 11284 126308 11340
rect 126364 11284 126374 11340
rect 126522 11284 126532 11340
rect 126588 11284 132747 11340
rect 133018 11284 133028 11340
rect 133084 11284 135940 11340
rect 135996 11284 136006 11340
rect 136714 11284 136724 11340
rect 136780 11284 144228 11340
rect 144284 11284 144294 11340
rect 146122 11284 146132 11340
rect 146188 11284 150052 11340
rect 150108 11284 150118 11340
rect 150378 11284 150388 11340
rect 150444 11284 159460 11340
rect 159516 11284 159526 11340
rect 162138 11284 162148 11340
rect 162204 11284 163828 11340
rect 163884 11284 166740 11340
rect 166796 11284 166806 11340
rect 167971 11284 183708 11340
rect 183866 11284 183876 11340
rect 183932 11284 194068 11340
rect 194124 11284 194134 11340
rect 103796 11228 103852 11284
rect 112980 11228 113036 11284
rect 167971 11228 168027 11284
rect 219200 11228 220000 11256
rect 48010 11172 48020 11228
rect 48076 11172 66276 11228
rect 66332 11172 66342 11228
rect 66490 11172 66500 11228
rect 66556 11172 68180 11228
rect 68236 11172 68246 11228
rect 68506 11172 68516 11228
rect 68572 11172 72660 11228
rect 72716 11172 72726 11228
rect 73434 11172 73444 11228
rect 73500 11172 73668 11228
rect 73724 11172 73734 11228
rect 73882 11172 73892 11228
rect 73948 11172 82347 11228
rect 82404 11172 82964 11228
rect 83020 11172 83030 11228
rect 83738 11172 83748 11228
rect 83804 11172 100212 11228
rect 100268 11172 100278 11228
rect 100426 11172 100436 11228
rect 100492 11172 100828 11228
rect 82404 11116 82460 11172
rect 100772 11116 100828 11172
rect 102452 11172 103852 11228
rect 104122 11172 104132 11228
rect 104188 11172 112756 11228
rect 112812 11172 112822 11228
rect 112980 11172 114436 11228
rect 114492 11172 114502 11228
rect 114762 11172 114772 11228
rect 114828 11172 129108 11228
rect 129164 11172 129174 11228
rect 129434 11172 129444 11228
rect 129500 11172 133868 11228
rect 134250 11172 134260 11228
rect 134316 11172 144340 11228
rect 144396 11172 144406 11228
rect 146234 11172 146244 11228
rect 146300 11172 152908 11228
rect 154522 11172 154532 11228
rect 154588 11172 158788 11228
rect 158844 11172 158854 11228
rect 159002 11172 159012 11228
rect 159068 11172 168027 11228
rect 175914 11172 175924 11228
rect 175980 11172 182868 11228
rect 182924 11172 182934 11228
rect 186330 11172 186340 11228
rect 186396 11172 197316 11228
rect 197372 11172 197382 11228
rect 219044 11172 220000 11228
rect 102452 11116 102508 11172
rect 133812 11116 133868 11172
rect 152852 11116 152908 11172
rect 14410 11060 14420 11116
rect 14476 11060 77924 11116
rect 77980 11060 77990 11116
rect 78138 11060 78148 11116
rect 78204 11004 78260 11116
rect 78362 11060 78372 11116
rect 78428 11060 78820 11116
rect 78876 11060 78886 11116
rect 79034 11060 79044 11116
rect 79100 11060 82460 11116
rect 82516 11060 92820 11116
rect 92876 11060 92886 11116
rect 93034 11060 93044 11116
rect 93100 11060 96852 11116
rect 96908 11060 96918 11116
rect 98186 11060 98196 11116
rect 98252 11060 100548 11116
rect 100604 11060 100614 11116
rect 100772 11060 102508 11116
rect 102666 11060 102676 11116
rect 102732 11060 112308 11116
rect 112364 11060 112374 11116
rect 113306 11060 113316 11116
rect 113372 11060 124180 11116
rect 124236 11060 124246 11116
rect 131002 11060 131012 11116
rect 131068 11060 131404 11116
rect 133550 11060 133588 11116
rect 133644 11060 133654 11116
rect 133812 11060 135044 11116
rect 135100 11060 135110 11116
rect 135258 11060 135268 11116
rect 135324 11060 135772 11116
rect 138282 11060 138292 11116
rect 138348 11060 143668 11116
rect 143724 11060 147924 11116
rect 147980 11060 147990 11116
rect 148698 11060 148708 11116
rect 148764 11060 151172 11116
rect 151228 11060 151238 11116
rect 152852 11060 154980 11116
rect 155036 11060 155046 11116
rect 156090 11060 156100 11116
rect 156156 11060 159236 11116
rect 159292 11060 159302 11116
rect 160906 11060 160916 11116
rect 160972 11060 161252 11116
rect 161308 11060 161318 11116
rect 162922 11060 162932 11116
rect 162988 11060 164892 11116
rect 166730 11060 166740 11116
rect 166796 11060 172788 11116
rect 172844 11060 179620 11116
rect 179676 11060 179686 11116
rect 179844 11060 187460 11116
rect 187516 11060 187526 11116
rect 187674 11060 187684 11116
rect 187740 11060 198324 11116
rect 198380 11060 198390 11116
rect 82516 11004 82572 11060
rect 10826 10948 10836 11004
rect 10892 10948 78036 11004
rect 78092 10948 78102 11004
rect 78204 10948 81900 11004
rect 82058 10948 82068 11004
rect 82124 10948 82572 11004
rect 83178 10948 83188 11004
rect 83244 10948 96740 11004
rect 96796 10948 96806 11004
rect 96964 10948 98420 11004
rect 98476 10948 98486 11004
rect 99194 10948 99204 11004
rect 99260 10948 103012 11004
rect 103068 10948 103078 11004
rect 103226 10948 103236 11004
rect 103292 10948 104468 11004
rect 104524 10948 104534 11004
rect 105578 10948 105588 11004
rect 105644 10948 113428 11004
rect 113484 10948 113494 11004
rect 113642 10948 113652 11004
rect 113708 10948 117348 11004
rect 117404 10948 117414 11004
rect 117562 10948 117572 11004
rect 117628 10948 120932 11004
rect 120988 10948 120998 11004
rect 121146 10948 121156 11004
rect 121212 10948 131124 11004
rect 131180 10948 131190 11004
rect 81844 10892 81900 10948
rect 96964 10892 97020 10948
rect 131348 10892 131404 11060
rect 135716 11004 135772 11060
rect 132122 10948 132132 11004
rect 132188 10948 135492 11004
rect 135548 10948 135558 11004
rect 135716 10948 139916 11004
rect 141082 10948 141092 11004
rect 141148 10948 147700 11004
rect 147756 10948 147766 11004
rect 150266 10948 150276 11004
rect 150332 10948 164612 11004
rect 164668 10948 164678 11004
rect 139860 10892 139916 10948
rect 164836 10892 164892 11060
rect 179844 11004 179900 11060
rect 166618 10948 166628 11004
rect 166684 10948 179900 11004
rect 180740 10948 187796 11004
rect 187852 10948 187862 11004
rect 189802 10948 189812 11004
rect 189868 10948 202356 11004
rect 202412 10948 202422 11004
rect 180740 10892 180796 10948
rect 219044 10892 219100 11172
rect 219200 11144 220000 11172
rect 13066 10836 13076 10892
rect 13132 10836 81620 10892
rect 81676 10836 81686 10892
rect 81844 10836 84924 10892
rect 85082 10836 85092 10892
rect 85148 10836 85988 10892
rect 86044 10836 86054 10892
rect 86174 10836 86212 10892
rect 86268 10836 86278 10892
rect 86426 10836 86436 10892
rect 86492 10836 91364 10892
rect 91420 10836 91430 10892
rect 92138 10836 92148 10892
rect 92204 10836 97020 10892
rect 98522 10836 98532 10892
rect 98588 10836 100548 10892
rect 100604 10836 100614 10892
rect 100762 10836 100772 10892
rect 100828 10836 102060 10892
rect 102218 10836 102228 10892
rect 102284 10836 107716 10892
rect 107772 10836 107782 10892
rect 107930 10836 107940 10892
rect 107996 10836 120708 10892
rect 120764 10836 120774 10892
rect 121034 10836 121044 10892
rect 121100 10836 124292 10892
rect 124348 10836 124358 10892
rect 124506 10836 124516 10892
rect 124572 10836 131292 10892
rect 131348 10836 133028 10892
rect 133084 10836 133094 10892
rect 133690 10836 133700 10892
rect 133756 10836 135380 10892
rect 135436 10836 135446 10892
rect 135594 10836 135604 10892
rect 135660 10836 139636 10892
rect 139692 10836 139702 10892
rect 139860 10836 141428 10892
rect 141484 10836 141494 10892
rect 142314 10836 142324 10892
rect 142380 10836 146916 10892
rect 146972 10836 146982 10892
rect 148922 10836 148932 10892
rect 148988 10836 151284 10892
rect 151340 10836 151350 10892
rect 152058 10836 152068 10892
rect 152124 10836 154644 10892
rect 154700 10836 154710 10892
rect 154970 10836 154980 10892
rect 155036 10836 158788 10892
rect 158844 10836 158854 10892
rect 159002 10836 159012 10892
rect 159068 10836 163380 10892
rect 163436 10836 163446 10892
rect 164836 10836 180796 10892
rect 180954 10836 180964 10892
rect 181020 10836 184324 10892
rect 184380 10836 184390 10892
rect 184538 10836 184548 10892
rect 184604 10836 188412 10892
rect 188570 10836 188580 10892
rect 188636 10836 202132 10892
rect 202188 10836 202198 10892
rect 219044 10836 219324 10892
rect 84868 10780 84924 10836
rect 102004 10780 102060 10836
rect 131236 10780 131292 10836
rect 188356 10780 188412 10836
rect 57642 10724 57652 10780
rect 57708 10724 77252 10780
rect 77308 10724 77318 10780
rect 77690 10724 77700 10780
rect 77756 10724 81508 10780
rect 81564 10724 81574 10780
rect 81722 10724 81732 10780
rect 81788 10724 84644 10780
rect 84700 10724 84710 10780
rect 84868 10724 86324 10780
rect 86380 10724 86390 10780
rect 86538 10724 86548 10780
rect 86604 10724 91812 10780
rect 91868 10724 91878 10780
rect 92026 10724 92036 10780
rect 92092 10724 96628 10780
rect 96684 10724 96694 10780
rect 96842 10724 96852 10780
rect 96908 10724 100044 10780
rect 100202 10724 100212 10780
rect 100268 10724 101220 10780
rect 101276 10724 101286 10780
rect 101434 10724 101444 10780
rect 101500 10724 101780 10780
rect 101836 10724 101846 10780
rect 102004 10724 103684 10780
rect 103740 10724 103750 10780
rect 104682 10724 104692 10780
rect 104748 10724 108836 10780
rect 108892 10724 108902 10780
rect 109060 10724 117124 10780
rect 117180 10724 117190 10780
rect 117338 10724 117348 10780
rect 117404 10724 126308 10780
rect 126364 10724 126374 10780
rect 131236 10724 131348 10780
rect 131404 10724 131414 10780
rect 131562 10724 131572 10780
rect 131628 10724 135828 10780
rect 135884 10724 135894 10780
rect 137722 10724 137732 10780
rect 137788 10724 146804 10780
rect 146860 10724 146870 10780
rect 147690 10724 147700 10780
rect 147756 10724 149716 10780
rect 149772 10724 149782 10780
rect 150276 10724 151508 10780
rect 151564 10724 151574 10780
rect 151722 10724 151732 10780
rect 151788 10724 183876 10780
rect 183932 10724 183942 10780
rect 185882 10724 185892 10780
rect 185948 10724 188300 10780
rect 188356 10724 198212 10780
rect 198268 10724 198278 10780
rect 99988 10668 100044 10724
rect 109060 10668 109116 10724
rect 150276 10668 150332 10724
rect 188244 10668 188300 10724
rect 14858 10612 14868 10668
rect 14924 10612 59556 10668
rect 59612 10612 59622 10668
rect 60778 10612 60788 10668
rect 60844 10612 67060 10668
rect 67116 10612 67126 10668
rect 67274 10612 67284 10668
rect 67340 10612 68404 10668
rect 68460 10612 68470 10668
rect 68730 10612 68740 10668
rect 68796 10612 70756 10668
rect 70812 10612 70822 10668
rect 70970 10612 70980 10668
rect 71036 10612 91140 10668
rect 91196 10612 91206 10668
rect 91354 10612 91364 10668
rect 91420 10612 99652 10668
rect 99708 10612 99718 10668
rect 99988 10612 100436 10668
rect 100492 10612 100502 10668
rect 100650 10612 100660 10668
rect 100716 10612 106204 10668
rect 108378 10612 108388 10668
rect 108444 10612 109116 10668
rect 109386 10612 109396 10668
rect 109452 10612 117684 10668
rect 117740 10612 117750 10668
rect 118010 10612 118020 10668
rect 118076 10612 120260 10668
rect 120316 10612 120326 10668
rect 120922 10612 120932 10668
rect 120988 10612 130452 10668
rect 130508 10612 130518 10668
rect 130862 10612 130900 10668
rect 130956 10612 130966 10668
rect 131674 10612 131684 10668
rect 131740 10612 139412 10668
rect 139468 10612 139478 10668
rect 139626 10612 139636 10668
rect 139692 10612 150332 10668
rect 151050 10612 151060 10668
rect 151116 10612 159012 10668
rect 159068 10612 159078 10668
rect 159226 10612 159236 10668
rect 159292 10612 178052 10668
rect 178108 10612 178118 10668
rect 178266 10612 178276 10668
rect 178332 10612 179396 10668
rect 179452 10612 188020 10668
rect 188076 10612 188086 10668
rect 188244 10612 200676 10668
rect 200732 10612 200742 10668
rect 53274 10500 53284 10556
rect 53340 10500 105924 10556
rect 105980 10500 105990 10556
rect 106148 10444 106204 10612
rect 106698 10500 106708 10556
rect 106764 10500 130004 10556
rect 130060 10500 130070 10556
rect 133886 10500 133924 10556
rect 133980 10500 133990 10556
rect 134138 10500 134148 10556
rect 134204 10500 146020 10556
rect 146076 10500 146086 10556
rect 147802 10500 147812 10556
rect 147868 10500 162148 10556
rect 162204 10500 162214 10556
rect 162362 10500 162372 10556
rect 162428 10500 164948 10556
rect 165004 10500 165014 10556
rect 165274 10500 165284 10556
rect 165340 10500 167636 10556
rect 167692 10500 167702 10556
rect 171658 10500 171668 10556
rect 171724 10500 191156 10556
rect 191212 10500 191222 10556
rect 25722 10388 25732 10444
rect 25788 10388 51828 10444
rect 51884 10388 51894 10444
rect 56298 10388 56308 10444
rect 56364 10388 56980 10444
rect 57036 10388 57046 10444
rect 62122 10388 62132 10444
rect 62188 10388 67620 10444
rect 67676 10388 67686 10444
rect 67834 10388 67844 10444
rect 67900 10388 68628 10444
rect 68684 10388 68694 10444
rect 68954 10388 68964 10444
rect 69020 10388 103124 10444
rect 103180 10388 103190 10444
rect 103348 10388 105812 10444
rect 105868 10388 105878 10444
rect 106148 10388 111244 10444
rect 111626 10388 111636 10444
rect 111692 10388 116228 10444
rect 116284 10388 116294 10444
rect 116666 10388 116676 10444
rect 116732 10388 117348 10444
rect 117404 10388 117414 10444
rect 117562 10388 117572 10444
rect 117628 10388 117684 10444
rect 117740 10388 117750 10444
rect 118234 10388 118244 10444
rect 118300 10388 126532 10444
rect 126588 10388 126598 10444
rect 129210 10388 129220 10444
rect 129276 10388 129556 10444
rect 129612 10388 129622 10444
rect 129770 10388 129780 10444
rect 129836 10388 133140 10444
rect 133196 10388 133206 10444
rect 133578 10388 133588 10444
rect 133644 10388 134036 10444
rect 134092 10388 134102 10444
rect 134222 10388 134260 10444
rect 134316 10388 134326 10444
rect 134474 10388 134484 10444
rect 134540 10388 139748 10444
rect 139804 10388 139814 10444
rect 140970 10388 140980 10444
rect 141036 10388 145796 10444
rect 145852 10388 145862 10444
rect 146570 10388 146580 10444
rect 146636 10388 147252 10444
rect 147308 10388 149716 10444
rect 149772 10388 149782 10444
rect 152394 10388 152404 10444
rect 152460 10388 153188 10444
rect 153244 10388 153254 10444
rect 153402 10388 153412 10444
rect 153468 10388 156212 10444
rect 156268 10388 156278 10444
rect 156426 10388 156436 10444
rect 156492 10388 159124 10444
rect 159180 10388 159190 10444
rect 161130 10388 161140 10444
rect 161196 10388 179787 10444
rect 183418 10388 183428 10444
rect 183484 10388 194292 10444
rect 194348 10388 194358 10444
rect 103348 10332 103404 10388
rect 111188 10332 111244 10388
rect 179731 10332 179787 10388
rect 28746 10276 28756 10332
rect 28812 10276 44436 10332
rect 44492 10276 44502 10332
rect 47338 10276 47348 10332
rect 47404 10276 48020 10332
rect 48076 10276 48086 10332
rect 48850 10276 48860 10332
rect 48916 10276 49140 10332
rect 49196 10276 49206 10332
rect 50810 10276 50820 10332
rect 50876 10276 51604 10332
rect 51660 10276 53396 10332
rect 53452 10276 53462 10332
rect 54170 10276 54180 10332
rect 54236 10276 66500 10332
rect 66556 10276 66566 10332
rect 66724 10276 78372 10332
rect 78428 10276 78438 10332
rect 78876 10276 82292 10332
rect 82348 10276 82358 10332
rect 82516 10276 83524 10332
rect 83580 10276 83590 10332
rect 83738 10276 83748 10332
rect 83804 10276 94836 10332
rect 94892 10276 94902 10332
rect 97850 10276 97860 10332
rect 97916 10276 103404 10332
rect 103562 10276 103572 10332
rect 103628 10276 104244 10332
rect 104300 10276 104310 10332
rect 106474 10276 106484 10332
rect 106540 10276 110964 10332
rect 111020 10276 111030 10332
rect 111188 10276 125860 10332
rect 125916 10276 125926 10332
rect 126074 10276 126084 10332
rect 126140 10276 130900 10332
rect 130956 10276 130966 10332
rect 131338 10276 131348 10332
rect 131404 10276 132132 10332
rect 132188 10276 132198 10332
rect 134362 10276 134372 10332
rect 134428 10276 141204 10332
rect 141260 10276 141270 10332
rect 141418 10276 141428 10332
rect 141484 10276 164836 10332
rect 164892 10276 164902 10332
rect 166590 10276 166628 10332
rect 166684 10276 166694 10332
rect 167850 10276 167860 10332
rect 167916 10276 168868 10332
rect 168924 10276 168934 10332
rect 173114 10276 173124 10332
rect 173180 10276 177548 10332
rect 179731 10276 180964 10332
rect 181020 10276 181030 10332
rect 181122 10276 181132 10332
rect 181188 10276 184492 10332
rect 189690 10276 189700 10332
rect 189756 10276 203307 10332
rect 66724 10220 66780 10276
rect 78876 10220 78932 10276
rect 82516 10220 82572 10276
rect 177492 10220 177548 10276
rect 184436 10220 184492 10276
rect 203251 10220 203307 10276
rect 28366 10164 28376 10220
rect 28432 10164 28480 10220
rect 28536 10164 28584 10220
rect 28640 10164 28650 10220
rect 32666 10164 32676 10220
rect 32732 10164 66780 10220
rect 66938 10164 66948 10220
rect 67004 10164 68964 10220
rect 69020 10164 69030 10220
rect 69290 10164 69300 10220
rect 69356 10164 77812 10220
rect 77868 10164 77878 10220
rect 78250 10164 78260 10220
rect 78316 10164 78932 10220
rect 79034 10164 79044 10220
rect 79100 10164 79380 10220
rect 79436 10164 79446 10220
rect 79594 10164 79604 10220
rect 79660 10164 80500 10220
rect 80556 10164 80566 10220
rect 80938 10164 80948 10220
rect 81004 10164 82180 10220
rect 82236 10164 82246 10220
rect 82394 10164 82404 10220
rect 82460 10164 82572 10220
rect 82694 10164 82704 10220
rect 82760 10164 82808 10220
rect 82864 10164 82912 10220
rect 82968 10164 82978 10220
rect 83178 10164 83188 10220
rect 83244 10164 91476 10220
rect 91532 10164 91542 10220
rect 91690 10164 91700 10220
rect 91756 10164 96068 10220
rect 96124 10164 96134 10220
rect 97290 10164 97300 10220
rect 97356 10164 98868 10220
rect 98924 10164 98934 10220
rect 99082 10164 99092 10220
rect 99148 10164 99876 10220
rect 99932 10164 99942 10220
rect 100090 10164 100100 10220
rect 100156 10164 103012 10220
rect 103068 10164 103078 10220
rect 103226 10164 103236 10220
rect 103292 10164 113988 10220
rect 114044 10164 114054 10220
rect 114156 10164 114884 10220
rect 114940 10164 114950 10220
rect 115434 10164 115444 10220
rect 115500 10164 119812 10220
rect 119868 10164 119878 10220
rect 120026 10164 120036 10220
rect 120092 10164 121044 10220
rect 121100 10164 121110 10220
rect 121258 10164 121268 10220
rect 121324 10164 125748 10220
rect 125804 10164 125814 10220
rect 127306 10164 127316 10220
rect 127372 10164 130900 10220
rect 130956 10164 130966 10220
rect 132906 10164 132916 10220
rect 132972 10164 136500 10220
rect 136556 10164 136566 10220
rect 137022 10164 137032 10220
rect 137088 10164 137136 10220
rect 137192 10164 137240 10220
rect 137296 10164 137306 10220
rect 137610 10164 137620 10220
rect 137676 10164 141540 10220
rect 141596 10164 141606 10220
rect 142426 10164 142436 10220
rect 142492 10164 146580 10220
rect 146636 10164 146646 10220
rect 146794 10164 146804 10220
rect 146860 10164 148428 10220
rect 148484 10164 148494 10220
rect 149146 10164 149156 10220
rect 149212 10164 153916 10220
rect 156202 10164 156212 10220
rect 156268 10164 157556 10220
rect 157612 10164 157622 10220
rect 157770 10164 157780 10220
rect 157836 10164 161476 10220
rect 161532 10164 161542 10220
rect 162810 10164 162820 10220
rect 162876 10164 164780 10220
rect 164938 10164 164948 10220
rect 165004 10164 168700 10220
rect 168756 10164 168766 10220
rect 169092 10164 177268 10220
rect 177324 10164 177334 10220
rect 177492 10164 183764 10220
rect 183820 10164 183830 10220
rect 184436 10164 190932 10220
rect 190988 10164 190998 10220
rect 191350 10164 191360 10220
rect 191416 10164 191464 10220
rect 191520 10164 191568 10220
rect 191624 10164 191634 10220
rect 203251 10164 211764 10220
rect 211820 10164 211830 10220
rect 114156 10108 114212 10164
rect 153860 10108 153916 10164
rect 164724 10108 164780 10164
rect 169092 10108 169148 10164
rect 177268 10108 177324 10164
rect 219268 10108 219324 10836
rect 16174 10052 16212 10108
rect 16268 10052 16278 10108
rect 26702 10052 26740 10108
rect 26796 10052 26806 10108
rect 36782 10052 36820 10108
rect 36876 10052 36886 10108
rect 41962 10052 41972 10108
rect 42028 10052 42644 10108
rect 42700 10052 42710 10108
rect 44426 10052 44436 10108
rect 44492 10052 51940 10108
rect 51996 10052 52006 10108
rect 52154 10052 52164 10108
rect 52220 10052 52780 10108
rect 52836 10052 54796 10108
rect 57194 10052 57204 10108
rect 57260 10052 60788 10108
rect 60844 10052 60854 10108
rect 62906 10052 62916 10108
rect 62972 10052 73444 10108
rect 73500 10052 73510 10108
rect 73658 10052 73668 10108
rect 73724 10052 75012 10108
rect 75068 10052 75078 10108
rect 75226 10052 75236 10108
rect 75292 10052 76468 10108
rect 76524 10052 76534 10108
rect 76794 10052 76804 10108
rect 76860 10052 78372 10108
rect 78428 10052 78438 10108
rect 78586 10052 78596 10108
rect 78652 10052 78820 10108
rect 78876 10052 78932 10108
rect 78988 10052 78998 10108
rect 79258 10052 79268 10108
rect 79324 10052 80724 10108
rect 80780 10052 80790 10108
rect 81386 10052 81396 10108
rect 81452 10052 83188 10108
rect 83244 10052 83254 10108
rect 83412 10052 85876 10108
rect 85932 10052 85942 10108
rect 86090 10052 86100 10108
rect 86156 10052 86194 10108
rect 86762 10052 86772 10108
rect 86828 10052 94276 10108
rect 94332 10052 94342 10108
rect 94490 10052 94500 10108
rect 94556 10052 97300 10108
rect 97356 10052 97366 10108
rect 97524 10052 98532 10108
rect 98588 10052 98598 10108
rect 98914 10052 98924 10108
rect 98980 10052 103796 10108
rect 103852 10052 103862 10108
rect 104010 10052 104020 10108
rect 104076 10052 105812 10108
rect 105868 10052 105878 10108
rect 106026 10052 106036 10108
rect 106092 10052 112532 10108
rect 112588 10052 112598 10108
rect 112746 10052 112756 10108
rect 112812 10052 114212 10108
rect 114426 10052 114436 10108
rect 114492 10052 115556 10108
rect 115612 10052 115622 10108
rect 115770 10052 115780 10108
rect 115836 10052 118356 10108
rect 118412 10052 118422 10108
rect 118570 10052 118580 10108
rect 118636 10052 129108 10108
rect 129164 10052 129174 10108
rect 131450 10052 131460 10108
rect 131516 10052 132020 10108
rect 132076 10052 132086 10108
rect 134250 10052 134260 10108
rect 134316 10052 139468 10108
rect 140746 10052 140756 10108
rect 140812 10052 141428 10108
rect 141484 10052 141494 10108
rect 144451 10052 147532 10108
rect 147588 10052 147598 10108
rect 147802 10052 147812 10108
rect 147868 10052 150724 10108
rect 150780 10052 151452 10108
rect 151508 10052 151518 10108
rect 152170 10052 152180 10108
rect 152236 10052 153412 10108
rect 153468 10052 153478 10108
rect 153860 10052 154588 10108
rect 157882 10052 157892 10108
rect 157948 10052 164668 10108
rect 164724 10052 167860 10108
rect 167916 10052 169148 10108
rect 169204 10052 171388 10108
rect 177268 10052 183652 10108
rect 183708 10052 183718 10108
rect 184314 10052 184324 10108
rect 184380 10052 190596 10108
rect 190652 10052 190662 10108
rect 197306 10052 197316 10108
rect 197372 10052 204260 10108
rect 204316 10052 204326 10108
rect 208170 10052 208180 10108
rect 208236 10052 219324 10108
rect 54740 9996 54796 10052
rect 83412 9996 83468 10052
rect 97524 9996 97580 10052
rect 137060 9996 137116 10052
rect 139412 9996 139468 10052
rect 144451 9996 144507 10052
rect 154532 9996 154588 10052
rect 164612 9996 164668 10052
rect 22362 9940 22372 9996
rect 22428 9940 54516 9996
rect 54572 9940 54582 9996
rect 54740 9940 67004 9996
rect 67162 9940 67172 9996
rect 67228 9940 72100 9996
rect 72156 9940 72166 9996
rect 72436 9940 77028 9996
rect 77084 9940 77094 9996
rect 77578 9940 77588 9996
rect 77644 9940 77700 9996
rect 77756 9940 77766 9996
rect 77914 9940 77924 9996
rect 77980 9940 78260 9996
rect 78316 9940 78326 9996
rect 78698 9940 78708 9996
rect 78764 9940 81284 9996
rect 81340 9940 81350 9996
rect 82282 9940 82292 9996
rect 82348 9940 83468 9996
rect 84298 9940 84308 9996
rect 84364 9940 87668 9996
rect 87724 9940 87734 9996
rect 87882 9940 87892 9996
rect 87948 9940 88900 9996
rect 88956 9940 88966 9996
rect 89114 9940 89124 9996
rect 89180 9940 90916 9996
rect 91018 9940 91028 9996
rect 91084 9940 97580 9996
rect 97738 9940 97748 9996
rect 97804 9940 103460 9996
rect 103516 9940 103526 9996
rect 103674 9940 103684 9996
rect 103740 9940 106316 9996
rect 106474 9940 106484 9996
rect 106540 9940 110180 9996
rect 110236 9940 110246 9996
rect 110394 9940 110404 9996
rect 110460 9940 115780 9996
rect 115836 9940 115846 9996
rect 115994 9940 116004 9996
rect 116060 9940 116900 9996
rect 116956 9940 116966 9996
rect 117124 9940 121604 9996
rect 121660 9940 121670 9996
rect 121818 9940 121828 9996
rect 121884 9940 132916 9996
rect 132972 9940 132982 9996
rect 133130 9940 133140 9996
rect 133196 9940 136724 9996
rect 136780 9940 136790 9996
rect 137050 9940 137060 9996
rect 137116 9940 137126 9996
rect 137386 9940 137396 9996
rect 137452 9940 138012 9996
rect 139412 9940 141708 9996
rect 141764 9940 141774 9996
rect 142762 9940 142772 9996
rect 142828 9940 144507 9996
rect 146132 9940 149380 9996
rect 149436 9940 149446 9996
rect 151050 9940 151060 9996
rect 151116 9940 152852 9996
rect 152908 9940 152918 9996
rect 154532 9940 154644 9996
rect 154700 9940 155372 9996
rect 155428 9940 155438 9996
rect 164042 9940 164052 9996
rect 164108 9940 164556 9996
rect 164612 9940 166292 9996
rect 166348 9940 166358 9996
rect 66948 9884 67004 9940
rect 13738 9828 13748 9884
rect 13804 9828 61460 9884
rect 61516 9828 61526 9884
rect 66948 9828 68964 9884
rect 69020 9828 69030 9884
rect 69178 9828 69188 9884
rect 69244 9828 72212 9884
rect 72268 9828 72278 9884
rect 72436 9772 72492 9940
rect 90860 9884 90916 9940
rect 106260 9884 106316 9940
rect 72650 9828 72660 9884
rect 72716 9828 90468 9884
rect 90524 9828 90534 9884
rect 90654 9828 90692 9884
rect 90748 9828 90758 9884
rect 90860 9828 106036 9884
rect 106092 9828 106102 9884
rect 106260 9828 108836 9884
rect 108892 9828 108902 9884
rect 109050 9828 109060 9884
rect 109116 9828 111188 9884
rect 111244 9828 111254 9884
rect 112970 9828 112980 9884
rect 113036 9828 116788 9884
rect 116844 9828 116854 9884
rect 117124 9772 117180 9940
rect 137956 9884 138012 9940
rect 146132 9884 146188 9940
rect 164500 9884 164556 9940
rect 169204 9884 169260 10052
rect 171332 9996 171388 10052
rect 171332 9940 173292 9996
rect 173348 9940 173358 9996
rect 178042 9940 178052 9996
rect 178108 9940 179060 9996
rect 179116 9940 179126 9996
rect 179731 9940 184772 9996
rect 184828 9940 184838 9996
rect 191370 9940 191380 9996
rect 191436 9940 204036 9996
rect 204092 9940 204102 9996
rect 179731 9884 179787 9940
rect 117450 9828 117460 9884
rect 117516 9828 122724 9884
rect 122780 9828 122790 9884
rect 125626 9828 125636 9884
rect 125692 9828 133308 9884
rect 134138 9828 134148 9884
rect 134204 9828 134932 9884
rect 134988 9828 137788 9884
rect 137844 9828 137854 9884
rect 137956 9828 139412 9884
rect 139468 9828 139478 9884
rect 142426 9828 142436 9884
rect 142492 9828 146188 9884
rect 148138 9828 148148 9884
rect 148204 9828 149772 9884
rect 149828 9828 149838 9884
rect 150266 9828 150276 9884
rect 150332 9828 150948 9884
rect 151004 9828 151014 9884
rect 151162 9828 151172 9884
rect 151228 9828 158004 9884
rect 158060 9828 158070 9884
rect 159338 9828 159348 9884
rect 159404 9828 164332 9884
rect 164388 9828 164398 9884
rect 164500 9828 169260 9884
rect 174682 9828 174692 9884
rect 174748 9828 179787 9884
rect 182718 9828 182756 9884
rect 182812 9828 182822 9884
rect 184986 9828 184996 9884
rect 185108 9828 185118 9884
rect 186442 9828 186452 9884
rect 186508 9828 192948 9884
rect 193004 9828 193014 9884
rect 198202 9828 198212 9884
rect 198268 9828 198492 9884
rect 198548 9828 198558 9884
rect 200330 9828 200340 9884
rect 200452 9828 203308 9884
rect 203364 9828 203374 9884
rect 210970 9828 210980 9884
rect 211036 9828 216580 9884
rect 216636 9828 216646 9884
rect 133252 9772 133308 9828
rect 6682 9716 6692 9772
rect 6748 9716 8316 9772
rect 8372 9716 11060 9772
rect 11116 9716 11126 9772
rect 15586 9716 15596 9772
rect 15652 9716 50427 9772
rect 53554 9716 53564 9772
rect 53620 9716 55188 9772
rect 55244 9716 55254 9772
rect 55402 9716 55412 9772
rect 55468 9716 56588 9772
rect 56644 9716 58660 9772
rect 58716 9716 58726 9772
rect 60554 9716 60564 9772
rect 60620 9716 72492 9772
rect 72762 9716 72772 9772
rect 72828 9716 77140 9772
rect 77196 9716 77206 9772
rect 77354 9716 77364 9772
rect 77420 9716 83188 9772
rect 83244 9716 83254 9772
rect 83402 9716 83412 9772
rect 83468 9716 91028 9772
rect 91084 9716 91094 9772
rect 91242 9716 91252 9772
rect 91308 9716 99316 9772
rect 99372 9716 99382 9772
rect 99866 9716 99876 9772
rect 99932 9716 102788 9772
rect 102844 9716 102854 9772
rect 102946 9716 102956 9772
rect 103012 9716 103684 9772
rect 103740 9716 103750 9772
rect 104234 9716 104244 9772
rect 104300 9716 105140 9772
rect 105196 9716 105206 9772
rect 105914 9716 105924 9772
rect 105980 9716 117180 9772
rect 117562 9716 117572 9772
rect 117628 9716 118580 9772
rect 118636 9716 118646 9772
rect 118794 9716 118804 9772
rect 118860 9716 119924 9772
rect 119980 9716 119990 9772
rect 120530 9716 120540 9772
rect 120596 9716 121044 9772
rect 121100 9716 121110 9772
rect 121258 9716 121268 9772
rect 121324 9716 131796 9772
rect 131852 9716 131862 9772
rect 133252 9716 135268 9772
rect 135324 9716 135334 9772
rect 135482 9716 135492 9772
rect 135548 9716 140980 9772
rect 141036 9716 141046 9772
rect 142762 9716 142772 9772
rect 142828 9716 142884 9772
rect 142940 9716 142950 9772
rect 143098 9716 143108 9772
rect 143164 9716 144956 9772
rect 145012 9716 145022 9772
rect 145674 9716 145684 9772
rect 145740 9716 150388 9772
rect 150444 9716 150454 9772
rect 150612 9716 157780 9772
rect 157836 9716 157846 9772
rect 158666 9716 158676 9772
rect 158732 9716 159628 9772
rect 159684 9716 160804 9772
rect 160860 9716 161588 9772
rect 161644 9716 163716 9772
rect 163772 9716 166460 9772
rect 166516 9716 166526 9772
rect 170090 9716 170100 9772
rect 170156 9716 174188 9772
rect 174244 9716 182084 9772
rect 182140 9716 185164 9772
rect 192126 9716 192164 9772
rect 192220 9716 192230 9772
rect 194702 9716 194740 9772
rect 194796 9716 201292 9772
rect 201348 9716 201358 9772
rect 204446 9716 204484 9772
rect 204540 9716 208516 9772
rect 208572 9716 208582 9772
rect 210746 9716 210756 9772
rect 210812 9716 217308 9772
rect 217364 9716 217374 9772
rect 50371 9660 50427 9716
rect 150612 9660 150668 9716
rect 185108 9660 185164 9716
rect 8866 9604 8876 9660
rect 8932 9604 10164 9660
rect 10220 9604 10230 9660
rect 43166 9604 43204 9660
rect 43260 9604 43270 9660
rect 45210 9604 45220 9660
rect 45276 9604 46060 9660
rect 46172 9604 46182 9660
rect 46666 9604 46676 9660
rect 46732 9604 47068 9660
rect 47124 9604 47134 9660
rect 50371 9604 69300 9660
rect 69356 9604 69366 9660
rect 69514 9604 69524 9660
rect 69580 9604 72996 9660
rect 73052 9604 73062 9660
rect 73210 9604 73220 9660
rect 73276 9604 76020 9660
rect 76076 9604 76086 9660
rect 76234 9604 76244 9660
rect 76300 9604 77252 9660
rect 77308 9604 77318 9660
rect 78138 9604 78148 9660
rect 78204 9604 79492 9660
rect 79548 9604 79558 9660
rect 79818 9604 79828 9660
rect 79884 9604 81060 9660
rect 81116 9604 81396 9660
rect 81452 9604 81462 9660
rect 81610 9604 81620 9660
rect 81676 9604 83076 9660
rect 83132 9604 83916 9660
rect 83972 9604 83982 9660
rect 84074 9604 84084 9660
rect 84140 9604 85540 9660
rect 85596 9604 85606 9660
rect 85922 9604 85932 9660
rect 85988 9604 86436 9660
rect 86492 9604 86502 9660
rect 87322 9604 87332 9660
rect 87388 9604 88676 9660
rect 88732 9604 88742 9660
rect 88890 9604 88900 9660
rect 88956 9604 93044 9660
rect 93100 9604 93110 9660
rect 97402 9604 97412 9660
rect 97468 9604 107492 9660
rect 107548 9604 107558 9660
rect 108154 9604 108164 9660
rect 108220 9604 114772 9660
rect 114828 9604 114838 9660
rect 114996 9604 124628 9660
rect 124684 9604 124694 9660
rect 124842 9604 124852 9660
rect 124908 9604 144228 9660
rect 144284 9604 144294 9660
rect 146122 9604 146132 9660
rect 146188 9604 148876 9660
rect 148932 9604 148942 9660
rect 149034 9604 149044 9660
rect 149100 9604 150668 9660
rect 151274 9604 151284 9660
rect 151340 9604 152516 9660
rect 152572 9604 152582 9660
rect 152842 9604 152852 9660
rect 152908 9604 166628 9660
rect 166684 9604 166694 9660
rect 169306 9604 169316 9660
rect 169372 9604 181020 9660
rect 181076 9604 181086 9660
rect 185098 9604 185108 9660
rect 185164 9604 186004 9660
rect 186060 9604 186676 9660
rect 186732 9604 186742 9660
rect 187786 9604 187796 9660
rect 187852 9604 188244 9660
rect 188300 9604 188310 9660
rect 188468 9604 189924 9660
rect 189980 9604 189990 9660
rect 191818 9604 191828 9660
rect 191884 9604 195636 9660
rect 195692 9604 195972 9660
rect 196028 9604 196038 9660
rect 197726 9604 197764 9660
rect 197820 9604 197830 9660
rect 197978 9604 197988 9660
rect 198044 9604 202860 9660
rect 202916 9604 202926 9660
rect 204698 9604 204708 9660
rect 204764 9604 205828 9660
rect 205884 9604 205894 9660
rect 206164 9604 212268 9660
rect 212324 9604 212334 9660
rect 23370 9492 23380 9548
rect 23436 9492 25228 9548
rect 25284 9492 50708 9548
rect 50764 9492 50774 9548
rect 56410 9492 56420 9548
rect 56476 9492 57036 9548
rect 57092 9492 87556 9548
rect 87612 9492 87622 9548
rect 87882 9492 87892 9548
rect 87948 9492 91252 9548
rect 91308 9492 91318 9548
rect 91466 9492 91476 9548
rect 91532 9492 91700 9548
rect 91756 9492 91766 9548
rect 92026 9492 92036 9548
rect 92092 9492 100660 9548
rect 100716 9492 100726 9548
rect 100874 9492 100884 9548
rect 100940 9492 101500 9548
rect 101882 9492 101892 9548
rect 101948 9492 102228 9548
rect 102284 9492 102294 9548
rect 102442 9492 102452 9548
rect 102508 9492 110964 9548
rect 111020 9492 111030 9548
rect 111178 9492 111188 9548
rect 111244 9492 114772 9548
rect 114828 9492 114838 9548
rect 101444 9436 101500 9492
rect 114996 9436 115052 9604
rect 188468 9548 188524 9604
rect 206164 9548 206220 9604
rect 115322 9492 115332 9548
rect 115388 9492 120036 9548
rect 120092 9492 120102 9548
rect 120250 9492 120260 9548
rect 120316 9492 125748 9548
rect 125804 9492 125814 9548
rect 128548 9492 178164 9548
rect 178220 9492 178230 9548
rect 182858 9492 182868 9548
rect 182924 9492 188524 9548
rect 189914 9492 189924 9548
rect 189980 9492 192780 9548
rect 192836 9492 199948 9548
rect 200004 9492 200396 9548
rect 200452 9492 200462 9548
rect 205706 9492 205716 9548
rect 205772 9492 206220 9548
rect 206378 9492 206388 9548
rect 206444 9492 214620 9548
rect 214676 9492 214686 9548
rect 11946 9380 11956 9436
rect 12012 9380 12572 9436
rect 12628 9380 50988 9436
rect 55530 9380 55540 9436
rect 55596 9380 55644 9436
rect 55700 9380 55748 9436
rect 55804 9380 55814 9436
rect 62131 9380 83132 9436
rect 83290 9380 83300 9436
rect 83356 9380 84420 9436
rect 84476 9380 84486 9436
rect 84634 9380 84644 9436
rect 84700 9380 89124 9436
rect 89180 9380 89190 9436
rect 89450 9380 89460 9436
rect 89516 9380 90244 9436
rect 90300 9380 90310 9436
rect 90458 9380 90468 9436
rect 90524 9380 98924 9436
rect 99082 9380 99092 9436
rect 99148 9380 99652 9436
rect 99764 9380 99774 9436
rect 99978 9380 99988 9436
rect 100044 9380 101220 9436
rect 101276 9380 101286 9436
rect 101444 9380 104356 9436
rect 104412 9380 104422 9436
rect 104570 9380 104580 9436
rect 104636 9380 109060 9436
rect 109116 9380 109126 9436
rect 109274 9380 109284 9436
rect 109340 9380 109396 9436
rect 109452 9380 109462 9436
rect 109858 9380 109868 9436
rect 109924 9380 109972 9436
rect 110028 9380 110076 9436
rect 110132 9380 110142 9436
rect 110842 9380 110852 9436
rect 110908 9380 115052 9436
rect 115210 9380 115220 9436
rect 115276 9380 117964 9436
rect 118234 9380 118244 9436
rect 118300 9380 118356 9436
rect 118412 9380 118422 9436
rect 119018 9380 119028 9436
rect 119084 9380 128380 9436
rect 128436 9380 128446 9436
rect 50932 9324 50988 9380
rect 62131 9324 62187 9380
rect 83076 9324 83132 9380
rect 98868 9324 98924 9380
rect 117908 9324 117964 9380
rect 128548 9324 128604 9492
rect 19898 9268 19908 9324
rect 19964 9268 20636 9324
rect 20692 9268 21700 9324
rect 21756 9268 21766 9324
rect 42522 9268 42532 9324
rect 42588 9268 43932 9324
rect 43988 9268 43998 9324
rect 44090 9268 44100 9324
rect 44156 9268 44548 9324
rect 44604 9268 44614 9324
rect 49914 9268 49924 9324
rect 49980 9268 50540 9324
rect 50596 9268 50606 9324
rect 50932 9268 62187 9324
rect 66378 9268 66388 9324
rect 66444 9268 67508 9324
rect 67564 9268 67574 9324
rect 69934 9268 69972 9324
rect 70028 9268 70038 9324
rect 70186 9268 70196 9324
rect 70252 9268 71204 9324
rect 71260 9268 71270 9324
rect 72538 9268 72548 9324
rect 72604 9268 78372 9324
rect 78428 9268 78438 9324
rect 78642 9268 78652 9324
rect 78708 9268 79940 9324
rect 79996 9268 80006 9324
rect 80108 9268 81844 9324
rect 81900 9268 81910 9324
rect 82068 9268 83020 9324
rect 83076 9268 98644 9324
rect 98700 9268 98710 9324
rect 98868 9268 100660 9324
rect 100716 9268 100726 9324
rect 101210 9268 101220 9324
rect 101276 9268 115780 9324
rect 115836 9268 115846 9324
rect 116666 9268 116676 9324
rect 116732 9268 117684 9324
rect 117740 9268 117750 9324
rect 117908 9268 119364 9324
rect 119420 9268 119430 9324
rect 119578 9268 119588 9324
rect 119644 9268 119682 9324
rect 120026 9268 120036 9324
rect 120092 9268 120708 9324
rect 120764 9268 120774 9324
rect 120922 9268 120932 9324
rect 120988 9268 123732 9324
rect 123788 9268 123798 9324
rect 123946 9268 123956 9324
rect 124012 9268 128604 9324
rect 128660 9380 131236 9436
rect 131292 9380 131302 9436
rect 133354 9380 133364 9436
rect 133420 9380 134932 9436
rect 134988 9380 134998 9436
rect 135258 9380 135268 9436
rect 135324 9380 137956 9436
rect 138012 9380 138022 9436
rect 140970 9380 140980 9436
rect 141036 9380 142772 9436
rect 142828 9380 142838 9436
rect 144442 9380 144452 9436
rect 144508 9380 149492 9436
rect 149548 9380 149558 9436
rect 150378 9380 150388 9436
rect 150444 9380 156324 9436
rect 156380 9380 156390 9436
rect 157210 9380 157220 9436
rect 157276 9380 161308 9436
rect 161364 9380 161374 9436
rect 164186 9380 164196 9436
rect 164252 9380 164300 9436
rect 164356 9380 164404 9436
rect 164460 9380 164470 9436
rect 164612 9380 181860 9436
rect 181916 9380 181926 9436
rect 182746 9380 182756 9436
rect 182812 9380 182980 9436
rect 183036 9380 183046 9436
rect 183754 9380 183764 9436
rect 183820 9380 199892 9436
rect 199948 9380 199958 9436
rect 202682 9380 202692 9436
rect 202748 9380 212660 9436
rect 212716 9380 215516 9436
rect 215572 9380 215582 9436
rect 80108 9212 80164 9268
rect 82068 9212 82124 9268
rect 82964 9212 83020 9268
rect 128660 9212 128716 9380
rect 164612 9324 164668 9380
rect 131114 9268 131124 9324
rect 131180 9268 164668 9324
rect 166450 9268 166460 9324
rect 166516 9268 166852 9324
rect 166908 9268 166918 9324
rect 167971 9268 185556 9324
rect 185612 9268 185622 9324
rect 185780 9268 191044 9324
rect 191100 9268 191110 9324
rect 191491 9268 194124 9324
rect 194954 9268 194964 9324
rect 195020 9268 201684 9324
rect 201740 9268 212996 9324
rect 213052 9268 214788 9324
rect 214844 9268 214854 9324
rect 215226 9268 215236 9324
rect 215292 9268 216020 9324
rect 216076 9268 216086 9324
rect 167971 9212 168027 9268
rect 185780 9212 185836 9268
rect 15082 9156 15092 9212
rect 15148 9156 15596 9212
rect 15652 9156 15662 9212
rect 17770 9156 17780 9212
rect 17836 9156 18508 9212
rect 18564 9156 50427 9212
rect 54842 9156 54852 9212
rect 54908 9156 57316 9212
rect 57372 9156 57382 9212
rect 57540 9156 61012 9212
rect 61068 9156 61078 9212
rect 61226 9156 61236 9212
rect 61292 9156 61964 9212
rect 62020 9156 71204 9212
rect 71260 9156 71270 9212
rect 71418 9156 71428 9212
rect 71484 9156 73668 9212
rect 73724 9156 73734 9212
rect 74106 9156 74116 9212
rect 74172 9156 74844 9212
rect 74900 9156 74910 9212
rect 75002 9156 75012 9212
rect 75068 9156 78820 9212
rect 78876 9156 78886 9212
rect 79146 9156 79156 9212
rect 79212 9156 80164 9212
rect 80602 9156 80612 9212
rect 80668 9156 82124 9212
rect 82254 9156 82292 9212
rect 82348 9156 82358 9212
rect 82506 9156 82516 9212
rect 82572 9156 82610 9212
rect 82964 9156 85540 9212
rect 85596 9156 85606 9212
rect 85754 9156 85764 9212
rect 85820 9156 87220 9212
rect 87276 9156 87286 9212
rect 87434 9156 87444 9212
rect 87500 9156 87724 9212
rect 87780 9156 87790 9212
rect 89226 9156 89236 9212
rect 89292 9156 92036 9212
rect 92092 9156 92102 9212
rect 92250 9156 92260 9212
rect 92316 9156 110740 9212
rect 110796 9156 110806 9212
rect 110954 9156 110964 9212
rect 111020 9156 116004 9212
rect 116060 9156 116070 9212
rect 116218 9156 116228 9212
rect 116284 9156 116900 9212
rect 116956 9156 116966 9212
rect 117114 9156 117124 9212
rect 117180 9156 119644 9212
rect 119802 9156 119812 9212
rect 119868 9156 121268 9212
rect 121324 9156 121334 9212
rect 121594 9156 121604 9212
rect 121660 9156 128716 9212
rect 129994 9156 130004 9212
rect 130060 9156 130340 9212
rect 130396 9156 130406 9212
rect 131002 9156 131012 9212
rect 131068 9156 135940 9212
rect 135996 9156 136006 9212
rect 137386 9156 137396 9212
rect 137452 9156 140308 9212
rect 140364 9156 140374 9212
rect 140746 9156 140756 9212
rect 140812 9156 143780 9212
rect 143836 9156 144676 9212
rect 144732 9156 144742 9212
rect 145002 9156 145012 9212
rect 145068 9156 168027 9212
rect 168970 9156 168980 9212
rect 169036 9156 174244 9212
rect 174300 9156 174310 9212
rect 178154 9156 178164 9212
rect 178220 9156 178276 9212
rect 178332 9156 178342 9212
rect 180776 9156 180852 9212
rect 180908 9156 184324 9212
rect 184380 9156 185836 9212
rect 186666 9156 186676 9212
rect 186732 9156 188692 9212
rect 188748 9156 189924 9212
rect 189980 9156 189990 9212
rect 190894 9156 190932 9212
rect 190988 9156 190998 9212
rect 50371 9100 50427 9156
rect 57540 9100 57596 9156
rect 119588 9100 119644 9156
rect 191491 9100 191547 9268
rect 194068 9212 194124 9268
rect 193806 9156 193844 9212
rect 193900 9156 193910 9212
rect 194068 9156 195188 9212
rect 195244 9156 195254 9212
rect 195374 9156 195412 9212
rect 195468 9156 195478 9212
rect 197978 9156 197988 9212
rect 198100 9156 198110 9212
rect 199098 9156 199108 9212
rect 199164 9156 202692 9212
rect 202748 9156 202758 9212
rect 206490 9156 206500 9212
rect 206556 9156 212548 9212
rect 212604 9156 212614 9212
rect 212762 9156 212772 9212
rect 212828 9156 216748 9212
rect 216804 9156 216814 9212
rect 8978 9044 8988 9100
rect 9044 9044 10052 9100
rect 10108 9044 10118 9100
rect 42858 9044 42868 9100
rect 42924 9044 43484 9100
rect 43540 9044 43550 9100
rect 46834 9044 46844 9100
rect 46900 9044 47348 9100
rect 47404 9044 47414 9100
rect 50371 9044 57596 9100
rect 58818 9044 58828 9100
rect 58884 9044 60228 9100
rect 60284 9044 60294 9100
rect 60442 9044 60452 9100
rect 60508 9044 101668 9100
rect 101724 9044 101734 9100
rect 101882 9044 101892 9100
rect 101948 9044 103012 9100
rect 103068 9044 103078 9100
rect 103236 9044 110404 9100
rect 110460 9044 110470 9100
rect 110618 9044 110628 9100
rect 110684 9044 110852 9100
rect 110908 9044 110918 9100
rect 111178 9044 111188 9100
rect 111244 9044 119532 9100
rect 119588 9044 123396 9100
rect 123452 9044 123462 9100
rect 124618 9044 124628 9100
rect 124684 9044 132468 9100
rect 132524 9044 132534 9100
rect 133466 9044 133476 9100
rect 133532 9044 133924 9100
rect 133980 9044 134092 9100
rect 134148 9044 135268 9100
rect 135324 9044 135996 9100
rect 138506 9044 138516 9100
rect 138572 9044 149604 9100
rect 149660 9044 149670 9100
rect 150378 9044 150388 9100
rect 150444 9044 158340 9100
rect 158396 9044 158406 9100
rect 158554 9044 158564 9100
rect 158620 9044 161756 9100
rect 161812 9044 161822 9100
rect 166058 9044 166068 9100
rect 166124 9044 170828 9100
rect 170884 9044 170894 9100
rect 170986 9044 170996 9100
rect 171052 9044 171090 9100
rect 173310 9044 173348 9100
rect 173404 9044 173414 9100
rect 182522 9044 182532 9100
rect 182588 9044 191547 9100
rect 193050 9044 193060 9100
rect 193116 9044 211204 9100
rect 211260 9044 211270 9100
rect 211418 9044 211428 9100
rect 211484 9044 216300 9100
rect 216356 9044 216366 9100
rect 14074 8932 14084 8988
rect 14140 8932 16044 8988
rect 16100 8932 16110 8988
rect 25610 8932 25620 8988
rect 25676 8932 26348 8988
rect 26460 8932 26470 8988
rect 48234 8932 48244 8988
rect 48300 8932 49308 8988
rect 49364 8932 52276 8988
rect 52332 8932 52342 8988
rect 52490 8932 52500 8988
rect 52556 8932 57204 8988
rect 57260 8932 57270 8988
rect 57418 8932 57428 8988
rect 57484 8932 57988 8988
rect 58044 8932 58828 8988
rect 59378 8932 59388 8988
rect 59444 8932 60340 8988
rect 60396 8932 60406 8988
rect 64922 8932 64932 8988
rect 64988 8932 65324 8988
rect 65380 8932 77980 8988
rect 78194 8932 78204 8988
rect 78260 8932 79268 8988
rect 79324 8932 79334 8988
rect 79482 8932 79492 8988
rect 79548 8932 80500 8988
rect 80556 8932 80566 8988
rect 80714 8932 80724 8988
rect 80780 8932 81060 8988
rect 81116 8932 81126 8988
rect 81284 8932 81900 8988
rect 82170 8932 82180 8988
rect 82236 8932 84252 8988
rect 84308 8932 84868 8988
rect 84924 8932 84934 8988
rect 85082 8932 85092 8988
rect 85148 8932 85428 8988
rect 85484 8932 85494 8988
rect 85642 8932 85652 8988
rect 85708 8932 88396 8988
rect 90906 8932 90916 8988
rect 90972 8932 94220 8988
rect 95330 8932 95340 8988
rect 95396 8932 95956 8988
rect 96012 8932 96022 8988
rect 98522 8932 98532 8988
rect 98588 8932 102900 8988
rect 102956 8932 102966 8988
rect 58772 8876 58828 8932
rect 77924 8876 77980 8932
rect 81284 8876 81340 8932
rect 81844 8876 81900 8932
rect 13626 8820 13636 8876
rect 13692 8820 58268 8876
rect 58324 8820 58334 8876
rect 58772 8820 66724 8876
rect 66780 8820 66790 8876
rect 67050 8820 67060 8876
rect 67116 8820 70420 8876
rect 70476 8820 70486 8876
rect 70578 8820 70588 8876
rect 70644 8820 72772 8876
rect 72828 8820 72838 8876
rect 72986 8820 72996 8876
rect 73052 8820 77812 8876
rect 77924 8820 81340 8876
rect 81498 8820 81508 8876
rect 81564 8820 81788 8876
rect 81844 8820 88116 8876
rect 88172 8820 88182 8876
rect 77756 8764 77812 8820
rect 81732 8764 81788 8820
rect 88340 8764 88396 8932
rect 94164 8876 94220 8932
rect 103236 8876 103292 9044
rect 119476 8988 119532 9044
rect 135940 8988 135996 9044
rect 103450 8932 103460 8988
rect 103516 8932 118132 8988
rect 118188 8932 118198 8988
rect 118682 8932 118692 8988
rect 118748 8932 119252 8988
rect 119308 8932 119318 8988
rect 119476 8932 126980 8988
rect 127036 8932 127046 8988
rect 127194 8932 127204 8988
rect 127260 8932 132636 8988
rect 132804 8932 134260 8988
rect 134316 8932 135772 8988
rect 135828 8932 135838 8988
rect 135930 8932 135940 8988
rect 135996 8932 138292 8988
rect 138348 8932 139748 8988
rect 139804 8932 140308 8988
rect 140364 8932 140756 8988
rect 140812 8932 140822 8988
rect 143882 8932 143892 8988
rect 143948 8932 168980 8988
rect 169036 8932 169046 8988
rect 169194 8932 169204 8988
rect 169260 8932 183428 8988
rect 183484 8932 183494 8988
rect 183698 8932 183708 8988
rect 183764 8932 195524 8988
rect 195580 8932 195590 8988
rect 195962 8932 195972 8988
rect 196028 8932 199388 8988
rect 200386 8932 200396 8988
rect 200452 8932 201740 8988
rect 201796 8932 201806 8988
rect 201898 8932 201908 8988
rect 201964 8932 206388 8988
rect 206444 8932 206454 8988
rect 208394 8932 208404 8988
rect 208460 8932 213948 8988
rect 214004 8932 214014 8988
rect 215562 8932 215572 8988
rect 215628 8932 216580 8988
rect 216636 8932 216646 8988
rect 132580 8876 132860 8932
rect 88666 8820 88676 8876
rect 88732 8820 90636 8876
rect 90794 8820 90804 8876
rect 90860 8820 93940 8876
rect 93996 8820 94006 8876
rect 94164 8820 103292 8876
rect 103450 8820 103460 8876
rect 103516 8820 106596 8876
rect 106652 8820 106662 8876
rect 107482 8820 107492 8876
rect 107548 8820 127988 8876
rect 128044 8820 128054 8876
rect 134026 8820 134036 8876
rect 134092 8820 139524 8876
rect 139580 8820 139590 8876
rect 139748 8820 144452 8876
rect 144508 8820 144518 8876
rect 144666 8820 144676 8876
rect 144732 8820 146020 8876
rect 146076 8820 146580 8876
rect 146636 8820 147420 8876
rect 147476 8820 148820 8876
rect 148876 8820 148886 8876
rect 149044 8820 181524 8876
rect 181580 8820 181590 8876
rect 186106 8820 186116 8876
rect 186172 8820 197988 8876
rect 198044 8820 198054 8876
rect 90580 8764 90636 8820
rect 139748 8764 139804 8820
rect 149044 8764 149100 8820
rect 199332 8764 199388 8932
rect 201282 8820 201292 8876
rect 201348 8820 214116 8876
rect 214172 8820 214182 8876
rect 219200 8764 220000 8792
rect 21914 8708 21924 8764
rect 21980 8708 22484 8764
rect 22540 8708 77588 8764
rect 77644 8708 77654 8764
rect 77756 8708 79716 8764
rect 79772 8708 79782 8764
rect 79930 8708 79940 8764
rect 79996 8708 80034 8764
rect 80490 8708 80500 8764
rect 80556 8708 81564 8764
rect 81732 8708 84700 8764
rect 84756 8708 84766 8764
rect 84858 8708 84868 8764
rect 84924 8708 86212 8764
rect 86268 8708 86278 8764
rect 86426 8708 86436 8764
rect 86492 8708 88116 8764
rect 88172 8708 88182 8764
rect 88340 8708 90412 8764
rect 90468 8708 90478 8764
rect 90580 8708 118468 8764
rect 118524 8708 118534 8764
rect 119354 8708 119364 8764
rect 119420 8708 124852 8764
rect 124908 8708 124918 8764
rect 127082 8708 127092 8764
rect 127148 8708 133364 8764
rect 133420 8708 133430 8764
rect 133690 8708 133700 8764
rect 133756 8708 135604 8764
rect 135660 8708 135670 8764
rect 136266 8708 136276 8764
rect 136332 8708 139804 8764
rect 140186 8708 140196 8764
rect 140252 8708 140980 8764
rect 141036 8708 141046 8764
rect 141754 8708 141764 8764
rect 141820 8708 149100 8764
rect 149258 8708 149268 8764
rect 149324 8708 172900 8764
rect 172956 8708 172966 8764
rect 178042 8708 178052 8764
rect 178108 8708 178500 8764
rect 178556 8708 185052 8764
rect 188010 8708 188020 8764
rect 188076 8708 193172 8764
rect 193228 8708 193238 8764
rect 193834 8708 193844 8764
rect 193900 8708 199108 8764
rect 199164 8708 199174 8764
rect 199332 8708 203307 8764
rect 212538 8708 212548 8764
rect 212604 8708 215180 8764
rect 81508 8652 81564 8708
rect 28366 8596 28376 8652
rect 28432 8596 28480 8652
rect 28536 8596 28584 8652
rect 28640 8596 28650 8652
rect 48234 8596 48244 8652
rect 48300 8596 48804 8652
rect 48860 8596 48870 8652
rect 51940 8596 60564 8652
rect 60620 8596 60630 8652
rect 60778 8596 60788 8652
rect 60844 8596 70196 8652
rect 70252 8596 70262 8652
rect 70410 8596 70420 8652
rect 70476 8596 77812 8652
rect 77868 8596 77878 8652
rect 77970 8596 77980 8652
rect 78036 8596 79436 8652
rect 79492 8596 79502 8652
rect 79706 8596 79716 8652
rect 79772 8596 81284 8652
rect 81340 8596 81350 8652
rect 81508 8596 82516 8652
rect 82572 8596 82582 8652
rect 82694 8596 82704 8652
rect 82760 8596 82808 8652
rect 82864 8596 82912 8652
rect 82968 8596 82978 8652
rect 83066 8596 83076 8652
rect 83132 8596 83748 8652
rect 83804 8596 83814 8652
rect 83962 8596 83972 8652
rect 84028 8596 85652 8652
rect 85708 8596 85718 8652
rect 85978 8596 85988 8652
rect 86044 8596 87108 8652
rect 87164 8596 87174 8652
rect 87322 8596 87332 8652
rect 87388 8596 88732 8652
rect 88890 8596 88900 8652
rect 88956 8596 91700 8652
rect 91756 8596 91766 8652
rect 92596 8596 99876 8652
rect 99932 8596 99942 8652
rect 100426 8596 100436 8652
rect 100492 8596 102452 8652
rect 102508 8596 102518 8652
rect 102666 8596 102676 8652
rect 102732 8596 106372 8652
rect 106428 8596 106438 8652
rect 106586 8596 106596 8652
rect 106652 8596 108892 8652
rect 109162 8596 109172 8652
rect 109228 8596 115220 8652
rect 115276 8596 115286 8652
rect 115434 8596 115444 8652
rect 115500 8596 115538 8652
rect 115770 8596 115780 8652
rect 115836 8596 117852 8652
rect 118122 8596 118132 8652
rect 118188 8596 120372 8652
rect 120428 8596 120438 8652
rect 120698 8596 120708 8652
rect 120764 8596 122164 8652
rect 122220 8596 122230 8652
rect 122378 8596 122388 8652
rect 122444 8596 123508 8652
rect 123564 8596 123574 8652
rect 123722 8596 123732 8652
rect 123788 8596 130676 8652
rect 130732 8596 130742 8652
rect 131114 8596 131124 8652
rect 131180 8596 133364 8652
rect 133420 8596 135156 8652
rect 135212 8596 135222 8652
rect 137022 8596 137032 8652
rect 137088 8596 137136 8652
rect 137192 8596 137240 8652
rect 137296 8596 137306 8652
rect 139626 8596 139636 8652
rect 139692 8596 183540 8652
rect 183596 8596 183606 8652
rect 51940 8540 51996 8596
rect 88676 8540 88732 8596
rect 92596 8540 92652 8596
rect 108836 8540 108892 8596
rect 117796 8540 117852 8596
rect 184996 8540 185052 8708
rect 203251 8652 203307 8708
rect 190820 8596 191212 8652
rect 191350 8596 191360 8652
rect 191416 8596 191464 8652
rect 191520 8596 191568 8652
rect 191624 8596 191634 8652
rect 196746 8596 196756 8652
rect 196812 8596 199444 8652
rect 199500 8596 201908 8652
rect 201964 8596 201974 8652
rect 203251 8596 212212 8652
rect 212268 8596 213500 8652
rect 213556 8596 213566 8652
rect 190820 8540 190876 8596
rect 30090 8484 30100 8540
rect 30156 8484 51996 8540
rect 52154 8484 52164 8540
rect 52220 8484 55972 8540
rect 56028 8484 56038 8540
rect 56420 8484 60452 8540
rect 60508 8484 60518 8540
rect 60666 8484 60676 8540
rect 60732 8484 72772 8540
rect 72828 8484 72838 8540
rect 72986 8484 72996 8540
rect 73052 8484 78484 8540
rect 78540 8484 78550 8540
rect 78708 8484 86436 8540
rect 86492 8484 86502 8540
rect 86650 8484 86660 8540
rect 86716 8484 87276 8540
rect 87434 8484 87444 8540
rect 87500 8484 88452 8540
rect 88508 8484 88518 8540
rect 88676 8484 91196 8540
rect 91252 8484 91262 8540
rect 91354 8484 91364 8540
rect 91420 8484 92652 8540
rect 93258 8484 93268 8540
rect 93324 8484 95284 8540
rect 95340 8484 95350 8540
rect 96282 8484 96292 8540
rect 96348 8484 96964 8540
rect 97020 8484 97030 8540
rect 98980 8484 102452 8540
rect 102508 8484 102518 8540
rect 103674 8484 103684 8540
rect 103740 8484 108612 8540
rect 108668 8484 108678 8540
rect 108836 8484 117572 8540
rect 117628 8484 117638 8540
rect 117796 8484 121156 8540
rect 121212 8484 121222 8540
rect 121324 8484 122500 8540
rect 122556 8484 122566 8540
rect 124058 8484 124068 8540
rect 124124 8484 126532 8540
rect 126588 8484 126598 8540
rect 126970 8484 126980 8540
rect 127036 8484 138516 8540
rect 138572 8484 138582 8540
rect 138842 8484 138852 8540
rect 138908 8484 139748 8540
rect 139804 8484 139814 8540
rect 141082 8484 141092 8540
rect 141148 8484 142996 8540
rect 143052 8484 143062 8540
rect 144666 8484 144676 8540
rect 144732 8484 148484 8540
rect 148540 8484 148550 8540
rect 148698 8484 148708 8540
rect 148764 8484 151116 8540
rect 151172 8484 151182 8540
rect 151386 8484 151396 8540
rect 151452 8484 151844 8540
rect 151900 8484 152292 8540
rect 152348 8484 153076 8540
rect 153132 8484 153142 8540
rect 153300 8484 157444 8540
rect 157500 8484 157510 8540
rect 157770 8484 157780 8540
rect 157836 8484 168756 8540
rect 168812 8484 168822 8540
rect 170426 8484 170436 8540
rect 170492 8484 171668 8540
rect 171724 8484 171734 8540
rect 173012 8484 181300 8540
rect 181356 8484 181366 8540
rect 181850 8484 181860 8540
rect 181916 8484 182756 8540
rect 182812 8484 182822 8540
rect 184996 8484 190876 8540
rect 191156 8540 191212 8596
rect 215124 8540 215180 8708
rect 219044 8708 220000 8764
rect 191156 8484 193732 8540
rect 193788 8484 193798 8540
rect 197530 8484 197540 8540
rect 197596 8484 200116 8540
rect 200172 8484 214396 8540
rect 214452 8484 214462 8540
rect 215114 8484 215124 8540
rect 215180 8484 215684 8540
rect 215740 8484 215750 8540
rect 56420 8428 56476 8484
rect 78708 8428 78764 8484
rect 87220 8428 87276 8484
rect 98980 8428 99036 8484
rect 121324 8428 121380 8484
rect 153300 8428 153356 8484
rect 9706 8372 9716 8428
rect 9772 8372 56476 8428
rect 58986 8372 58996 8428
rect 59052 8372 59444 8428
rect 59500 8372 63252 8428
rect 63308 8372 63318 8428
rect 63466 8372 63476 8428
rect 63532 8372 65604 8428
rect 65660 8372 65670 8428
rect 66826 8372 66836 8428
rect 66892 8372 67788 8428
rect 67946 8372 67956 8428
rect 68012 8372 69748 8428
rect 69804 8372 69814 8428
rect 70308 8372 72100 8428
rect 72156 8372 72166 8428
rect 72650 8372 72660 8428
rect 72716 8372 74676 8428
rect 74732 8372 74742 8428
rect 74890 8372 74900 8428
rect 74956 8372 78764 8428
rect 78820 8372 85932 8428
rect 85988 8372 85998 8428
rect 86090 8372 86100 8428
rect 86156 8372 86772 8428
rect 86828 8372 86838 8428
rect 87220 8372 99036 8428
rect 99194 8372 99204 8428
rect 99260 8372 100436 8428
rect 100492 8372 100502 8428
rect 100650 8372 100660 8428
rect 100716 8372 105700 8428
rect 105756 8372 105766 8428
rect 105924 8372 116004 8428
rect 116060 8372 116070 8428
rect 116218 8372 116228 8428
rect 116284 8372 116732 8428
rect 117002 8372 117012 8428
rect 117068 8372 118244 8428
rect 118300 8372 118310 8428
rect 118794 8372 118804 8428
rect 118860 8372 121380 8428
rect 121492 8372 124852 8428
rect 124908 8372 124918 8428
rect 125066 8372 125076 8428
rect 125132 8372 126700 8428
rect 127950 8372 127988 8428
rect 128044 8372 128054 8428
rect 128212 8372 132916 8428
rect 132972 8372 132982 8428
rect 135370 8372 135380 8428
rect 135436 8372 142828 8428
rect 143658 8372 143668 8428
rect 143724 8372 145460 8428
rect 145516 8372 145526 8428
rect 145674 8372 145684 8428
rect 145740 8372 149380 8428
rect 149436 8372 149446 8428
rect 149594 8372 149604 8428
rect 149660 8372 150052 8428
rect 150108 8372 150500 8428
rect 150556 8372 150566 8428
rect 150938 8372 150948 8428
rect 151004 8372 152740 8428
rect 152796 8372 152806 8428
rect 152954 8372 152964 8428
rect 153020 8372 153356 8428
rect 153962 8372 153972 8428
rect 154028 8372 156100 8428
rect 156156 8372 156166 8428
rect 157780 8372 158564 8428
rect 158620 8372 158630 8428
rect 158788 8372 170324 8428
rect 170380 8372 170390 8428
rect 67732 8316 67788 8372
rect 70308 8316 70364 8372
rect 78820 8316 78876 8372
rect 105924 8316 105980 8372
rect 10238 8260 10276 8316
rect 10332 8260 10342 8316
rect 12842 8260 12852 8316
rect 12908 8260 13580 8316
rect 13636 8260 13646 8316
rect 43194 8260 43204 8316
rect 43260 8260 64260 8316
rect 64316 8260 64326 8316
rect 65706 8260 65716 8316
rect 65772 8260 66556 8316
rect 66612 8260 66948 8316
rect 67004 8260 67014 8316
rect 67732 8260 70364 8316
rect 70522 8260 70532 8316
rect 70588 8260 74340 8316
rect 74396 8260 74406 8316
rect 74890 8260 74900 8316
rect 74956 8260 76804 8316
rect 76860 8260 76870 8316
rect 77130 8260 77140 8316
rect 77196 8260 78876 8316
rect 79034 8260 79044 8316
rect 79100 8260 79268 8316
rect 79324 8260 79334 8316
rect 79482 8260 79492 8316
rect 79548 8260 81844 8316
rect 81900 8260 81910 8316
rect 82058 8260 82068 8316
rect 82124 8260 85316 8316
rect 85372 8260 85382 8316
rect 85530 8260 85540 8316
rect 85596 8260 87780 8316
rect 88498 8260 88508 8316
rect 88564 8260 89460 8316
rect 89516 8260 89526 8316
rect 89870 8260 89908 8316
rect 89964 8260 89974 8316
rect 90132 8260 99540 8316
rect 99596 8260 99606 8316
rect 100090 8260 100100 8316
rect 100156 8260 100548 8316
rect 100604 8260 100614 8316
rect 100762 8260 100772 8316
rect 100828 8260 101220 8316
rect 101276 8260 101286 8316
rect 101434 8260 101444 8316
rect 101500 8260 103908 8316
rect 103964 8260 103974 8316
rect 104122 8260 104132 8316
rect 104188 8260 105980 8316
rect 107258 8260 107268 8316
rect 107324 8260 107884 8316
rect 107940 8260 107950 8316
rect 108276 8260 109172 8316
rect 109228 8260 109620 8316
rect 109676 8260 109686 8316
rect 110394 8260 110404 8316
rect 110516 8260 110526 8316
rect 110730 8260 110740 8316
rect 110796 8260 116452 8316
rect 116508 8260 116518 8316
rect 87724 8204 87780 8260
rect 90132 8204 90188 8260
rect 108276 8204 108332 8260
rect 116676 8204 116732 8372
rect 121492 8316 121548 8372
rect 126644 8316 126700 8372
rect 128212 8316 128268 8372
rect 117114 8260 117124 8316
rect 117180 8260 117460 8316
rect 117516 8260 117526 8316
rect 117674 8260 117684 8316
rect 117740 8260 121548 8316
rect 121706 8260 121716 8316
rect 121772 8260 121828 8316
rect 121884 8260 121894 8316
rect 124730 8260 124740 8316
rect 124796 8260 125972 8316
rect 126028 8260 126038 8316
rect 126634 8260 126644 8316
rect 126700 8260 126710 8316
rect 127642 8260 127652 8316
rect 127708 8260 128268 8316
rect 128426 8260 128436 8316
rect 128492 8260 133700 8316
rect 133756 8260 133766 8316
rect 134810 8260 134820 8316
rect 134876 8260 137620 8316
rect 137676 8260 137686 8316
rect 142772 8204 142828 8372
rect 157780 8316 157836 8372
rect 158788 8316 158844 8372
rect 173012 8316 173068 8484
rect 219044 8428 219100 8708
rect 219200 8680 220000 8708
rect 144442 8260 144452 8316
rect 144508 8260 144564 8316
rect 144620 8260 144630 8316
rect 145226 8260 145236 8316
rect 145292 8260 147532 8316
rect 147588 8260 147598 8316
rect 148474 8260 148484 8316
rect 148540 8260 152852 8316
rect 152908 8260 152918 8316
rect 153188 8260 157836 8316
rect 158330 8260 158340 8316
rect 158396 8260 158844 8316
rect 160570 8260 160580 8316
rect 160636 8260 166964 8316
rect 167020 8260 167030 8316
rect 167850 8260 167860 8316
rect 167916 8260 169092 8316
rect 169148 8260 169158 8316
rect 169530 8260 169540 8316
rect 169596 8260 170772 8316
rect 170828 8260 173068 8316
rect 173796 8372 180404 8428
rect 180460 8372 180470 8428
rect 181290 8372 181300 8428
rect 181356 8372 190708 8428
rect 190764 8372 190774 8428
rect 191034 8372 191044 8428
rect 191100 8372 194796 8428
rect 153188 8204 153244 8260
rect 173796 8204 173852 8372
rect 194740 8316 194796 8372
rect 197316 8372 198940 8428
rect 198996 8372 199006 8428
rect 219044 8372 219324 8428
rect 197316 8316 197372 8372
rect 219268 8316 219324 8372
rect 175018 8260 175028 8316
rect 175084 8260 183652 8316
rect 183708 8260 183718 8316
rect 185070 8260 185108 8316
rect 185164 8260 185174 8316
rect 187562 8260 187572 8316
rect 187684 8260 187694 8316
rect 194740 8260 197316 8316
rect 197372 8260 197382 8316
rect 197530 8260 197540 8316
rect 197596 8260 197634 8316
rect 199882 8260 199892 8316
rect 199948 8260 206556 8316
rect 206714 8260 206724 8316
rect 206780 8260 209188 8316
rect 209244 8260 209254 8316
rect 209850 8260 209860 8316
rect 209916 8260 219324 8316
rect 206500 8204 206556 8260
rect 26618 8148 26628 8204
rect 26684 8148 27468 8204
rect 27524 8148 27534 8204
rect 29530 8148 29540 8204
rect 29596 8148 30324 8204
rect 30380 8148 30390 8204
rect 31546 8148 31556 8204
rect 31612 8148 32340 8204
rect 32396 8148 32406 8204
rect 34906 8148 34916 8204
rect 34972 8148 35756 8204
rect 35812 8148 35822 8204
rect 36362 8148 36372 8204
rect 36428 8148 36932 8204
rect 36988 8148 36998 8204
rect 38611 8148 50427 8204
rect 51818 8148 51828 8204
rect 51884 8148 60004 8204
rect 60060 8148 60070 8204
rect 60498 8148 60508 8204
rect 60564 8148 63252 8204
rect 63308 8148 63318 8204
rect 66042 8148 66052 8204
rect 66108 8148 69412 8204
rect 69468 8148 69478 8204
rect 70634 8148 70644 8204
rect 70700 8148 71204 8204
rect 71260 8148 71270 8204
rect 71418 8148 71428 8204
rect 71484 8148 71988 8204
rect 72044 8148 72054 8204
rect 72426 8148 72436 8204
rect 72492 8148 81284 8204
rect 81340 8148 81350 8204
rect 81722 8148 81732 8204
rect 81788 8148 81844 8204
rect 81900 8148 81910 8204
rect 82282 8148 82292 8204
rect 82348 8148 84532 8204
rect 84588 8148 84598 8204
rect 84746 8148 84756 8204
rect 84812 8148 87556 8204
rect 87612 8148 87622 8204
rect 87724 8148 90188 8204
rect 90346 8148 90356 8204
rect 90412 8148 93268 8204
rect 93324 8148 93334 8204
rect 94714 8148 94724 8204
rect 94780 8148 98644 8204
rect 98700 8148 98710 8204
rect 98858 8148 98868 8204
rect 98924 8148 108332 8204
rect 108602 8148 108612 8204
rect 108668 8148 112980 8204
rect 113036 8148 113046 8204
rect 113642 8148 113652 8204
rect 113708 8148 116452 8204
rect 116508 8148 116518 8204
rect 116676 8148 117908 8204
rect 117964 8148 117974 8204
rect 118122 8148 118132 8204
rect 118188 8148 120260 8204
rect 120316 8148 120326 8204
rect 120810 8148 120820 8204
rect 120876 8148 123340 8204
rect 123396 8148 123406 8204
rect 126410 8148 126420 8204
rect 126476 8148 129444 8204
rect 129500 8148 129510 8204
rect 132346 8148 132356 8204
rect 132412 8148 133252 8204
rect 133308 8148 133318 8204
rect 134922 8148 134932 8204
rect 134988 8148 141092 8204
rect 141148 8148 141158 8204
rect 142772 8148 144788 8204
rect 144844 8148 144854 8204
rect 145002 8148 145012 8204
rect 145068 8148 145124 8204
rect 145180 8148 146020 8204
rect 146076 8148 146086 8204
rect 146346 8148 146356 8204
rect 146412 8148 150164 8204
rect 150220 8148 150230 8204
rect 150658 8148 150668 8204
rect 150724 8148 151396 8204
rect 151452 8148 151462 8204
rect 151890 8148 151900 8204
rect 151956 8148 152628 8204
rect 152684 8148 153244 8204
rect 155978 8148 155988 8204
rect 156044 8148 160692 8204
rect 160748 8148 160758 8204
rect 166618 8148 166628 8204
rect 166684 8148 173852 8204
rect 177594 8148 177604 8204
rect 177660 8148 187516 8204
rect 187572 8148 187582 8204
rect 188458 8148 188468 8204
rect 188524 8148 202188 8204
rect 202244 8148 202254 8204
rect 203028 8148 203924 8204
rect 203980 8148 203990 8204
rect 206500 8148 206948 8204
rect 207004 8148 214508 8204
rect 214564 8148 214574 8204
rect 38611 8092 38667 8148
rect 50371 8092 50427 8148
rect 203028 8092 203084 8148
rect 11610 8036 11620 8092
rect 11676 8036 13916 8092
rect 14028 8036 14038 8092
rect 16650 8036 16660 8092
rect 16716 8036 19180 8092
rect 19236 8036 19348 8092
rect 19404 8036 19414 8092
rect 25050 8036 25060 8092
rect 25116 8036 25452 8092
rect 25508 8036 38667 8092
rect 47272 8036 47348 8092
rect 47404 8036 48580 8092
rect 48636 8036 48646 8092
rect 50371 8036 62187 8092
rect 62570 8036 62580 8092
rect 62636 8036 74900 8092
rect 74956 8036 74966 8092
rect 75114 8036 75124 8092
rect 75180 8036 77476 8092
rect 77532 8036 77542 8092
rect 77914 8036 77924 8092
rect 77980 8036 78708 8092
rect 78764 8036 78774 8092
rect 78866 8036 78876 8092
rect 78932 8036 80052 8092
rect 80108 8036 80118 8092
rect 80378 8036 80388 8092
rect 80444 8036 80948 8092
rect 81004 8036 81014 8092
rect 81274 8036 81284 8092
rect 81340 8036 82180 8092
rect 82236 8036 82246 8092
rect 82394 8036 82404 8092
rect 82460 8036 83972 8092
rect 84028 8036 84038 8092
rect 84410 8036 84420 8092
rect 84476 8036 87668 8092
rect 87724 8036 87734 8092
rect 89226 8036 89236 8092
rect 89292 8036 91084 8092
rect 91140 8036 91150 8092
rect 91242 8036 91252 8092
rect 91308 8036 93268 8092
rect 93324 8036 93334 8092
rect 95722 8036 95732 8092
rect 95788 8036 96404 8092
rect 96460 8036 96470 8092
rect 96954 8036 96964 8092
rect 97020 8036 101220 8092
rect 101276 8036 101286 8092
rect 101434 8036 101444 8092
rect 101500 8036 101668 8092
rect 101770 8036 101780 8092
rect 101836 8036 102228 8092
rect 102284 8036 102294 8092
rect 102554 8036 102564 8092
rect 102620 8036 104076 8092
rect 104132 8036 104142 8092
rect 104794 8036 104804 8092
rect 104860 8036 110740 8092
rect 110796 8036 110806 8092
rect 110898 8036 110908 8092
rect 110964 8036 111076 8092
rect 111132 8036 111142 8092
rect 111290 8036 111300 8092
rect 111356 8036 112028 8092
rect 112298 8036 112308 8092
rect 112364 8036 112532 8092
rect 112588 8036 112598 8092
rect 113082 8036 113092 8092
rect 113148 8036 118244 8092
rect 118300 8036 118310 8092
rect 118458 8036 118468 8092
rect 118524 8036 119364 8092
rect 119420 8036 119430 8092
rect 119802 8036 119812 8092
rect 119868 8036 121492 8092
rect 121548 8036 121558 8092
rect 122042 8036 122052 8092
rect 122108 8036 123228 8092
rect 123284 8036 123294 8092
rect 123386 8036 123396 8092
rect 123452 8036 127092 8092
rect 127148 8036 127158 8092
rect 127530 8036 127540 8092
rect 127596 8036 132916 8092
rect 132972 8036 132982 8092
rect 133130 8036 133140 8092
rect 133196 8036 135828 8092
rect 135884 8036 135894 8092
rect 136490 8036 136500 8092
rect 136556 8036 136948 8092
rect 137004 8036 137508 8092
rect 137564 8036 137574 8092
rect 137946 8036 137956 8092
rect 138012 8036 144564 8092
rect 144620 8036 144630 8092
rect 144778 8036 144788 8092
rect 144844 8036 156267 8092
rect 158554 8036 158564 8092
rect 158620 8036 173404 8092
rect 173460 8036 173470 8092
rect 174990 8036 175028 8092
rect 175084 8036 175094 8092
rect 175924 8036 181076 8092
rect 181132 8036 181142 8092
rect 181290 8036 181300 8092
rect 181356 8036 191324 8092
rect 191380 8036 191390 8092
rect 193050 8036 193060 8092
rect 193116 8036 194348 8092
rect 202010 8036 202020 8092
rect 202076 8036 203084 8092
rect 203140 8036 203150 8092
rect 203251 8036 206052 8092
rect 206108 8036 206118 8092
rect 211866 8036 211876 8092
rect 211932 8036 212268 8092
rect 212324 8036 212334 8092
rect 212706 8036 212716 8092
rect 212772 8036 216300 8092
rect 216412 8036 216422 8092
rect 62131 7980 62187 8036
rect 101612 7980 101668 8036
rect 111972 7980 112028 8036
rect 156211 7980 156267 8036
rect 175924 7980 175980 8036
rect 194292 7980 194348 8036
rect 203251 7980 203307 8036
rect 74 7924 84 7980
rect 140 7924 364 7980
rect 23370 7924 23380 7980
rect 23436 7924 25900 7980
rect 26012 7924 26022 7980
rect 40730 7924 40740 7980
rect 40796 7924 53620 7980
rect 53676 7924 53686 7980
rect 54030 7924 54068 7980
rect 54124 7924 54134 7980
rect 56634 7924 56644 7980
rect 56700 7924 57428 7980
rect 57484 7924 60676 7980
rect 60732 7924 60742 7980
rect 62131 7924 70532 7980
rect 70588 7924 70598 7980
rect 72202 7924 72212 7980
rect 72268 7924 77252 7980
rect 77308 7924 77318 7980
rect 77466 7924 77476 7980
rect 77532 7924 77588 7980
rect 77644 7924 77654 7980
rect 77802 7924 77812 7980
rect 77868 7924 84084 7980
rect 84140 7924 84150 7980
rect 84298 7924 84308 7980
rect 84364 7924 85092 7980
rect 85148 7924 85158 7980
rect 85250 7924 85260 7980
rect 85316 7924 85820 7980
rect 85876 7924 86548 7980
rect 86604 7924 86614 7980
rect 86874 7924 86884 7980
rect 86940 7924 87220 7980
rect 87276 7924 87286 7980
rect 87546 7924 87556 7980
rect 87612 7924 89068 7980
rect 89124 7924 89572 7980
rect 89628 7924 89638 7980
rect 90132 7924 90804 7980
rect 90860 7924 90870 7980
rect 91018 7924 91028 7980
rect 91084 7924 91924 7980
rect 91980 7924 91990 7980
rect 95386 7924 95396 7980
rect 95452 7924 96068 7980
rect 96124 7924 96852 7980
rect 96908 7924 96918 7980
rect 97626 7924 97636 7980
rect 97692 7924 101444 7980
rect 101500 7924 101510 7980
rect 101612 7924 107492 7980
rect 107548 7924 107558 7980
rect 107706 7924 107716 7980
rect 107772 7924 111748 7980
rect 111804 7924 111814 7980
rect 111972 7924 113876 7980
rect 113932 7924 113942 7980
rect 114100 7924 117404 7980
rect 118570 7924 118580 7980
rect 118636 7924 120596 7980
rect 120652 7924 120662 7980
rect 120922 7924 120932 7980
rect 120988 7924 131628 7980
rect 132458 7924 132468 7980
rect 132524 7924 134484 7980
rect 134540 7924 134550 7980
rect 134810 7924 134820 7980
rect 134876 7924 141204 7980
rect 141260 7924 141270 7980
rect 141866 7924 141876 7980
rect 141932 7924 142996 7980
rect 143052 7924 143062 7980
rect 144218 7924 144228 7980
rect 144284 7924 147700 7980
rect 147756 7924 147766 7980
rect 147914 7924 147924 7980
rect 147980 7924 150388 7980
rect 150444 7924 150454 7980
rect 156211 7924 162932 7980
rect 162988 7924 162998 7980
rect 166394 7924 166404 7980
rect 166460 7924 166964 7980
rect 167020 7924 167030 7980
rect 172218 7924 172228 7980
rect 172284 7924 175980 7980
rect 179731 7924 193060 7980
rect 193116 7924 193126 7980
rect 194292 7924 203307 7980
rect 203634 7924 203644 7980
rect 203756 7924 203766 7980
rect 203914 7924 203924 7980
rect 203980 7924 213612 7980
rect 213668 7924 213678 7980
rect 308 7756 364 7924
rect 90132 7868 90188 7924
rect 114100 7868 114156 7924
rect 117348 7868 117404 7924
rect 131572 7868 131628 7924
rect 179731 7868 179787 7924
rect 55530 7812 55540 7868
rect 55596 7812 55644 7868
rect 55700 7812 55748 7868
rect 55804 7812 55814 7868
rect 58426 7812 58436 7868
rect 58492 7812 60452 7868
rect 60508 7812 88396 7868
rect 88452 7812 88462 7868
rect 88564 7812 90188 7868
rect 90458 7812 90468 7868
rect 90524 7812 99204 7868
rect 99260 7812 99270 7868
rect 99866 7812 99876 7868
rect 99932 7812 102900 7868
rect 102956 7812 102966 7868
rect 103338 7812 103348 7868
rect 103404 7812 104132 7868
rect 104188 7812 104198 7868
rect 108266 7812 108276 7868
rect 108332 7812 109788 7868
rect 109858 7812 109868 7868
rect 109924 7812 109972 7868
rect 110028 7812 110076 7868
rect 110132 7812 110142 7868
rect 110292 7812 113652 7868
rect 113708 7812 113718 7868
rect 113876 7812 114156 7868
rect 114314 7812 114324 7868
rect 114380 7812 116676 7868
rect 116732 7812 116742 7868
rect 116890 7812 116900 7868
rect 116956 7812 117124 7868
rect 117180 7812 117190 7868
rect 117348 7812 119476 7868
rect 119532 7812 119542 7868
rect 119914 7812 119924 7868
rect 119980 7812 127204 7868
rect 127260 7812 127270 7868
rect 128426 7812 128436 7868
rect 128492 7812 129052 7868
rect 129108 7812 129118 7868
rect 129210 7812 129220 7868
rect 129276 7812 131067 7868
rect 131572 7812 137956 7868
rect 138012 7812 138022 7868
rect 138628 7812 148708 7868
rect 148764 7812 148774 7868
rect 149370 7812 149380 7868
rect 149436 7812 157780 7868
rect 157836 7812 157846 7868
rect 158004 7812 163268 7868
rect 163324 7812 163334 7868
rect 164186 7812 164196 7868
rect 164252 7812 164300 7868
rect 164356 7812 164404 7868
rect 164460 7812 164470 7868
rect 166282 7812 166292 7868
rect 166348 7812 174412 7868
rect 174794 7812 174804 7868
rect 174860 7812 179787 7868
rect 181066 7812 181076 7868
rect 181132 7812 184996 7868
rect 185052 7812 185062 7868
rect 187338 7812 187348 7868
rect 187404 7812 200564 7868
rect 200620 7812 200630 7868
rect 203251 7812 208404 7868
rect 208460 7812 208470 7868
rect 210970 7812 210980 7868
rect 211036 7812 212716 7868
rect 212772 7812 212782 7868
rect 88564 7756 88620 7812
rect 109732 7756 109788 7812
rect 110292 7756 110348 7812
rect 113876 7756 113932 7812
rect 131011 7756 131067 7812
rect 138628 7756 138684 7812
rect 158004 7756 158060 7812
rect 308 7700 924 7756
rect 21466 7700 21476 7756
rect 21532 7700 56868 7756
rect 56924 7700 56934 7756
rect 57530 7700 57540 7756
rect 57596 7700 58324 7756
rect 58380 7700 58390 7756
rect 58650 7700 58660 7756
rect 58716 7700 59332 7756
rect 59388 7700 60788 7756
rect 60844 7700 60854 7756
rect 62906 7700 62916 7756
rect 62972 7700 63420 7756
rect 63476 7700 66724 7756
rect 66780 7700 66790 7756
rect 67050 7700 67060 7756
rect 67116 7700 67900 7756
rect 67956 7700 68964 7756
rect 69020 7700 69030 7756
rect 69514 7700 69524 7756
rect 69580 7700 85708 7756
rect 85764 7700 85774 7756
rect 85866 7700 85876 7756
rect 85932 7700 88004 7756
rect 88060 7700 88070 7756
rect 88228 7700 88620 7756
rect 90346 7700 90356 7756
rect 90412 7700 91532 7756
rect 91588 7700 91598 7756
rect 91690 7700 91700 7756
rect 91756 7700 109508 7756
rect 109564 7700 109574 7756
rect 109732 7700 110348 7756
rect 111066 7700 111076 7756
rect 111132 7700 113932 7756
rect 114090 7700 114100 7756
rect 114156 7700 114324 7756
rect 114380 7700 114390 7756
rect 114762 7700 114772 7756
rect 114828 7700 115108 7756
rect 115164 7700 115174 7756
rect 115322 7700 115332 7756
rect 115388 7700 120036 7756
rect 120092 7700 120102 7756
rect 120250 7700 120260 7756
rect 120316 7700 126868 7756
rect 126924 7700 126934 7756
rect 127082 7700 127092 7756
rect 127148 7700 128436 7756
rect 128492 7700 128502 7756
rect 129434 7700 129444 7756
rect 129500 7700 130396 7756
rect 130452 7700 130462 7756
rect 131011 7700 132804 7756
rect 132860 7700 132870 7756
rect 133354 7700 133364 7756
rect 133420 7700 136220 7756
rect 136826 7700 136836 7756
rect 136892 7700 138684 7756
rect 141194 7700 141204 7756
rect 141260 7700 142548 7756
rect 142604 7700 142614 7756
rect 142762 7700 142772 7756
rect 142828 7700 154196 7756
rect 154252 7700 154262 7756
rect 155978 7700 155988 7756
rect 156044 7700 156548 7756
rect 156604 7700 156614 7756
rect 156884 7700 158060 7756
rect 162586 7700 162596 7756
rect 162652 7700 167860 7756
rect 167916 7700 167926 7756
rect 0 7532 800 7560
rect 868 7532 924 7700
rect 88228 7644 88284 7700
rect 136164 7644 136220 7700
rect 156884 7644 156940 7700
rect 174356 7644 174412 7812
rect 203251 7756 203307 7812
rect 177678 7700 177716 7756
rect 177772 7700 177782 7756
rect 182942 7700 182980 7756
rect 183036 7700 183046 7756
rect 188906 7700 188916 7756
rect 188972 7700 190820 7756
rect 190876 7700 190886 7756
rect 191706 7700 191716 7756
rect 191772 7700 196028 7756
rect 196084 7700 196094 7756
rect 196410 7700 196420 7756
rect 196476 7700 203307 7756
rect 207498 7700 207508 7756
rect 207564 7700 214396 7756
rect 214452 7700 214462 7756
rect 8922 7588 8932 7644
rect 8988 7588 9548 7644
rect 9604 7588 20187 7644
rect 42158 7588 42196 7644
rect 42252 7588 42262 7644
rect 46190 7588 46228 7644
rect 46284 7588 46294 7644
rect 47114 7588 47124 7644
rect 47180 7588 62580 7644
rect 62636 7588 62646 7644
rect 63802 7588 63812 7644
rect 63868 7588 71764 7644
rect 71820 7588 71830 7644
rect 71978 7588 71988 7644
rect 72044 7588 74116 7644
rect 74172 7588 74182 7644
rect 74330 7588 74340 7644
rect 74396 7588 79436 7644
rect 79492 7588 79502 7644
rect 79706 7588 79716 7644
rect 79772 7588 83076 7644
rect 83132 7588 83142 7644
rect 83290 7588 83300 7644
rect 83356 7588 83972 7644
rect 84028 7588 84038 7644
rect 84410 7588 84420 7644
rect 84476 7588 86100 7644
rect 86156 7588 86166 7644
rect 86426 7588 86436 7644
rect 86492 7588 88284 7644
rect 88666 7588 88676 7644
rect 88732 7588 91812 7644
rect 91868 7588 91878 7644
rect 95610 7588 95620 7644
rect 95676 7588 106148 7644
rect 106204 7588 106214 7644
rect 106362 7588 106372 7644
rect 106428 7588 113204 7644
rect 113260 7588 113270 7644
rect 113754 7588 113764 7644
rect 113820 7588 115220 7644
rect 115276 7588 115286 7644
rect 115546 7588 115556 7644
rect 115612 7588 115948 7644
rect 116004 7588 117628 7644
rect 117786 7588 117796 7644
rect 117852 7588 118692 7644
rect 118748 7588 118758 7644
rect 119018 7588 119028 7644
rect 119084 7588 119364 7644
rect 119420 7588 119430 7644
rect 119690 7588 119700 7644
rect 119756 7588 134260 7644
rect 134316 7588 134326 7644
rect 134586 7588 134596 7644
rect 134652 7588 135996 7644
rect 136052 7588 136062 7644
rect 136164 7588 139524 7644
rect 139580 7588 139590 7644
rect 139738 7588 139748 7644
rect 139804 7588 143556 7644
rect 143612 7588 143622 7644
rect 143714 7588 143724 7644
rect 143780 7588 144228 7644
rect 144284 7588 144294 7644
rect 144778 7588 144788 7644
rect 144844 7588 146916 7644
rect 146972 7588 146982 7644
rect 147140 7588 148820 7644
rect 148876 7588 148886 7644
rect 149034 7588 149044 7644
rect 149100 7588 153300 7644
rect 153356 7588 153366 7644
rect 155978 7588 155988 7644
rect 156044 7588 156940 7644
rect 157098 7588 157108 7644
rect 157164 7588 158564 7644
rect 158620 7588 158630 7644
rect 159450 7588 159460 7644
rect 159516 7588 161364 7644
rect 161420 7588 161430 7644
rect 164266 7588 164276 7644
rect 164332 7588 167748 7644
rect 167804 7588 167814 7644
rect 174346 7588 174356 7644
rect 174412 7588 175980 7644
rect 176138 7588 176148 7644
rect 176204 7588 182532 7644
rect 182588 7588 182598 7644
rect 190810 7588 190820 7644
rect 190876 7588 190932 7644
rect 190988 7588 190998 7644
rect 192266 7588 192276 7644
rect 192332 7588 193788 7644
rect 193844 7588 193854 7644
rect 195122 7588 195132 7644
rect 195188 7588 196420 7644
rect 196476 7588 196486 7644
rect 196634 7588 196644 7644
rect 196700 7588 196924 7644
rect 196980 7588 196990 7644
rect 209850 7588 209860 7644
rect 209916 7588 215292 7644
rect 215348 7588 215358 7644
rect 20131 7532 20187 7588
rect 117572 7532 117628 7588
rect 147140 7532 147196 7588
rect 175924 7532 175980 7588
rect 0 7476 924 7532
rect 12730 7476 12740 7532
rect 12796 7476 13748 7532
rect 13804 7476 13814 7532
rect 20131 7476 68348 7532
rect 68404 7476 68414 7532
rect 68506 7476 68516 7532
rect 68572 7476 71148 7532
rect 71306 7476 71316 7532
rect 71372 7476 73892 7532
rect 73948 7476 73958 7532
rect 74452 7476 75236 7532
rect 75338 7476 75348 7532
rect 75404 7476 78260 7532
rect 78316 7476 78326 7532
rect 78474 7476 78484 7532
rect 78540 7476 85036 7532
rect 86090 7476 86100 7532
rect 86156 7476 86884 7532
rect 86940 7476 86950 7532
rect 88106 7476 88116 7532
rect 88172 7476 91028 7532
rect 91084 7476 91094 7532
rect 91242 7476 91252 7532
rect 91308 7476 99876 7532
rect 99932 7476 99942 7532
rect 100090 7476 100100 7532
rect 100156 7476 103460 7532
rect 103516 7476 103526 7532
rect 104122 7476 104132 7532
rect 104188 7476 104972 7532
rect 105028 7476 105038 7532
rect 105130 7476 105140 7532
rect 105196 7476 117348 7532
rect 117404 7476 117414 7532
rect 117572 7476 118020 7532
rect 118076 7476 118086 7532
rect 118234 7476 118244 7532
rect 118300 7476 125412 7532
rect 125468 7476 125478 7532
rect 127082 7476 127092 7532
rect 127148 7476 133644 7532
rect 133802 7476 133812 7532
rect 133868 7476 146020 7532
rect 146076 7476 146086 7532
rect 146234 7476 146244 7532
rect 146300 7476 147196 7532
rect 147550 7476 147588 7532
rect 147644 7476 147654 7532
rect 147914 7476 147924 7532
rect 147980 7476 149996 7532
rect 150052 7476 150062 7532
rect 150154 7476 150164 7532
rect 150220 7476 150724 7532
rect 150780 7476 150790 7532
rect 152730 7476 152740 7532
rect 152796 7476 161476 7532
rect 161532 7476 161542 7532
rect 163594 7476 163604 7532
rect 163660 7476 165452 7532
rect 167850 7476 167860 7532
rect 167916 7476 175756 7532
rect 175812 7476 175822 7532
rect 175924 7476 192836 7532
rect 192892 7476 192902 7532
rect 197988 7476 199612 7532
rect 199668 7476 199678 7532
rect 199770 7476 199780 7532
rect 199836 7476 203924 7532
rect 203980 7476 203990 7532
rect 206042 7476 206052 7532
rect 206108 7476 213948 7532
rect 214004 7476 214014 7532
rect 0 7448 800 7476
rect 10322 7364 10332 7420
rect 10388 7364 10948 7420
rect 11004 7364 11014 7420
rect 15866 7364 15876 7420
rect 15932 7364 18060 7420
rect 18116 7364 18228 7420
rect 18284 7364 18294 7420
rect 18610 7364 18620 7420
rect 18676 7364 59780 7420
rect 59836 7364 59846 7420
rect 59994 7364 60004 7420
rect 60060 7364 62804 7420
rect 62860 7364 62870 7420
rect 63018 7364 63028 7420
rect 63084 7364 63868 7420
rect 63924 7364 63934 7420
rect 64586 7364 64596 7420
rect 64652 7364 67956 7420
rect 68012 7364 68022 7420
rect 68114 7364 68124 7420
rect 68180 7364 70868 7420
rect 70924 7364 70934 7420
rect 71092 7308 71148 7476
rect 74452 7420 74508 7476
rect 75180 7420 75236 7476
rect 84980 7420 85036 7476
rect 133588 7420 133644 7476
rect 165396 7420 165452 7476
rect 197988 7420 198044 7476
rect 71418 7364 71428 7420
rect 71484 7364 74508 7420
rect 74666 7364 74676 7420
rect 74732 7364 75012 7420
rect 75068 7364 75078 7420
rect 75180 7364 75796 7420
rect 75852 7364 75862 7420
rect 76066 7364 76076 7420
rect 76132 7364 80052 7420
rect 80108 7364 80118 7420
rect 80266 7364 80276 7420
rect 80332 7364 83748 7420
rect 83804 7364 84756 7420
rect 84812 7364 84822 7420
rect 84980 7364 91476 7420
rect 91532 7364 91542 7420
rect 91690 7364 91700 7420
rect 91756 7364 97524 7420
rect 97580 7364 97590 7420
rect 97682 7364 97692 7420
rect 97804 7364 99092 7420
rect 99148 7364 99158 7420
rect 99418 7364 99428 7420
rect 99484 7364 102340 7420
rect 102396 7364 102406 7420
rect 102666 7364 102676 7420
rect 102732 7364 103628 7420
rect 103786 7364 103796 7420
rect 103852 7364 115052 7420
rect 115210 7364 115220 7420
rect 115276 7364 118468 7420
rect 118524 7364 118534 7420
rect 118906 7364 118916 7420
rect 118972 7364 119700 7420
rect 119756 7364 119766 7420
rect 119914 7364 119924 7420
rect 119980 7364 121324 7420
rect 121380 7364 121390 7420
rect 121594 7364 121604 7420
rect 121660 7364 121716 7420
rect 121772 7364 122836 7420
rect 122892 7364 122902 7420
rect 123060 7364 127876 7420
rect 127932 7364 127942 7420
rect 128258 7364 128268 7420
rect 128324 7364 130228 7420
rect 130284 7364 130294 7420
rect 130442 7364 130452 7420
rect 130508 7364 133364 7420
rect 133420 7364 133430 7420
rect 133588 7364 138180 7420
rect 138236 7364 138246 7420
rect 140410 7364 140420 7420
rect 140476 7364 142156 7420
rect 142426 7364 142436 7420
rect 142492 7364 144956 7420
rect 145562 7364 145572 7420
rect 145628 7364 149268 7420
rect 149324 7364 149334 7420
rect 149594 7364 149604 7420
rect 149660 7364 154084 7420
rect 154140 7364 154150 7420
rect 154410 7364 154420 7420
rect 154476 7364 164836 7420
rect 164892 7364 164902 7420
rect 165396 7364 182980 7420
rect 183036 7364 183046 7420
rect 190586 7364 190596 7420
rect 190652 7364 198044 7420
rect 198202 7364 198212 7420
rect 198268 7364 199164 7420
rect 199220 7364 199230 7420
rect 201562 7364 201572 7420
rect 201628 7364 202636 7420
rect 202692 7364 202702 7420
rect 203522 7364 203532 7420
rect 203588 7364 203924 7420
rect 203980 7364 210980 7420
rect 211036 7364 211046 7420
rect 211184 7364 211204 7420
rect 211316 7364 212324 7420
rect 212380 7364 212390 7420
rect 214386 7364 214396 7420
rect 214508 7364 214518 7420
rect 103572 7308 103628 7364
rect 114996 7308 115052 7364
rect 123060 7308 123116 7364
rect 142100 7308 142156 7364
rect 144900 7308 144956 7364
rect 7914 7252 7924 7308
rect 7980 7252 8764 7308
rect 8820 7252 8830 7308
rect 16874 7252 16884 7308
rect 16940 7252 17612 7308
rect 17668 7252 58044 7308
rect 58100 7252 58110 7308
rect 58314 7252 58324 7308
rect 58380 7252 60900 7308
rect 60956 7252 60966 7308
rect 62346 7252 62356 7308
rect 62412 7252 69524 7308
rect 69580 7252 69590 7308
rect 69738 7252 69748 7308
rect 69804 7252 70587 7308
rect 71092 7252 71988 7308
rect 72044 7252 72054 7308
rect 72314 7252 72324 7308
rect 72380 7252 73892 7308
rect 73948 7252 73958 7308
rect 74554 7252 74564 7308
rect 74620 7252 75628 7308
rect 75684 7252 75694 7308
rect 75898 7252 75908 7308
rect 75964 7252 77924 7308
rect 77980 7252 77990 7308
rect 78138 7252 78148 7308
rect 78204 7252 78708 7308
rect 78764 7252 78774 7308
rect 78866 7252 78876 7308
rect 78988 7252 80164 7308
rect 80220 7252 80230 7308
rect 80490 7252 80500 7308
rect 80556 7252 80948 7308
rect 81004 7252 81014 7308
rect 81162 7252 81172 7308
rect 81228 7252 81266 7308
rect 81386 7252 81396 7308
rect 81452 7252 84027 7308
rect 84186 7252 84196 7308
rect 84252 7252 84420 7308
rect 84476 7252 84486 7308
rect 84858 7252 84868 7308
rect 84924 7252 85372 7308
rect 85428 7252 90244 7308
rect 90300 7252 90310 7308
rect 90458 7252 90468 7308
rect 90524 7252 103348 7308
rect 103404 7252 103414 7308
rect 103572 7252 105700 7308
rect 105756 7252 105766 7308
rect 106138 7252 106148 7308
rect 106204 7252 114324 7308
rect 114380 7252 114390 7308
rect 114996 7252 121044 7308
rect 121100 7252 121110 7308
rect 121258 7252 121268 7308
rect 121324 7252 121940 7308
rect 121996 7252 122006 7308
rect 122266 7252 122276 7308
rect 122332 7252 123116 7308
rect 125402 7252 125412 7308
rect 125468 7252 126812 7308
rect 126970 7252 126980 7308
rect 127036 7252 141876 7308
rect 141932 7252 141942 7308
rect 142100 7252 144676 7308
rect 144732 7252 144742 7308
rect 144900 7252 150052 7308
rect 150108 7252 150118 7308
rect 155418 7252 155428 7308
rect 155484 7252 160524 7308
rect 162922 7252 162932 7308
rect 162988 7252 168868 7308
rect 168924 7252 168934 7308
rect 172890 7252 172900 7308
rect 172956 7252 177940 7308
rect 177996 7252 178006 7308
rect 180170 7252 180180 7308
rect 180236 7252 191660 7308
rect 191716 7252 191726 7308
rect 193610 7252 193620 7308
rect 193676 7252 200004 7308
rect 200060 7252 200070 7308
rect 70531 7196 70587 7252
rect 83971 7196 84027 7252
rect 126756 7196 126812 7252
rect 160468 7196 160524 7252
rect 23034 7140 23044 7196
rect 23100 7140 25564 7196
rect 25676 7140 25686 7196
rect 28186 7140 28196 7196
rect 28252 7140 30604 7196
rect 30716 7140 30726 7196
rect 34010 7140 34020 7196
rect 34076 7140 34524 7196
rect 34636 7140 34646 7196
rect 44594 7140 44604 7196
rect 44716 7140 44726 7196
rect 50371 7140 69860 7196
rect 69916 7140 69926 7196
rect 70531 7140 72100 7196
rect 72156 7140 72166 7196
rect 72314 7140 72324 7196
rect 72380 7140 74788 7196
rect 74844 7140 74854 7196
rect 75002 7140 75012 7196
rect 75068 7140 76132 7196
rect 76188 7140 76198 7196
rect 76290 7140 76300 7196
rect 76356 7140 82292 7196
rect 82348 7140 82358 7196
rect 82506 7140 82516 7196
rect 82572 7140 83412 7196
rect 83468 7140 83478 7196
rect 83626 7140 83636 7196
rect 83692 7140 83730 7196
rect 83971 7140 91252 7196
rect 91308 7140 91318 7196
rect 91466 7140 91476 7196
rect 91532 7140 91588 7196
rect 91644 7140 91756 7196
rect 91812 7140 91822 7196
rect 91914 7140 91924 7196
rect 91980 7140 96852 7196
rect 96908 7140 96918 7196
rect 100426 7140 100436 7196
rect 100492 7140 100772 7196
rect 100828 7140 100838 7196
rect 100986 7140 100996 7196
rect 101052 7140 102004 7196
rect 102060 7140 102070 7196
rect 102218 7140 102228 7196
rect 102284 7140 103012 7196
rect 103068 7140 103078 7196
rect 103338 7140 103348 7196
rect 103404 7140 103908 7196
rect 103964 7140 103974 7196
rect 104122 7140 104132 7196
rect 104188 7140 115220 7196
rect 115276 7140 115286 7196
rect 115434 7140 115444 7196
rect 115500 7140 117460 7196
rect 117516 7140 117526 7196
rect 117674 7140 117684 7196
rect 117740 7140 121828 7196
rect 121884 7140 121894 7196
rect 122490 7140 122500 7196
rect 122556 7140 126084 7196
rect 126140 7140 126150 7196
rect 126756 7140 139860 7196
rect 139916 7140 139926 7196
rect 140522 7140 140532 7196
rect 140588 7140 142436 7196
rect 142492 7140 142502 7196
rect 142650 7140 142660 7196
rect 142716 7140 153748 7196
rect 153804 7140 153814 7196
rect 153972 7140 159460 7196
rect 159516 7140 159526 7196
rect 160468 7140 164612 7196
rect 164668 7140 164678 7196
rect 164826 7140 164836 7196
rect 164892 7140 180684 7196
rect 180740 7140 180750 7196
rect 182970 7140 182980 7196
rect 183036 7140 197820 7196
rect 197876 7140 197886 7196
rect 207722 7140 207732 7196
rect 207788 7140 210700 7196
rect 210756 7140 210766 7196
rect 50371 7084 50427 7140
rect 153972 7084 154028 7140
rect 28366 7028 28376 7084
rect 28432 7028 28480 7084
rect 28536 7028 28584 7084
rect 28640 7028 28650 7084
rect 38714 7028 38724 7084
rect 38780 7028 39788 7084
rect 39844 7028 50427 7084
rect 52658 7028 52668 7084
rect 52724 7028 79268 7084
rect 79324 7028 79334 7084
rect 79818 7028 79828 7084
rect 79884 7028 82460 7084
rect 82694 7028 82704 7084
rect 82760 7028 82808 7084
rect 82864 7028 82912 7084
rect 82968 7028 82978 7084
rect 83188 7028 84644 7084
rect 84700 7028 84710 7084
rect 84970 7028 84980 7084
rect 85036 7028 85764 7084
rect 85820 7028 85830 7084
rect 85978 7028 85988 7084
rect 86044 7028 87780 7084
rect 87836 7028 87846 7084
rect 87994 7028 88004 7084
rect 88060 7028 89404 7084
rect 90234 7028 90244 7084
rect 90300 7028 91252 7084
rect 91308 7028 91318 7084
rect 91466 7028 91476 7084
rect 91532 7028 103796 7084
rect 103852 7028 103862 7084
rect 104010 7028 104020 7084
rect 104076 7028 110852 7084
rect 110908 7028 110918 7084
rect 111626 7028 111636 7084
rect 111692 7028 120652 7084
rect 121146 7028 121156 7084
rect 121212 7028 121324 7084
rect 121380 7028 121390 7084
rect 121930 7028 121940 7084
rect 121996 7028 122948 7084
rect 123004 7028 123014 7084
rect 123274 7028 123284 7084
rect 123340 7028 127092 7084
rect 127148 7028 127158 7084
rect 129322 7028 129332 7084
rect 129388 7028 136836 7084
rect 136892 7028 136902 7084
rect 137022 7028 137032 7084
rect 137088 7028 137136 7084
rect 137192 7028 137240 7084
rect 137296 7028 137306 7084
rect 137498 7028 137508 7084
rect 137564 7028 144452 7084
rect 144508 7028 144518 7084
rect 144666 7028 144676 7084
rect 144732 7028 149044 7084
rect 149100 7028 149110 7084
rect 149482 7028 149492 7084
rect 149548 7028 154028 7084
rect 154186 7028 154196 7084
rect 154252 7028 169540 7084
rect 169596 7028 169606 7084
rect 173898 7028 173908 7084
rect 173964 7028 186564 7084
rect 186620 7028 186630 7084
rect 186778 7028 186788 7084
rect 186844 7028 188860 7084
rect 191350 7028 191360 7084
rect 191416 7028 191464 7084
rect 191520 7028 191568 7084
rect 191624 7028 191634 7084
rect 197530 7028 197540 7084
rect 197596 7028 214116 7084
rect 214172 7028 214182 7084
rect 82404 6972 82460 7028
rect 83188 6972 83244 7028
rect 89348 6972 89404 7028
rect 120596 6972 120652 7028
rect 188804 6972 188860 7028
rect 30594 6916 30604 6972
rect 30660 6916 67452 6972
rect 67946 6916 67956 6972
rect 68012 6916 69020 6972
rect 70522 6916 70532 6972
rect 70588 6916 75348 6972
rect 75404 6916 75414 6972
rect 75618 6916 75628 6972
rect 75684 6916 78148 6972
rect 78204 6916 78214 6972
rect 78316 6916 80052 6972
rect 80108 6916 80118 6972
rect 80378 6916 80388 6972
rect 80444 6916 82068 6972
rect 82124 6916 82134 6972
rect 82404 6916 83244 6972
rect 83402 6916 83412 6972
rect 83468 6916 83524 6972
rect 83580 6916 83590 6972
rect 84298 6916 84308 6972
rect 84364 6916 87444 6972
rect 87500 6916 87510 6972
rect 87658 6916 87668 6972
rect 87724 6916 88340 6972
rect 88396 6916 88406 6972
rect 88554 6916 88564 6972
rect 88620 6916 89124 6972
rect 89180 6916 89190 6972
rect 89348 6916 90580 6972
rect 90636 6916 90646 6972
rect 90738 6916 90748 6972
rect 90804 6916 91252 6972
rect 91308 6916 91318 6972
rect 91466 6916 91476 6972
rect 91532 6916 99316 6972
rect 99372 6916 99382 6972
rect 99530 6916 99540 6972
rect 99596 6916 100100 6972
rect 100156 6916 100166 6972
rect 100314 6916 100324 6972
rect 100380 6916 102788 6972
rect 102844 6916 102854 6972
rect 103002 6916 103012 6972
rect 103068 6916 105140 6972
rect 105196 6916 105206 6972
rect 105364 6916 106932 6972
rect 106988 6916 106998 6972
rect 107818 6916 107828 6972
rect 107884 6916 109172 6972
rect 109228 6916 109238 6972
rect 109386 6916 109396 6972
rect 109452 6916 120372 6972
rect 120428 6916 120438 6972
rect 120596 6916 122500 6972
rect 122556 6916 122566 6972
rect 122714 6916 122724 6972
rect 122780 6916 130452 6972
rect 130508 6916 130518 6972
rect 132570 6916 132580 6972
rect 132636 6916 134260 6972
rect 134316 6916 134326 6972
rect 135930 6916 135940 6972
rect 135996 6916 136108 6972
rect 136164 6916 136500 6972
rect 136556 6916 137620 6972
rect 137676 6916 137686 6972
rect 138170 6916 138180 6972
rect 138236 6916 142660 6972
rect 142716 6916 142726 6972
rect 142986 6916 142996 6972
rect 143052 6916 147812 6972
rect 147868 6916 147878 6972
rect 148810 6916 148820 6972
rect 148876 6916 149940 6972
rect 149996 6916 150006 6972
rect 152170 6916 152180 6972
rect 152236 6916 174804 6972
rect 174860 6916 174870 6972
rect 178826 6916 178836 6972
rect 178892 6916 186452 6972
rect 186508 6916 186518 6972
rect 187002 6916 187012 6972
rect 187068 6916 188748 6972
rect 188804 6916 193732 6972
rect 193788 6916 193798 6972
rect 195738 6916 195748 6972
rect 195804 6916 198324 6972
rect 198380 6916 203307 6972
rect 21690 6804 21700 6860
rect 21756 6804 48356 6860
rect 48412 6804 48422 6860
rect 51594 6804 51604 6860
rect 51660 6804 52556 6860
rect 52612 6804 52622 6860
rect 56746 6804 56756 6860
rect 56812 6804 58604 6860
rect 58660 6804 58670 6860
rect 58884 6804 62244 6860
rect 62300 6804 62310 6860
rect 62468 6804 66276 6860
rect 66332 6804 66342 6860
rect 66714 6804 66724 6860
rect 66780 6804 67172 6860
rect 67228 6804 67238 6860
rect 58884 6748 58940 6804
rect 62468 6748 62524 6804
rect 67396 6748 67452 6916
rect 67890 6804 67900 6860
rect 67956 6804 68740 6860
rect 68796 6804 68806 6860
rect 68964 6748 69020 6916
rect 78316 6860 78372 6916
rect 105364 6860 105420 6916
rect 188692 6860 188748 6916
rect 203251 6860 203307 6916
rect 69178 6804 69188 6860
rect 69244 6804 70140 6860
rect 70196 6804 74900 6860
rect 74956 6804 74966 6860
rect 75058 6804 75068 6860
rect 75124 6804 76020 6860
rect 76076 6804 76086 6860
rect 76234 6804 76244 6860
rect 76300 6804 78372 6860
rect 78586 6804 78596 6860
rect 78652 6804 79828 6860
rect 79884 6804 79894 6860
rect 80042 6804 80052 6860
rect 80108 6804 82180 6860
rect 82236 6804 82246 6860
rect 82618 6804 82628 6860
rect 82684 6804 84027 6860
rect 84186 6804 84196 6860
rect 84252 6804 86212 6860
rect 86268 6804 86278 6860
rect 86650 6804 86660 6860
rect 86716 6804 91588 6860
rect 91802 6804 91812 6860
rect 91868 6804 103628 6860
rect 103786 6804 103796 6860
rect 103852 6804 105420 6860
rect 105690 6804 105700 6860
rect 105756 6804 109508 6860
rect 109564 6804 109574 6860
rect 110170 6804 110180 6860
rect 110236 6804 111300 6860
rect 111356 6804 111366 6860
rect 112074 6804 112084 6860
rect 112140 6804 114212 6860
rect 114314 6804 114324 6860
rect 114380 6804 114660 6860
rect 114716 6804 114726 6860
rect 115098 6804 115108 6860
rect 115164 6804 115332 6860
rect 115388 6804 115398 6860
rect 115658 6804 115668 6860
rect 115724 6804 116564 6860
rect 116620 6804 116630 6860
rect 116788 6804 117124 6860
rect 117180 6804 117190 6860
rect 117450 6804 117460 6860
rect 117516 6804 134820 6860
rect 134876 6804 134886 6860
rect 135828 6804 139412 6860
rect 139468 6804 139478 6860
rect 139850 6804 139860 6860
rect 139916 6804 141764 6860
rect 141820 6804 141830 6860
rect 143210 6804 143220 6860
rect 143276 6804 143556 6860
rect 143612 6804 143622 6860
rect 143770 6804 143780 6860
rect 143836 6804 144564 6860
rect 144620 6804 144630 6860
rect 145114 6804 145124 6860
rect 145180 6804 145796 6860
rect 145852 6804 145862 6860
rect 147634 6804 147644 6860
rect 147700 6804 149156 6860
rect 149212 6804 149222 6860
rect 150276 6804 157108 6860
rect 157164 6804 157174 6860
rect 157322 6804 157332 6860
rect 157388 6804 176148 6860
rect 176204 6804 176214 6860
rect 179731 6804 181188 6860
rect 181244 6804 181254 6860
rect 182606 6804 182644 6860
rect 182700 6804 182710 6860
rect 185210 6804 185220 6860
rect 185276 6804 188468 6860
rect 188524 6804 188534 6860
rect 188692 6804 200788 6860
rect 200844 6804 200854 6860
rect 203251 6804 213108 6860
rect 213164 6804 213174 6860
rect 83971 6748 84027 6804
rect 91532 6748 91588 6804
rect 20010 6692 20020 6748
rect 20076 6692 21476 6748
rect 21532 6692 21542 6748
rect 43418 6692 43428 6748
rect 43484 6692 43932 6748
rect 43988 6692 43998 6748
rect 47394 6692 47404 6748
rect 47460 6692 49028 6748
rect 49084 6692 49094 6748
rect 51762 6692 51772 6748
rect 51828 6692 52164 6748
rect 52220 6692 52230 6748
rect 56970 6692 56980 6748
rect 57036 6692 58940 6748
rect 60452 6692 62524 6748
rect 62682 6692 62692 6748
rect 62748 6692 64148 6748
rect 64204 6692 64214 6748
rect 65818 6692 65828 6748
rect 65884 6692 67060 6748
rect 67116 6692 67126 6748
rect 67396 6692 68852 6748
rect 68964 6692 73668 6748
rect 73724 6692 73734 6748
rect 73891 6692 79100 6748
rect 79230 6692 79268 6748
rect 79324 6692 79334 6748
rect 79482 6692 79492 6748
rect 79548 6692 80388 6748
rect 80444 6692 80454 6748
rect 80602 6692 80612 6748
rect 80668 6692 82516 6748
rect 82572 6692 82582 6748
rect 82730 6692 82740 6748
rect 82796 6692 83748 6748
rect 83804 6692 83814 6748
rect 83971 6692 84532 6748
rect 84634 6692 84644 6748
rect 84700 6692 86884 6748
rect 86940 6692 86950 6748
rect 87098 6692 87108 6748
rect 87164 6692 87556 6748
rect 87612 6692 87622 6748
rect 87770 6692 87780 6748
rect 87836 6692 91364 6748
rect 91420 6692 91430 6748
rect 91532 6692 103236 6748
rect 103292 6692 103302 6748
rect 60452 6636 60508 6692
rect 68796 6636 68852 6692
rect 73891 6636 73947 6692
rect 79044 6636 79100 6692
rect 84476 6636 84532 6692
rect 103572 6636 103628 6804
rect 114156 6748 114212 6804
rect 116788 6748 116844 6804
rect 135828 6748 135884 6804
rect 150276 6748 150332 6804
rect 179731 6748 179787 6804
rect 104010 6692 104020 6748
rect 104076 6692 113988 6748
rect 114044 6692 114054 6748
rect 114156 6692 115556 6748
rect 115612 6692 115622 6748
rect 115770 6692 115780 6748
rect 115836 6692 116844 6748
rect 117002 6692 117012 6748
rect 117068 6692 117124 6748
rect 117180 6692 117190 6748
rect 117338 6692 117348 6748
rect 117404 6692 117796 6748
rect 117852 6692 117862 6748
rect 118122 6692 118132 6748
rect 118188 6692 118412 6748
rect 118468 6692 122276 6748
rect 122332 6692 122342 6748
rect 122490 6692 122500 6748
rect 122556 6692 129836 6748
rect 130778 6692 130788 6748
rect 130844 6692 135884 6748
rect 135940 6692 139468 6748
rect 140634 6692 140644 6748
rect 140700 6692 141316 6748
rect 141372 6692 141382 6748
rect 142772 6692 150332 6748
rect 150490 6692 150500 6748
rect 150556 6692 152907 6748
rect 153066 6692 153076 6748
rect 153132 6692 154700 6748
rect 155306 6692 155316 6748
rect 155372 6692 179787 6748
rect 181290 6692 181300 6748
rect 181356 6692 186900 6748
rect 186956 6692 186966 6748
rect 188234 6692 188244 6748
rect 188300 6692 190596 6748
rect 190652 6692 190662 6748
rect 191706 6692 191716 6748
rect 191828 6692 191838 6748
rect 194842 6692 194852 6748
rect 194908 6692 196420 6748
rect 196476 6692 196486 6748
rect 196634 6692 196644 6748
rect 196700 6692 198772 6748
rect 198828 6692 199780 6748
rect 199836 6692 199846 6748
rect 199994 6692 200004 6748
rect 200060 6692 211876 6748
rect 211932 6692 211942 6748
rect 16650 6580 16660 6636
rect 16716 6580 19236 6636
rect 19292 6580 19302 6636
rect 28690 6580 28700 6636
rect 28812 6580 28822 6636
rect 37818 6580 37828 6636
rect 37884 6580 39004 6636
rect 39060 6580 39070 6636
rect 43306 6580 43316 6636
rect 43372 6580 43820 6636
rect 43876 6580 43886 6636
rect 53834 6580 53844 6636
rect 53900 6580 54964 6636
rect 55020 6580 56588 6636
rect 56644 6580 56654 6636
rect 56858 6580 56868 6636
rect 56924 6580 60508 6636
rect 60666 6580 60676 6636
rect 60732 6580 63700 6636
rect 63756 6580 63766 6636
rect 66836 6580 68628 6636
rect 68684 6580 68694 6636
rect 68796 6580 73947 6636
rect 75170 6580 75180 6636
rect 75236 6580 78820 6636
rect 78876 6580 78886 6636
rect 79044 6580 80836 6636
rect 80892 6580 80902 6636
rect 81172 6580 82516 6636
rect 82572 6580 82582 6636
rect 83066 6580 83076 6636
rect 83132 6580 84308 6636
rect 84364 6580 84374 6636
rect 84476 6580 85876 6636
rect 85932 6580 85942 6636
rect 86202 6580 86212 6636
rect 86268 6580 87668 6636
rect 87724 6580 87734 6636
rect 87994 6580 88004 6636
rect 88060 6580 90580 6636
rect 90636 6580 90646 6636
rect 90850 6580 90860 6636
rect 90916 6580 102116 6636
rect 102172 6580 102182 6636
rect 102330 6580 102340 6636
rect 102396 6580 103124 6636
rect 103180 6580 103190 6636
rect 103572 6580 108276 6636
rect 108332 6580 108342 6636
rect 108490 6580 108500 6636
rect 108556 6580 110068 6636
rect 110124 6580 110134 6636
rect 110282 6580 110292 6636
rect 110348 6580 113652 6636
rect 113708 6580 113718 6636
rect 113876 6580 115780 6636
rect 115836 6580 115846 6636
rect 116554 6580 116564 6636
rect 116620 6580 117460 6636
rect 117516 6580 117526 6636
rect 117674 6580 117684 6636
rect 117740 6580 122276 6636
rect 122332 6580 122342 6636
rect 122490 6580 122500 6636
rect 122556 6580 124740 6636
rect 124796 6580 124806 6636
rect 124954 6580 124964 6636
rect 125020 6580 127036 6636
rect 128258 6580 128268 6636
rect 128324 6580 128548 6636
rect 128604 6580 129556 6636
rect 129612 6580 129622 6636
rect 66836 6524 66892 6580
rect 81172 6524 81228 6580
rect 113876 6524 113932 6580
rect 126980 6524 127036 6580
rect 12842 6468 12852 6524
rect 12908 6468 14028 6524
rect 14084 6468 14094 6524
rect 20682 6468 20692 6524
rect 20748 6468 21532 6524
rect 21588 6468 21598 6524
rect 24602 6468 24612 6524
rect 24668 6468 37716 6524
rect 37772 6468 37782 6524
rect 43642 6468 43652 6524
rect 43708 6468 44380 6524
rect 44436 6468 44446 6524
rect 52546 6468 52556 6524
rect 52612 6468 56420 6524
rect 56476 6468 56486 6524
rect 58986 6468 58996 6524
rect 59052 6468 59948 6524
rect 60004 6468 66892 6524
rect 67050 6468 67060 6524
rect 67116 6468 75740 6524
rect 75796 6468 75806 6524
rect 76906 6468 76916 6524
rect 76972 6468 78092 6524
rect 78148 6468 81228 6524
rect 81834 6468 81844 6524
rect 81900 6468 82292 6524
rect 82348 6468 82358 6524
rect 82506 6468 82516 6524
rect 82572 6468 84084 6524
rect 84140 6468 84150 6524
rect 84298 6468 84308 6524
rect 84364 6468 90468 6524
rect 90524 6468 90534 6524
rect 90682 6468 90692 6524
rect 90748 6468 92820 6524
rect 92876 6468 92886 6524
rect 93258 6468 93268 6524
rect 93324 6468 95844 6524
rect 95900 6468 95910 6524
rect 96058 6468 96068 6524
rect 96124 6468 98644 6524
rect 98700 6468 98710 6524
rect 100202 6468 100212 6524
rect 100268 6468 101052 6524
rect 101164 6468 101174 6524
rect 101322 6468 101332 6524
rect 101388 6468 101612 6524
rect 101668 6468 103124 6524
rect 103180 6468 103190 6524
rect 103348 6468 104692 6524
rect 104748 6468 104758 6524
rect 105018 6468 105028 6524
rect 105084 6468 105364 6524
rect 105420 6468 105430 6524
rect 105690 6468 105700 6524
rect 105756 6468 111300 6524
rect 111356 6468 111366 6524
rect 112186 6468 112196 6524
rect 112252 6468 113932 6524
rect 114090 6468 114100 6524
rect 114156 6468 117236 6524
rect 117292 6468 117302 6524
rect 117786 6468 117796 6524
rect 117852 6468 118020 6524
rect 118076 6468 118086 6524
rect 118570 6468 118580 6524
rect 118636 6468 119140 6524
rect 119196 6468 119206 6524
rect 119354 6468 119364 6524
rect 119420 6468 122164 6524
rect 122220 6468 122230 6524
rect 122490 6468 122500 6524
rect 122556 6468 123564 6524
rect 123620 6468 123630 6524
rect 123834 6468 123844 6524
rect 123900 6468 126924 6524
rect 126980 6468 129220 6524
rect 129276 6468 129286 6524
rect 103348 6412 103404 6468
rect 4442 6356 4452 6412
rect 4508 6356 26404 6412
rect 26460 6356 26470 6412
rect 34682 6356 34692 6412
rect 34748 6356 35084 6412
rect 35140 6356 70588 6412
rect 70644 6356 70654 6412
rect 72090 6356 72100 6412
rect 72156 6356 75796 6412
rect 76010 6356 76020 6412
rect 76076 6356 78484 6412
rect 78540 6356 78550 6412
rect 78698 6356 78708 6412
rect 78764 6356 80276 6412
rect 80332 6356 80342 6412
rect 80490 6356 80500 6412
rect 80556 6356 81956 6412
rect 82012 6356 82022 6412
rect 82170 6356 82180 6412
rect 82236 6356 83860 6412
rect 83916 6356 83926 6412
rect 84074 6356 84084 6412
rect 84140 6356 86212 6412
rect 86268 6356 86278 6412
rect 86538 6356 86548 6412
rect 86604 6356 90244 6412
rect 90300 6356 90310 6412
rect 90570 6356 90580 6412
rect 90636 6356 91420 6412
rect 91476 6356 98196 6412
rect 98252 6356 98262 6412
rect 98354 6356 98364 6412
rect 98420 6356 103404 6412
rect 103562 6356 103572 6412
rect 103628 6356 105700 6412
rect 105756 6356 105766 6412
rect 109171 6356 126644 6412
rect 126700 6356 126710 6412
rect 75740 6300 75796 6356
rect 109171 6300 109227 6356
rect 126868 6300 126924 6468
rect 129780 6412 129836 6692
rect 135940 6636 135996 6692
rect 139412 6636 139468 6692
rect 142772 6636 142828 6692
rect 152851 6636 152907 6692
rect 154644 6636 154700 6692
rect 130890 6580 130900 6636
rect 130956 6580 131404 6636
rect 131460 6580 131470 6636
rect 134250 6580 134260 6636
rect 134316 6580 135996 6636
rect 136266 6580 136276 6636
rect 136332 6580 138628 6636
rect 138684 6580 138694 6636
rect 139412 6580 142828 6636
rect 144106 6580 144116 6636
rect 144172 6580 145236 6636
rect 145292 6580 145302 6636
rect 146010 6580 146020 6636
rect 146076 6580 149380 6636
rect 149436 6580 149446 6636
rect 149594 6580 149604 6636
rect 149660 6580 151508 6636
rect 151564 6580 151574 6636
rect 151722 6580 151732 6636
rect 151788 6580 151826 6636
rect 152851 6580 153692 6636
rect 153748 6580 154420 6636
rect 154476 6580 154486 6636
rect 154644 6580 154980 6636
rect 155036 6580 155046 6636
rect 155530 6580 155540 6636
rect 155596 6580 157556 6636
rect 157612 6580 157622 6636
rect 160906 6580 160916 6636
rect 160972 6580 163828 6636
rect 163884 6580 163894 6636
rect 166814 6580 166852 6636
rect 166908 6580 166918 6636
rect 167598 6580 167636 6636
rect 167692 6580 167702 6636
rect 167971 6580 175140 6636
rect 175196 6580 175206 6636
rect 178266 6580 178276 6636
rect 178332 6580 178836 6636
rect 178892 6580 178902 6636
rect 179610 6580 179620 6636
rect 179732 6580 179742 6636
rect 179834 6580 179844 6636
rect 179900 6580 189588 6636
rect 189644 6580 189654 6636
rect 189802 6580 189812 6636
rect 189868 6580 196364 6636
rect 196420 6580 196430 6636
rect 196522 6580 196532 6636
rect 196588 6580 197260 6636
rect 197316 6580 197326 6636
rect 200862 6580 200900 6636
rect 200956 6580 200966 6636
rect 202570 6580 202580 6636
rect 202636 6580 203084 6636
rect 203140 6580 203150 6636
rect 206490 6580 206500 6636
rect 206556 6580 214508 6636
rect 214564 6580 214574 6636
rect 151732 6524 151788 6580
rect 167971 6524 168027 6580
rect 130778 6468 130788 6524
rect 130844 6468 131852 6524
rect 131908 6468 131918 6524
rect 132691 6468 142660 6524
rect 142716 6468 142726 6524
rect 144218 6468 144228 6524
rect 144284 6468 145012 6524
rect 145068 6468 145078 6524
rect 145450 6468 145460 6524
rect 145516 6468 147644 6524
rect 147700 6468 147710 6524
rect 149258 6468 149268 6524
rect 149324 6468 151116 6524
rect 151172 6468 151182 6524
rect 151732 6468 153524 6524
rect 153580 6468 153590 6524
rect 154298 6468 154308 6524
rect 154364 6468 156324 6524
rect 156380 6468 156390 6524
rect 156538 6468 156548 6524
rect 156604 6468 158228 6524
rect 158284 6468 158294 6524
rect 160626 6468 160636 6524
rect 160692 6468 161028 6524
rect 161084 6468 161094 6524
rect 161354 6468 161364 6524
rect 161420 6468 165004 6524
rect 165060 6468 165070 6524
rect 166282 6468 166292 6524
rect 166348 6468 168027 6524
rect 168634 6468 168644 6524
rect 168700 6468 170996 6524
rect 171052 6468 171062 6524
rect 171210 6468 171220 6524
rect 171276 6468 179732 6524
rect 179788 6468 179798 6524
rect 179946 6468 179956 6524
rect 180012 6468 192668 6524
rect 192724 6468 192734 6524
rect 192826 6468 192836 6524
rect 192892 6468 193564 6524
rect 193620 6468 193630 6524
rect 193722 6468 193732 6524
rect 193788 6468 195244 6524
rect 195300 6468 195310 6524
rect 199658 6468 199668 6524
rect 199724 6468 212268 6524
rect 212324 6468 212334 6524
rect 213322 6468 213332 6524
rect 213388 6468 213892 6524
rect 213948 6468 215404 6524
rect 215460 6468 215796 6524
rect 215852 6468 215862 6524
rect 132691 6412 132747 6468
rect 156548 6412 156604 6468
rect 129780 6356 132747 6412
rect 133018 6356 133028 6412
rect 133084 6356 138292 6412
rect 138348 6356 138358 6412
rect 138618 6356 138628 6412
rect 138684 6356 154532 6412
rect 154588 6356 154598 6412
rect 154690 6356 154700 6412
rect 154812 6356 154822 6412
rect 154970 6356 154980 6412
rect 155036 6356 156100 6412
rect 156156 6356 156604 6412
rect 156734 6356 156772 6412
rect 156828 6356 156838 6412
rect 157546 6356 157556 6412
rect 157612 6356 165172 6412
rect 165228 6356 165238 6412
rect 165834 6356 165844 6412
rect 165900 6356 173796 6412
rect 173852 6356 173862 6412
rect 174122 6356 174132 6412
rect 174188 6356 174468 6412
rect 174524 6356 174534 6412
rect 179162 6356 179172 6412
rect 179228 6356 182420 6412
rect 182476 6356 189364 6412
rect 189420 6356 189430 6412
rect 189578 6356 189588 6412
rect 189644 6356 192892 6412
rect 192948 6356 192958 6412
rect 193162 6356 193172 6412
rect 193228 6356 194796 6412
rect 194852 6356 194862 6412
rect 200890 6356 200900 6412
rect 200956 6356 214060 6412
rect 214116 6356 214126 6412
rect 219200 6300 220000 6328
rect 24378 6244 24388 6300
rect 24444 6244 25004 6300
rect 25060 6244 52444 6300
rect 55530 6244 55540 6300
rect 55596 6244 55644 6300
rect 55700 6244 55748 6300
rect 55804 6244 55814 6300
rect 57362 6244 57372 6300
rect 57484 6244 57494 6300
rect 58370 6244 58380 6300
rect 58492 6244 58502 6300
rect 59994 6244 60004 6300
rect 60060 6244 61740 6300
rect 61796 6244 62692 6300
rect 62748 6244 62758 6300
rect 66826 6244 66836 6300
rect 66892 6244 68180 6300
rect 68236 6244 68246 6300
rect 68338 6244 68348 6300
rect 68404 6244 70700 6300
rect 70756 6244 70766 6300
rect 70858 6244 70868 6300
rect 70924 6244 72940 6300
rect 73098 6244 73108 6300
rect 73164 6244 75572 6300
rect 75628 6244 75638 6300
rect 75740 6244 84980 6300
rect 85036 6244 85046 6300
rect 85642 6244 85652 6300
rect 85708 6244 91308 6300
rect 91466 6244 91476 6300
rect 91532 6244 109227 6300
rect 109508 6244 109620 6300
rect 109676 6244 109686 6300
rect 109858 6244 109868 6300
rect 109924 6244 109972 6300
rect 110028 6244 110076 6300
rect 110132 6244 110142 6300
rect 110292 6244 116228 6300
rect 116284 6244 116294 6300
rect 116554 6244 116564 6300
rect 116620 6244 119364 6300
rect 119420 6244 119430 6300
rect 119690 6244 119700 6300
rect 119756 6244 121828 6300
rect 121884 6244 121894 6300
rect 122154 6244 122164 6300
rect 122220 6244 122948 6300
rect 123004 6244 123014 6300
rect 123172 6244 124964 6300
rect 125020 6244 125030 6300
rect 126868 6244 133476 6300
rect 133532 6244 133542 6300
rect 134138 6244 134148 6300
rect 134204 6244 144004 6300
rect 144060 6244 144070 6300
rect 144442 6244 144452 6300
rect 144508 6244 146244 6300
rect 146300 6244 146310 6300
rect 148586 6244 148596 6300
rect 148652 6244 155988 6300
rect 156044 6244 156054 6300
rect 164186 6244 164196 6300
rect 164252 6244 164300 6300
rect 164356 6244 164404 6300
rect 164460 6244 164470 6300
rect 164602 6244 164612 6300
rect 164668 6244 168644 6300
rect 168700 6244 168710 6300
rect 168858 6244 168868 6300
rect 168924 6244 171892 6300
rect 171948 6244 171958 6300
rect 177930 6244 177940 6300
rect 177996 6244 189812 6300
rect 189868 6244 189878 6300
rect 191818 6244 191828 6300
rect 191884 6244 192220 6300
rect 192276 6244 192286 6300
rect 194272 6244 194292 6300
rect 194404 6244 197764 6300
rect 197820 6244 197830 6300
rect 203242 6244 203252 6300
rect 203308 6244 203924 6300
rect 203980 6244 213276 6300
rect 213332 6244 213342 6300
rect 52388 6188 52444 6244
rect 72884 6188 72940 6244
rect 91252 6188 91308 6244
rect 109508 6188 109564 6244
rect 110292 6188 110348 6244
rect 123172 6188 123228 6244
rect 213556 6188 213612 6300
rect 213668 6244 216020 6300
rect 216076 6244 216086 6300
rect 217354 6244 217364 6300
rect 217420 6244 220000 6300
rect 219200 6216 220000 6244
rect 27738 6132 27748 6188
rect 27804 6132 28364 6188
rect 28420 6132 38667 6188
rect 40058 6132 40068 6188
rect 40124 6132 43204 6188
rect 43260 6132 43270 6188
rect 48626 6132 48636 6188
rect 48692 6132 52332 6188
rect 52388 6132 62468 6188
rect 62524 6132 62534 6188
rect 66714 6132 66724 6188
rect 66780 6132 68628 6188
rect 68684 6132 68694 6188
rect 68786 6132 68796 6188
rect 68852 6132 71428 6188
rect 71484 6132 71494 6188
rect 72884 6132 83972 6188
rect 84028 6132 84038 6188
rect 84410 6132 84420 6188
rect 84476 6132 84868 6188
rect 84924 6132 84934 6188
rect 85194 6132 85204 6188
rect 85260 6132 86436 6188
rect 86492 6132 86502 6188
rect 86986 6132 86996 6188
rect 87052 6132 87332 6188
rect 87388 6132 87398 6188
rect 87546 6132 87556 6188
rect 87612 6132 88900 6188
rect 88956 6132 88966 6188
rect 89068 6132 90692 6188
rect 90748 6132 90758 6188
rect 91252 6132 92372 6188
rect 92428 6132 93828 6188
rect 93884 6132 93894 6188
rect 97402 6132 97412 6188
rect 97468 6132 98364 6188
rect 98420 6132 98430 6188
rect 98522 6132 98532 6188
rect 98588 6132 100100 6188
rect 100156 6132 100166 6188
rect 100650 6132 100660 6188
rect 100716 6132 109564 6188
rect 109722 6132 109732 6188
rect 109788 6132 110348 6188
rect 110506 6132 110516 6188
rect 110572 6132 111972 6188
rect 112028 6132 112038 6188
rect 112298 6132 112308 6188
rect 112364 6132 113204 6188
rect 113260 6132 113708 6188
rect 113764 6132 113774 6188
rect 113866 6132 113876 6188
rect 113932 6132 116004 6188
rect 116060 6132 116070 6188
rect 116330 6132 116340 6188
rect 116396 6132 123228 6188
rect 124394 6132 124404 6188
rect 124460 6132 129220 6188
rect 129276 6132 129286 6188
rect 129434 6132 129444 6188
rect 129500 6132 141764 6188
rect 141820 6132 141830 6188
rect 145338 6132 145348 6188
rect 145404 6132 146916 6188
rect 146972 6132 146982 6188
rect 149258 6132 149268 6188
rect 149324 6132 155484 6188
rect 38611 6076 38667 6132
rect 52276 6076 52332 6132
rect 89068 6076 89124 6132
rect 155428 6076 155484 6132
rect 156324 6132 158116 6188
rect 158172 6132 158182 6188
rect 158666 6132 158676 6188
rect 158732 6132 166404 6188
rect 166460 6132 166470 6188
rect 166618 6132 166628 6188
rect 166684 6132 173908 6188
rect 173964 6132 173974 6188
rect 177594 6132 177604 6188
rect 177660 6132 179620 6188
rect 179676 6132 179686 6188
rect 182298 6132 182308 6188
rect 182364 6132 182868 6188
rect 182924 6132 182934 6188
rect 183418 6132 183428 6188
rect 183484 6132 184772 6188
rect 184828 6132 199388 6188
rect 199444 6132 199454 6188
rect 209850 6132 209860 6188
rect 209916 6132 211988 6188
rect 212044 6132 212054 6188
rect 212538 6132 212548 6188
rect 212604 6132 213612 6188
rect 156324 6076 156380 6132
rect 8810 6020 8820 6076
rect 8876 6020 9548 6076
rect 9604 6020 9614 6076
rect 10658 6020 10668 6076
rect 10724 6020 12740 6076
rect 12796 6020 25676 6076
rect 30090 6020 30100 6076
rect 30156 6020 31947 6076
rect 33450 6020 33460 6076
rect 33516 6020 35532 6076
rect 35644 6020 35654 6076
rect 38611 6020 52052 6076
rect 52108 6020 52118 6076
rect 52276 6020 71932 6076
rect 71988 6020 71998 6076
rect 73322 6020 73332 6076
rect 73388 6020 76300 6076
rect 76458 6020 76468 6076
rect 76524 6020 82908 6076
rect 83178 6020 83188 6076
rect 83244 6020 89124 6076
rect 89786 6020 89796 6076
rect 89852 6020 120708 6076
rect 120764 6020 120774 6076
rect 120931 6020 122164 6076
rect 122220 6020 122230 6076
rect 122602 6020 122612 6076
rect 122668 6020 122948 6076
rect 123004 6020 123014 6076
rect 123498 6020 123508 6076
rect 123564 6020 130900 6076
rect 130956 6020 130966 6076
rect 131450 6020 131460 6076
rect 131516 6020 137732 6076
rect 137788 6020 137798 6076
rect 139402 6020 139412 6076
rect 139468 6020 144788 6076
rect 144844 6020 144854 6076
rect 145114 6020 145124 6076
rect 145180 6020 152852 6076
rect 152908 6020 152918 6076
rect 155428 6020 156380 6076
rect 156762 6020 156772 6076
rect 156828 6020 159236 6076
rect 159292 6020 159302 6076
rect 159450 6020 159460 6076
rect 159516 6020 166516 6076
rect 166572 6020 166582 6076
rect 166740 6020 169316 6076
rect 169372 6020 169382 6076
rect 170986 6020 170996 6076
rect 171052 6020 174692 6076
rect 174748 6020 174758 6076
rect 175102 6020 175140 6076
rect 175196 6020 175206 6076
rect 175466 6020 175476 6076
rect 175532 6020 179620 6076
rect 179676 6020 179686 6076
rect 180170 6020 180180 6076
rect 180236 6020 191212 6076
rect 191268 6020 191278 6076
rect 193274 6020 193284 6076
rect 193396 6020 193406 6076
rect 194842 6020 194852 6076
rect 194908 6020 195132 6076
rect 195188 6020 195198 6076
rect 195300 6020 197708 6076
rect 197764 6020 205716 6076
rect 205772 6020 205782 6076
rect 209626 6020 209636 6076
rect 209692 6020 214900 6076
rect 214956 6020 214966 6076
rect 25620 5964 25676 6020
rect 31891 5964 31947 6020
rect 24714 5908 24724 5964
rect 24780 5908 25452 5964
rect 25508 5908 25518 5964
rect 25620 5908 30100 5964
rect 30156 5908 30166 5964
rect 31891 5908 51828 5964
rect 51884 5908 51894 5964
rect 52154 5908 52164 5964
rect 52220 5908 69916 5964
rect 69972 5908 69982 5964
rect 70084 5908 73780 5964
rect 73836 5908 73846 5964
rect 73994 5908 74004 5964
rect 74060 5908 75460 5964
rect 75516 5908 75526 5964
rect 70084 5852 70140 5908
rect 76244 5852 76300 6020
rect 82852 5964 82908 6020
rect 120931 5964 120987 6020
rect 166740 5964 166796 6020
rect 195300 5964 195356 6020
rect 76458 5908 76468 5964
rect 76524 5908 77812 5964
rect 77868 5908 77878 5964
rect 78204 5908 82404 5964
rect 82460 5908 82470 5964
rect 82852 5908 84644 5964
rect 84700 5908 84710 5964
rect 84858 5908 84868 5964
rect 84924 5908 85540 5964
rect 85596 5908 85606 5964
rect 85754 5908 85764 5964
rect 85820 5908 99428 5964
rect 99484 5908 99494 5964
rect 100650 5908 100660 5964
rect 100716 5908 108500 5964
rect 108556 5908 108566 5964
rect 109610 5908 109620 5964
rect 109676 5908 109732 5964
rect 109788 5908 109798 5964
rect 110058 5908 110068 5964
rect 110124 5908 113764 5964
rect 113820 5908 113830 5964
rect 113988 5908 117012 5964
rect 117068 5908 117078 5964
rect 117674 5908 117684 5964
rect 117740 5908 118804 5964
rect 118860 5908 118870 5964
rect 119018 5908 119028 5964
rect 119084 5908 119122 5964
rect 119242 5908 119252 5964
rect 119308 5908 119756 5964
rect 119812 5908 120987 5964
rect 121258 5908 121268 5964
rect 121324 5908 121604 5964
rect 121660 5908 121670 5964
rect 121818 5908 121828 5964
rect 121884 5908 122612 5964
rect 122668 5908 122678 5964
rect 122826 5908 122836 5964
rect 122892 5908 129556 5964
rect 129612 5908 129622 5964
rect 130554 5908 130564 5964
rect 130620 5908 131068 5964
rect 131124 5908 131134 5964
rect 131226 5908 131236 5964
rect 131292 5908 135100 5964
rect 135156 5908 135166 5964
rect 135538 5908 135548 5964
rect 135604 5908 135940 5964
rect 135996 5908 136006 5964
rect 136602 5908 136612 5964
rect 136668 5908 139300 5964
rect 139356 5908 139366 5964
rect 140858 5908 140868 5964
rect 140924 5908 144676 5964
rect 144732 5908 144742 5964
rect 145226 5908 145236 5964
rect 145292 5908 165396 5964
rect 165452 5908 165462 5964
rect 166394 5908 166404 5964
rect 166460 5908 166796 5964
rect 167290 5908 167300 5964
rect 167356 5908 169204 5964
rect 169260 5908 169270 5964
rect 171098 5908 171108 5964
rect 171164 5908 173012 5964
rect 173068 5908 173078 5964
rect 174570 5908 174580 5964
rect 174636 5908 190484 5964
rect 190540 5908 190550 5964
rect 194506 5908 194516 5964
rect 194572 5908 195356 5964
rect 205482 5908 205492 5964
rect 205548 5908 214172 5964
rect 214228 5908 214238 5964
rect 78204 5852 78260 5908
rect 113988 5852 114044 5908
rect 16874 5796 16884 5852
rect 16940 5796 17500 5852
rect 17556 5796 41748 5852
rect 41804 5796 41814 5852
rect 41962 5796 41972 5852
rect 42028 5796 42364 5852
rect 42476 5796 42486 5852
rect 42746 5796 42756 5852
rect 42812 5796 43260 5852
rect 43316 5796 43326 5852
rect 46554 5796 46564 5852
rect 46620 5796 47068 5852
rect 47124 5796 47134 5852
rect 47236 5796 50372 5852
rect 50428 5796 50438 5852
rect 51034 5796 51044 5852
rect 51100 5796 51548 5852
rect 51660 5796 51670 5852
rect 52042 5796 52052 5852
rect 52108 5796 64596 5852
rect 64652 5796 64662 5852
rect 65594 5796 65604 5852
rect 65660 5796 67284 5852
rect 67340 5796 67350 5852
rect 67442 5796 67452 5852
rect 67508 5796 69412 5852
rect 69468 5796 69478 5852
rect 69626 5796 69636 5852
rect 69692 5796 70140 5852
rect 70298 5796 70308 5852
rect 70364 5796 73388 5852
rect 73546 5796 73556 5852
rect 73612 5796 75908 5852
rect 75964 5796 75974 5852
rect 76244 5796 78260 5852
rect 78586 5796 78596 5852
rect 78652 5796 81004 5852
rect 81498 5796 81508 5852
rect 81564 5796 83300 5852
rect 83356 5796 83366 5852
rect 83738 5796 83748 5852
rect 83804 5796 85204 5852
rect 85260 5796 85270 5852
rect 85418 5796 85428 5852
rect 85484 5796 85820 5852
rect 85876 5796 86996 5852
rect 87052 5796 87062 5852
rect 87210 5796 87220 5852
rect 87276 5796 87948 5852
rect 88004 5796 88564 5852
rect 88620 5796 88630 5852
rect 88778 5796 88788 5852
rect 88844 5796 89236 5852
rect 89292 5796 89302 5852
rect 89450 5796 89460 5852
rect 89516 5796 100436 5852
rect 100492 5796 100502 5852
rect 100650 5796 100660 5852
rect 100716 5796 101724 5852
rect 101780 5796 101790 5852
rect 102106 5796 102116 5852
rect 102172 5796 103236 5852
rect 103292 5796 103302 5852
rect 103674 5796 103684 5852
rect 103740 5796 104132 5852
rect 104188 5796 104198 5852
rect 104346 5796 104356 5852
rect 104412 5796 104468 5852
rect 104524 5796 104534 5852
rect 104906 5796 104916 5852
rect 104972 5796 114044 5852
rect 114202 5796 114212 5852
rect 114268 5796 115444 5852
rect 115500 5796 115510 5852
rect 115882 5796 115892 5852
rect 115948 5796 119364 5852
rect 119420 5796 119430 5852
rect 119914 5796 119924 5852
rect 119980 5796 120372 5852
rect 120428 5796 120438 5852
rect 120931 5796 123284 5852
rect 123340 5796 123350 5852
rect 126634 5796 126644 5852
rect 126700 5796 133140 5852
rect 133196 5796 133206 5852
rect 134250 5796 134260 5852
rect 134316 5796 137844 5852
rect 137900 5796 137910 5852
rect 138730 5796 138740 5852
rect 138796 5796 140980 5852
rect 141036 5796 141046 5852
rect 141194 5796 141204 5852
rect 141260 5796 144228 5852
rect 144284 5796 144294 5852
rect 144442 5796 144452 5852
rect 144508 5796 146244 5852
rect 146300 5796 146310 5852
rect 146906 5796 146916 5852
rect 146972 5796 150276 5852
rect 150332 5796 150342 5852
rect 150910 5796 150948 5852
rect 151004 5796 151014 5852
rect 151778 5796 151788 5852
rect 151844 5796 181300 5852
rect 181356 5796 181366 5852
rect 183194 5796 183204 5852
rect 183260 5796 183540 5852
rect 183596 5796 198492 5852
rect 198548 5796 198558 5852
rect 210298 5796 210308 5852
rect 210364 5796 210980 5852
rect 211036 5796 214620 5852
rect 214676 5796 214686 5852
rect 15866 5684 15876 5740
rect 15932 5684 18060 5740
rect 18172 5684 18182 5740
rect 32666 5684 32676 5740
rect 32732 5684 33460 5740
rect 33516 5684 33526 5740
rect 33842 5684 33852 5740
rect 33964 5684 33974 5740
rect 37706 5684 37716 5740
rect 37772 5684 47012 5740
rect 47068 5684 47078 5740
rect 47236 5628 47292 5796
rect 73332 5740 73388 5796
rect 80948 5740 81004 5796
rect 120931 5740 120987 5796
rect 50371 5684 69244 5740
rect 69300 5684 69310 5740
rect 69402 5684 69412 5740
rect 69468 5684 73108 5740
rect 73164 5684 73174 5740
rect 73332 5684 74788 5740
rect 74844 5684 74854 5740
rect 75002 5684 75012 5740
rect 75068 5684 80052 5740
rect 80108 5684 80118 5740
rect 80276 5684 80724 5740
rect 80780 5684 80790 5740
rect 80948 5684 82180 5740
rect 82236 5684 82246 5740
rect 82730 5684 82740 5740
rect 82796 5684 84476 5740
rect 84532 5684 84542 5740
rect 84634 5684 84644 5740
rect 84700 5684 87108 5740
rect 87164 5684 87174 5740
rect 87322 5684 87332 5740
rect 87388 5684 87780 5740
rect 87836 5684 87846 5740
rect 88116 5684 90468 5740
rect 90524 5684 90534 5740
rect 91186 5684 91196 5740
rect 91252 5684 98196 5740
rect 98252 5684 98262 5740
rect 98410 5684 98420 5740
rect 98476 5684 98980 5740
rect 99036 5684 99046 5740
rect 100762 5684 100772 5740
rect 100828 5684 105364 5740
rect 105420 5684 105430 5740
rect 105690 5684 105700 5740
rect 105756 5684 120987 5740
rect 121146 5684 121156 5740
rect 121212 5684 121828 5740
rect 121884 5684 121894 5740
rect 122266 5684 122276 5740
rect 122332 5684 133140 5740
rect 133196 5684 133206 5740
rect 135594 5684 135604 5740
rect 135660 5684 138068 5740
rect 138124 5684 138134 5740
rect 139402 5684 139412 5740
rect 139468 5684 156996 5740
rect 157052 5684 157062 5740
rect 157210 5684 157220 5740
rect 157276 5684 160580 5740
rect 160636 5684 160646 5740
rect 160738 5684 160748 5740
rect 160804 5684 186788 5740
rect 186844 5684 186854 5740
rect 187012 5684 191436 5740
rect 191492 5684 191502 5740
rect 197754 5684 197764 5740
rect 197820 5684 212548 5740
rect 212604 5684 212614 5740
rect 212762 5684 212772 5740
rect 212884 5684 212996 5740
rect 213052 5684 213062 5740
rect 50371 5628 50427 5684
rect 80276 5628 80332 5684
rect 18778 5572 18788 5628
rect 18844 5572 37100 5628
rect 38490 5572 38500 5628
rect 38556 5572 39228 5628
rect 39284 5572 40068 5628
rect 40124 5572 40134 5628
rect 41738 5572 41748 5628
rect 41804 5572 47292 5628
rect 47450 5572 47460 5628
rect 47516 5572 50427 5628
rect 52042 5572 52052 5628
rect 52108 5572 54180 5628
rect 54236 5572 54246 5628
rect 56186 5572 56196 5628
rect 56252 5572 73276 5628
rect 73332 5572 73342 5628
rect 73658 5572 73668 5628
rect 73724 5572 75572 5628
rect 75628 5572 75638 5628
rect 75786 5572 75796 5628
rect 75852 5572 78708 5628
rect 78764 5572 78774 5628
rect 78922 5572 78932 5628
rect 78988 5572 80332 5628
rect 80490 5572 80500 5628
rect 80556 5572 87892 5628
rect 87948 5572 87958 5628
rect 37044 5516 37100 5572
rect 88116 5516 88172 5684
rect 88330 5572 88340 5628
rect 88396 5572 89796 5628
rect 89852 5572 89862 5628
rect 90010 5572 90020 5628
rect 90076 5572 91700 5628
rect 91756 5572 91766 5628
rect 92250 5572 92260 5628
rect 92316 5572 92596 5628
rect 92652 5572 92662 5628
rect 95162 5572 95172 5628
rect 95228 5572 100044 5628
rect 100426 5572 100436 5628
rect 100492 5572 109508 5628
rect 109564 5572 109574 5628
rect 109722 5572 109732 5628
rect 109788 5572 118580 5628
rect 118636 5572 118646 5628
rect 119018 5572 119028 5628
rect 119084 5572 123508 5628
rect 123564 5572 123574 5628
rect 123722 5572 123732 5628
rect 123788 5572 131012 5628
rect 131068 5572 131078 5628
rect 132514 5572 132524 5628
rect 132580 5572 134260 5628
rect 134316 5572 134326 5628
rect 137498 5572 137508 5628
rect 137564 5572 144788 5628
rect 144844 5572 144854 5628
rect 145002 5572 145012 5628
rect 145068 5572 145348 5628
rect 145404 5572 145414 5628
rect 145674 5572 145684 5628
rect 145740 5572 155652 5628
rect 155708 5572 155718 5628
rect 155978 5572 155988 5628
rect 156044 5572 161140 5628
rect 161196 5572 161206 5628
rect 161466 5572 161476 5628
rect 161532 5572 166628 5628
rect 166684 5572 166694 5628
rect 166954 5572 166964 5628
rect 167020 5572 169484 5628
rect 169540 5572 169550 5628
rect 173786 5572 173796 5628
rect 173852 5572 184772 5628
rect 184828 5572 184838 5628
rect 99988 5516 100044 5572
rect 187012 5516 187068 5684
rect 187898 5572 187908 5628
rect 187964 5572 188020 5628
rect 188076 5572 188086 5628
rect 188654 5572 188692 5628
rect 188748 5572 188758 5628
rect 202010 5572 202020 5628
rect 202076 5572 203140 5628
rect 203196 5572 213444 5628
rect 213500 5572 213724 5628
rect 213780 5572 213790 5628
rect 28366 5460 28376 5516
rect 28432 5460 28480 5516
rect 28536 5460 28584 5516
rect 28640 5460 28650 5516
rect 31770 5460 31780 5516
rect 31836 5460 33908 5516
rect 33964 5460 33974 5516
rect 37044 5460 57204 5516
rect 57260 5460 57270 5516
rect 57418 5460 57428 5516
rect 57484 5460 73220 5516
rect 73276 5460 73286 5516
rect 73434 5460 73444 5516
rect 73500 5460 75012 5516
rect 75068 5460 75078 5516
rect 75170 5460 75180 5516
rect 75236 5460 81396 5516
rect 81452 5460 81462 5516
rect 81610 5460 81620 5516
rect 81676 5460 82516 5516
rect 82572 5460 82582 5516
rect 82694 5460 82704 5516
rect 82760 5460 82808 5516
rect 82864 5460 82912 5516
rect 82968 5460 82978 5516
rect 83514 5460 83524 5516
rect 83580 5460 83916 5516
rect 83972 5460 83982 5516
rect 84466 5460 84476 5516
rect 84532 5460 88172 5516
rect 88340 5460 97972 5516
rect 98028 5460 98038 5516
rect 98186 5460 98196 5516
rect 98252 5460 99428 5516
rect 99484 5460 99494 5516
rect 99988 5460 101444 5516
rect 101500 5460 101510 5516
rect 101658 5460 101668 5516
rect 101724 5460 102340 5516
rect 102396 5460 102406 5516
rect 102666 5460 102676 5516
rect 102732 5460 110292 5516
rect 110348 5460 110358 5516
rect 111962 5460 111972 5516
rect 112028 5460 114212 5516
rect 114268 5460 114278 5516
rect 114650 5460 114660 5516
rect 114716 5460 123004 5516
rect 123162 5460 123172 5516
rect 123228 5460 133028 5516
rect 133084 5460 133094 5516
rect 137022 5460 137032 5516
rect 137088 5460 137136 5516
rect 137192 5460 137240 5516
rect 137296 5460 137306 5516
rect 137498 5460 137508 5516
rect 137564 5460 137620 5516
rect 137676 5460 137686 5516
rect 137834 5460 137844 5516
rect 137900 5460 141372 5516
rect 142146 5460 142156 5516
rect 142212 5460 161140 5516
rect 161196 5460 161206 5516
rect 162250 5460 162260 5516
rect 162316 5460 163828 5516
rect 163884 5460 163894 5516
rect 166170 5460 166180 5516
rect 166236 5460 167076 5516
rect 167132 5460 167142 5516
rect 167850 5460 167860 5516
rect 167916 5460 176484 5516
rect 176540 5460 187068 5516
rect 191350 5460 191360 5516
rect 191416 5460 191464 5516
rect 191520 5460 191568 5516
rect 191624 5460 191634 5516
rect 193050 5460 193060 5516
rect 193116 5460 203307 5516
rect 210746 5460 210756 5516
rect 210812 5460 213892 5516
rect 213948 5460 213958 5516
rect 88340 5404 88396 5460
rect 122948 5404 123004 5460
rect 141316 5404 141372 5460
rect 203251 5404 203307 5460
rect 25442 5348 25452 5404
rect 25508 5348 57092 5404
rect 57148 5348 57158 5404
rect 58650 5348 58660 5404
rect 58716 5348 60508 5404
rect 60564 5348 72828 5404
rect 72772 5292 72828 5348
rect 73556 5348 84308 5404
rect 84364 5348 84374 5404
rect 84522 5348 84532 5404
rect 84588 5348 85204 5404
rect 85260 5348 85270 5404
rect 85418 5348 85428 5404
rect 85484 5348 88396 5404
rect 88554 5348 88564 5404
rect 88620 5348 92372 5404
rect 92428 5348 92438 5404
rect 93930 5348 93940 5404
rect 93996 5348 94780 5404
rect 94836 5348 122724 5404
rect 122780 5348 122790 5404
rect 122948 5348 129332 5404
rect 129388 5348 129398 5404
rect 129546 5348 129556 5404
rect 129612 5348 131236 5404
rect 131292 5348 131302 5404
rect 134250 5348 134260 5404
rect 134316 5348 141092 5404
rect 141148 5348 141158 5404
rect 141316 5348 143780 5404
rect 143836 5348 143846 5404
rect 143994 5348 144004 5404
rect 144060 5348 149716 5404
rect 149772 5348 149782 5404
rect 150266 5348 150276 5404
rect 150332 5348 152012 5404
rect 152618 5348 152628 5404
rect 152684 5348 160748 5404
rect 160804 5348 160814 5404
rect 162474 5348 162484 5404
rect 162540 5348 167188 5404
rect 167244 5348 167254 5404
rect 169474 5348 169484 5404
rect 169540 5348 170100 5404
rect 170156 5348 170166 5404
rect 171658 5348 171668 5404
rect 171724 5348 177492 5404
rect 177548 5348 177558 5404
rect 177930 5348 177940 5404
rect 177996 5348 178164 5404
rect 178220 5348 181300 5404
rect 181356 5348 181366 5404
rect 184314 5348 184324 5404
rect 184380 5348 194404 5404
rect 194460 5348 194470 5404
rect 203251 5348 209860 5404
rect 209916 5348 209926 5404
rect 211278 5348 211316 5404
rect 211372 5348 215068 5404
rect 215124 5348 216468 5404
rect 216524 5348 216534 5404
rect 73556 5292 73612 5348
rect 151956 5292 152012 5348
rect 14074 5236 14084 5292
rect 14140 5236 68180 5292
rect 68236 5236 68246 5292
rect 68394 5236 68404 5292
rect 68460 5236 70868 5292
rect 70924 5236 70934 5292
rect 71754 5236 71764 5292
rect 71820 5236 72548 5292
rect 72604 5236 72614 5292
rect 72772 5236 73612 5292
rect 73770 5236 73780 5292
rect 73836 5236 91476 5292
rect 91532 5236 91542 5292
rect 91690 5236 91700 5292
rect 91756 5236 95284 5292
rect 95340 5236 95350 5292
rect 96292 5236 100996 5292
rect 101052 5236 101062 5292
rect 101210 5236 101220 5292
rect 101276 5236 103012 5292
rect 103068 5236 103078 5292
rect 103226 5236 103236 5292
rect 103292 5236 107380 5292
rect 107436 5236 107446 5292
rect 107594 5236 107604 5292
rect 107660 5236 113204 5292
rect 113260 5236 113270 5292
rect 113418 5236 113428 5292
rect 113484 5236 114156 5292
rect 114212 5236 116676 5292
rect 116732 5236 116742 5292
rect 117338 5236 117348 5292
rect 117404 5236 119028 5292
rect 119084 5236 119094 5292
rect 119242 5236 119252 5292
rect 119308 5236 121716 5292
rect 121772 5236 121782 5292
rect 122602 5236 122612 5292
rect 122668 5236 128548 5292
rect 128604 5236 128614 5292
rect 128762 5236 128772 5292
rect 128828 5236 129444 5292
rect 129500 5236 129510 5292
rect 129658 5236 129668 5292
rect 129724 5236 131348 5292
rect 131404 5236 131414 5292
rect 132346 5236 132356 5292
rect 132412 5236 134148 5292
rect 134204 5236 134214 5292
rect 136388 5236 138628 5292
rect 138684 5236 138694 5292
rect 139178 5236 139188 5292
rect 139244 5236 142380 5292
rect 142538 5236 142548 5292
rect 142604 5236 144452 5292
rect 144508 5236 144518 5292
rect 144676 5236 145684 5292
rect 145740 5236 145750 5292
rect 145898 5236 145908 5292
rect 145964 5236 151788 5292
rect 151844 5236 151854 5292
rect 151956 5236 159348 5292
rect 159404 5236 159414 5292
rect 159562 5236 159572 5292
rect 159628 5236 164500 5292
rect 164556 5236 164566 5292
rect 165386 5236 165396 5292
rect 165452 5236 183708 5292
rect 183764 5236 183774 5292
rect 187898 5236 187908 5292
rect 187964 5236 201684 5292
rect 201740 5236 201750 5292
rect 19198 5124 19236 5180
rect 19292 5124 19302 5180
rect 20458 5124 20468 5180
rect 20524 5124 21700 5180
rect 21756 5124 21766 5180
rect 23006 5124 23044 5180
rect 23100 5124 23110 5180
rect 43866 5124 43876 5180
rect 43932 5124 50427 5180
rect 55738 5124 55748 5180
rect 55804 5124 55972 5180
rect 56028 5124 56038 5180
rect 56186 5124 56196 5180
rect 56252 5124 57428 5180
rect 57484 5124 57494 5180
rect 58650 5124 58660 5180
rect 58716 5124 60676 5180
rect 60732 5124 60742 5180
rect 63802 5124 63812 5180
rect 63868 5124 73332 5180
rect 73388 5124 73398 5180
rect 73556 5124 78708 5180
rect 78764 5124 78774 5180
rect 79034 5124 79044 5180
rect 79100 5124 79716 5180
rect 79772 5124 79782 5180
rect 80042 5124 80052 5180
rect 80108 5124 82292 5180
rect 82348 5124 82358 5180
rect 83178 5124 83188 5180
rect 83244 5124 84924 5180
rect 84980 5124 84990 5180
rect 85082 5124 85092 5180
rect 85148 5124 86212 5180
rect 86268 5124 86278 5180
rect 87434 5124 87444 5180
rect 87500 5124 89908 5180
rect 89964 5124 89974 5180
rect 90570 5124 90580 5180
rect 90636 5124 91196 5180
rect 91252 5124 91262 5180
rect 91354 5124 91364 5180
rect 91420 5124 91924 5180
rect 91980 5124 91990 5180
rect 92250 5124 92260 5180
rect 92316 5124 96068 5180
rect 96124 5124 96134 5180
rect 50371 5068 50427 5124
rect 73556 5068 73612 5124
rect 96292 5068 96348 5236
rect 136388 5180 136444 5236
rect 142324 5180 142380 5236
rect 144676 5180 144732 5236
rect 97402 5124 97412 5180
rect 97468 5124 98028 5180
rect 98084 5124 104020 5180
rect 104076 5124 104086 5180
rect 106698 5124 106708 5180
rect 106764 5124 107548 5180
rect 107604 5124 136444 5180
rect 136602 5124 136612 5180
rect 136668 5124 142156 5180
rect 142212 5124 142222 5180
rect 142324 5124 144732 5180
rect 145114 5124 145124 5180
rect 145180 5124 158676 5180
rect 158732 5124 158742 5180
rect 159450 5124 159460 5180
rect 159516 5124 166292 5180
rect 166348 5124 166358 5180
rect 166730 5124 166740 5180
rect 166796 5124 167636 5180
rect 167692 5124 167702 5180
rect 175914 5124 175924 5180
rect 175980 5124 177716 5180
rect 177772 5124 177782 5180
rect 178042 5124 178052 5180
rect 178108 5124 181636 5180
rect 181692 5124 181702 5180
rect 189354 5124 189364 5180
rect 189420 5124 205492 5180
rect 205548 5124 205558 5180
rect 21102 5012 21140 5068
rect 21196 5012 21206 5068
rect 23342 5012 23380 5068
rect 23436 5012 23446 5068
rect 24378 5012 24388 5068
rect 24444 5012 25228 5068
rect 25284 5012 25294 5068
rect 49774 5012 49812 5068
rect 49868 5012 49878 5068
rect 50371 5012 71204 5068
rect 71260 5012 71270 5068
rect 71418 5012 71428 5068
rect 71484 5012 73612 5068
rect 73882 5012 73892 5068
rect 73948 5012 75180 5068
rect 75236 5012 75246 5068
rect 75348 5012 77140 5068
rect 77196 5012 77206 5068
rect 77354 5012 77364 5068
rect 77420 5012 86660 5068
rect 86716 5012 86726 5068
rect 87098 5012 87108 5068
rect 87164 5012 87948 5068
rect 88004 5012 88014 5068
rect 88218 5012 88228 5068
rect 88284 5012 90020 5068
rect 90076 5012 90086 5068
rect 90234 5012 90244 5068
rect 90300 5012 96348 5068
rect 96954 5012 96964 5068
rect 97020 5012 98868 5068
rect 98924 5012 98934 5068
rect 99194 5012 99204 5068
rect 99260 5012 101556 5068
rect 101612 5012 101622 5068
rect 101770 5012 101780 5068
rect 101836 5012 110068 5068
rect 110124 5012 110134 5068
rect 110282 5012 110292 5068
rect 110348 5012 111468 5068
rect 111524 5012 111534 5068
rect 112634 5012 112644 5068
rect 112700 5012 115668 5068
rect 115724 5012 115734 5068
rect 115882 5012 115892 5068
rect 115948 5012 135268 5068
rect 135324 5012 135334 5068
rect 140634 5012 140644 5068
rect 140700 5012 147644 5068
rect 148530 5012 148540 5068
rect 148652 5012 148662 5068
rect 149426 5012 149436 5068
rect 149492 5012 154532 5068
rect 154588 5012 154598 5068
rect 157434 5012 157444 5068
rect 157500 5012 159012 5068
rect 159068 5012 159078 5068
rect 159338 5012 159348 5068
rect 159404 5012 162988 5068
rect 164042 5012 164052 5068
rect 164108 5012 185220 5068
rect 185276 5012 185286 5068
rect 188906 5012 188916 5068
rect 189028 5012 189038 5068
rect 189130 5012 189140 5068
rect 189196 5012 205604 5068
rect 205660 5012 205670 5068
rect 207778 5012 207788 5068
rect 207844 5012 210532 5068
rect 210588 5012 212268 5068
rect 75348 4956 75404 5012
rect 8698 4900 8708 4956
rect 8764 4900 9548 4956
rect 9660 4900 9670 4956
rect 10546 4900 10556 4956
rect 10612 4900 11620 4956
rect 11676 4900 11686 4956
rect 15754 4900 15764 4956
rect 15820 4900 16380 4956
rect 16492 4900 16502 4956
rect 28298 4900 28308 4956
rect 28364 4900 29148 4956
rect 29204 4900 29214 4956
rect 35018 4900 35028 4956
rect 35084 4900 35644 4956
rect 35756 4900 35766 4956
rect 38611 4900 56196 4956
rect 56252 4900 56262 4956
rect 56578 4900 56588 4956
rect 56700 4900 56710 4956
rect 57978 4900 57988 4956
rect 58044 4900 66836 4956
rect 66892 4900 66902 4956
rect 67050 4900 67060 4956
rect 67116 4900 68404 4956
rect 68460 4900 68470 4956
rect 68954 4900 68964 4956
rect 69020 4900 69748 4956
rect 69804 4900 69814 4956
rect 70074 4900 70084 4956
rect 70140 4900 70868 4956
rect 70924 4900 70934 4956
rect 71194 4900 71204 4956
rect 71260 4900 72828 4956
rect 73658 4900 73668 4956
rect 73724 4900 74284 4956
rect 74778 4900 74788 4956
rect 74844 4900 75404 4956
rect 76794 4900 76804 4956
rect 76860 4900 78484 4956
rect 78540 4900 78550 4956
rect 79258 4900 79268 4956
rect 79324 4900 80108 4956
rect 80164 4900 80174 4956
rect 80378 4900 80388 4956
rect 80444 4900 80836 4956
rect 80892 4900 80902 4956
rect 81274 4900 81284 4956
rect 81340 4900 81956 4956
rect 82012 4900 82022 4956
rect 82170 4900 82180 4956
rect 82236 4900 83636 4956
rect 83692 4900 83702 4956
rect 83962 4900 83972 4956
rect 84028 4900 84532 4956
rect 84588 4900 84598 4956
rect 84914 4900 84924 4956
rect 84980 4900 85764 4956
rect 85820 4900 85830 4956
rect 85978 4900 85988 4956
rect 86044 4900 89572 4956
rect 89628 4900 89638 4956
rect 89898 4900 89908 4956
rect 89964 4900 91700 4956
rect 91756 4900 91766 4956
rect 91914 4900 91924 4956
rect 91980 4900 97076 4956
rect 97132 4900 97142 4956
rect 97290 4900 97300 4956
rect 97356 4900 100100 4956
rect 100156 4900 100166 4956
rect 100314 4900 100324 4956
rect 100380 4900 101332 4956
rect 101388 4900 110516 4956
rect 110572 4900 110582 4956
rect 110954 4900 110964 4956
rect 111020 4900 112532 4956
rect 112588 4900 112598 4956
rect 113194 4900 113204 4956
rect 113260 4900 116452 4956
rect 116508 4900 116518 4956
rect 116666 4900 116676 4956
rect 116732 4900 118804 4956
rect 118860 4900 118870 4956
rect 119018 4900 119028 4956
rect 119084 4900 121156 4956
rect 121212 4900 121222 4956
rect 121370 4900 121380 4956
rect 121436 4900 121604 4956
rect 121660 4900 121670 4956
rect 121818 4900 121828 4956
rect 121884 4900 123116 4956
rect 123274 4900 123284 4956
rect 123340 4900 126532 4956
rect 126588 4900 126598 4956
rect 126746 4900 126756 4956
rect 126812 4900 133588 4956
rect 133644 4900 133654 4956
rect 133802 4900 133812 4956
rect 133868 4900 135604 4956
rect 135660 4900 135670 4956
rect 135930 4900 135940 4956
rect 135996 4900 139412 4956
rect 139468 4900 139478 4956
rect 140522 4900 140532 4956
rect 140588 4900 141596 4956
rect 141652 4900 141662 4956
rect 141754 4900 141764 4956
rect 141820 4900 147084 4956
rect 147140 4900 147150 4956
rect 147588 4900 147644 5012
rect 162932 4956 162988 5012
rect 212212 4956 212268 5012
rect 147700 4900 151060 4956
rect 151116 4900 151126 4956
rect 152842 4900 152852 4956
rect 152908 4900 154476 4956
rect 154532 4900 154542 4956
rect 154634 4900 154644 4956
rect 154700 4900 156436 4956
rect 156492 4900 156502 4956
rect 161354 4900 161364 4956
rect 161420 4900 162484 4956
rect 162540 4900 162550 4956
rect 162932 4900 165452 4956
rect 165508 4900 165518 4956
rect 166282 4900 166292 4956
rect 166348 4900 168868 4956
rect 168924 4900 168934 4956
rect 173002 4900 173012 4956
rect 173068 4900 179396 4956
rect 179452 4900 179462 4956
rect 180058 4900 180068 4956
rect 180124 4900 189756 4956
rect 189812 4900 189822 4956
rect 190026 4900 190036 4956
rect 190092 4900 190652 4956
rect 190708 4900 190718 4956
rect 191930 4900 191940 4956
rect 191996 4900 192444 4956
rect 192500 4900 192510 4956
rect 193162 4900 193172 4956
rect 193228 4900 193676 4956
rect 193732 4900 193742 4956
rect 194842 4900 194852 4956
rect 194908 4900 195468 4956
rect 195524 4900 195534 4956
rect 195636 4900 200900 4956
rect 200956 4900 200966 4956
rect 207890 4900 207900 4956
rect 207956 4900 208740 4956
rect 208796 4900 208806 4956
rect 209962 4900 209972 4956
rect 210028 4900 211596 4956
rect 211652 4900 211662 4956
rect 211754 4900 211764 4956
rect 211820 4900 212044 4956
rect 212100 4900 212110 4956
rect 212212 4900 214620 4956
rect 214676 4900 214686 4956
rect 215058 4900 215068 4956
rect 215124 4900 216132 4956
rect 216188 4900 216198 4956
rect 3770 4788 3780 4844
rect 3836 4788 23044 4844
rect 23100 4788 23110 4844
rect 38611 4732 38667 4900
rect 72772 4844 72828 4900
rect 74228 4844 74284 4900
rect 123060 4844 123116 4900
rect 195636 4844 195692 4900
rect 43082 4788 43092 4844
rect 43148 4788 43708 4844
rect 43764 4788 45108 4844
rect 45164 4788 45174 4844
rect 48346 4788 48356 4844
rect 48412 4788 49644 4844
rect 49700 4788 49710 4844
rect 52266 4788 52276 4844
rect 52332 4788 54516 4844
rect 54572 4788 54582 4844
rect 55412 4788 56140 4844
rect 63466 4788 63476 4844
rect 63532 4788 64428 4844
rect 64484 4788 67284 4844
rect 67340 4788 67350 4844
rect 67610 4788 67620 4844
rect 67676 4788 69524 4844
rect 69580 4788 69590 4844
rect 71988 4788 72548 4844
rect 72604 4788 72614 4844
rect 72772 4788 74004 4844
rect 74060 4788 74070 4844
rect 74228 4788 82068 4844
rect 82124 4788 82134 4844
rect 82394 4788 82404 4844
rect 82460 4788 102788 4844
rect 102844 4788 102854 4844
rect 103002 4788 103012 4844
rect 103068 4788 112084 4844
rect 112140 4788 112150 4844
rect 112410 4788 112420 4844
rect 112476 4788 119868 4844
rect 120026 4788 120036 4844
rect 120092 4788 122836 4844
rect 122892 4788 122902 4844
rect 123060 4788 127204 4844
rect 127260 4788 127270 4844
rect 129994 4788 130004 4844
rect 130060 4788 132356 4844
rect 132412 4788 132422 4844
rect 132570 4788 132580 4844
rect 132636 4788 133420 4844
rect 133476 4788 137396 4844
rect 137452 4788 137462 4844
rect 137946 4788 137956 4844
rect 138012 4788 139412 4844
rect 139468 4788 139478 4844
rect 140970 4788 140980 4844
rect 141036 4788 142828 4844
rect 142884 4788 144228 4844
rect 144284 4788 144294 4844
rect 144442 4788 144452 4844
rect 144508 4788 144676 4844
rect 144732 4788 144742 4844
rect 144890 4788 144900 4844
rect 144956 4788 146020 4844
rect 146076 4788 148876 4844
rect 148932 4788 148942 4844
rect 149482 4788 149492 4844
rect 149548 4788 149940 4844
rect 149996 4788 153132 4844
rect 153188 4788 153198 4844
rect 153300 4788 180180 4844
rect 180236 4788 180246 4844
rect 180394 4788 180404 4844
rect 180460 4788 181132 4844
rect 181188 4788 181198 4844
rect 182158 4788 182196 4844
rect 182252 4788 182262 4844
rect 183316 4788 185332 4844
rect 185388 4788 185398 4844
rect 185556 4788 192892 4844
rect 192948 4788 192958 4844
rect 193050 4788 193060 4844
rect 193116 4788 195692 4844
rect 196644 4788 201796 4844
rect 201852 4788 201862 4844
rect 209850 4788 209860 4844
rect 209916 4788 211092 4844
rect 211148 4788 215516 4844
rect 215572 4788 215582 4844
rect 5002 4676 5012 4732
rect 5068 4676 26964 4732
rect 27020 4676 27030 4732
rect 33450 4676 33460 4732
rect 33516 4676 38667 4732
rect 41850 4676 41860 4732
rect 41916 4676 44324 4732
rect 44380 4676 44772 4732
rect 44828 4676 44838 4732
rect 52042 4676 52052 4732
rect 52108 4676 52724 4732
rect 52780 4676 52790 4732
rect 54618 4676 54628 4732
rect 54684 4676 55188 4732
rect 55244 4676 55254 4732
rect 55412 4620 55468 4788
rect 56084 4732 56140 4788
rect 71988 4732 72044 4788
rect 119812 4732 119868 4788
rect 153300 4732 153356 4788
rect 183316 4732 183372 4788
rect 55530 4676 55540 4732
rect 55596 4676 55644 4732
rect 55700 4676 55748 4732
rect 55804 4676 55814 4732
rect 56084 4676 60228 4732
rect 60284 4676 60294 4732
rect 65258 4676 65268 4732
rect 65324 4676 72044 4732
rect 72202 4676 72212 4732
rect 72268 4676 82292 4732
rect 82348 4676 82358 4732
rect 83038 4676 83076 4732
rect 83132 4676 83142 4732
rect 83290 4676 83300 4732
rect 83356 4676 84980 4732
rect 85036 4676 85046 4732
rect 85418 4676 85428 4732
rect 85484 4676 90804 4732
rect 90860 4676 90870 4732
rect 91018 4676 91028 4732
rect 91084 4676 96180 4732
rect 96236 4676 96246 4732
rect 96394 4676 96404 4732
rect 96460 4676 98644 4732
rect 98700 4676 98710 4732
rect 99194 4676 99204 4732
rect 99260 4676 101780 4732
rect 101836 4676 101846 4732
rect 101994 4676 102004 4732
rect 102060 4676 107492 4732
rect 107548 4676 107558 4732
rect 107706 4676 107716 4732
rect 107772 4676 109396 4732
rect 109452 4676 109462 4732
rect 109858 4676 109868 4732
rect 109924 4676 109972 4732
rect 110028 4676 110076 4732
rect 110132 4676 110142 4732
rect 110506 4676 110516 4732
rect 110572 4676 112644 4732
rect 112700 4676 112710 4732
rect 112858 4676 112868 4732
rect 112924 4676 119588 4732
rect 119644 4676 119654 4732
rect 119812 4676 126756 4732
rect 126812 4676 126822 4732
rect 126970 4676 126980 4732
rect 127036 4676 135660 4732
rect 136490 4676 136500 4732
rect 136556 4676 137116 4732
rect 137172 4676 137182 4732
rect 137274 4676 137284 4732
rect 137340 4676 138964 4732
rect 139020 4676 141148 4732
rect 141204 4676 141214 4732
rect 142650 4676 142660 4732
rect 142716 4676 146692 4732
rect 146748 4676 146758 4732
rect 146906 4676 146916 4732
rect 146972 4676 149772 4732
rect 149828 4676 149838 4732
rect 150042 4676 150052 4732
rect 150108 4676 152292 4732
rect 152348 4676 152358 4732
rect 152618 4676 152628 4732
rect 152684 4676 153356 4732
rect 153514 4676 153524 4732
rect 153636 4676 153646 4732
rect 153738 4676 153748 4732
rect 153804 4676 154644 4732
rect 154700 4676 154710 4732
rect 155978 4676 155988 4732
rect 156044 4676 163604 4732
rect 163660 4676 163670 4732
rect 164186 4676 164196 4732
rect 164252 4676 164300 4732
rect 164356 4676 164404 4732
rect 164460 4676 164470 4732
rect 165106 4676 165116 4732
rect 165228 4676 165238 4732
rect 167962 4676 167972 4732
rect 168028 4676 172564 4732
rect 172620 4676 172630 4732
rect 175812 4676 183372 4732
rect 11498 4564 11508 4620
rect 11564 4564 13300 4620
rect 13356 4564 13366 4620
rect 20131 4564 30884 4620
rect 30940 4564 30950 4620
rect 46890 4564 46900 4620
rect 46956 4564 48748 4620
rect 48804 4564 55468 4620
rect 56186 4564 56196 4620
rect 56252 4564 64820 4620
rect 64876 4564 64886 4620
rect 66826 4564 66836 4620
rect 66892 4564 74116 4620
rect 74172 4564 74182 4620
rect 74330 4564 74340 4620
rect 74396 4564 76692 4620
rect 76748 4564 77700 4620
rect 77756 4564 77766 4620
rect 78250 4564 78260 4620
rect 78316 4564 79716 4620
rect 79772 4564 79782 4620
rect 80490 4564 80500 4620
rect 80556 4564 85652 4620
rect 85708 4564 85718 4620
rect 85866 4564 85876 4620
rect 85932 4564 86212 4620
rect 86268 4564 86278 4620
rect 86538 4564 86548 4620
rect 86604 4564 86996 4620
rect 87052 4564 87062 4620
rect 87434 4564 87444 4620
rect 87500 4564 92708 4620
rect 92764 4564 92774 4620
rect 93370 4564 93380 4620
rect 93436 4564 97188 4620
rect 97244 4564 97254 4620
rect 97402 4564 97412 4620
rect 97468 4564 101892 4620
rect 101948 4564 101958 4620
rect 102106 4564 102116 4620
rect 102172 4564 108724 4620
rect 108780 4564 108790 4620
rect 110618 4564 110628 4620
rect 110684 4564 114772 4620
rect 114828 4564 114838 4620
rect 115546 4564 115556 4620
rect 115612 4564 116116 4620
rect 116172 4564 116182 4620
rect 116330 4564 116340 4620
rect 116396 4564 116434 4620
rect 116554 4564 116564 4620
rect 116620 4564 124292 4620
rect 124348 4564 124358 4620
rect 126756 4564 132132 4620
rect 132188 4564 132198 4620
rect 20131 4508 20187 4564
rect 126756 4508 126812 4564
rect 135604 4508 135660 4676
rect 135818 4564 135828 4620
rect 135884 4564 139188 4620
rect 139244 4564 139254 4620
rect 139402 4564 139412 4620
rect 139468 4564 143612 4620
rect 143668 4564 143678 4620
rect 143770 4564 143780 4620
rect 143836 4564 145572 4620
rect 145628 4564 145638 4620
rect 149594 4564 149604 4620
rect 149660 4564 151284 4620
rect 151340 4564 151350 4620
rect 151498 4564 151508 4620
rect 151564 4564 161364 4620
rect 161420 4564 161430 4620
rect 161690 4564 161700 4620
rect 161756 4564 174356 4620
rect 174412 4564 174422 4620
rect 175812 4508 175868 4676
rect 185556 4620 185612 4788
rect 196644 4732 196700 4788
rect 185770 4676 185780 4732
rect 185836 4676 196700 4732
rect 197838 4676 197876 4732
rect 197932 4676 197942 4732
rect 198426 4676 198436 4732
rect 198492 4676 200284 4732
rect 200340 4676 200350 4732
rect 203251 4676 203756 4732
rect 203812 4676 203822 4732
rect 208562 4676 208572 4732
rect 208628 4676 215068 4732
rect 215124 4676 215134 4732
rect 178714 4564 178724 4620
rect 178780 4564 185612 4620
rect 189214 4564 189252 4620
rect 189308 4564 189318 4620
rect 189550 4564 189588 4620
rect 189644 4564 189654 4620
rect 189914 4564 189924 4620
rect 189980 4564 191996 4620
rect 192052 4564 192062 4620
rect 192154 4564 192164 4620
rect 192220 4564 202020 4620
rect 202076 4564 202086 4620
rect 203251 4508 203307 4676
rect 204586 4564 204596 4620
rect 204652 4564 213724 4620
rect 213780 4564 215236 4620
rect 215292 4564 215302 4620
rect 12954 4452 12964 4508
rect 13020 4452 20187 4508
rect 35914 4452 35924 4508
rect 35980 4452 67956 4508
rect 68012 4452 68022 4508
rect 69066 4452 69076 4508
rect 69132 4452 79492 4508
rect 79548 4452 79558 4508
rect 79706 4452 79716 4508
rect 79772 4452 89572 4508
rect 89628 4452 89638 4508
rect 89796 4452 91252 4508
rect 91308 4452 91318 4508
rect 91420 4452 99147 4508
rect 99418 4452 99428 4508
rect 99484 4452 117460 4508
rect 117516 4452 117526 4508
rect 117898 4452 117908 4508
rect 117964 4452 118132 4508
rect 118188 4452 118198 4508
rect 118346 4452 118356 4508
rect 118412 4452 126812 4508
rect 131002 4452 131012 4508
rect 131068 4452 133476 4508
rect 133532 4452 133542 4508
rect 133690 4452 133700 4508
rect 133756 4452 134372 4508
rect 134428 4452 134438 4508
rect 135604 4452 139860 4508
rect 139916 4452 139926 4508
rect 140970 4452 140980 4508
rect 141036 4452 142996 4508
rect 143052 4452 143062 4508
rect 144330 4452 144340 4508
rect 144396 4452 147700 4508
rect 147756 4452 147766 4508
rect 149482 4452 149492 4508
rect 149548 4452 152852 4508
rect 152908 4452 152918 4508
rect 153290 4452 153300 4508
rect 153356 4452 154868 4508
rect 154924 4452 154934 4508
rect 155642 4452 155652 4508
rect 155708 4452 156100 4508
rect 156156 4452 164556 4508
rect 164612 4452 164622 4508
rect 164714 4452 164724 4508
rect 164780 4452 167860 4508
rect 167916 4452 167926 4508
rect 171994 4452 172004 4508
rect 172060 4452 175868 4508
rect 176932 4452 191100 4508
rect 191156 4452 191166 4508
rect 191370 4452 191380 4508
rect 191436 4452 203307 4508
rect 205594 4452 205604 4508
rect 205660 4452 214172 4508
rect 214228 4452 214238 4508
rect 89796 4396 89852 4452
rect 91420 4396 91476 4452
rect 99091 4396 99147 4452
rect 176932 4396 176988 4452
rect 55290 4340 55300 4396
rect 55356 4340 72548 4396
rect 72604 4340 72614 4396
rect 72762 4340 72772 4396
rect 72828 4340 76468 4396
rect 76524 4340 76534 4396
rect 76682 4340 76692 4396
rect 76748 4340 78260 4396
rect 78316 4340 78326 4396
rect 78474 4340 78484 4396
rect 78540 4340 79044 4396
rect 79100 4340 79110 4396
rect 79818 4340 79828 4396
rect 79884 4340 80052 4396
rect 80108 4340 80118 4396
rect 80500 4340 84308 4396
rect 84364 4340 84374 4396
rect 84606 4340 84644 4396
rect 84700 4340 84710 4396
rect 84868 4340 85988 4396
rect 86044 4340 86054 4396
rect 86538 4340 86548 4396
rect 86604 4340 87668 4396
rect 87724 4340 87734 4396
rect 87882 4340 87892 4396
rect 87948 4340 88900 4396
rect 88956 4340 88966 4396
rect 89114 4340 89124 4396
rect 89180 4340 89852 4396
rect 90010 4340 90020 4396
rect 90076 4340 91476 4396
rect 91690 4340 91700 4396
rect 91756 4340 98700 4396
rect 99091 4340 100212 4396
rect 100268 4340 100278 4396
rect 100538 4340 100548 4396
rect 100604 4340 101220 4396
rect 101276 4340 101286 4396
rect 101434 4340 101444 4396
rect 101500 4340 110516 4396
rect 110572 4340 110582 4396
rect 110730 4340 110740 4396
rect 110796 4340 114324 4396
rect 114380 4340 114390 4396
rect 115658 4340 115668 4396
rect 115724 4340 119812 4396
rect 119868 4340 119878 4396
rect 120138 4340 120148 4396
rect 120204 4340 120372 4396
rect 120428 4340 120438 4396
rect 120586 4340 120596 4396
rect 120652 4340 125412 4396
rect 125468 4340 125478 4396
rect 125626 4340 125636 4396
rect 125692 4340 142772 4396
rect 142828 4340 142838 4396
rect 142996 4340 147252 4396
rect 147308 4340 147318 4396
rect 147466 4340 147476 4396
rect 147532 4340 151956 4396
rect 152012 4340 152022 4396
rect 152282 4340 152292 4396
rect 152348 4340 156380 4396
rect 156538 4340 156548 4396
rect 156604 4340 162596 4396
rect 162652 4340 162662 4396
rect 162810 4340 162820 4396
rect 162876 4340 166964 4396
rect 167020 4340 167030 4396
rect 168970 4340 168980 4396
rect 169036 4340 176932 4396
rect 176988 4340 176998 4396
rect 177146 4340 177156 4396
rect 177212 4340 180404 4396
rect 180460 4340 180470 4396
rect 180618 4340 180628 4396
rect 180684 4340 182980 4396
rect 183036 4340 196364 4396
rect 196420 4340 196430 4396
rect 197754 4340 197764 4396
rect 197820 4340 212492 4396
rect 212548 4340 212558 4396
rect 80500 4284 80556 4340
rect 84868 4284 84924 4340
rect 98644 4284 98700 4340
rect 142996 4284 143052 4340
rect 156324 4284 156380 4340
rect 30314 4228 30324 4284
rect 30380 4228 39396 4284
rect 39452 4228 39462 4284
rect 40170 4228 40180 4284
rect 40236 4228 54964 4284
rect 55020 4228 55030 4284
rect 55178 4228 55188 4284
rect 55244 4228 58772 4284
rect 58828 4228 58838 4284
rect 59108 4228 66612 4284
rect 66668 4228 66678 4284
rect 66836 4228 71428 4284
rect 71484 4228 71494 4284
rect 72090 4228 72100 4284
rect 72156 4228 74228 4284
rect 74284 4228 74294 4284
rect 74442 4228 74452 4284
rect 74508 4228 75908 4284
rect 75964 4228 75974 4284
rect 76122 4228 76132 4284
rect 76188 4228 80556 4284
rect 80714 4228 80724 4284
rect 80780 4228 81620 4284
rect 81676 4228 81686 4284
rect 82170 4228 82180 4284
rect 82236 4228 82964 4284
rect 83020 4228 83030 4284
rect 83514 4228 83524 4284
rect 83580 4228 84924 4284
rect 85530 4228 85540 4284
rect 85596 4228 91420 4284
rect 92138 4228 92148 4284
rect 92204 4228 95284 4284
rect 95340 4228 96404 4284
rect 96460 4228 96470 4284
rect 96730 4228 96740 4284
rect 96796 4228 97188 4284
rect 97244 4228 97254 4284
rect 98644 4228 102340 4284
rect 102396 4228 102406 4284
rect 102554 4228 102564 4284
rect 102620 4228 111524 4284
rect 111580 4228 111590 4284
rect 113082 4228 113092 4284
rect 113148 4228 113540 4284
rect 113596 4228 113606 4284
rect 114090 4228 114100 4284
rect 114156 4228 119364 4284
rect 119420 4228 119430 4284
rect 119578 4228 119588 4284
rect 119644 4228 140980 4284
rect 141036 4228 141046 4284
rect 141194 4228 141204 4284
rect 141260 4228 143052 4284
rect 144340 4228 145348 4284
rect 145404 4228 145414 4284
rect 145562 4228 145572 4284
rect 145628 4228 147700 4284
rect 147756 4228 147766 4284
rect 151050 4228 151060 4284
rect 151116 4228 156100 4284
rect 156156 4228 156166 4284
rect 156324 4228 159460 4284
rect 159516 4228 159526 4284
rect 159898 4228 159908 4284
rect 159964 4228 170436 4284
rect 170492 4228 170502 4284
rect 178238 4228 178276 4284
rect 178332 4228 178342 4284
rect 185994 4228 186004 4284
rect 186060 4228 186340 4284
rect 186396 4228 191492 4284
rect 191548 4228 191558 4284
rect 191706 4228 191716 4284
rect 191772 4228 195636 4284
rect 195692 4228 195702 4284
rect 10042 4116 10052 4172
rect 10108 4116 58884 4172
rect 58940 4116 58950 4172
rect 59108 4060 59164 4228
rect 66836 4172 66892 4228
rect 91364 4172 91420 4228
rect 144340 4172 144396 4228
rect 197764 4172 197820 4340
rect 201674 4228 201684 4284
rect 201740 4228 213220 4284
rect 213276 4228 213286 4284
rect 59434 4116 59444 4172
rect 59500 4116 62580 4172
rect 62636 4116 62646 4172
rect 62794 4116 62804 4172
rect 62860 4116 66892 4172
rect 66948 4116 69188 4172
rect 69244 4116 69254 4172
rect 69412 4116 78036 4172
rect 78092 4116 78102 4172
rect 78250 4116 78260 4172
rect 78316 4116 78354 4172
rect 78820 4116 79716 4172
rect 79772 4116 79782 4172
rect 80042 4116 80052 4172
rect 80108 4116 81508 4172
rect 81564 4116 81574 4172
rect 81834 4116 81844 4172
rect 81900 4116 90020 4172
rect 90076 4116 90086 4172
rect 91364 4116 95564 4172
rect 95722 4116 95732 4172
rect 95788 4116 115444 4172
rect 115500 4116 115510 4172
rect 115658 4116 115668 4172
rect 115724 4116 119924 4172
rect 119980 4116 119990 4172
rect 120138 4116 120148 4172
rect 120204 4116 120764 4172
rect 121258 4116 121268 4172
rect 121324 4116 123956 4172
rect 124012 4116 124022 4172
rect 124142 4116 124180 4172
rect 124236 4116 124246 4172
rect 124394 4116 124404 4172
rect 124460 4116 128100 4172
rect 128156 4116 128166 4172
rect 131002 4116 131012 4172
rect 131068 4116 139412 4172
rect 139468 4116 139478 4172
rect 139626 4116 139636 4172
rect 139692 4116 140644 4172
rect 140700 4116 140710 4172
rect 140858 4116 140868 4172
rect 140924 4116 144396 4172
rect 146458 4116 146468 4172
rect 146524 4116 153076 4172
rect 153132 4116 153142 4172
rect 154410 4116 154420 4172
rect 154476 4116 156548 4172
rect 156604 4116 156614 4172
rect 156762 4116 156772 4172
rect 156828 4116 158676 4172
rect 158732 4116 158742 4172
rect 159226 4116 159236 4172
rect 159292 4116 166516 4172
rect 166572 4116 166582 4172
rect 166740 4116 175028 4172
rect 175084 4116 175094 4172
rect 176698 4116 176708 4172
rect 176764 4116 181860 4172
rect 181916 4116 194516 4172
rect 194572 4116 194582 4172
rect 195290 4116 195300 4172
rect 195356 4116 197820 4172
rect 203802 4116 203812 4172
rect 203868 4116 213108 4172
rect 213164 4116 213174 4172
rect 66948 4060 67004 4116
rect 13290 4004 13300 4060
rect 13356 4004 42196 4060
rect 42252 4004 42262 4060
rect 44436 4004 56196 4060
rect 56252 4004 56262 4060
rect 56970 4004 56980 4060
rect 57036 4004 57092 4060
rect 57148 4004 57158 4060
rect 57306 4004 57316 4060
rect 57372 4004 59164 4060
rect 60666 4004 60676 4060
rect 60732 4004 66276 4060
rect 66332 4004 66342 4060
rect 66490 4004 66500 4060
rect 66556 4004 67004 4060
rect 67386 4004 67396 4060
rect 67452 4004 68292 4060
rect 68348 4004 68358 4060
rect 44436 3948 44492 4004
rect 69412 3948 69468 4116
rect 70746 4004 70756 4060
rect 70812 4004 73108 4060
rect 73164 4004 73174 4060
rect 73322 4004 73332 4060
rect 73388 4004 73556 4060
rect 73612 4004 73622 4060
rect 73994 4004 74004 4060
rect 74060 4004 77364 4060
rect 77420 4004 77430 4060
rect 77802 4004 77812 4060
rect 77868 4004 78596 4060
rect 78652 4004 78662 4060
rect 78820 3948 78876 4116
rect 95508 4060 95564 4116
rect 120708 4060 120764 4116
rect 166740 4060 166796 4116
rect 79370 4004 79380 4060
rect 79436 4004 84196 4060
rect 84252 4004 84262 4060
rect 84410 4004 84420 4060
rect 84476 4004 85876 4060
rect 85932 4004 85942 4060
rect 86426 4004 86436 4060
rect 86492 4004 86660 4060
rect 86716 4004 86726 4060
rect 86874 4004 86884 4060
rect 86940 4004 88340 4060
rect 88396 4004 88406 4060
rect 88890 4004 88900 4060
rect 88956 4004 95172 4060
rect 95228 4004 95238 4060
rect 95508 4004 96740 4060
rect 96796 4004 96806 4060
rect 96954 4004 96964 4060
rect 97020 4004 97412 4060
rect 97468 4004 97478 4060
rect 97626 4004 97636 4060
rect 97692 4004 99540 4060
rect 99596 4004 99606 4060
rect 99978 4004 99988 4060
rect 100044 4004 100940 4060
rect 101210 4004 101220 4060
rect 101276 4004 109172 4060
rect 109228 4004 109238 4060
rect 110282 4004 110292 4060
rect 110348 4004 112756 4060
rect 112812 4004 112822 4060
rect 112970 4004 112980 4060
rect 113036 4004 118468 4060
rect 118524 4004 118534 4060
rect 119354 4004 119364 4060
rect 119420 4004 119924 4060
rect 119980 4004 119990 4060
rect 120138 4004 120148 4060
rect 120204 4004 120260 4060
rect 120316 4004 120326 4060
rect 120708 4004 121156 4060
rect 121212 4004 121222 4060
rect 121370 4004 121380 4060
rect 121436 4004 126980 4060
rect 127036 4004 127046 4060
rect 127194 4004 127204 4060
rect 127260 4004 132244 4060
rect 132300 4004 132310 4060
rect 134138 4004 134148 4060
rect 134204 4004 134596 4060
rect 134652 4004 134662 4060
rect 134810 4004 134820 4060
rect 134876 4004 144228 4060
rect 144284 4004 144294 4060
rect 147466 4004 147476 4060
rect 147532 4004 155316 4060
rect 155372 4004 155382 4060
rect 156211 4004 156660 4060
rect 156716 4004 156726 4060
rect 157434 4004 157444 4060
rect 157500 4004 166796 4060
rect 166954 4004 166964 4060
rect 167020 4004 168644 4060
rect 168700 4004 168710 4060
rect 169194 4004 169204 4060
rect 169260 4004 175924 4060
rect 175980 4004 175990 4060
rect 187450 4004 187460 4060
rect 187516 4004 191268 4060
rect 191324 4004 191334 4060
rect 191482 4004 191492 4060
rect 191548 4004 192052 4060
rect 192108 4004 192118 4060
rect 192266 4004 192276 4060
rect 192332 4004 194292 4060
rect 194348 4004 194358 4060
rect 100884 3948 100940 4004
rect 156211 3948 156267 4004
rect 29194 3892 29204 3948
rect 29260 3892 44492 3948
rect 50362 3892 50372 3948
rect 50428 3892 52388 3948
rect 52444 3892 52454 3948
rect 52714 3892 52724 3948
rect 52780 3892 61684 3948
rect 61740 3892 61750 3948
rect 62570 3892 62580 3948
rect 62636 3892 65268 3948
rect 65324 3892 65334 3948
rect 65482 3892 65492 3948
rect 65548 3892 69468 3948
rect 69626 3892 69636 3948
rect 69692 3892 75796 3948
rect 77018 3892 77028 3948
rect 77084 3892 77140 3948
rect 77196 3892 77206 3948
rect 77354 3892 77364 3948
rect 77420 3892 77700 3948
rect 77756 3892 77766 3948
rect 77914 3892 77924 3948
rect 77980 3892 78876 3948
rect 79146 3892 79156 3948
rect 79212 3892 100660 3948
rect 100716 3892 100726 3948
rect 100884 3892 101108 3948
rect 101164 3892 101174 3948
rect 101322 3892 101332 3948
rect 101388 3892 103460 3948
rect 103516 3892 103526 3948
rect 103786 3892 103796 3948
rect 103852 3892 105028 3948
rect 105084 3892 105094 3948
rect 106922 3892 106932 3948
rect 106988 3892 115556 3948
rect 115612 3892 115622 3948
rect 115770 3892 115780 3948
rect 115836 3892 134260 3948
rect 134316 3892 134326 3948
rect 134484 3892 141204 3948
rect 141260 3892 141270 3948
rect 141530 3892 141540 3948
rect 141596 3892 146580 3948
rect 146636 3892 146646 3948
rect 147354 3892 147364 3948
rect 147420 3892 152180 3948
rect 152236 3892 152246 3948
rect 152506 3892 152516 3948
rect 152572 3892 152852 3948
rect 152908 3892 152918 3948
rect 153066 3892 153076 3948
rect 153132 3892 156267 3948
rect 157546 3892 157556 3948
rect 157612 3892 162820 3948
rect 162876 3892 162886 3948
rect 165162 3892 165172 3948
rect 165228 3892 173124 3948
rect 173180 3892 173190 3948
rect 175242 3892 175252 3948
rect 175308 3892 178724 3948
rect 178780 3892 178790 3948
rect 180170 3892 180180 3948
rect 180236 3892 188020 3948
rect 188076 3892 191380 3948
rect 191436 3892 191446 3948
rect 191706 3892 191716 3948
rect 191772 3892 200676 3948
rect 200732 3892 200742 3948
rect 75740 3836 75796 3892
rect 134484 3836 134540 3892
rect 219200 3836 220000 3864
rect 53834 3780 53844 3836
rect 53900 3780 55076 3836
rect 55132 3780 55142 3836
rect 55290 3780 55300 3836
rect 55356 3780 60340 3836
rect 60396 3780 60406 3836
rect 66686 3780 66724 3836
rect 66780 3780 66790 3836
rect 67022 3780 67060 3836
rect 67116 3780 67126 3836
rect 67274 3780 67284 3836
rect 67340 3780 70532 3836
rect 70588 3780 70598 3836
rect 70746 3780 70756 3836
rect 70812 3780 74676 3836
rect 74732 3780 74742 3836
rect 75310 3780 75348 3836
rect 75404 3780 75414 3836
rect 75740 3780 79044 3836
rect 79100 3780 79110 3836
rect 79370 3780 79380 3836
rect 79436 3780 80276 3836
rect 80332 3780 80342 3836
rect 80714 3780 80724 3836
rect 80780 3780 84420 3836
rect 84476 3780 84486 3836
rect 84634 3780 84644 3836
rect 84700 3780 85428 3836
rect 85484 3780 85494 3836
rect 85642 3780 85652 3836
rect 85708 3780 86548 3836
rect 86604 3780 86614 3836
rect 86874 3780 86884 3836
rect 86940 3780 88340 3836
rect 88396 3780 88406 3836
rect 88554 3780 88564 3836
rect 88620 3780 89348 3836
rect 89404 3780 89414 3836
rect 89562 3780 89572 3836
rect 89628 3780 91588 3836
rect 91644 3780 96964 3836
rect 97020 3780 97030 3836
rect 100762 3780 100772 3836
rect 100828 3780 108948 3836
rect 109004 3780 109014 3836
rect 109162 3780 109172 3836
rect 109228 3780 114996 3836
rect 115052 3780 115062 3836
rect 115210 3780 115220 3836
rect 115276 3780 115314 3836
rect 116078 3780 116116 3836
rect 116172 3780 116182 3836
rect 116330 3780 116340 3836
rect 116396 3780 118524 3836
rect 118682 3780 118692 3836
rect 118748 3780 119252 3836
rect 119308 3780 119318 3836
rect 119690 3780 119700 3836
rect 119756 3780 125636 3836
rect 125692 3780 125702 3836
rect 125850 3780 125860 3836
rect 125916 3780 129556 3836
rect 129612 3780 129622 3836
rect 131982 3780 132020 3836
rect 132076 3780 132086 3836
rect 132682 3780 132692 3836
rect 132748 3780 134540 3836
rect 136154 3780 136164 3836
rect 136220 3780 142772 3836
rect 142828 3780 142838 3836
rect 144442 3780 144452 3836
rect 144508 3780 146916 3836
rect 146972 3780 146982 3836
rect 150388 3780 152964 3836
rect 153020 3780 153030 3836
rect 153178 3780 153188 3836
rect 153244 3780 155092 3836
rect 155148 3780 155158 3836
rect 156202 3780 156212 3836
rect 156268 3780 186564 3836
rect 186620 3780 186630 3836
rect 189466 3780 189476 3836
rect 189532 3780 194068 3836
rect 194124 3780 194134 3836
rect 194926 3780 194964 3836
rect 195020 3780 195030 3836
rect 209598 3780 209636 3836
rect 209692 3780 209702 3836
rect 214890 3780 214900 3836
rect 214956 3780 220000 3836
rect 118468 3724 118524 3780
rect 49690 3668 49700 3724
rect 49756 3668 63700 3724
rect 63756 3668 63766 3724
rect 63924 3668 72996 3724
rect 73052 3668 73062 3724
rect 73210 3668 73220 3724
rect 73276 3668 80948 3724
rect 81004 3668 81014 3724
rect 81162 3668 81172 3724
rect 81228 3668 82516 3724
rect 82572 3668 82582 3724
rect 82730 3668 82740 3724
rect 82796 3668 83188 3724
rect 83244 3668 83254 3724
rect 83402 3668 83412 3724
rect 83468 3668 97748 3724
rect 97804 3668 97814 3724
rect 97962 3668 97972 3724
rect 98028 3668 99204 3724
rect 99260 3668 99270 3724
rect 99754 3668 99764 3724
rect 99820 3668 101444 3724
rect 101500 3668 101510 3724
rect 101658 3668 101668 3724
rect 101724 3668 110628 3724
rect 110684 3668 110694 3724
rect 110842 3668 110852 3724
rect 110908 3668 118244 3724
rect 118300 3668 118310 3724
rect 118468 3668 123060 3724
rect 123116 3668 123126 3724
rect 123274 3668 123284 3724
rect 123340 3668 136724 3724
rect 136780 3668 136790 3724
rect 137386 3668 137396 3724
rect 137452 3668 139524 3724
rect 139580 3668 139590 3724
rect 139738 3668 139748 3724
rect 139804 3668 141428 3724
rect 141484 3668 141494 3724
rect 142202 3668 142212 3724
rect 142268 3668 144004 3724
rect 144060 3668 144070 3724
rect 144218 3668 144228 3724
rect 144284 3668 146132 3724
rect 146188 3668 146198 3724
rect 146682 3668 146692 3724
rect 146748 3668 148708 3724
rect 148764 3668 148774 3724
rect 25274 3556 25284 3612
rect 25340 3556 50372 3612
rect 50428 3556 50438 3612
rect 50586 3556 50596 3612
rect 50652 3556 57316 3612
rect 57372 3556 57382 3612
rect 61674 3556 61684 3612
rect 61740 3556 63700 3612
rect 63756 3556 63766 3612
rect 63924 3500 63980 3668
rect 150388 3612 150444 3780
rect 219200 3752 220000 3780
rect 151050 3668 151060 3724
rect 151116 3668 153188 3724
rect 153244 3668 153254 3724
rect 154298 3668 154308 3724
rect 154364 3668 162820 3724
rect 162876 3668 162886 3724
rect 163034 3668 163044 3724
rect 163100 3668 166740 3724
rect 166796 3668 166806 3724
rect 167066 3668 167076 3724
rect 167132 3668 168420 3724
rect 168476 3668 168486 3724
rect 173226 3668 173236 3724
rect 173292 3668 205716 3724
rect 205772 3668 205782 3724
rect 65370 3556 65380 3612
rect 65436 3556 68404 3612
rect 68460 3556 68470 3612
rect 68618 3556 68628 3612
rect 68684 3556 69188 3612
rect 69244 3556 69254 3612
rect 70074 3556 70084 3612
rect 70140 3556 72772 3612
rect 72828 3556 72838 3612
rect 73210 3556 73220 3612
rect 73276 3556 74788 3612
rect 74844 3556 74854 3612
rect 75002 3556 75012 3612
rect 75068 3556 78260 3612
rect 78316 3556 78326 3612
rect 78428 3556 79156 3612
rect 79212 3556 79222 3612
rect 79370 3556 79380 3612
rect 79436 3556 79474 3612
rect 79930 3556 79940 3612
rect 79996 3556 81956 3612
rect 82012 3556 82022 3612
rect 82842 3556 82852 3612
rect 82908 3556 84084 3612
rect 84140 3556 84150 3612
rect 84298 3556 84308 3612
rect 84364 3556 95620 3612
rect 95676 3556 95686 3612
rect 96058 3556 96068 3612
rect 96124 3556 98084 3612
rect 98140 3556 98150 3612
rect 99054 3556 99092 3612
rect 99148 3556 99158 3612
rect 99866 3556 99876 3612
rect 99932 3556 102116 3612
rect 102172 3556 102182 3612
rect 102666 3556 102676 3612
rect 102732 3556 102844 3612
rect 103450 3556 103460 3612
rect 103516 3556 112420 3612
rect 112476 3556 112486 3612
rect 112634 3556 112644 3612
rect 112700 3556 113652 3612
rect 113708 3556 113718 3612
rect 113876 3556 120428 3612
rect 120698 3556 120708 3612
rect 120764 3556 122388 3612
rect 122444 3556 122454 3612
rect 122938 3556 122948 3612
rect 123004 3556 127707 3612
rect 78428 3500 78484 3556
rect 102788 3500 102844 3556
rect 113876 3500 113932 3556
rect 31210 3444 31220 3500
rect 31276 3444 55300 3500
rect 55356 3444 55366 3500
rect 56196 3444 61908 3500
rect 61964 3444 61974 3500
rect 63028 3444 63980 3500
rect 67274 3444 67284 3500
rect 67340 3444 72884 3500
rect 72940 3444 72950 3500
rect 73098 3444 73108 3500
rect 73164 3444 76692 3500
rect 76748 3444 76758 3500
rect 77242 3444 77252 3500
rect 77308 3444 77644 3500
rect 77774 3444 77812 3500
rect 77868 3444 77878 3500
rect 78026 3444 78036 3500
rect 78092 3444 78484 3500
rect 78586 3444 78596 3500
rect 78652 3444 78932 3500
rect 78988 3444 78998 3500
rect 79146 3444 79156 3500
rect 79212 3444 80388 3500
rect 80444 3444 80454 3500
rect 80602 3444 80612 3500
rect 80668 3444 81396 3500
rect 81452 3444 81462 3500
rect 81722 3444 81732 3500
rect 81788 3444 82068 3500
rect 82124 3444 82134 3500
rect 82618 3444 82628 3500
rect 82684 3444 83524 3500
rect 83580 3444 83590 3500
rect 83738 3444 83748 3500
rect 83804 3444 89012 3500
rect 89068 3444 89078 3500
rect 89226 3444 89236 3500
rect 89292 3444 91364 3500
rect 91420 3444 91430 3500
rect 91578 3444 91588 3500
rect 91644 3444 92316 3500
rect 92474 3444 92484 3500
rect 92540 3444 100716 3500
rect 100874 3444 100884 3500
rect 100940 3444 102564 3500
rect 102620 3444 102630 3500
rect 102788 3444 112980 3500
rect 113036 3444 113046 3500
rect 113194 3444 113204 3500
rect 113260 3444 113932 3500
rect 113988 3444 114772 3500
rect 114828 3444 114838 3500
rect 115182 3444 115220 3500
rect 115276 3444 115286 3500
rect 115658 3444 115668 3500
rect 115724 3444 118020 3500
rect 118076 3444 118086 3500
rect 118346 3444 118356 3500
rect 118412 3444 120148 3500
rect 120204 3444 120214 3500
rect 56196 3388 56252 3444
rect 8698 3332 8708 3388
rect 8764 3332 11172 3388
rect 11228 3332 11238 3388
rect 30650 3332 30660 3388
rect 30716 3332 56252 3388
rect 62244 3332 62804 3388
rect 62860 3332 62870 3388
rect 62244 3276 62300 3332
rect 32442 3220 32452 3276
rect 32508 3220 55300 3276
rect 55356 3220 55366 3276
rect 56186 3220 56196 3276
rect 56252 3220 58772 3276
rect 58828 3220 58838 3276
rect 60330 3220 60340 3276
rect 60396 3220 62300 3276
rect 63028 3164 63084 3444
rect 77588 3388 77644 3444
rect 92260 3388 92316 3444
rect 100660 3388 100716 3444
rect 113988 3388 114044 3444
rect 120372 3388 120428 3556
rect 127651 3500 127707 3556
rect 132468 3556 137844 3612
rect 137900 3556 137910 3612
rect 138618 3556 138628 3612
rect 138684 3556 142548 3612
rect 142604 3556 142614 3612
rect 142762 3556 142772 3612
rect 142828 3556 150444 3612
rect 151050 3556 151060 3612
rect 151116 3556 172676 3612
rect 172732 3556 172742 3612
rect 176138 3556 176148 3612
rect 176204 3556 179787 3612
rect 181290 3556 181300 3612
rect 181356 3556 195860 3612
rect 195916 3556 195926 3612
rect 132468 3500 132524 3556
rect 120586 3444 120596 3500
rect 120652 3444 122444 3500
rect 122602 3444 122612 3500
rect 122668 3444 127428 3500
rect 127484 3444 127494 3500
rect 127651 3444 132524 3500
rect 132682 3444 132692 3500
rect 132748 3444 134036 3500
rect 134092 3444 134102 3500
rect 134250 3444 134260 3500
rect 134316 3444 135212 3500
rect 122388 3388 122444 3444
rect 66154 3332 66164 3388
rect 66220 3332 71876 3388
rect 71932 3332 71942 3388
rect 72762 3332 72772 3388
rect 72828 3332 73500 3388
rect 73658 3332 73668 3388
rect 73724 3332 74900 3388
rect 74956 3332 74966 3388
rect 75180 3332 76804 3388
rect 76860 3332 76870 3388
rect 77588 3332 84252 3388
rect 84410 3332 84420 3388
rect 84476 3332 88900 3388
rect 88956 3332 88966 3388
rect 89124 3332 92036 3388
rect 92092 3332 92102 3388
rect 92260 3332 100604 3388
rect 100660 3332 100996 3388
rect 101052 3332 101062 3388
rect 101322 3332 101332 3388
rect 101388 3332 102676 3388
rect 102732 3332 102742 3388
rect 102890 3332 102900 3388
rect 102956 3332 104468 3388
rect 104524 3332 104534 3388
rect 105476 3332 110404 3388
rect 110460 3332 110470 3388
rect 112298 3332 112308 3388
rect 112364 3332 112756 3388
rect 112812 3332 112822 3388
rect 113502 3332 113540 3388
rect 113596 3332 113606 3388
rect 113754 3332 113764 3388
rect 113820 3332 114044 3388
rect 114314 3332 114324 3388
rect 114380 3332 115108 3388
rect 115164 3332 115174 3388
rect 115434 3332 115444 3388
rect 115500 3332 118020 3388
rect 118076 3332 118086 3388
rect 118234 3332 118244 3388
rect 118300 3332 119140 3388
rect 119196 3332 119206 3388
rect 120372 3332 121604 3388
rect 121660 3332 121670 3388
rect 122388 3332 134484 3388
rect 134540 3332 134550 3388
rect 73444 3276 73500 3332
rect 75180 3276 75236 3332
rect 84196 3276 84252 3332
rect 89124 3276 89180 3332
rect 100548 3276 100604 3332
rect 105476 3276 105532 3332
rect 63690 3220 63700 3276
rect 63756 3220 67172 3276
rect 67228 3220 67238 3276
rect 67386 3220 67396 3276
rect 67452 3220 69972 3276
rect 70028 3220 70038 3276
rect 70186 3220 70196 3276
rect 70252 3220 72884 3276
rect 72940 3220 72950 3276
rect 73444 3220 74340 3276
rect 74396 3220 74406 3276
rect 74554 3220 74564 3276
rect 74620 3220 75236 3276
rect 75338 3220 75348 3276
rect 75404 3220 75572 3276
rect 75628 3220 75638 3276
rect 75786 3220 75796 3276
rect 75852 3220 77476 3276
rect 77532 3220 77542 3276
rect 77690 3220 77700 3276
rect 77756 3220 78260 3276
rect 78316 3220 78326 3276
rect 78474 3220 78484 3276
rect 78540 3220 81284 3276
rect 81340 3220 81350 3276
rect 81498 3220 81508 3276
rect 81564 3220 82740 3276
rect 82796 3220 82806 3276
rect 82954 3220 82964 3276
rect 83020 3220 83972 3276
rect 84028 3220 84038 3276
rect 84196 3220 89180 3276
rect 89786 3220 89796 3276
rect 89852 3220 96292 3276
rect 96348 3220 96358 3276
rect 97850 3220 97860 3276
rect 97916 3220 100212 3276
rect 100268 3220 100278 3276
rect 100548 3220 102004 3276
rect 102060 3220 102070 3276
rect 102666 3220 102676 3276
rect 102732 3220 105532 3276
rect 105690 3220 105700 3276
rect 105756 3220 107380 3276
rect 107436 3220 107446 3276
rect 107594 3220 107604 3276
rect 107660 3220 109060 3276
rect 109116 3220 109126 3276
rect 109274 3220 109284 3276
rect 109340 3220 112644 3276
rect 112700 3220 112710 3276
rect 112858 3220 112868 3276
rect 112924 3220 114716 3276
rect 114874 3220 114884 3276
rect 114940 3220 117236 3276
rect 117292 3220 117302 3276
rect 117562 3220 117572 3276
rect 117628 3220 120260 3276
rect 120316 3220 120326 3276
rect 121146 3220 121156 3276
rect 121212 3220 123284 3276
rect 123340 3220 123350 3276
rect 126756 3220 132244 3276
rect 132300 3220 132310 3276
rect 132570 3220 132580 3276
rect 132636 3220 133700 3276
rect 133756 3220 133766 3276
rect 134138 3220 134148 3276
rect 134204 3220 134820 3276
rect 134876 3220 134886 3276
rect 114660 3164 114716 3220
rect 126756 3164 126812 3220
rect 135156 3164 135212 3444
rect 138068 3444 139636 3500
rect 139692 3444 139702 3500
rect 140298 3444 140308 3500
rect 140364 3444 140756 3500
rect 140812 3444 140822 3500
rect 140970 3444 140980 3500
rect 141036 3444 141316 3500
rect 141372 3444 141382 3500
rect 141754 3444 141764 3500
rect 141820 3444 141830 3500
rect 142762 3444 142772 3500
rect 142828 3444 150948 3500
rect 151004 3444 151014 3500
rect 153178 3444 153188 3500
rect 153244 3444 178836 3500
rect 178892 3444 178902 3500
rect 138068 3388 138124 3444
rect 141764 3388 141820 3444
rect 179731 3388 179787 3556
rect 182634 3444 182644 3500
rect 182700 3444 196756 3500
rect 196812 3444 196822 3500
rect 135706 3332 135716 3388
rect 135772 3332 138124 3388
rect 138506 3332 138516 3388
rect 138572 3332 140644 3388
rect 140700 3332 140710 3388
rect 140858 3332 140868 3388
rect 140924 3332 141540 3388
rect 141596 3332 141606 3388
rect 141764 3332 147700 3388
rect 147756 3332 147766 3388
rect 150154 3332 150164 3388
rect 150220 3332 154476 3388
rect 154634 3332 154644 3388
rect 154700 3332 156492 3388
rect 159674 3332 159684 3388
rect 159740 3332 167076 3388
rect 167132 3332 167142 3388
rect 168634 3332 168644 3388
rect 168700 3332 178948 3388
rect 179004 3332 179014 3388
rect 179731 3332 188804 3388
rect 188860 3332 188870 3388
rect 190138 3332 190148 3388
rect 190204 3332 193116 3388
rect 194058 3332 194068 3388
rect 194124 3332 212660 3388
rect 212716 3332 212726 3388
rect 154420 3276 154476 3332
rect 156436 3276 156492 3332
rect 193060 3276 193116 3332
rect 135370 3220 135380 3276
rect 135436 3220 136052 3276
rect 136108 3220 136500 3276
rect 136556 3220 136566 3276
rect 136714 3220 136724 3276
rect 136780 3220 141764 3276
rect 141820 3220 141830 3276
rect 144218 3220 144228 3276
rect 144284 3220 147812 3276
rect 147868 3220 147878 3276
rect 149482 3220 149492 3276
rect 149548 3220 153020 3276
rect 154420 3220 156212 3276
rect 156268 3220 156278 3276
rect 156436 3220 160468 3276
rect 160524 3220 160534 3276
rect 161130 3220 161140 3276
rect 161196 3220 166404 3276
rect 166460 3220 166470 3276
rect 178042 3220 178052 3276
rect 178108 3220 179396 3276
rect 179452 3220 179620 3276
rect 179676 3220 179686 3276
rect 179946 3220 179956 3276
rect 180012 3220 184660 3276
rect 184716 3220 184726 3276
rect 184996 3220 186900 3276
rect 186956 3220 186966 3276
rect 187310 3220 187348 3276
rect 187404 3220 187414 3276
rect 187786 3220 187796 3276
rect 187852 3220 190932 3276
rect 190988 3220 190998 3276
rect 193060 3220 193956 3276
rect 194012 3220 194022 3276
rect 152964 3164 153020 3220
rect 184996 3164 185052 3220
rect 24490 3108 24500 3164
rect 24556 3108 52500 3164
rect 52556 3108 52566 3164
rect 52714 3108 52724 3164
rect 52780 3108 60004 3164
rect 60060 3108 60070 3164
rect 60218 3108 60228 3164
rect 60284 3108 63084 3164
rect 63914 3108 63924 3164
rect 63980 3108 66052 3164
rect 66108 3108 66118 3164
rect 66266 3108 66276 3164
rect 66332 3108 70532 3164
rect 70588 3108 70598 3164
rect 70746 3108 70756 3164
rect 70812 3108 91476 3164
rect 91532 3108 91542 3164
rect 91700 3108 100660 3164
rect 100716 3108 100726 3164
rect 101098 3108 101108 3164
rect 101164 3108 101220 3164
rect 101276 3108 101286 3164
rect 101546 3108 101556 3164
rect 101612 3108 102452 3164
rect 102508 3108 102518 3164
rect 102890 3108 102900 3164
rect 102956 3108 109172 3164
rect 109228 3108 109238 3164
rect 109396 3108 112308 3164
rect 112364 3108 112374 3164
rect 112522 3108 112532 3164
rect 112588 3108 113428 3164
rect 113484 3108 113494 3164
rect 113642 3108 113652 3164
rect 113708 3108 114604 3164
rect 114660 3108 117124 3164
rect 117180 3108 117190 3164
rect 117338 3108 117348 3164
rect 117404 3108 126812 3164
rect 126868 3108 131460 3164
rect 131516 3108 131526 3164
rect 131674 3108 131684 3164
rect 131740 3108 134596 3164
rect 134652 3108 134662 3164
rect 135156 3108 139636 3164
rect 139692 3108 139702 3164
rect 139850 3108 139860 3164
rect 139916 3108 140532 3164
rect 140588 3108 140598 3164
rect 140746 3108 140756 3164
rect 140812 3108 146244 3164
rect 146300 3108 146310 3164
rect 147690 3108 147700 3164
rect 147756 3108 152907 3164
rect 152964 3108 154532 3164
rect 154588 3108 154598 3164
rect 154746 3108 154756 3164
rect 154812 3108 161140 3164
rect 161196 3108 161206 3164
rect 161354 3108 161364 3164
rect 161420 3108 162260 3164
rect 162316 3108 162326 3164
rect 162474 3108 162484 3164
rect 162540 3108 168756 3164
rect 168812 3108 168822 3164
rect 175914 3108 175924 3164
rect 175980 3108 180068 3164
rect 180124 3108 180134 3164
rect 180282 3108 180292 3164
rect 180348 3108 180964 3164
rect 181020 3108 182140 3164
rect 184202 3108 184212 3164
rect 184268 3108 185052 3164
rect 185210 3108 185220 3164
rect 185276 3108 194740 3164
rect 194796 3108 194806 3164
rect 91700 3052 91756 3108
rect 109396 3052 109452 3108
rect 114548 3052 114604 3108
rect 126868 3052 126924 3108
rect 152851 3052 152907 3108
rect 182084 3052 182140 3108
rect 14186 2996 14196 3052
rect 14252 2996 41748 3052
rect 41804 2996 41814 3052
rect 45098 2996 45108 3052
rect 45164 2996 52780 3052
rect 28186 2884 28196 2940
rect 28252 2884 49588 2940
rect 49644 2884 49654 2940
rect 52724 2828 52780 2996
rect 55076 2996 57092 3052
rect 57148 2996 57158 3052
rect 57418 2996 57428 3052
rect 57484 2996 60116 3052
rect 60172 2996 60182 3052
rect 60890 2996 60900 3052
rect 60956 2996 64148 3052
rect 64204 2996 64214 3052
rect 64698 2996 64708 3052
rect 64764 2996 65772 3052
rect 66938 2996 66948 3052
rect 67004 2996 70756 3052
rect 70812 2996 70822 3052
rect 71642 2996 71652 3052
rect 71708 2996 75012 3052
rect 75068 2996 75078 3052
rect 75180 2996 76692 3052
rect 76748 2996 76758 3052
rect 76906 2996 76916 3052
rect 76972 2996 79940 3052
rect 79996 2996 80006 3052
rect 80154 2996 80164 3052
rect 80220 2996 82516 3052
rect 82572 2996 82582 3052
rect 83178 2996 83188 3052
rect 83244 2996 85428 3052
rect 85484 2996 85494 3052
rect 85642 2996 85652 3052
rect 85708 2996 86212 3052
rect 86268 2996 86278 3052
rect 86426 2996 86436 3052
rect 86492 2996 89684 3052
rect 89740 2996 89750 3052
rect 90570 2996 90580 3052
rect 90636 2996 91756 3052
rect 91914 2996 91924 3052
rect 91980 2996 94164 3052
rect 94220 2996 94230 3052
rect 94378 2996 94388 3052
rect 94444 2996 100996 3052
rect 101052 2996 101062 3052
rect 102330 2996 102340 3052
rect 102396 2996 109452 3052
rect 109610 2996 109620 3052
rect 109676 2996 110404 3052
rect 110460 2996 110470 3052
rect 110618 2996 110628 3052
rect 110684 2996 110740 3052
rect 110796 2996 110806 3052
rect 110954 2996 110964 3052
rect 111020 2996 112196 3052
rect 112252 2996 112262 3052
rect 112410 2996 112420 3052
rect 112476 2996 114324 3052
rect 114380 2996 114390 3052
rect 114548 2996 114772 3052
rect 114828 2996 114838 3052
rect 114986 2996 114996 3052
rect 115052 2996 118468 3052
rect 118524 2996 118534 3052
rect 119018 2996 119028 3052
rect 119084 2996 125636 3052
rect 125692 2996 125702 3052
rect 125850 2996 125860 3052
rect 125916 2996 126924 3052
rect 127082 2996 127092 3052
rect 127148 2996 132468 3052
rect 132524 2996 132534 3052
rect 132681 2996 132691 3052
rect 132747 2996 152628 3052
rect 152684 2996 152694 3052
rect 152851 2996 167076 3052
rect 167132 2996 167142 3052
rect 174122 2996 174132 3052
rect 174188 2996 181860 3052
rect 181916 2996 181926 3052
rect 182084 2996 184268 3052
rect 184398 2996 184436 3052
rect 184492 2996 184502 3052
rect 184771 2996 191716 3052
rect 191772 2996 191782 3052
rect 192266 2996 192276 3052
rect 192332 2996 202468 3052
rect 202524 2996 202534 3052
rect 55076 2940 55132 2996
rect 65716 2940 65772 2996
rect 75180 2940 75236 2996
rect 184212 2940 184268 2996
rect 184771 2940 184827 2996
rect 52938 2884 52948 2940
rect 53004 2884 55132 2940
rect 55290 2884 55300 2940
rect 55356 2884 62580 2940
rect 62636 2884 62646 2940
rect 65716 2884 72324 2940
rect 72380 2884 72390 2940
rect 73434 2884 73444 2940
rect 73500 2884 75236 2940
rect 75348 2884 83860 2940
rect 83916 2884 83926 2940
rect 84074 2884 84084 2940
rect 84140 2884 87668 2940
rect 87724 2884 87734 2940
rect 87882 2884 87892 2940
rect 87948 2884 88788 2940
rect 88844 2884 88854 2940
rect 89002 2884 89012 2940
rect 89068 2884 104132 2940
rect 104188 2884 104198 2940
rect 104346 2884 104356 2940
rect 104412 2884 108724 2940
rect 108780 2884 108790 2940
rect 109050 2884 109060 2940
rect 109116 2884 114548 2940
rect 114604 2884 114614 2940
rect 115098 2884 115108 2940
rect 115164 2884 121044 2940
rect 121100 2884 121110 2940
rect 121258 2884 121268 2940
rect 121324 2884 129332 2940
rect 129388 2884 129398 2940
rect 131898 2884 131908 2940
rect 131964 2884 134148 2940
rect 134204 2884 134214 2940
rect 134586 2884 134596 2940
rect 134652 2884 135492 2940
rect 135548 2884 135558 2940
rect 135818 2884 135828 2940
rect 135884 2884 139076 2940
rect 139132 2884 139142 2940
rect 139402 2884 139412 2940
rect 139468 2884 146020 2940
rect 146076 2884 146086 2940
rect 150042 2884 150052 2940
rect 150108 2884 183092 2940
rect 183148 2884 183158 2940
rect 184212 2884 184827 2940
rect 185854 2884 185892 2940
rect 185948 2884 185958 2940
rect 186106 2884 186116 2940
rect 186172 2884 188916 2940
rect 188972 2884 188982 2940
rect 190026 2884 190036 2940
rect 190092 2884 194068 2940
rect 194124 2884 194134 2940
rect 75348 2828 75404 2884
rect 26954 2772 26964 2828
rect 27020 2772 45892 2828
rect 45948 2772 45958 2828
rect 52724 2772 67060 2828
rect 67116 2772 67126 2828
rect 68394 2772 68404 2828
rect 68460 2772 75404 2828
rect 75674 2772 75684 2828
rect 75740 2772 82404 2828
rect 82460 2772 82470 2828
rect 82618 2772 82628 2828
rect 82684 2772 82852 2828
rect 82908 2772 82918 2828
rect 83178 2772 83188 2828
rect 83244 2772 83636 2828
rect 83692 2772 83702 2828
rect 83962 2772 83972 2828
rect 84028 2772 88676 2828
rect 88732 2772 88742 2828
rect 88890 2772 88900 2828
rect 88956 2772 102228 2828
rect 102284 2772 102294 2828
rect 102666 2772 102676 2828
rect 102732 2772 109620 2828
rect 109676 2772 109686 2828
rect 110282 2772 110292 2828
rect 110348 2772 114436 2828
rect 114492 2772 114502 2828
rect 114884 2772 115164 2828
rect 115322 2772 115332 2828
rect 115388 2772 116900 2828
rect 116956 2772 116966 2828
rect 117226 2772 117236 2828
rect 117292 2772 119028 2828
rect 119084 2772 119094 2828
rect 119466 2772 119476 2828
rect 119532 2772 121828 2828
rect 121884 2772 121894 2828
rect 122154 2772 122164 2828
rect 122220 2772 128772 2828
rect 128828 2772 128838 2828
rect 130890 2772 130900 2828
rect 130956 2772 132692 2828
rect 132748 2772 132758 2828
rect 133018 2772 133028 2828
rect 133084 2772 134036 2828
rect 134092 2772 134102 2828
rect 134250 2772 134260 2828
rect 134316 2772 142548 2828
rect 142604 2772 142614 2828
rect 142762 2772 142772 2828
rect 142828 2772 149268 2828
rect 149324 2772 149334 2828
rect 150266 2772 150276 2828
rect 150332 2772 162484 2828
rect 162540 2772 162550 2828
rect 162670 2772 162708 2828
rect 162764 2772 162774 2828
rect 166282 2772 166292 2828
rect 166348 2772 178220 2828
rect 178378 2772 178388 2828
rect 178444 2772 186004 2828
rect 186060 2772 186070 2828
rect 186218 2772 186228 2828
rect 186284 2772 187628 2828
rect 190586 2772 190596 2828
rect 190652 2772 200676 2828
rect 200732 2772 200742 2828
rect 114884 2716 114940 2772
rect 14746 2660 14756 2716
rect 14812 2660 45220 2716
rect 45276 2660 45286 2716
rect 56970 2660 56980 2716
rect 57036 2660 57316 2716
rect 57372 2660 57382 2716
rect 59882 2660 59892 2716
rect 59948 2660 70084 2716
rect 70140 2660 70150 2716
rect 70298 2660 70308 2716
rect 70364 2660 73332 2716
rect 73388 2660 73398 2716
rect 73546 2660 73556 2716
rect 73612 2660 85764 2716
rect 85820 2660 85830 2716
rect 85978 2660 85988 2716
rect 86044 2660 87108 2716
rect 87164 2660 87174 2716
rect 87658 2660 87668 2716
rect 87724 2660 92372 2716
rect 92428 2660 92438 2716
rect 92586 2660 92596 2716
rect 92652 2660 97524 2716
rect 97580 2660 97590 2716
rect 100426 2660 100436 2716
rect 100492 2660 101052 2716
rect 101434 2660 101444 2716
rect 101500 2660 104356 2716
rect 104412 2660 104422 2716
rect 106586 2660 106596 2716
rect 106652 2660 107492 2716
rect 107548 2660 107558 2716
rect 107706 2660 107716 2716
rect 107772 2660 114940 2716
rect 115108 2716 115164 2772
rect 178164 2716 178220 2772
rect 187572 2716 187628 2772
rect 115108 2660 121380 2716
rect 121482 2660 121492 2716
rect 121548 2660 125860 2716
rect 125916 2660 125926 2716
rect 126074 2660 126084 2716
rect 126140 2660 127652 2716
rect 127708 2660 127718 2716
rect 132122 2660 132132 2716
rect 132188 2660 132692 2716
rect 132748 2660 132758 2716
rect 132906 2660 132916 2716
rect 132972 2660 138516 2716
rect 138572 2660 138582 2716
rect 139626 2660 139636 2716
rect 139692 2660 140756 2716
rect 140812 2660 140822 2716
rect 146010 2660 146020 2716
rect 146076 2660 150164 2716
rect 150220 2660 150230 2716
rect 150612 2660 155988 2716
rect 156044 2660 156054 2716
rect 156201 2660 156211 2716
rect 156267 2660 174132 2716
rect 174188 2660 174198 2716
rect 174346 2660 174356 2716
rect 174412 2660 174450 2716
rect 178164 2660 187348 2716
rect 187404 2660 187414 2716
rect 187572 2660 199780 2716
rect 199836 2660 199846 2716
rect 0 2604 800 2632
rect 100996 2604 101052 2660
rect 121324 2604 121380 2660
rect 150612 2604 150668 2660
rect 0 2548 10276 2604
rect 10332 2548 10342 2604
rect 15418 2548 15428 2604
rect 15484 2548 46564 2604
rect 46620 2548 46630 2604
rect 50698 2548 50708 2604
rect 50764 2548 59668 2604
rect 59724 2548 59734 2604
rect 62458 2548 62468 2604
rect 62524 2548 67004 2604
rect 67162 2548 67172 2604
rect 67228 2548 68628 2604
rect 68684 2548 68694 2604
rect 69066 2548 69076 2604
rect 69132 2548 73947 2604
rect 74330 2548 74340 2604
rect 74396 2548 75684 2604
rect 75740 2548 75750 2604
rect 75898 2548 75908 2604
rect 75964 2548 77924 2604
rect 77980 2548 77990 2604
rect 78810 2548 78820 2604
rect 78876 2548 84644 2604
rect 84700 2548 84710 2604
rect 84858 2548 84868 2604
rect 84924 2548 98644 2604
rect 98700 2548 98710 2604
rect 99278 2548 99316 2604
rect 99372 2548 99382 2604
rect 99540 2548 99764 2604
rect 99820 2548 99830 2604
rect 99978 2548 99988 2604
rect 100044 2548 100772 2604
rect 100828 2548 100838 2604
rect 100996 2548 103348 2604
rect 103404 2548 103414 2604
rect 103674 2548 103684 2604
rect 103740 2548 108388 2604
rect 108444 2548 108454 2604
rect 109050 2548 109060 2604
rect 109116 2548 114772 2604
rect 114828 2548 114838 2604
rect 114996 2548 117684 2604
rect 117740 2548 117750 2604
rect 117898 2548 117908 2604
rect 117964 2548 118002 2604
rect 118122 2548 118132 2604
rect 118188 2548 118916 2604
rect 118972 2548 118982 2604
rect 119914 2548 119924 2604
rect 119980 2548 121156 2604
rect 121212 2548 121222 2604
rect 121324 2548 122164 2604
rect 122220 2548 122230 2604
rect 123050 2548 123060 2604
rect 123116 2548 137732 2604
rect 137788 2548 137798 2604
rect 138170 2548 138180 2604
rect 138236 2548 148260 2604
rect 148316 2548 148326 2604
rect 148484 2548 150668 2604
rect 153178 2548 153188 2604
rect 153244 2548 186340 2604
rect 186396 2548 186406 2604
rect 187002 2548 187012 2604
rect 187068 2548 197540 2604
rect 197596 2548 197606 2604
rect 0 2520 800 2548
rect 66948 2492 67004 2548
rect 73891 2492 73947 2548
rect 99540 2492 99596 2548
rect 114996 2492 115052 2548
rect 148484 2492 148540 2548
rect 16538 2436 16548 2492
rect 16604 2436 50484 2492
rect 50540 2436 50550 2492
rect 54954 2436 54964 2492
rect 55020 2436 59892 2492
rect 59948 2436 59958 2492
rect 60106 2436 60116 2492
rect 60172 2436 61572 2492
rect 61628 2436 61638 2492
rect 61898 2436 61908 2492
rect 61964 2436 65380 2492
rect 65436 2436 65446 2492
rect 66948 2436 67452 2492
rect 67610 2436 67620 2492
rect 67676 2436 71316 2492
rect 71372 2436 71382 2492
rect 71530 2436 71540 2492
rect 71596 2436 72660 2492
rect 72716 2436 72726 2492
rect 73098 2436 73108 2492
rect 73164 2436 73668 2492
rect 73724 2436 73734 2492
rect 73891 2436 86884 2492
rect 86940 2436 86950 2492
rect 87098 2436 87108 2492
rect 87164 2436 90412 2492
rect 90570 2436 90580 2492
rect 90636 2436 96068 2492
rect 96124 2436 96134 2492
rect 96282 2436 96292 2492
rect 96348 2436 99596 2492
rect 99754 2436 99764 2492
rect 99820 2436 101668 2492
rect 101724 2436 101734 2492
rect 102442 2436 102452 2492
rect 102508 2436 106596 2492
rect 106652 2436 106662 2492
rect 106810 2436 106820 2492
rect 106876 2436 111972 2492
rect 112028 2436 112038 2492
rect 112186 2436 112196 2492
rect 112252 2436 115052 2492
rect 115108 2436 125412 2492
rect 125468 2436 125478 2492
rect 125626 2436 125636 2492
rect 125692 2436 127764 2492
rect 127820 2436 127830 2492
rect 127988 2436 145684 2492
rect 145740 2436 145750 2492
rect 147578 2436 147588 2492
rect 147644 2436 148540 2492
rect 149482 2436 149492 2492
rect 149548 2436 152628 2492
rect 152684 2436 152694 2492
rect 154410 2436 154420 2492
rect 154476 2436 154532 2492
rect 154588 2436 154598 2492
rect 154746 2436 154756 2492
rect 154812 2436 155876 2492
rect 155932 2436 155942 2492
rect 156100 2436 178388 2492
rect 178444 2436 178454 2492
rect 179022 2436 179060 2492
rect 179116 2436 179126 2492
rect 179274 2436 179284 2492
rect 179340 2436 180292 2492
rect 180348 2436 180358 2492
rect 183054 2436 183092 2492
rect 183148 2436 183158 2492
rect 184538 2436 184548 2492
rect 184604 2436 185444 2492
rect 185500 2436 186228 2492
rect 186284 2436 186294 2492
rect 186442 2436 186452 2492
rect 186508 2436 189252 2492
rect 189308 2436 189318 2492
rect 189466 2436 189476 2492
rect 189532 2436 201572 2492
rect 201628 2436 201638 2492
rect 67396 2380 67452 2436
rect 90356 2380 90412 2436
rect 115108 2380 115164 2436
rect 127988 2380 128044 2436
rect 156100 2380 156156 2436
rect 37594 2324 37604 2380
rect 37660 2324 52948 2380
rect 53004 2324 53014 2380
rect 53162 2324 53172 2380
rect 53228 2324 56980 2380
rect 57036 2324 57046 2380
rect 57204 2324 61796 2380
rect 61852 2324 61862 2380
rect 62010 2324 62020 2380
rect 62076 2324 65492 2380
rect 65548 2324 65558 2380
rect 67396 2324 68740 2380
rect 68796 2324 72436 2380
rect 72492 2324 72502 2380
rect 72650 2324 72660 2380
rect 72716 2324 79828 2380
rect 79884 2324 79894 2380
rect 80798 2324 80836 2380
rect 80892 2324 80902 2380
rect 81162 2324 81172 2380
rect 81228 2324 81396 2380
rect 81452 2324 81462 2380
rect 81610 2324 81620 2380
rect 81676 2324 82068 2380
rect 82124 2324 82134 2380
rect 82282 2324 82292 2380
rect 82348 2324 90132 2380
rect 90188 2324 90198 2380
rect 90356 2324 92596 2380
rect 92652 2324 92662 2380
rect 94154 2324 94164 2380
rect 94220 2324 102340 2380
rect 102396 2324 102406 2380
rect 102564 2324 103180 2380
rect 103338 2324 103348 2380
rect 103404 2324 103684 2380
rect 103740 2324 103750 2380
rect 103898 2324 103908 2380
rect 103964 2324 108948 2380
rect 109004 2324 109014 2380
rect 109161 2324 109171 2380
rect 109227 2324 115164 2380
rect 115546 2324 115556 2380
rect 115612 2324 117236 2380
rect 117292 2324 117302 2380
rect 117450 2324 117460 2380
rect 117516 2324 118356 2380
rect 118412 2324 118422 2380
rect 118570 2324 118580 2380
rect 118636 2324 120372 2380
rect 120428 2324 120438 2380
rect 120586 2324 120596 2380
rect 120652 2324 120820 2380
rect 120876 2324 120886 2380
rect 121594 2324 121604 2380
rect 121660 2324 122052 2380
rect 122108 2324 122118 2380
rect 122602 2324 122612 2380
rect 122668 2324 128044 2380
rect 129546 2324 129556 2380
rect 129612 2324 133364 2380
rect 133420 2324 133430 2380
rect 134222 2324 134260 2380
rect 134316 2324 134326 2380
rect 134586 2324 134596 2380
rect 134652 2324 136388 2380
rect 136444 2324 136454 2380
rect 137722 2324 137732 2380
rect 137788 2324 140980 2380
rect 141036 2324 141046 2380
rect 141530 2324 141540 2380
rect 141596 2324 150612 2380
rect 150668 2324 150678 2380
rect 152506 2324 152516 2380
rect 152572 2324 156156 2380
rect 157770 2324 157780 2380
rect 157836 2324 161028 2380
rect 161084 2324 161094 2380
rect 161241 2324 161251 2380
rect 161307 2324 165732 2380
rect 165788 2324 165798 2380
rect 167066 2324 167076 2380
rect 167132 2324 173124 2380
rect 173180 2324 173190 2380
rect 174906 2324 174916 2380
rect 174972 2324 186676 2380
rect 186732 2324 186742 2380
rect 187562 2324 187572 2380
rect 187628 2324 190372 2380
rect 190428 2324 190438 2380
rect 190586 2324 190596 2380
rect 190652 2324 198100 2380
rect 198156 2324 198166 2380
rect 57204 2268 57260 2324
rect 102564 2268 102620 2324
rect 103124 2268 103180 2324
rect 41626 2212 41636 2268
rect 41692 2212 53508 2268
rect 53564 2212 53574 2268
rect 56858 2212 56868 2268
rect 56924 2212 57260 2268
rect 58650 2212 58660 2268
rect 58716 2212 61292 2268
rect 62121 2212 62131 2268
rect 62187 2212 62412 2268
rect 62570 2212 62580 2268
rect 62636 2212 67620 2268
rect 67676 2212 67686 2268
rect 67834 2212 67844 2268
rect 67900 2212 75236 2268
rect 75292 2212 75302 2268
rect 75562 2212 75572 2268
rect 75628 2212 82068 2268
rect 82124 2212 82134 2268
rect 82291 2212 83636 2268
rect 83692 2212 83702 2268
rect 83850 2212 83860 2268
rect 83916 2212 85764 2268
rect 85820 2212 85830 2268
rect 85978 2212 85988 2268
rect 86044 2212 87220 2268
rect 87276 2212 87286 2268
rect 87434 2212 87444 2268
rect 87500 2212 88788 2268
rect 88844 2212 88854 2268
rect 89226 2212 89236 2268
rect 89292 2212 93940 2268
rect 93996 2212 94006 2268
rect 95610 2212 95620 2268
rect 95676 2212 95732 2268
rect 95788 2212 95798 2268
rect 95946 2212 95956 2268
rect 96012 2212 98196 2268
rect 98252 2212 98262 2268
rect 99530 2212 99540 2268
rect 99596 2212 101556 2268
rect 101612 2212 101622 2268
rect 101770 2212 101780 2268
rect 101836 2212 102620 2268
rect 102862 2212 102900 2268
rect 102956 2212 102966 2268
rect 103124 2212 104244 2268
rect 104300 2212 104310 2268
rect 104458 2212 104468 2268
rect 104524 2212 113204 2268
rect 113260 2212 113270 2268
rect 113642 2212 113652 2268
rect 113708 2212 114100 2268
rect 114156 2212 114166 2268
rect 114314 2212 114324 2268
rect 114380 2212 119140 2268
rect 119196 2212 119206 2268
rect 119354 2212 119364 2268
rect 119420 2212 120932 2268
rect 120988 2212 120998 2268
rect 121146 2212 121156 2268
rect 121212 2212 122500 2268
rect 122556 2212 122566 2268
rect 123834 2212 123844 2268
rect 123900 2212 132804 2268
rect 132860 2212 132870 2268
rect 133028 2212 134148 2268
rect 134204 2212 134214 2268
rect 134474 2212 134484 2268
rect 134540 2212 136276 2268
rect 136332 2212 136342 2268
rect 136714 2212 136724 2268
rect 136780 2212 139860 2268
rect 139916 2212 139926 2268
rect 140074 2212 140084 2268
rect 140140 2212 150052 2268
rect 150108 2212 150118 2268
rect 151162 2212 151172 2268
rect 151228 2212 152852 2268
rect 152908 2212 152918 2268
rect 153822 2212 153860 2268
rect 153916 2212 153926 2268
rect 156211 2212 177996 2268
rect 178154 2212 178164 2268
rect 178220 2212 193844 2268
rect 193900 2212 193910 2268
rect 203550 2212 203588 2268
rect 203644 2212 203654 2268
rect 61236 2156 61292 2212
rect 62356 2156 62412 2212
rect 82291 2156 82347 2212
rect 133028 2156 133084 2212
rect 156211 2156 156267 2212
rect 177940 2156 177996 2212
rect 45882 2100 45892 2156
rect 45948 2100 57988 2156
rect 58044 2100 58054 2156
rect 61236 2100 62132 2156
rect 62188 2100 62198 2156
rect 62356 2100 64708 2156
rect 64764 2100 64774 2156
rect 64932 2100 68292 2156
rect 68348 2100 68358 2156
rect 69626 2100 69636 2156
rect 69692 2100 71932 2156
rect 72090 2100 72100 2156
rect 72156 2100 73220 2156
rect 73276 2100 73286 2156
rect 73434 2100 73444 2156
rect 73500 2100 75012 2156
rect 75068 2100 75078 2156
rect 75226 2100 75236 2156
rect 75292 2100 77700 2156
rect 77756 2100 77766 2156
rect 77914 2100 77924 2156
rect 77980 2100 82347 2156
rect 82506 2100 82516 2156
rect 82572 2100 83076 2156
rect 83132 2100 83142 2156
rect 83402 2100 83412 2156
rect 83468 2100 84868 2156
rect 84924 2100 84934 2156
rect 85194 2100 85204 2156
rect 85260 2100 86100 2156
rect 86156 2100 86166 2156
rect 86314 2100 86324 2156
rect 86380 2100 90244 2156
rect 90300 2100 90310 2156
rect 91130 2100 91140 2156
rect 91196 2100 91924 2156
rect 91980 2100 91990 2156
rect 92138 2100 92148 2156
rect 92204 2100 94388 2156
rect 94444 2100 94454 2156
rect 94602 2100 94612 2156
rect 94668 2100 96292 2156
rect 96348 2100 96358 2156
rect 96506 2100 96516 2156
rect 96572 2100 96610 2156
rect 97626 2100 97636 2156
rect 97692 2100 113316 2156
rect 113372 2100 113382 2156
rect 113530 2100 113540 2156
rect 113596 2100 117236 2156
rect 117292 2100 117302 2156
rect 117562 2100 117572 2156
rect 117628 2100 127652 2156
rect 127708 2100 127718 2156
rect 127866 2100 127876 2156
rect 127932 2100 133084 2156
rect 133242 2100 133252 2156
rect 133308 2100 137732 2156
rect 137788 2100 137798 2156
rect 141530 2100 141540 2156
rect 141596 2100 144900 2156
rect 144956 2100 144966 2156
rect 148922 2100 148932 2156
rect 148988 2100 156267 2156
rect 159114 2100 159124 2156
rect 159180 2100 161028 2156
rect 161084 2100 161094 2156
rect 161251 2100 177716 2156
rect 177772 2100 177782 2156
rect 177940 2100 179284 2156
rect 179340 2100 179350 2156
rect 184874 2100 184884 2156
rect 184940 2100 187460 2156
rect 187516 2100 187526 2156
rect 188654 2100 188692 2156
rect 188748 2100 188758 2156
rect 188906 2100 188916 2156
rect 188972 2100 198884 2156
rect 198940 2100 198950 2156
rect 64932 2044 64988 2100
rect 71876 2044 71932 2100
rect 96516 2044 96572 2100
rect 161251 2044 161307 2100
rect 43306 1988 43316 2044
rect 43372 1988 56980 2044
rect 57036 1988 57046 2044
rect 57866 1988 57876 2044
rect 57932 1988 60788 2044
rect 60844 1988 60854 2044
rect 61786 1988 61796 2044
rect 61852 1988 64988 2044
rect 65146 1988 65156 2044
rect 65212 1988 71652 2044
rect 71708 1988 71718 2044
rect 71876 1988 75460 2044
rect 75516 1988 75526 2044
rect 75674 1988 75684 2044
rect 75740 1988 76468 2044
rect 76524 1988 76534 2044
rect 76682 1988 76692 2044
rect 76748 1988 81396 2044
rect 81452 1988 81462 2044
rect 81722 1988 81732 2044
rect 81788 1988 94276 2044
rect 94332 1988 94342 2044
rect 94490 1988 94500 2044
rect 94556 1988 96572 2044
rect 98858 1988 98868 2044
rect 98924 1988 101332 2044
rect 101388 1988 101398 2044
rect 101546 1988 101556 2044
rect 101612 1988 101650 2044
rect 101994 1988 102004 2044
rect 102060 1988 108388 2044
rect 108444 1988 108454 2044
rect 108602 1988 108612 2044
rect 108668 1988 109732 2044
rect 109788 1988 109798 2044
rect 109946 1988 109956 2044
rect 110012 1988 113316 2044
rect 113372 1988 113382 2044
rect 113614 1988 113652 2044
rect 113708 1988 113718 2044
rect 113866 1988 113876 2044
rect 113932 1988 114604 2044
rect 114762 1988 114772 2044
rect 114828 1988 120932 2044
rect 120988 1988 120998 2044
rect 121146 1988 121156 2044
rect 121212 1988 124796 2044
rect 125850 1988 125860 2044
rect 125916 1988 133196 2044
rect 133354 1988 133364 2044
rect 133420 1988 147924 2044
rect 147980 1988 147990 2044
rect 150042 1988 150052 2044
rect 150108 1988 150724 2044
rect 150780 1988 150790 2044
rect 151050 1988 151060 2044
rect 151116 1988 161307 2044
rect 162250 1988 162260 2044
rect 162316 1988 165172 2044
rect 165228 1988 165238 2044
rect 165386 1988 165396 2044
rect 165452 1988 168084 2044
rect 168140 1988 168150 2044
rect 172890 1988 172900 2044
rect 172956 1988 178164 2044
rect 178220 1988 178230 2044
rect 178826 1988 178836 2044
rect 178892 1988 210756 2044
rect 210812 1988 210822 2044
rect 114548 1932 114604 1988
rect 48346 1876 48356 1932
rect 48412 1876 52724 1932
rect 52780 1876 52790 1932
rect 56186 1876 56196 1932
rect 56252 1876 60116 1932
rect 60172 1876 60182 1932
rect 62430 1876 62468 1932
rect 62524 1876 62534 1932
rect 62766 1876 62804 1932
rect 62860 1876 62870 1932
rect 65258 1876 65268 1932
rect 65324 1876 74396 1932
rect 74526 1876 74564 1932
rect 74620 1876 74630 1932
rect 75450 1876 75460 1932
rect 75516 1876 80724 1932
rect 80780 1876 80790 1932
rect 80938 1876 80948 1932
rect 81004 1876 81956 1932
rect 82012 1876 82022 1932
rect 82282 1876 82292 1932
rect 82348 1876 84308 1932
rect 84410 1876 84420 1932
rect 84476 1876 85540 1932
rect 85596 1876 85606 1932
rect 85754 1876 85764 1932
rect 85820 1876 89516 1932
rect 89674 1876 89684 1932
rect 89740 1876 114324 1932
rect 114380 1876 114390 1932
rect 114548 1876 115164 1932
rect 115434 1876 115444 1932
rect 115500 1876 118356 1932
rect 118412 1876 118422 1932
rect 119354 1876 119364 1932
rect 119420 1876 123844 1932
rect 123900 1876 123910 1932
rect 74340 1820 74396 1876
rect 84252 1820 84308 1876
rect 89460 1820 89516 1876
rect 115108 1820 115164 1876
rect 124740 1820 124796 1988
rect 133140 1932 133196 1988
rect 125850 1876 125860 1932
rect 125916 1876 133084 1932
rect 133140 1876 136164 1932
rect 136220 1876 136230 1932
rect 136378 1876 136388 1932
rect 136444 1876 143444 1932
rect 143500 1876 143510 1932
rect 144451 1876 147364 1932
rect 147420 1876 147430 1932
rect 148250 1876 148260 1932
rect 148316 1876 150836 1932
rect 150892 1876 150902 1932
rect 151050 1876 151060 1932
rect 151116 1876 151508 1932
rect 151564 1876 151574 1932
rect 151722 1876 151732 1932
rect 151788 1876 154420 1932
rect 154476 1876 154486 1932
rect 155978 1876 155988 1932
rect 156044 1876 159572 1932
rect 159628 1876 159638 1932
rect 162362 1876 162372 1932
rect 162428 1876 164724 1932
rect 164780 1876 164790 1932
rect 164938 1876 164948 1932
rect 165004 1876 167748 1932
rect 167804 1876 167814 1932
rect 167962 1876 167972 1932
rect 168028 1876 189700 1932
rect 189756 1876 189766 1932
rect 189914 1876 189924 1932
rect 189980 1876 201908 1932
rect 201964 1876 201974 1932
rect 133028 1820 133084 1876
rect 55626 1764 55636 1820
rect 55692 1764 60676 1820
rect 60732 1764 60742 1820
rect 65370 1764 65380 1820
rect 65436 1764 69076 1820
rect 69132 1764 69142 1820
rect 70858 1764 70868 1820
rect 70924 1764 72996 1820
rect 73052 1764 73062 1820
rect 74340 1764 83972 1820
rect 84028 1764 84038 1820
rect 84252 1764 88452 1820
rect 88508 1764 88518 1820
rect 88666 1764 88676 1820
rect 88732 1764 89236 1820
rect 89292 1764 89302 1820
rect 89460 1764 93380 1820
rect 93436 1764 93446 1820
rect 94042 1764 94052 1820
rect 94108 1764 96236 1820
rect 96618 1764 96628 1820
rect 96684 1764 97412 1820
rect 97468 1764 97478 1820
rect 97626 1764 97636 1820
rect 97692 1764 99652 1820
rect 99708 1764 99718 1820
rect 99866 1764 99876 1820
rect 99932 1764 102788 1820
rect 102844 1764 102854 1820
rect 103002 1764 103012 1820
rect 103068 1764 109004 1820
rect 109162 1764 109172 1820
rect 109228 1764 114772 1820
rect 114828 1764 114838 1820
rect 115108 1764 115668 1820
rect 115724 1764 115734 1820
rect 115882 1764 115892 1820
rect 115948 1764 121044 1820
rect 121100 1764 121110 1820
rect 121258 1764 121268 1820
rect 121324 1764 124516 1820
rect 124572 1764 124582 1820
rect 124740 1764 128212 1820
rect 128268 1764 128278 1820
rect 129322 1764 129332 1820
rect 129388 1764 132804 1820
rect 132860 1764 132870 1820
rect 133028 1764 138180 1820
rect 138236 1764 138246 1820
rect 96180 1708 96236 1764
rect 108948 1708 109004 1764
rect 144451 1708 144507 1876
rect 145786 1764 145796 1820
rect 145852 1764 152404 1820
rect 152460 1764 152470 1820
rect 154634 1764 154644 1820
rect 154700 1764 157780 1820
rect 157836 1764 157846 1820
rect 162810 1764 162820 1820
rect 162876 1764 188468 1820
rect 188524 1764 188534 1820
rect 188682 1764 188692 1820
rect 188748 1764 191716 1820
rect 191772 1764 191782 1820
rect 26394 1652 26404 1708
rect 26460 1652 53004 1708
rect 53162 1652 53172 1708
rect 53228 1652 54628 1708
rect 54684 1652 54694 1708
rect 56410 1652 56420 1708
rect 56476 1652 57428 1708
rect 57484 1652 57494 1708
rect 60442 1652 60452 1708
rect 60508 1652 75236 1708
rect 75292 1652 75302 1708
rect 75450 1652 75460 1708
rect 75516 1652 79716 1708
rect 79772 1652 79782 1708
rect 80042 1652 80052 1708
rect 80108 1652 81172 1708
rect 81228 1652 81238 1708
rect 81386 1652 81396 1708
rect 81452 1652 85428 1708
rect 85484 1652 85494 1708
rect 85642 1652 85652 1708
rect 85708 1652 86884 1708
rect 86940 1652 86950 1708
rect 88330 1652 88340 1708
rect 88396 1652 95956 1708
rect 96012 1652 96022 1708
rect 96180 1652 99764 1708
rect 99820 1652 99830 1708
rect 100090 1652 100100 1708
rect 100156 1652 101220 1708
rect 101276 1652 101286 1708
rect 103114 1652 103124 1708
rect 103180 1652 108388 1708
rect 108444 1652 108454 1708
rect 108948 1652 114996 1708
rect 115052 1652 115062 1708
rect 115220 1652 118748 1708
rect 118906 1652 118916 1708
rect 118972 1652 120932 1708
rect 120988 1652 120998 1708
rect 121156 1652 126924 1708
rect 127194 1652 127204 1708
rect 127260 1652 131796 1708
rect 131852 1652 131862 1708
rect 132010 1652 132020 1708
rect 132076 1652 132804 1708
rect 132860 1652 132870 1708
rect 133018 1652 133028 1708
rect 133084 1652 133700 1708
rect 133756 1652 133766 1708
rect 133914 1652 133924 1708
rect 133980 1652 134820 1708
rect 134876 1652 134886 1708
rect 135044 1652 136164 1708
rect 136220 1652 136230 1708
rect 138506 1652 138516 1708
rect 138572 1652 144507 1708
rect 147354 1652 147364 1708
rect 147420 1652 147924 1708
rect 147980 1652 147990 1708
rect 150238 1652 150276 1708
rect 150332 1652 150342 1708
rect 150714 1652 150724 1708
rect 150780 1652 155988 1708
rect 156044 1652 156054 1708
rect 8250 1540 8260 1596
rect 8316 1540 9940 1596
rect 9996 1540 10006 1596
rect 11050 1540 11060 1596
rect 11116 1540 14420 1596
rect 14476 1540 14486 1596
rect 17742 1540 17780 1596
rect 17836 1540 17846 1596
rect 22670 1540 22708 1596
rect 22764 1540 22774 1596
rect 28718 1540 28756 1596
rect 28812 1540 28822 1596
rect 29950 1540 29988 1596
rect 30044 1540 30054 1596
rect 34206 1540 34244 1596
rect 34300 1540 34310 1596
rect 35438 1540 35476 1596
rect 35532 1540 35542 1596
rect 44762 1540 44772 1596
rect 44828 1540 46452 1596
rect 46508 1540 46518 1596
rect 47674 1540 47684 1596
rect 47740 1540 52164 1596
rect 52220 1540 52230 1596
rect 52948 1484 53004 1652
rect 115220 1596 115276 1652
rect 118692 1596 118748 1652
rect 121156 1596 121212 1652
rect 126868 1596 126924 1652
rect 55066 1540 55076 1596
rect 55132 1540 55972 1596
rect 56028 1540 56038 1596
rect 62121 1540 62131 1596
rect 62187 1540 62244 1596
rect 62300 1540 62310 1596
rect 62458 1540 62468 1596
rect 62524 1540 65940 1596
rect 65996 1540 66006 1596
rect 66266 1540 66276 1596
rect 66332 1540 71540 1596
rect 71596 1540 71606 1596
rect 71754 1540 71764 1596
rect 71820 1540 90356 1596
rect 90412 1540 90422 1596
rect 90570 1540 90580 1596
rect 90636 1540 100492 1596
rect 100650 1540 100660 1596
rect 100716 1540 102452 1596
rect 102508 1540 102518 1596
rect 104010 1540 104020 1596
rect 104076 1540 108668 1596
rect 108826 1540 108836 1596
rect 108892 1540 110292 1596
rect 110348 1540 110358 1596
rect 111514 1540 111524 1596
rect 111580 1540 115276 1596
rect 115546 1540 115556 1596
rect 115612 1540 115892 1596
rect 115948 1540 115958 1596
rect 116106 1540 116116 1596
rect 116172 1540 116564 1596
rect 116620 1540 116630 1596
rect 117786 1540 117796 1596
rect 117852 1540 118020 1596
rect 118076 1540 118086 1596
rect 118430 1540 118468 1596
rect 118524 1540 118534 1596
rect 118692 1540 120484 1596
rect 120540 1540 120550 1596
rect 120698 1540 120708 1596
rect 120764 1540 121212 1596
rect 121268 1540 124628 1596
rect 124684 1540 124694 1596
rect 126868 1540 132747 1596
rect 132906 1540 132916 1596
rect 132972 1540 134372 1596
rect 134428 1540 134438 1596
rect 100436 1484 100492 1540
rect 108612 1484 108668 1540
rect 121268 1484 121324 1540
rect 132691 1484 132747 1540
rect 135044 1484 135100 1652
rect 156211 1596 156268 1708
rect 156426 1652 156436 1708
rect 156492 1652 194628 1708
rect 194684 1652 194694 1708
rect 196410 1652 196420 1708
rect 196476 1652 197932 1708
rect 135706 1540 135716 1596
rect 135772 1540 142436 1596
rect 142492 1540 142502 1596
rect 143406 1540 143444 1596
rect 143500 1540 143510 1596
rect 143966 1540 144004 1596
rect 144060 1540 144070 1596
rect 144442 1540 144452 1596
rect 144508 1540 145012 1596
rect 145068 1540 145078 1596
rect 145198 1540 145236 1596
rect 145292 1540 145302 1596
rect 146122 1540 146132 1596
rect 146188 1540 154308 1596
rect 154364 1540 154374 1596
rect 154532 1540 159684 1596
rect 159740 1540 159750 1596
rect 160458 1540 160468 1596
rect 160524 1540 162708 1596
rect 162764 1540 162774 1596
rect 162922 1540 162932 1596
rect 162988 1540 163156 1596
rect 163212 1540 163222 1596
rect 164714 1540 164724 1596
rect 164780 1540 164836 1596
rect 164892 1540 164902 1596
rect 166478 1540 166516 1596
rect 166572 1540 166582 1596
rect 167402 1540 167412 1596
rect 167468 1540 170212 1596
rect 170268 1540 170278 1596
rect 175102 1540 175140 1596
rect 175196 1540 175206 1596
rect 179358 1540 179396 1596
rect 179452 1540 179462 1596
rect 180394 1540 180404 1596
rect 180460 1540 181188 1596
rect 181244 1540 181254 1596
rect 186078 1540 186116 1596
rect 186172 1540 186182 1596
rect 187870 1540 187908 1596
rect 187964 1540 187974 1596
rect 189102 1540 189140 1596
rect 189196 1540 189206 1596
rect 196410 1540 196420 1596
rect 196476 1540 197652 1596
rect 197708 1540 197718 1596
rect 154532 1484 154588 1540
rect 197876 1484 197932 1652
rect 199406 1540 199444 1596
rect 199500 1540 199510 1596
rect 200078 1540 200116 1596
rect 200172 1540 200182 1596
rect 204334 1540 204372 1596
rect 204428 1540 204438 1596
rect 211614 1540 211652 1596
rect 211708 1540 211718 1596
rect 8138 1428 8148 1484
rect 8204 1428 10500 1484
rect 10556 1428 10566 1484
rect 11722 1428 11732 1484
rect 11788 1428 19348 1484
rect 19404 1428 19414 1484
rect 25134 1428 25172 1484
rect 25228 1428 25238 1484
rect 39050 1428 39060 1484
rect 39116 1428 45892 1484
rect 45948 1428 45958 1484
rect 49466 1428 49476 1484
rect 49532 1428 49700 1484
rect 49756 1428 49766 1484
rect 52948 1428 59780 1484
rect 59836 1428 59846 1484
rect 60330 1428 60340 1484
rect 60396 1428 70532 1484
rect 70588 1428 70598 1484
rect 71950 1428 71988 1484
rect 72044 1428 72054 1484
rect 72324 1428 74900 1484
rect 74956 1428 74966 1484
rect 75180 1428 76244 1484
rect 76300 1428 76310 1484
rect 76458 1428 76468 1484
rect 76524 1428 77252 1484
rect 77308 1428 77318 1484
rect 77466 1428 77476 1484
rect 77532 1428 79324 1484
rect 79454 1428 79492 1484
rect 79548 1428 79558 1484
rect 79706 1428 79716 1484
rect 79772 1428 86996 1484
rect 87052 1428 87062 1484
rect 87210 1428 87220 1484
rect 87276 1428 87780 1484
rect 87994 1428 88004 1484
rect 88060 1428 88676 1484
rect 88732 1428 88742 1484
rect 88890 1428 88900 1484
rect 88956 1428 100380 1484
rect 100436 1428 108556 1484
rect 108612 1428 120820 1484
rect 120876 1428 120886 1484
rect 121034 1428 121044 1484
rect 121100 1428 121324 1484
rect 121594 1428 121604 1484
rect 121660 1428 122108 1484
rect 122490 1428 122500 1484
rect 122556 1428 129332 1484
rect 129388 1428 129398 1484
rect 132691 1428 135100 1484
rect 135594 1428 135604 1484
rect 135660 1428 138628 1484
rect 138684 1428 138694 1484
rect 138964 1428 141652 1484
rect 141708 1428 141718 1484
rect 142202 1428 142212 1484
rect 142268 1428 144340 1484
rect 144396 1428 144406 1484
rect 144666 1428 144676 1484
rect 144732 1428 147924 1484
rect 147980 1428 147990 1484
rect 148260 1428 152180 1484
rect 152236 1428 152246 1484
rect 152842 1428 152852 1484
rect 152908 1428 154588 1484
rect 154858 1428 154868 1484
rect 154924 1428 164500 1484
rect 164556 1428 164566 1484
rect 164714 1428 164724 1484
rect 164780 1428 167748 1484
rect 167804 1428 167814 1484
rect 180590 1428 180628 1484
rect 180684 1428 180694 1484
rect 190586 1428 190596 1484
rect 190652 1428 196532 1484
rect 196588 1428 196598 1484
rect 197876 1428 201908 1484
rect 201964 1428 201974 1484
rect 209738 1428 209748 1484
rect 209804 1428 219044 1484
rect 219100 1428 219110 1484
rect 8026 1316 8036 1372
rect 8092 1316 11956 1372
rect 12012 1316 12022 1372
rect 25610 1316 25620 1372
rect 25676 1316 43988 1372
rect 44044 1316 44054 1372
rect 44212 1316 45220 1372
rect 45276 1316 45286 1372
rect 48906 1316 48916 1372
rect 48972 1316 53620 1372
rect 53676 1316 53686 1372
rect 53844 1316 62244 1372
rect 62300 1316 62310 1372
rect 62570 1316 62580 1372
rect 62636 1316 66836 1372
rect 66892 1316 66902 1372
rect 67050 1316 67060 1372
rect 67116 1316 72100 1372
rect 72156 1316 72166 1372
rect 44212 1260 44268 1316
rect 9258 1204 9268 1260
rect 9324 1204 11396 1260
rect 11452 1204 11462 1260
rect 33646 1204 33684 1260
rect 33740 1204 33750 1260
rect 35578 1204 35588 1260
rect 35644 1204 44268 1260
rect 44426 1204 44436 1260
rect 44492 1204 50596 1260
rect 50652 1204 50662 1260
rect 53844 1148 53900 1316
rect 72324 1260 72380 1428
rect 75180 1372 75236 1428
rect 79268 1372 79324 1428
rect 87724 1372 87780 1428
rect 100324 1372 100380 1428
rect 108500 1372 108556 1428
rect 122052 1372 122108 1428
rect 138964 1372 139020 1428
rect 148260 1372 148316 1428
rect 219200 1372 220000 1400
rect 72538 1316 72548 1372
rect 72604 1316 75236 1372
rect 75338 1316 75348 1372
rect 75404 1316 76692 1372
rect 76748 1316 76758 1372
rect 77018 1316 77028 1372
rect 77084 1316 78708 1372
rect 78764 1316 78774 1372
rect 78922 1316 78932 1372
rect 78988 1316 79044 1372
rect 79100 1316 79110 1372
rect 79268 1316 79940 1372
rect 79996 1316 80006 1372
rect 80154 1316 80164 1372
rect 80220 1316 82628 1372
rect 82684 1316 82694 1372
rect 82842 1316 82852 1372
rect 82908 1316 85652 1372
rect 85708 1316 85718 1372
rect 85876 1316 87556 1372
rect 87612 1316 87622 1372
rect 87724 1316 88844 1372
rect 89002 1316 89012 1372
rect 89068 1316 89796 1372
rect 89852 1316 89862 1372
rect 90570 1316 90580 1372
rect 90636 1316 99204 1372
rect 99260 1316 99270 1372
rect 99418 1316 99428 1372
rect 99484 1316 99522 1372
rect 100324 1316 100996 1372
rect 101052 1316 101062 1372
rect 101210 1316 101220 1372
rect 101276 1316 108276 1372
rect 108332 1316 108342 1372
rect 108500 1316 109060 1372
rect 109116 1316 109126 1372
rect 109274 1316 109284 1372
rect 109340 1316 111412 1372
rect 111468 1316 111478 1372
rect 111626 1316 111636 1372
rect 111692 1316 120260 1372
rect 120316 1316 120326 1372
rect 120670 1316 120708 1372
rect 120764 1316 120774 1372
rect 122052 1316 123284 1372
rect 123340 1316 123350 1372
rect 123498 1316 123508 1372
rect 123564 1316 126084 1372
rect 126140 1316 126150 1372
rect 126298 1316 126308 1372
rect 126364 1316 132972 1372
rect 135006 1316 135044 1372
rect 135100 1316 135110 1372
rect 137162 1316 137172 1372
rect 137228 1316 139020 1372
rect 139402 1316 139412 1372
rect 139468 1316 148316 1372
rect 150154 1316 150164 1372
rect 150220 1316 156100 1372
rect 156156 1316 156166 1372
rect 163482 1316 163492 1372
rect 163548 1316 166180 1372
rect 166236 1316 166246 1372
rect 172666 1316 172676 1372
rect 172732 1316 201684 1372
rect 201740 1316 201750 1372
rect 203251 1316 205828 1372
rect 205884 1316 205894 1372
rect 211054 1316 211092 1372
rect 211148 1316 211158 1372
rect 214442 1316 214452 1372
rect 214508 1316 220000 1372
rect 85876 1260 85932 1316
rect 88788 1260 88844 1316
rect 132916 1260 132972 1316
rect 203251 1260 203307 1316
rect 219200 1288 220000 1316
rect 59182 1204 59220 1260
rect 59276 1204 59286 1260
rect 60442 1204 60452 1260
rect 60508 1204 61908 1260
rect 61964 1204 61974 1260
rect 62122 1204 62132 1260
rect 62188 1204 62198 1260
rect 62570 1204 62580 1260
rect 62636 1204 68068 1260
rect 68124 1204 68134 1260
rect 68506 1204 68516 1260
rect 68572 1204 72380 1260
rect 72538 1204 72548 1260
rect 72604 1204 74508 1260
rect 74890 1204 74900 1260
rect 74956 1204 85932 1260
rect 86986 1204 86996 1260
rect 87052 1204 88564 1260
rect 88620 1204 88630 1260
rect 88788 1204 89908 1260
rect 89964 1204 89974 1260
rect 90346 1204 90356 1260
rect 90412 1204 99988 1260
rect 100044 1204 100054 1260
rect 100202 1204 100212 1260
rect 100268 1204 105812 1260
rect 105868 1204 105878 1260
rect 106026 1204 106036 1260
rect 106092 1204 108836 1260
rect 108892 1204 108902 1260
rect 109386 1204 109396 1260
rect 109452 1204 113988 1260
rect 114044 1204 114054 1260
rect 114202 1204 114212 1260
rect 114268 1204 116788 1260
rect 116844 1204 116854 1260
rect 117002 1204 117012 1260
rect 117068 1204 117106 1260
rect 117562 1204 117572 1260
rect 117628 1204 125748 1260
rect 125804 1204 125814 1260
rect 125962 1204 125972 1260
rect 126028 1204 127540 1260
rect 127596 1204 127606 1260
rect 132682 1204 132692 1260
rect 132748 1204 132860 1260
rect 132916 1204 135828 1260
rect 135884 1204 135894 1260
rect 138058 1204 138068 1260
rect 138124 1204 144004 1260
rect 144060 1204 144070 1260
rect 144228 1204 150164 1260
rect 150220 1204 150230 1260
rect 150378 1204 150388 1260
rect 150444 1204 152740 1260
rect 152796 1204 152806 1260
rect 164154 1204 164164 1260
rect 164220 1204 181412 1260
rect 181468 1204 181478 1260
rect 197316 1204 203307 1260
rect 208282 1204 208292 1260
rect 208348 1204 209860 1260
rect 209916 1204 209926 1260
rect 62131 1148 62187 1204
rect 74452 1148 74508 1204
rect 132804 1148 132860 1204
rect 144228 1148 144284 1204
rect 10126 1092 10164 1148
rect 10220 1092 10230 1148
rect 12282 1092 12292 1148
rect 12348 1092 26852 1148
rect 26908 1092 26918 1148
rect 30650 1092 30660 1148
rect 30716 1092 44660 1148
rect 44716 1092 44726 1148
rect 50110 1092 50148 1148
rect 50204 1092 50214 1148
rect 50362 1092 50372 1148
rect 50428 1092 53900 1148
rect 54058 1092 54068 1148
rect 54124 1092 62187 1148
rect 63924 1092 70532 1148
rect 70588 1092 70598 1148
rect 70746 1092 70756 1148
rect 70812 1092 74116 1148
rect 74172 1092 74182 1148
rect 74452 1092 87220 1148
rect 87276 1092 87286 1148
rect 87434 1092 87444 1148
rect 87500 1092 90580 1148
rect 90636 1092 90646 1148
rect 91018 1092 91028 1148
rect 91084 1092 92372 1148
rect 92428 1092 92438 1148
rect 94042 1092 94052 1148
rect 94108 1092 103236 1148
rect 103292 1092 103302 1148
rect 103460 1092 109620 1148
rect 109676 1092 109686 1148
rect 109834 1092 109844 1148
rect 109900 1092 110740 1148
rect 110796 1092 110806 1148
rect 110954 1092 110964 1148
rect 111020 1092 125860 1148
rect 125916 1092 125926 1148
rect 126186 1092 126196 1148
rect 126252 1092 126980 1148
rect 127036 1092 127046 1148
rect 127418 1092 127428 1148
rect 127484 1092 130564 1148
rect 130620 1092 130630 1148
rect 132804 1092 140308 1148
rect 140364 1092 140374 1148
rect 142874 1092 142884 1148
rect 142940 1092 144284 1148
rect 144452 1092 168644 1148
rect 168700 1092 168710 1148
rect 170874 1092 170884 1148
rect 170940 1092 190596 1148
rect 190652 1092 190662 1148
rect 192798 1092 192836 1148
rect 192892 1092 192902 1148
rect 63924 1036 63980 1092
rect 103460 1036 103516 1092
rect 144452 1036 144508 1092
rect 18414 980 18452 1036
rect 18508 980 18518 1036
rect 19226 980 19236 1036
rect 19292 980 39172 1036
rect 39228 980 39238 1036
rect 39386 980 39396 1036
rect 39452 980 63980 1036
rect 64138 980 64148 1036
rect 64204 980 65380 1036
rect 65436 980 65446 1036
rect 68954 980 68964 1036
rect 69020 980 76020 1036
rect 76076 980 76086 1036
rect 76682 980 76692 1036
rect 76748 980 80724 1036
rect 80780 980 80790 1036
rect 80938 980 80948 1036
rect 81004 980 84420 1036
rect 84476 980 84486 1036
rect 84746 980 84756 1036
rect 84812 980 85540 1036
rect 85596 980 85606 1036
rect 85754 980 85764 1036
rect 85820 980 87108 1036
rect 87164 980 87174 1036
rect 87322 980 87332 1036
rect 87388 980 96292 1036
rect 96348 980 96358 1036
rect 97402 980 97412 1036
rect 97468 980 97524 1036
rect 97580 980 97590 1036
rect 97738 980 97748 1036
rect 97804 980 100436 1036
rect 100492 980 100502 1036
rect 100762 980 100772 1036
rect 100828 980 103516 1036
rect 103674 980 103684 1036
rect 103740 980 105924 1036
rect 105980 980 105990 1036
rect 106138 980 106148 1036
rect 106204 980 106242 1036
rect 106362 980 106372 1036
rect 106428 980 106466 1036
rect 106596 980 107996 1036
rect 108154 980 108164 1036
rect 108220 980 110068 1036
rect 110124 980 110134 1036
rect 110282 980 110292 1036
rect 110348 980 116116 1036
rect 116172 980 116182 1036
rect 116442 980 116452 1036
rect 116508 980 119252 1036
rect 119308 980 119318 1036
rect 119466 980 119476 1036
rect 119532 980 119700 1036
rect 119756 980 119766 1036
rect 119914 980 119924 1036
rect 119980 980 137172 1036
rect 137228 980 137238 1036
rect 138292 980 144508 1036
rect 144666 980 144676 1036
rect 144732 980 144956 1036
rect 147662 980 147700 1036
rect 147756 980 147766 1036
rect 147914 980 147924 1036
rect 147980 980 152852 1036
rect 152908 980 152918 1036
rect 153710 980 153748 1036
rect 153804 980 153814 1036
rect 153962 980 153972 1036
rect 154028 980 173067 1036
rect 174458 980 174468 1036
rect 174524 980 194068 1036
rect 194124 980 194134 1036
rect 195150 980 195188 1036
rect 195244 980 195254 1036
rect 197054 980 197092 1036
rect 197148 980 197158 1036
rect 106596 924 106652 980
rect 746 868 756 924
rect 812 868 822 924
rect 1278 868 1316 924
rect 1372 868 1382 924
rect 1950 868 1988 924
rect 2044 868 2054 924
rect 2510 868 2548 924
rect 2604 868 2614 924
rect 3210 868 3220 924
rect 3276 868 3286 924
rect 15950 868 15988 924
rect 16044 868 16054 924
rect 18890 868 18900 924
rect 18956 868 18966 924
rect 19646 868 19684 924
rect 19740 868 19750 924
rect 31891 868 39732 924
rect 39788 868 39798 924
rect 40366 868 40404 924
rect 40460 868 40470 924
rect 40926 868 40964 924
rect 41020 868 41030 924
rect 68292 868 75236 924
rect 75292 868 75302 924
rect 75450 868 75460 924
rect 75516 868 76020 924
rect 76076 868 76086 924
rect 76206 868 76244 924
rect 76300 868 76310 924
rect 76570 868 76580 924
rect 76636 868 80164 924
rect 80220 868 80230 924
rect 80378 868 80388 924
rect 80444 868 81172 924
rect 81228 868 81238 924
rect 81386 868 81396 924
rect 81452 868 81508 924
rect 81564 868 81574 924
rect 81722 868 81732 924
rect 81788 868 81844 924
rect 81900 868 81910 924
rect 82170 868 82180 924
rect 82236 868 82852 924
rect 82908 868 82918 924
rect 83066 868 83076 924
rect 83132 868 106652 924
rect 107940 924 107996 980
rect 107940 868 123844 924
rect 123900 868 123910 924
rect 125850 868 125860 924
rect 125916 868 133924 924
rect 133980 868 133990 924
rect 756 700 812 868
rect 3220 812 3276 868
rect 18900 812 18956 868
rect 31891 812 31947 868
rect 3220 756 18956 812
rect 19338 756 19348 812
rect 19404 756 31947 812
rect 39386 756 39396 812
rect 39452 756 44436 812
rect 44492 756 44502 812
rect 44650 756 44660 812
rect 44716 756 50372 812
rect 50428 756 50438 812
rect 50586 756 50596 812
rect 50652 756 66164 812
rect 66220 756 66230 812
rect 68292 700 68348 868
rect 138292 812 138348 980
rect 144900 924 144956 980
rect 138506 868 138516 924
rect 138572 868 144452 924
rect 144508 868 144518 924
rect 144900 868 151172 924
rect 151228 868 151238 924
rect 151918 868 151956 924
rect 152012 868 152022 924
rect 161251 868 162820 924
rect 162876 868 162886 924
rect 171406 868 171444 924
rect 171500 868 171510 924
rect 161251 812 161307 868
rect 756 644 22932 700
rect 22988 644 22998 700
rect 29642 644 29652 700
rect 29708 644 50484 700
rect 50540 644 50550 700
rect 52042 644 52052 700
rect 52108 644 56812 700
rect 57082 644 57092 700
rect 57148 644 68348 700
rect 68404 756 72548 812
rect 72604 756 72614 812
rect 74106 756 74116 812
rect 74172 756 75348 812
rect 75404 756 75414 812
rect 76020 756 76692 812
rect 76748 756 76758 812
rect 77242 756 77252 812
rect 77308 756 81060 812
rect 81116 756 81126 812
rect 81498 756 81508 812
rect 81564 756 81956 812
rect 82012 756 82022 812
rect 82282 756 82292 812
rect 82348 756 107492 812
rect 107548 756 107558 812
rect 107716 756 108052 812
rect 108108 756 108118 812
rect 108266 756 108276 812
rect 108332 756 112084 812
rect 112140 756 112150 812
rect 112298 756 112308 812
rect 112364 756 138348 812
rect 142538 756 142548 812
rect 142604 756 161307 812
rect 173011 812 173067 980
rect 197316 924 197372 1204
rect 197530 1092 197540 1148
rect 197596 1092 214116 1148
rect 214172 1092 214182 1148
rect 216346 1092 216356 1148
rect 216412 1092 219604 1148
rect 219660 1092 219670 1148
rect 197642 980 197652 1036
rect 197708 980 201348 1036
rect 201404 980 201414 1036
rect 201562 980 201572 1036
rect 201628 980 212324 1036
rect 212380 980 212390 1036
rect 173898 868 173908 924
rect 173964 868 197372 924
rect 202990 868 203028 924
rect 203084 868 203094 924
rect 203251 868 203812 924
rect 203868 868 203878 924
rect 205566 868 205604 924
rect 205660 868 205670 924
rect 206798 868 206836 924
rect 206892 868 206902 924
rect 212846 868 212884 924
rect 212940 868 212950 924
rect 217102 868 217140 924
rect 217196 868 217206 924
rect 203251 812 203307 868
rect 173011 756 203307 812
rect 204138 756 204148 812
rect 204204 756 204214 812
rect 6570 532 6580 588
rect 6636 532 31444 588
rect 31500 532 31510 588
rect 46666 532 46676 588
rect 46732 532 50427 588
rect 52126 532 52164 588
rect 52220 532 52230 588
rect 50371 476 50427 532
rect 56756 476 56812 644
rect 68404 588 68460 756
rect 76020 700 76076 756
rect 107716 700 107772 756
rect 204148 700 204204 756
rect 74778 644 74788 700
rect 74844 644 76076 700
rect 76234 644 76244 700
rect 76300 644 76804 700
rect 76860 644 76870 700
rect 77130 644 77140 700
rect 77196 644 78596 700
rect 78652 644 78662 700
rect 79258 644 79268 700
rect 79324 644 80388 700
rect 80444 644 80454 700
rect 80714 644 80724 700
rect 80780 644 107772 700
rect 107930 644 107940 700
rect 107996 644 117012 700
rect 117068 644 117078 700
rect 117562 644 117572 700
rect 117628 644 118916 700
rect 118972 644 118982 700
rect 119130 644 119140 700
rect 119196 644 121716 700
rect 121772 644 121782 700
rect 123498 644 123508 700
rect 123564 644 134596 700
rect 134652 644 134662 700
rect 141306 644 141316 700
rect 141372 644 144452 700
rect 144508 644 144518 700
rect 144666 644 144676 700
rect 144732 644 144742 700
rect 145002 644 145012 700
rect 145068 644 191828 700
rect 191884 644 191894 700
rect 194058 644 194068 700
rect 194124 644 204204 700
rect 144676 588 144732 644
rect 56970 532 56980 588
rect 57036 532 68460 588
rect 68730 532 68740 588
rect 68796 532 76972 588
rect 77130 532 77140 588
rect 77196 532 124180 588
rect 124236 532 124246 588
rect 125290 532 125300 588
rect 125356 532 132020 588
rect 132076 532 132086 588
rect 134474 532 134484 588
rect 134540 532 144732 588
rect 144890 532 144900 588
rect 144956 532 150388 588
rect 150444 532 150454 588
rect 151050 532 151060 588
rect 151116 532 214340 588
rect 214396 532 214406 588
rect 13962 420 13972 476
rect 14028 420 41188 476
rect 41244 420 41254 476
rect 49886 420 49924 476
rect 49980 420 49990 476
rect 50371 420 56532 476
rect 56588 420 56598 476
rect 56756 420 57428 476
rect 57484 420 57494 476
rect 59770 420 59780 476
rect 59836 420 72324 476
rect 72380 420 72390 476
rect 72538 420 72548 476
rect 72604 420 76580 476
rect 76636 420 76646 476
rect 76916 364 76972 532
rect 77242 420 77252 476
rect 77308 420 79044 476
rect 79100 420 79110 476
rect 79268 420 80052 476
rect 80108 420 80118 476
rect 80266 420 80276 476
rect 80332 420 81340 476
rect 81610 420 81620 476
rect 81676 420 91700 476
rect 91756 420 91766 476
rect 97290 420 97300 476
rect 97356 420 97412 476
rect 97468 420 97478 476
rect 98130 420 98140 476
rect 98196 420 100548 476
rect 100604 420 100614 476
rect 100762 420 100772 476
rect 100828 420 102004 476
rect 102060 420 102070 476
rect 102218 420 102228 476
rect 102284 420 109844 476
rect 109900 420 109910 476
rect 110058 420 110068 476
rect 110124 420 116228 476
rect 116284 420 116294 476
rect 116452 420 117572 476
rect 117628 420 117638 476
rect 117786 420 117796 476
rect 117852 420 120820 476
rect 120876 420 120886 476
rect 121930 420 121940 476
rect 121996 420 124740 476
rect 124796 420 124806 476
rect 124964 420 130788 476
rect 130844 420 130854 476
rect 131114 420 131124 476
rect 131180 420 138516 476
rect 138572 420 138582 476
rect 141978 420 141988 476
rect 142044 420 217364 476
rect 217420 420 217430 476
rect 79268 364 79324 420
rect 81284 364 81340 420
rect 116452 364 116508 420
rect 124964 364 125020 420
rect 7802 308 7812 364
rect 7868 308 35812 364
rect 35868 308 35878 364
rect 44202 308 44212 364
rect 44268 308 57764 364
rect 57820 308 57830 364
rect 59658 308 59668 364
rect 59724 308 76692 364
rect 76748 308 76758 364
rect 76916 308 79324 364
rect 79594 308 79604 364
rect 79660 308 81060 364
rect 81116 308 81126 364
rect 81284 308 83300 364
rect 83356 308 83366 364
rect 83514 308 83524 364
rect 83580 308 85764 364
rect 85820 308 85830 364
rect 85978 308 85988 364
rect 86044 308 86660 364
rect 86716 308 86726 364
rect 86874 308 86884 364
rect 86940 308 97300 364
rect 97356 308 97366 364
rect 99194 308 99204 364
rect 99260 308 103012 364
rect 103068 308 103078 364
rect 103226 308 103236 364
rect 103292 308 110852 364
rect 110908 308 110918 364
rect 111066 308 111076 364
rect 111132 308 116508 364
rect 116666 308 116676 364
rect 116732 308 121044 364
rect 121100 308 121110 364
rect 121258 308 121268 364
rect 121324 308 125020 364
rect 127530 308 127540 364
rect 127596 308 204708 364
rect 204764 308 204774 364
rect 522 196 532 252
rect 588 196 19908 252
rect 19964 196 19974 252
rect 20682 196 20692 252
rect 20748 196 52052 252
rect 52108 196 52118 252
rect 52266 196 52276 252
rect 52332 196 60564 252
rect 60620 196 60630 252
rect 71866 196 71876 252
rect 71932 196 205828 252
rect 205884 196 205894 252
rect 19226 84 19236 140
rect 19292 84 63588 140
rect 63644 84 63654 140
rect 65930 84 65940 140
rect 65996 84 207620 140
rect 207676 84 207686 140
<< via3 >>
rect 102452 14868 102508 14924
rect 103012 14868 103068 14924
rect 115444 14868 115500 14924
rect 120932 14868 120988 14924
rect 151620 14868 151676 14924
rect 70196 14756 70252 14812
rect 71652 14756 71708 14812
rect 77588 14756 77644 14812
rect 80836 14756 80892 14812
rect 82180 14756 82236 14812
rect 98308 14756 98364 14812
rect 111412 14756 111468 14812
rect 81284 14644 81340 14700
rect 100660 14644 100716 14700
rect 103908 14644 103964 14700
rect 121044 14644 121100 14700
rect 121268 14644 121324 14700
rect 124628 14644 124684 14700
rect 151060 14644 151116 14700
rect 153076 14644 153132 14700
rect 153524 14644 153580 14700
rect 156100 14644 156156 14700
rect 65604 14532 65660 14588
rect 77924 14532 77980 14588
rect 78148 14532 78204 14588
rect 79604 14532 79660 14588
rect 80388 14532 80444 14588
rect 80612 14532 80668 14588
rect 92596 14532 92652 14588
rect 92820 14532 92876 14588
rect 98308 14532 98364 14588
rect 98532 14532 98588 14588
rect 102788 14532 102844 14588
rect 113988 14532 114044 14588
rect 120372 14532 120428 14588
rect 149380 14532 149436 14588
rect 82068 14420 82124 14476
rect 82292 14420 82348 14476
rect 82628 14420 82684 14476
rect 114996 14420 115052 14476
rect 118804 14420 118860 14476
rect 119364 14420 119420 14476
rect 119924 14420 119980 14476
rect 120484 14420 120540 14476
rect 124404 14420 124460 14476
rect 124628 14420 124684 14476
rect 156212 14420 156268 14476
rect 156436 14420 156492 14476
rect 70084 14308 70140 14364
rect 77476 14308 77532 14364
rect 114212 14308 114268 14364
rect 120708 14308 120764 14364
rect 121044 14308 121100 14364
rect 139412 14308 139468 14364
rect 156772 14308 156828 14364
rect 182756 14308 182812 14364
rect 77588 14196 77644 14252
rect 78148 14196 78204 14252
rect 79492 14196 79548 14252
rect 79716 14196 79772 14252
rect 103348 14196 103404 14252
rect 116340 14196 116396 14252
rect 116564 14196 116620 14252
rect 117236 14196 117292 14252
rect 117796 14196 117852 14252
rect 118356 14196 118412 14252
rect 142660 14196 142716 14252
rect 149268 14196 149324 14252
rect 151284 14196 151340 14252
rect 152740 14196 152796 14252
rect 153076 14196 153132 14252
rect 158676 14196 158732 14252
rect 21476 14084 21532 14140
rect 69636 14084 69692 14140
rect 79044 14084 79100 14140
rect 79604 14084 79660 14140
rect 80612 14084 80668 14140
rect 80836 14084 80892 14140
rect 124516 14084 124572 14140
rect 124740 14084 124796 14140
rect 154084 14084 154140 14140
rect 14868 13972 14924 14028
rect 17780 13972 17836 14028
rect 77700 13972 77756 14028
rect 78708 13972 78764 14028
rect 81284 13972 81340 14028
rect 92372 13972 92428 14028
rect 92596 13972 92652 14028
rect 97300 13972 97356 14028
rect 115444 13972 115500 14028
rect 116004 13972 116060 14028
rect 134036 13972 134092 14028
rect 134260 13972 134316 14028
rect 151172 13972 151228 14028
rect 156436 13972 156492 14028
rect 159460 13972 159516 14028
rect 162708 13972 162764 14028
rect 166852 13972 166908 14028
rect 191156 13972 191212 14028
rect 25060 13860 25116 13916
rect 61460 13860 61516 13916
rect 73108 13860 73164 13916
rect 74676 13860 74732 13916
rect 77140 13860 77196 13916
rect 77364 13860 77420 13916
rect 81732 13860 81788 13916
rect 82292 13860 82348 13916
rect 92484 13860 92540 13916
rect 99876 13860 99932 13916
rect 114772 13860 114828 13916
rect 117908 13860 117964 13916
rect 118132 13860 118188 13916
rect 118804 13860 118860 13916
rect 119700 13860 119756 13916
rect 126980 13860 127036 13916
rect 138068 13860 138124 13916
rect 139524 13860 139580 13916
rect 158340 13860 158396 13916
rect 172452 13860 172508 13916
rect 174468 13860 174524 13916
rect 193396 13860 193452 13916
rect 57092 13748 57148 13804
rect 74228 13748 74284 13804
rect 82852 13748 82908 13804
rect 83076 13748 83132 13804
rect 120596 13748 120652 13804
rect 120820 13748 120876 13804
rect 124292 13748 124348 13804
rect 155876 13748 155932 13804
rect 183204 13748 183260 13804
rect 65604 13636 65660 13692
rect 65940 13636 65996 13692
rect 67732 13636 67788 13692
rect 81844 13636 81900 13692
rect 82068 13636 82124 13692
rect 92484 13636 92540 13692
rect 102788 13636 102844 13692
rect 116452 13636 116508 13692
rect 146020 13636 146076 13692
rect 147924 13636 147980 13692
rect 148148 13636 148204 13692
rect 174020 13636 174076 13692
rect 10500 13524 10556 13580
rect 64036 13524 64092 13580
rect 68068 13524 68124 13580
rect 68292 13524 68348 13580
rect 83188 13524 83244 13580
rect 83412 13524 83468 13580
rect 83972 13524 84028 13580
rect 85204 13524 85260 13580
rect 91252 13524 91308 13580
rect 97076 13524 97132 13580
rect 97300 13524 97356 13580
rect 103796 13524 103852 13580
rect 119476 13524 119532 13580
rect 120372 13524 120428 13580
rect 120596 13524 120652 13580
rect 162260 13524 162316 13580
rect 173572 13524 173628 13580
rect 25732 13412 25788 13468
rect 53844 13412 53900 13468
rect 63924 13412 63980 13468
rect 77588 13412 77644 13468
rect 77812 13412 77868 13468
rect 117796 13412 117852 13468
rect 124740 13412 124796 13468
rect 136500 13412 136556 13468
rect 137956 13412 138012 13468
rect 148148 13412 148204 13468
rect 148372 13412 148428 13468
rect 152292 13412 152348 13468
rect 167972 13412 168028 13468
rect 187572 13412 187628 13468
rect 82740 13300 82796 13356
rect 83300 13300 83356 13356
rect 103236 13300 103292 13356
rect 149828 13300 149884 13356
rect 165396 13300 165452 13356
rect 172452 13300 172508 13356
rect 211652 13300 211708 13356
rect 18452 13188 18508 13244
rect 53060 13188 53116 13244
rect 68068 13188 68124 13244
rect 73780 13188 73836 13244
rect 77476 13188 77532 13244
rect 133476 13188 133532 13244
rect 134260 13188 134316 13244
rect 135604 13188 135660 13244
rect 146916 13188 146972 13244
rect 161028 13188 161084 13244
rect 162596 13188 162652 13244
rect 164948 13188 165004 13244
rect 73220 13076 73276 13132
rect 73444 13076 73500 13132
rect 77588 13076 77644 13132
rect 80724 13076 80780 13132
rect 81060 13076 81116 13132
rect 83524 13076 83580 13132
rect 83748 13076 83804 13132
rect 84644 13076 84700 13132
rect 84868 13076 84924 13132
rect 85204 13076 85260 13132
rect 86996 13076 87052 13132
rect 103012 13076 103068 13132
rect 119924 13076 119980 13132
rect 132692 13076 132748 13132
rect 149156 13076 149212 13132
rect 149492 13076 149548 13132
rect 154308 13076 154364 13132
rect 27972 12964 28028 13020
rect 34468 12964 34524 13020
rect 64036 12964 64092 13020
rect 77140 12964 77196 13020
rect 77924 12964 77980 13020
rect 78932 12964 78988 13020
rect 91252 12964 91308 13020
rect 103236 12964 103292 13020
rect 103572 12964 103628 13020
rect 104132 12964 104188 13020
rect 109620 12964 109676 13020
rect 122724 12964 122780 13020
rect 146916 12964 146972 13020
rect 148932 12964 148988 13020
rect 165396 12964 165452 13020
rect 165732 12964 165788 13020
rect 185332 12964 185388 13020
rect 195524 12964 195580 13020
rect 56196 12852 56252 12908
rect 73780 12852 73836 12908
rect 75236 12852 75292 12908
rect 103684 12852 103740 12908
rect 103908 12852 103964 12908
rect 104692 12852 104748 12908
rect 114324 12852 114380 12908
rect 114548 12852 114604 12908
rect 119140 12852 119196 12908
rect 119364 12852 119420 12908
rect 137620 12852 137676 12908
rect 142436 12852 142492 12908
rect 142772 12852 142828 12908
rect 152852 12852 152908 12908
rect 162148 12852 162204 12908
rect 173796 12852 173852 12908
rect 196532 12852 196588 12908
rect 27188 12740 27244 12796
rect 77812 12740 77868 12796
rect 78820 12740 78876 12796
rect 80500 12740 80556 12796
rect 80836 12740 80892 12796
rect 91700 12740 91756 12796
rect 102564 12740 102620 12796
rect 102788 12740 102844 12796
rect 120932 12740 120988 12796
rect 149156 12740 149212 12796
rect 149492 12740 149548 12796
rect 150948 12740 151004 12796
rect 173684 12740 173740 12796
rect 69524 12628 69580 12684
rect 73108 12628 73164 12684
rect 77924 12628 77980 12684
rect 94948 12628 95004 12684
rect 96068 12628 96124 12684
rect 102004 12628 102060 12684
rect 102340 12628 102396 12684
rect 114772 12628 114828 12684
rect 114996 12628 115052 12684
rect 137620 12628 137676 12684
rect 137844 12628 137900 12684
rect 149268 12628 149324 12684
rect 149940 12628 149996 12684
rect 151284 12628 151340 12684
rect 174020 12628 174076 12684
rect 174244 12628 174300 12684
rect 180852 12628 180908 12684
rect 193844 12628 193900 12684
rect 200900 12628 200956 12684
rect 30100 12516 30156 12572
rect 68852 12516 68908 12572
rect 69076 12516 69132 12572
rect 78148 12516 78204 12572
rect 78372 12516 78428 12572
rect 78932 12516 78988 12572
rect 80052 12516 80108 12572
rect 80388 12516 80444 12572
rect 81284 12516 81340 12572
rect 81732 12516 81788 12572
rect 84308 12516 84364 12572
rect 84756 12516 84812 12572
rect 86548 12516 86604 12572
rect 91700 12516 91756 12572
rect 111748 12516 111804 12572
rect 114436 12516 114492 12572
rect 120708 12516 120764 12572
rect 148708 12516 148764 12572
rect 195412 12516 195468 12572
rect 63252 12404 63308 12460
rect 69748 12404 69804 12460
rect 69972 12404 70028 12460
rect 73556 12404 73612 12460
rect 74004 12404 74060 12460
rect 77364 12404 77420 12460
rect 80276 12404 80332 12460
rect 81508 12404 81564 12460
rect 83300 12404 83356 12460
rect 97636 12404 97692 12460
rect 99876 12404 99932 12460
rect 102116 12404 102172 12460
rect 114548 12404 114604 12460
rect 114772 12404 114828 12460
rect 119028 12404 119084 12460
rect 119364 12404 119420 12460
rect 122724 12404 122780 12460
rect 125524 12404 125580 12460
rect 126532 12404 126588 12460
rect 154084 12404 154140 12460
rect 154308 12404 154364 12460
rect 155764 12404 155820 12460
rect 156212 12404 156268 12460
rect 55412 12292 55468 12348
rect 55636 12292 55692 12348
rect 158676 12404 158732 12460
rect 164276 12404 164332 12460
rect 166516 12404 166572 12460
rect 174244 12404 174300 12460
rect 174468 12404 174524 12460
rect 193844 12404 193900 12460
rect 70084 12292 70140 12348
rect 70308 12292 70364 12348
rect 78484 12292 78540 12348
rect 79828 12292 79884 12348
rect 83412 12292 83468 12348
rect 83748 12292 83804 12348
rect 83972 12292 84028 12348
rect 84644 12292 84700 12348
rect 84868 12292 84924 12348
rect 89460 12292 89516 12348
rect 103908 12292 103964 12348
rect 104468 12292 104524 12348
rect 113652 12292 113708 12348
rect 114212 12292 114268 12348
rect 116788 12292 116844 12348
rect 117908 12292 117964 12348
rect 121044 12292 121100 12348
rect 130788 12292 130844 12348
rect 138292 12292 138348 12348
rect 160580 12292 160636 12348
rect 162708 12292 162764 12348
rect 171220 12292 171276 12348
rect 172228 12292 172284 12348
rect 180852 12292 180908 12348
rect 187012 12292 187068 12348
rect 56196 12180 56252 12236
rect 67508 12180 67564 12236
rect 71988 12180 72044 12236
rect 73556 12180 73612 12236
rect 79940 12180 79996 12236
rect 80388 12180 80444 12236
rect 89012 12180 89068 12236
rect 90356 12180 90412 12236
rect 97636 12180 97692 12236
rect 98084 12180 98140 12236
rect 99092 12180 99148 12236
rect 102564 12180 102620 12236
rect 103012 12180 103068 12236
rect 109396 12180 109452 12236
rect 120260 12180 120316 12236
rect 120596 12180 120652 12236
rect 125524 12180 125580 12236
rect 125748 12180 125804 12236
rect 131460 12180 131516 12236
rect 132468 12180 132524 12236
rect 141204 12180 141260 12236
rect 156212 12180 156268 12236
rect 178836 12180 178892 12236
rect 212996 12180 213052 12236
rect 55412 12068 55468 12124
rect 63476 12068 63532 12124
rect 63700 12068 63756 12124
rect 68852 12068 68908 12124
rect 74116 12068 74172 12124
rect 80836 12068 80892 12124
rect 81172 12068 81228 12124
rect 98980 12068 99036 12124
rect 106148 12068 106204 12124
rect 114100 12068 114156 12124
rect 114324 12068 114380 12124
rect 115668 12068 115724 12124
rect 115892 12068 115948 12124
rect 117348 12068 117404 12124
rect 118244 12068 118300 12124
rect 162036 12068 162092 12124
rect 164276 12068 164332 12124
rect 164500 12068 164556 12124
rect 194852 12068 194908 12124
rect 197764 12068 197820 12124
rect 75012 11956 75068 12012
rect 80276 11956 80332 12012
rect 80500 11956 80556 12012
rect 82292 11956 82348 12012
rect 82516 11956 82572 12012
rect 89236 11956 89292 12012
rect 97748 11956 97804 12012
rect 108724 11956 108780 12012
rect 108948 11956 109004 12012
rect 109284 11956 109340 12012
rect 115220 11956 115276 12012
rect 138180 11956 138236 12012
rect 147476 11956 147532 12012
rect 149044 11956 149100 12012
rect 149380 11956 149436 12012
rect 162148 11956 162204 12012
rect 162484 11956 162540 12012
rect 163716 11956 163772 12012
rect 166292 11956 166348 12012
rect 166516 11956 166572 12012
rect 75124 11844 75180 11900
rect 78708 11844 78764 11900
rect 79044 11844 79100 11900
rect 82068 11844 82124 11900
rect 84532 11844 84588 11900
rect 95284 11844 95340 11900
rect 98868 11844 98924 11900
rect 104244 11844 104300 11900
rect 107492 11844 107548 11900
rect 116340 11844 116396 11900
rect 119252 11844 119308 11900
rect 121380 11844 121436 11900
rect 126308 11844 126364 11900
rect 131460 11844 131516 11900
rect 135492 11844 135548 11900
rect 141316 11844 141372 11900
rect 141540 11844 141596 11900
rect 146132 11844 146188 11900
rect 148036 11844 148092 11900
rect 149156 11844 149212 11900
rect 151172 11844 151228 11900
rect 153524 11844 153580 11900
rect 168868 11844 168924 11900
rect 172564 11844 172620 11900
rect 57092 11732 57148 11788
rect 57764 11732 57820 11788
rect 62132 11732 62188 11788
rect 65380 11732 65436 11788
rect 67172 11732 67228 11788
rect 67508 11732 67564 11788
rect 74116 11732 74172 11788
rect 77700 11732 77756 11788
rect 77924 11732 77980 11788
rect 96068 11732 96124 11788
rect 97076 11732 97132 11788
rect 100436 11732 100492 11788
rect 106148 11732 106204 11788
rect 113316 11732 113372 11788
rect 117124 11732 117180 11788
rect 119364 11732 119420 11788
rect 120932 11732 120988 11788
rect 122276 11732 122332 11788
rect 122500 11732 122556 11788
rect 132692 11732 132748 11788
rect 137732 11732 137788 11788
rect 173796 11844 173852 11900
rect 187012 11844 187068 11900
rect 198436 11844 198492 11900
rect 206948 11844 207004 11900
rect 154868 11732 154924 11788
rect 155092 11732 155148 11788
rect 174468 11732 174524 11788
rect 55748 11620 55804 11676
rect 66612 11620 66668 11676
rect 66836 11620 66892 11676
rect 67396 11620 67452 11676
rect 68180 11620 68236 11676
rect 69524 11620 69580 11676
rect 69748 11620 69804 11676
rect 77252 11620 77308 11676
rect 102340 11620 102396 11676
rect 103012 11620 103068 11676
rect 112756 11620 112812 11676
rect 116004 11620 116060 11676
rect 116228 11620 116284 11676
rect 116788 11620 116844 11676
rect 119924 11620 119980 11676
rect 120148 11620 120204 11676
rect 134260 11620 134316 11676
rect 156212 11620 156268 11676
rect 158564 11620 158620 11676
rect 158788 11620 158844 11676
rect 162260 11620 162316 11676
rect 182980 11620 183036 11676
rect 51716 11508 51772 11564
rect 56196 11508 56252 11564
rect 57092 11508 57148 11564
rect 103460 11508 103516 11564
rect 107940 11508 107996 11564
rect 109060 11508 109116 11564
rect 110964 11508 111020 11564
rect 112532 11508 112588 11564
rect 113988 11508 114044 11564
rect 114324 11508 114380 11564
rect 115780 11508 115836 11564
rect 116340 11508 116396 11564
rect 116564 11508 116620 11564
rect 117684 11508 117740 11564
rect 126532 11508 126588 11564
rect 140756 11508 140812 11564
rect 152740 11508 152796 11564
rect 168532 11508 168588 11564
rect 170996 11508 171052 11564
rect 191716 11508 191772 11564
rect 63924 11396 63980 11452
rect 66836 11396 66892 11452
rect 67172 11396 67228 11452
rect 82068 11396 82124 11452
rect 82964 11396 83020 11452
rect 83300 11396 83356 11452
rect 83524 11396 83580 11452
rect 84084 11396 84140 11452
rect 88564 11396 88620 11452
rect 88788 11396 88844 11452
rect 92708 11396 92764 11452
rect 99092 11396 99148 11452
rect 99316 11396 99372 11452
rect 113540 11396 113596 11452
rect 118580 11396 118636 11452
rect 119140 11396 119196 11452
rect 138628 11396 138684 11452
rect 141316 11396 141372 11452
rect 146020 11396 146076 11452
rect 164836 11396 164892 11452
rect 183428 11396 183484 11452
rect 189812 11396 189868 11452
rect 51716 11284 51772 11340
rect 51940 11284 51996 11340
rect 55300 11284 55356 11340
rect 56196 11284 56252 11340
rect 65044 11284 65100 11340
rect 69412 11284 69468 11340
rect 79828 11284 79884 11340
rect 80388 11284 80444 11340
rect 81956 11284 82012 11340
rect 82516 11284 82572 11340
rect 91140 11284 91196 11340
rect 102676 11284 102732 11340
rect 103572 11284 103628 11340
rect 104804 11284 104860 11340
rect 105028 11284 105084 11340
rect 109508 11284 109564 11340
rect 111076 11284 111132 11340
rect 116228 11284 116284 11340
rect 118804 11284 118860 11340
rect 126308 11284 126364 11340
rect 126532 11284 126588 11340
rect 133028 11284 133084 11340
rect 135940 11284 135996 11340
rect 136724 11284 136780 11340
rect 144228 11284 144284 11340
rect 162148 11284 162204 11340
rect 166740 11284 166796 11340
rect 68516 11172 68572 11228
rect 73668 11172 73724 11228
rect 83748 11172 83804 11228
rect 104132 11172 104188 11228
rect 114772 11172 114828 11228
rect 129444 11172 129500 11228
rect 144340 11172 144396 11228
rect 146244 11172 146300 11228
rect 158788 11172 158844 11228
rect 159012 11172 159068 11228
rect 182868 11172 182924 11228
rect 197316 11172 197372 11228
rect 77924 11060 77980 11116
rect 78372 11060 78428 11116
rect 79044 11060 79100 11116
rect 96852 11060 96908 11116
rect 102676 11060 102732 11116
rect 131012 11060 131068 11116
rect 133588 11060 133644 11116
rect 138292 11060 138348 11116
rect 154980 11060 155036 11116
rect 156100 11060 156156 11116
rect 160916 11060 160972 11116
rect 166740 11060 166796 11116
rect 179620 11060 179676 11116
rect 187460 11060 187516 11116
rect 82068 10948 82124 11004
rect 83188 10948 83244 11004
rect 103012 10948 103068 11004
rect 103236 10948 103292 11004
rect 113652 10948 113708 11004
rect 117572 10948 117628 11004
rect 121156 10948 121212 11004
rect 131124 10948 131180 11004
rect 132132 10948 132188 11004
rect 141092 10948 141148 11004
rect 164612 10948 164668 11004
rect 166628 10948 166684 11004
rect 187796 10948 187852 11004
rect 81620 10836 81676 10892
rect 86212 10836 86268 10892
rect 92148 10836 92204 10892
rect 98532 10836 98588 10892
rect 100548 10836 100604 10892
rect 102228 10836 102284 10892
rect 107716 10836 107772 10892
rect 107940 10836 107996 10892
rect 124516 10836 124572 10892
rect 133028 10836 133084 10892
rect 133700 10836 133756 10892
rect 139636 10836 139692 10892
rect 141428 10836 141484 10892
rect 148932 10836 148988 10892
rect 151284 10836 151340 10892
rect 154980 10836 155036 10892
rect 163380 10836 163436 10892
rect 180964 10836 181020 10892
rect 184324 10836 184380 10892
rect 77700 10724 77756 10780
rect 81508 10724 81564 10780
rect 86324 10724 86380 10780
rect 92036 10724 92092 10780
rect 101220 10724 101276 10780
rect 101780 10724 101836 10780
rect 103684 10724 103740 10780
rect 104692 10724 104748 10780
rect 117348 10724 117404 10780
rect 126308 10724 126364 10780
rect 137732 10724 137788 10780
rect 147700 10724 147756 10780
rect 149716 10724 149772 10780
rect 151508 10724 151564 10780
rect 59556 10612 59612 10668
rect 68404 10612 68460 10668
rect 68740 10612 68796 10668
rect 70756 10612 70812 10668
rect 100660 10612 100716 10668
rect 108388 10612 108444 10668
rect 118020 10612 118076 10668
rect 130900 10612 130956 10668
rect 139636 10612 139692 10668
rect 151060 10612 151116 10668
rect 159012 10612 159068 10668
rect 188020 10612 188076 10668
rect 105924 10500 105980 10556
rect 106708 10500 106764 10556
rect 133924 10500 133980 10556
rect 146020 10500 146076 10556
rect 162148 10500 162204 10556
rect 164948 10500 165004 10556
rect 56980 10388 57036 10444
rect 62132 10388 62188 10444
rect 68628 10388 68684 10444
rect 103124 10388 103180 10444
rect 116228 10388 116284 10444
rect 117348 10388 117404 10444
rect 117684 10388 117740 10444
rect 118244 10388 118300 10444
rect 129780 10388 129836 10444
rect 134260 10388 134316 10444
rect 139748 10388 139804 10444
rect 140980 10388 141036 10444
rect 145796 10388 145852 10444
rect 153188 10388 153244 10444
rect 161140 10388 161196 10444
rect 183428 10388 183484 10444
rect 194292 10388 194348 10444
rect 28756 10276 28812 10332
rect 44436 10276 44492 10332
rect 49140 10276 49196 10332
rect 53396 10276 53452 10332
rect 83524 10276 83580 10332
rect 97860 10276 97916 10332
rect 103572 10276 103628 10332
rect 104244 10276 104300 10332
rect 110964 10276 111020 10332
rect 126084 10276 126140 10332
rect 130900 10276 130956 10332
rect 141428 10276 141484 10332
rect 164836 10276 164892 10332
rect 166628 10276 166684 10332
rect 167860 10276 167916 10332
rect 173124 10276 173180 10332
rect 180964 10276 181020 10332
rect 28376 10164 28432 10220
rect 28480 10164 28536 10220
rect 28584 10164 28640 10220
rect 66948 10164 67004 10220
rect 77812 10164 77868 10220
rect 78260 10164 78316 10220
rect 79380 10164 79436 10220
rect 80500 10164 80556 10220
rect 80948 10164 81004 10220
rect 82404 10164 82460 10220
rect 82704 10164 82760 10220
rect 82808 10164 82864 10220
rect 82912 10164 82968 10220
rect 91700 10164 91756 10220
rect 96068 10164 96124 10220
rect 97300 10164 97356 10220
rect 98868 10164 98924 10220
rect 99092 10164 99148 10220
rect 100100 10164 100156 10220
rect 103012 10164 103068 10220
rect 103236 10164 103292 10220
rect 114884 10164 114940 10220
rect 115444 10164 115500 10220
rect 120036 10164 120092 10220
rect 121044 10164 121100 10220
rect 121268 10164 121324 10220
rect 125748 10164 125804 10220
rect 137032 10164 137088 10220
rect 137136 10164 137192 10220
rect 137240 10164 137296 10220
rect 149156 10164 149212 10220
rect 156212 10164 156268 10220
rect 157556 10164 157612 10220
rect 162820 10164 162876 10220
rect 164948 10164 165004 10220
rect 183764 10164 183820 10220
rect 190932 10164 190988 10220
rect 191360 10164 191416 10220
rect 191464 10164 191520 10220
rect 191568 10164 191624 10220
rect 16212 10052 16268 10108
rect 26740 10052 26796 10108
rect 36820 10052 36876 10108
rect 44436 10052 44492 10108
rect 51940 10052 51996 10108
rect 57204 10052 57260 10108
rect 62916 10052 62972 10108
rect 73444 10052 73500 10108
rect 73668 10052 73724 10108
rect 75012 10052 75068 10108
rect 76468 10052 76524 10108
rect 78820 10052 78876 10108
rect 80724 10052 80780 10108
rect 81396 10052 81452 10108
rect 83188 10052 83244 10108
rect 85876 10052 85932 10108
rect 86100 10052 86156 10108
rect 94500 10052 94556 10108
rect 105812 10052 105868 10108
rect 106036 10052 106092 10108
rect 112756 10052 112812 10108
rect 114436 10052 114492 10108
rect 118356 10052 118412 10108
rect 134260 10052 134316 10108
rect 141428 10052 141484 10108
rect 147812 10052 147868 10108
rect 152180 10052 152236 10108
rect 153412 10052 153468 10108
rect 157892 10052 157948 10108
rect 184324 10052 184380 10108
rect 190596 10052 190652 10108
rect 197316 10052 197372 10108
rect 77028 9940 77084 9996
rect 77700 9940 77756 9996
rect 77924 9940 77980 9996
rect 78708 9940 78764 9996
rect 82292 9940 82348 9996
rect 87892 9940 87948 9996
rect 89124 9940 89180 9996
rect 91028 9940 91084 9996
rect 97748 9940 97804 9996
rect 103684 9940 103740 9996
rect 106484 9940 106540 9996
rect 110404 9940 110460 9996
rect 115780 9940 115836 9996
rect 121604 9940 121660 9996
rect 121828 9940 121884 9996
rect 142772 9940 142828 9996
rect 152852 9940 152908 9996
rect 166292 9940 166348 9996
rect 61460 9828 61516 9884
rect 68964 9828 69020 9884
rect 72212 9828 72268 9884
rect 90468 9828 90524 9884
rect 90692 9828 90748 9884
rect 106036 9828 106092 9884
rect 111188 9828 111244 9884
rect 112980 9828 113036 9884
rect 116788 9828 116844 9884
rect 178052 9940 178108 9996
rect 122724 9828 122780 9884
rect 134148 9828 134204 9884
rect 139412 9828 139468 9884
rect 142436 9828 142492 9884
rect 158004 9828 158060 9884
rect 174692 9828 174748 9884
rect 182756 9828 182812 9884
rect 184996 9828 185052 9884
rect 186452 9828 186508 9884
rect 198212 9828 198268 9884
rect 200340 9828 200396 9884
rect 58660 9716 58716 9772
rect 77364 9716 77420 9772
rect 83188 9716 83244 9772
rect 83412 9716 83468 9772
rect 91028 9716 91084 9772
rect 99316 9716 99372 9772
rect 99876 9716 99932 9772
rect 102788 9716 102844 9772
rect 104244 9716 104300 9772
rect 105924 9716 105980 9772
rect 117572 9716 117628 9772
rect 119924 9716 119980 9772
rect 135268 9716 135324 9772
rect 140980 9716 141036 9772
rect 142772 9716 142828 9772
rect 145684 9716 145740 9772
rect 157780 9716 157836 9772
rect 192164 9716 192220 9772
rect 194740 9716 194796 9772
rect 204484 9716 204540 9772
rect 10164 9604 10220 9660
rect 43204 9604 43260 9660
rect 46116 9604 46172 9660
rect 69524 9604 69580 9660
rect 72996 9604 73052 9660
rect 76244 9604 76300 9660
rect 77252 9604 77308 9660
rect 78148 9604 78204 9660
rect 79492 9604 79548 9660
rect 83076 9604 83132 9660
rect 85540 9604 85596 9660
rect 93044 9604 93100 9660
rect 107492 9604 107548 9660
rect 114772 9604 114828 9660
rect 124628 9604 124684 9660
rect 124852 9604 124908 9660
rect 144228 9604 144284 9660
rect 146132 9604 146188 9660
rect 149044 9604 149100 9660
rect 151284 9604 151340 9660
rect 152852 9604 152908 9660
rect 188244 9604 188300 9660
rect 189924 9604 189980 9660
rect 197764 9604 197820 9660
rect 197988 9604 198044 9660
rect 91476 9492 91532 9548
rect 92036 9492 92092 9548
rect 100660 9492 100716 9548
rect 101892 9492 101948 9548
rect 102452 9492 102508 9548
rect 111188 9492 111244 9548
rect 120036 9492 120092 9548
rect 182868 9492 182924 9548
rect 205716 9492 205772 9548
rect 206388 9492 206444 9548
rect 55540 9380 55596 9436
rect 55644 9380 55700 9436
rect 55748 9380 55804 9436
rect 83300 9380 83356 9436
rect 84420 9380 84476 9436
rect 89124 9380 89180 9436
rect 89460 9380 89516 9436
rect 90244 9380 90300 9436
rect 90468 9380 90524 9436
rect 99652 9380 99708 9436
rect 99988 9380 100044 9436
rect 104580 9380 104636 9436
rect 109060 9380 109116 9436
rect 109396 9380 109452 9436
rect 109868 9380 109924 9436
rect 109972 9380 110028 9436
rect 110076 9380 110132 9436
rect 110852 9380 110908 9436
rect 118244 9380 118300 9436
rect 119028 9380 119084 9436
rect 21700 9268 21756 9324
rect 44548 9268 44604 9324
rect 69972 9268 70028 9324
rect 72548 9268 72604 9324
rect 78372 9268 78428 9324
rect 79940 9268 79996 9324
rect 81844 9268 81900 9324
rect 98644 9268 98700 9324
rect 100660 9268 100716 9324
rect 101220 9268 101276 9324
rect 115780 9268 115836 9324
rect 117684 9268 117740 9324
rect 119364 9268 119420 9324
rect 119588 9268 119644 9324
rect 120036 9268 120092 9324
rect 120708 9268 120764 9324
rect 133364 9380 133420 9436
rect 135268 9380 135324 9436
rect 142772 9380 142828 9436
rect 144452 9380 144508 9436
rect 149492 9380 149548 9436
rect 150388 9380 150444 9436
rect 164196 9380 164252 9436
rect 164300 9380 164356 9436
rect 164404 9380 164460 9436
rect 182980 9380 183036 9436
rect 183764 9380 183820 9436
rect 199892 9380 199948 9436
rect 191044 9268 191100 9324
rect 71204 9156 71260 9212
rect 71428 9156 71484 9212
rect 75012 9156 75068 9212
rect 78820 9156 78876 9212
rect 82292 9156 82348 9212
rect 82516 9156 82572 9212
rect 85764 9156 85820 9212
rect 89236 9156 89292 9212
rect 92036 9156 92092 9212
rect 92260 9156 92316 9212
rect 110740 9156 110796 9212
rect 116004 9156 116060 9212
rect 116900 9156 116956 9212
rect 117124 9156 117180 9212
rect 121268 9156 121324 9212
rect 121604 9156 121660 9212
rect 131012 9156 131068 9212
rect 135940 9156 135996 9212
rect 140308 9156 140364 9212
rect 168980 9156 169036 9212
rect 178164 9156 178220 9212
rect 180852 9156 180908 9212
rect 190932 9156 190988 9212
rect 193844 9156 193900 9212
rect 195412 9156 195468 9212
rect 197988 9156 198044 9212
rect 212548 9156 212604 9212
rect 10052 9044 10108 9100
rect 47348 9044 47404 9100
rect 60228 9044 60284 9100
rect 103012 9044 103068 9100
rect 110404 9044 110460 9100
rect 110852 9044 110908 9100
rect 124628 9044 124684 9100
rect 132468 9044 132524 9100
rect 138516 9044 138572 9100
rect 158340 9044 158396 9100
rect 170996 9044 171052 9100
rect 173348 9044 173404 9100
rect 26404 8932 26460 8988
rect 52276 8932 52332 8988
rect 57204 8932 57260 8988
rect 60340 8932 60396 8988
rect 80500 8932 80556 8988
rect 84868 8932 84924 8988
rect 85092 8932 85148 8988
rect 85428 8932 85484 8988
rect 90916 8932 90972 8988
rect 66724 8820 66780 8876
rect 67060 8820 67116 8876
rect 70420 8820 70476 8876
rect 72772 8820 72828 8876
rect 72996 8820 73052 8876
rect 118132 8932 118188 8988
rect 118692 8932 118748 8988
rect 126980 8932 127036 8988
rect 127204 8932 127260 8988
rect 168980 8932 169036 8988
rect 201908 8932 201964 8988
rect 206388 8932 206444 8988
rect 208404 8932 208460 8988
rect 88676 8820 88732 8876
rect 90804 8820 90860 8876
rect 103460 8820 103516 8876
rect 106596 8820 106652 8876
rect 107492 8820 107548 8876
rect 127988 8820 128044 8876
rect 134036 8820 134092 8876
rect 79716 8708 79772 8764
rect 79940 8708 79996 8764
rect 80500 8708 80556 8764
rect 86436 8708 86492 8764
rect 88116 8708 88172 8764
rect 118468 8708 118524 8764
rect 119364 8708 119420 8764
rect 133364 8708 133420 8764
rect 135604 8708 135660 8764
rect 141764 8708 141820 8764
rect 172900 8708 172956 8764
rect 188020 8708 188076 8764
rect 193172 8708 193228 8764
rect 212548 8708 212604 8764
rect 28376 8596 28432 8652
rect 28480 8596 28536 8652
rect 28584 8596 28640 8652
rect 70420 8596 70476 8652
rect 77812 8596 77868 8652
rect 81284 8596 81340 8652
rect 82704 8596 82760 8652
rect 82808 8596 82864 8652
rect 82912 8596 82968 8652
rect 83748 8596 83804 8652
rect 83972 8596 84028 8652
rect 85988 8596 86044 8652
rect 87108 8596 87164 8652
rect 87332 8596 87388 8652
rect 91700 8596 91756 8652
rect 102452 8596 102508 8652
rect 102676 8596 102732 8652
rect 106372 8596 106428 8652
rect 106596 8596 106652 8652
rect 109172 8596 109228 8652
rect 115444 8596 115500 8652
rect 118132 8596 118188 8652
rect 123508 8596 123564 8652
rect 131124 8596 131180 8652
rect 137032 8596 137088 8652
rect 137136 8596 137192 8652
rect 137240 8596 137296 8652
rect 191360 8596 191416 8652
rect 191464 8596 191520 8652
rect 191568 8596 191624 8652
rect 199444 8596 199500 8652
rect 201908 8596 201964 8652
rect 30100 8484 30156 8540
rect 55972 8484 56028 8540
rect 60676 8484 60732 8540
rect 72996 8484 73052 8540
rect 78484 8484 78540 8540
rect 86660 8484 86716 8540
rect 87444 8484 87500 8540
rect 91364 8484 91420 8540
rect 95284 8484 95340 8540
rect 96964 8484 97020 8540
rect 103684 8484 103740 8540
rect 108612 8484 108668 8540
rect 126980 8484 127036 8540
rect 138516 8484 138572 8540
rect 139748 8484 139804 8540
rect 144676 8484 144732 8540
rect 148484 8484 148540 8540
rect 157444 8484 157500 8540
rect 170436 8484 170492 8540
rect 181300 8484 181356 8540
rect 181860 8484 181916 8540
rect 193732 8484 193788 8540
rect 200116 8484 200172 8540
rect 63252 8372 63308 8428
rect 63476 8372 63532 8428
rect 72660 8372 72716 8428
rect 74900 8372 74956 8428
rect 86772 8372 86828 8428
rect 99204 8372 99260 8428
rect 100436 8372 100492 8428
rect 100660 8372 100716 8428
rect 118244 8372 118300 8428
rect 118804 8372 118860 8428
rect 124852 8372 124908 8428
rect 127988 8372 128044 8428
rect 145460 8372 145516 8428
rect 149380 8372 149436 8428
rect 152740 8372 152796 8428
rect 156100 8372 156156 8428
rect 10276 8260 10332 8316
rect 66948 8260 67004 8316
rect 70532 8260 70588 8316
rect 74340 8260 74396 8316
rect 79044 8260 79100 8316
rect 79492 8260 79548 8316
rect 85540 8260 85596 8316
rect 89460 8260 89516 8316
rect 89908 8260 89964 8316
rect 104132 8260 104188 8316
rect 110404 8260 110460 8316
rect 110740 8260 110796 8316
rect 117124 8260 117180 8316
rect 117684 8260 117740 8316
rect 121828 8260 121884 8316
rect 128436 8260 128492 8316
rect 133700 8260 133756 8316
rect 144564 8260 144620 8316
rect 148484 8260 148540 8316
rect 152852 8260 152908 8316
rect 158340 8260 158396 8316
rect 167860 8260 167916 8316
rect 191044 8372 191100 8428
rect 185108 8260 185164 8316
rect 187572 8260 187628 8316
rect 197540 8260 197596 8316
rect 199892 8260 199948 8316
rect 60004 8148 60060 8204
rect 72436 8148 72492 8204
rect 81844 8148 81900 8204
rect 82292 8148 82348 8204
rect 84532 8148 84588 8204
rect 84756 8148 84812 8204
rect 93268 8148 93324 8204
rect 98644 8148 98700 8204
rect 98868 8148 98924 8204
rect 108612 8148 108668 8204
rect 112980 8148 113036 8204
rect 116452 8148 116508 8204
rect 117908 8148 117964 8204
rect 120260 8148 120316 8204
rect 120820 8148 120876 8204
rect 129444 8148 129500 8204
rect 134932 8148 134988 8204
rect 145012 8148 145068 8204
rect 146020 8148 146076 8204
rect 13972 8036 14028 8092
rect 19348 8036 19404 8092
rect 47348 8036 47404 8092
rect 48580 8036 48636 8092
rect 62580 8036 62636 8092
rect 74900 8036 74956 8092
rect 75124 8036 75180 8092
rect 78708 8036 78764 8092
rect 80948 8036 81004 8092
rect 81284 8036 81340 8092
rect 82404 8036 82460 8092
rect 83972 8036 84028 8092
rect 91252 8036 91308 8092
rect 96964 8036 97020 8092
rect 101220 8036 101276 8092
rect 101444 8036 101500 8092
rect 102228 8036 102284 8092
rect 104804 8036 104860 8092
rect 111076 8036 111132 8092
rect 111300 8036 111356 8092
rect 112308 8036 112364 8092
rect 118244 8036 118300 8092
rect 119812 8036 119868 8092
rect 121492 8036 121548 8092
rect 123396 8036 123452 8092
rect 127092 8036 127148 8092
rect 132916 8036 132972 8092
rect 135828 8036 135884 8092
rect 136500 8036 136556 8092
rect 137508 8036 137564 8092
rect 137956 8036 138012 8092
rect 144788 8036 144844 8092
rect 175028 8036 175084 8092
rect 181076 8036 181132 8092
rect 181300 8036 181356 8092
rect 193060 8036 193116 8092
rect 216356 8036 216412 8092
rect 25956 7924 26012 7980
rect 53620 7924 53676 7980
rect 54068 7924 54124 7980
rect 57428 7924 57484 7980
rect 60676 7924 60732 7980
rect 70532 7924 70588 7980
rect 77252 7924 77308 7980
rect 77476 7924 77532 7980
rect 84308 7924 84364 7980
rect 85092 7924 85148 7980
rect 86884 7924 86940 7980
rect 87220 7924 87276 7980
rect 91028 7924 91084 7980
rect 91924 7924 91980 7980
rect 96852 7924 96908 7980
rect 107492 7924 107548 7980
rect 107716 7924 107772 7980
rect 113876 7924 113932 7980
rect 120596 7924 120652 7980
rect 120932 7924 120988 7980
rect 134820 7924 134876 7980
rect 141204 7924 141260 7980
rect 142996 7924 143052 7980
rect 144228 7924 144284 7980
rect 147700 7924 147756 7980
rect 147924 7924 147980 7980
rect 150388 7924 150444 7980
rect 162932 7924 162988 7980
rect 166404 7924 166460 7980
rect 203700 7924 203756 7980
rect 203924 7924 203980 7980
rect 55540 7812 55596 7868
rect 55644 7812 55700 7868
rect 55748 7812 55804 7868
rect 60452 7812 60508 7868
rect 90468 7812 90524 7868
rect 102900 7812 102956 7868
rect 104132 7812 104188 7868
rect 108276 7812 108332 7868
rect 109868 7812 109924 7868
rect 109972 7812 110028 7868
rect 110076 7812 110132 7868
rect 114324 7812 114380 7868
rect 116676 7812 116732 7868
rect 117124 7812 117180 7868
rect 119476 7812 119532 7868
rect 127204 7812 127260 7868
rect 129220 7812 129276 7868
rect 137956 7812 138012 7868
rect 149380 7812 149436 7868
rect 157780 7812 157836 7868
rect 164196 7812 164252 7868
rect 164300 7812 164356 7868
rect 164404 7812 164460 7868
rect 166292 7812 166348 7868
rect 181076 7812 181132 7868
rect 208404 7812 208460 7868
rect 60788 7700 60844 7756
rect 85876 7700 85932 7756
rect 91700 7700 91756 7756
rect 114100 7700 114156 7756
rect 115108 7700 115164 7756
rect 115332 7700 115388 7756
rect 120036 7700 120092 7756
rect 126868 7700 126924 7756
rect 127092 7700 127148 7756
rect 128436 7700 128492 7756
rect 133364 7700 133420 7756
rect 136836 7700 136892 7756
rect 141204 7700 141260 7756
rect 142548 7700 142604 7756
rect 142772 7700 142828 7756
rect 154196 7700 154252 7756
rect 155988 7700 156044 7756
rect 156548 7700 156604 7756
rect 167860 7700 167916 7756
rect 177716 7700 177772 7756
rect 182980 7700 183036 7756
rect 188916 7700 188972 7756
rect 191716 7700 191772 7756
rect 196420 7700 196476 7756
rect 42196 7588 42252 7644
rect 46228 7588 46284 7644
rect 62580 7588 62636 7644
rect 63812 7588 63868 7644
rect 71988 7588 72044 7644
rect 74340 7588 74396 7644
rect 79716 7588 79772 7644
rect 83076 7588 83132 7644
rect 83972 7588 84028 7644
rect 91812 7588 91868 7644
rect 106148 7588 106204 7644
rect 106372 7588 106428 7644
rect 115220 7588 115276 7644
rect 117796 7588 117852 7644
rect 118692 7588 118748 7644
rect 119364 7588 119420 7644
rect 134260 7588 134316 7644
rect 139524 7588 139580 7644
rect 139748 7588 139804 7644
rect 143556 7588 143612 7644
rect 146916 7588 146972 7644
rect 148820 7588 148876 7644
rect 149044 7588 149100 7644
rect 157108 7588 157164 7644
rect 176148 7588 176204 7644
rect 190820 7588 190876 7644
rect 196644 7588 196700 7644
rect 68516 7476 68572 7532
rect 71316 7476 71372 7532
rect 75348 7476 75404 7532
rect 78260 7476 78316 7532
rect 78484 7476 78540 7532
rect 86100 7476 86156 7532
rect 86884 7476 86940 7532
rect 91028 7476 91084 7532
rect 99876 7476 99932 7532
rect 103460 7476 103516 7532
rect 105140 7476 105196 7532
rect 117348 7476 117404 7532
rect 118244 7476 118300 7532
rect 127092 7476 127148 7532
rect 146020 7476 146076 7532
rect 147588 7476 147644 7532
rect 152740 7476 152796 7532
rect 192836 7476 192892 7532
rect 203924 7476 203980 7532
rect 18228 7364 18284 7420
rect 60004 7364 60060 7420
rect 62804 7364 62860 7420
rect 64596 7364 64652 7420
rect 67956 7364 68012 7420
rect 75796 7364 75852 7420
rect 80052 7364 80108 7420
rect 83748 7364 83804 7420
rect 84756 7364 84812 7420
rect 91476 7364 91532 7420
rect 91700 7364 91756 7420
rect 97748 7364 97804 7420
rect 99428 7364 99484 7420
rect 102340 7364 102396 7420
rect 103796 7364 103852 7420
rect 115220 7364 115276 7420
rect 118468 7364 118524 7420
rect 121604 7364 121660 7420
rect 133364 7364 133420 7420
rect 138180 7364 138236 7420
rect 142436 7364 142492 7420
rect 149268 7364 149324 7420
rect 149604 7364 149660 7420
rect 154084 7364 154140 7420
rect 198212 7364 198268 7420
rect 201572 7364 201628 7420
rect 211204 7364 211260 7420
rect 214452 7364 214508 7420
rect 69748 7252 69804 7308
rect 71988 7252 72044 7308
rect 72324 7252 72380 7308
rect 73892 7252 73948 7308
rect 75908 7252 75964 7308
rect 78148 7252 78204 7308
rect 78932 7252 78988 7308
rect 80948 7252 81004 7308
rect 81172 7252 81228 7308
rect 81396 7252 81452 7308
rect 84196 7252 84252 7308
rect 90244 7252 90300 7308
rect 105700 7252 105756 7308
rect 106148 7252 106204 7308
rect 114324 7252 114380 7308
rect 121268 7252 121324 7308
rect 126980 7252 127036 7308
rect 144676 7252 144732 7308
rect 150052 7252 150108 7308
rect 162932 7252 162988 7308
rect 172900 7252 172956 7308
rect 177940 7252 177996 7308
rect 200004 7252 200060 7308
rect 25620 7140 25676 7196
rect 30660 7140 30716 7196
rect 34580 7140 34636 7196
rect 44660 7140 44716 7196
rect 72100 7140 72156 7196
rect 75012 7140 75068 7196
rect 76132 7140 76188 7196
rect 82516 7140 82572 7196
rect 83412 7140 83468 7196
rect 83636 7140 83692 7196
rect 91588 7140 91644 7196
rect 91924 7140 91980 7196
rect 100436 7140 100492 7196
rect 100996 7140 101052 7196
rect 102004 7140 102060 7196
rect 102228 7140 102284 7196
rect 103348 7140 103404 7196
rect 103908 7140 103964 7196
rect 115220 7140 115276 7196
rect 115444 7140 115500 7196
rect 117684 7140 117740 7196
rect 121828 7140 121884 7196
rect 122500 7140 122556 7196
rect 126084 7140 126140 7196
rect 140532 7140 140588 7196
rect 142436 7140 142492 7196
rect 142660 7140 142716 7196
rect 28376 7028 28432 7084
rect 28480 7028 28536 7084
rect 28584 7028 28640 7084
rect 82704 7028 82760 7084
rect 82808 7028 82864 7084
rect 82912 7028 82968 7084
rect 84644 7028 84700 7084
rect 85988 7028 86044 7084
rect 88004 7028 88060 7084
rect 90244 7028 90300 7084
rect 91252 7028 91308 7084
rect 91476 7028 91532 7084
rect 103796 7028 103852 7084
rect 110852 7028 110908 7084
rect 121156 7028 121212 7084
rect 121940 7028 121996 7084
rect 127092 7028 127148 7084
rect 129332 7028 129388 7084
rect 136836 7028 136892 7084
rect 137032 7028 137088 7084
rect 137136 7028 137192 7084
rect 137240 7028 137296 7084
rect 144452 7028 144508 7084
rect 149044 7028 149100 7084
rect 149492 7028 149548 7084
rect 154196 7028 154252 7084
rect 173908 7028 173964 7084
rect 186788 7028 186844 7084
rect 191360 7028 191416 7084
rect 191464 7028 191520 7084
rect 191568 7028 191624 7084
rect 67956 6916 68012 6972
rect 75348 6916 75404 6972
rect 78148 6916 78204 6972
rect 80388 6916 80444 6972
rect 82068 6916 82124 6972
rect 83524 6916 83580 6972
rect 87444 6916 87500 6972
rect 88564 6916 88620 6972
rect 90580 6916 90636 6972
rect 99540 6916 99596 6972
rect 100324 6916 100380 6972
rect 105140 6916 105196 6972
rect 106932 6916 106988 6972
rect 109396 6916 109452 6972
rect 122500 6916 122556 6972
rect 122724 6916 122780 6972
rect 134260 6916 134316 6972
rect 135940 6916 135996 6972
rect 137620 6916 137676 6972
rect 138180 6916 138236 6972
rect 149940 6916 149996 6972
rect 178836 6916 178892 6972
rect 186452 6916 186508 6972
rect 68740 6804 68796 6860
rect 69188 6804 69244 6860
rect 74900 6804 74956 6860
rect 76244 6804 76300 6860
rect 80052 6804 80108 6860
rect 82180 6804 82236 6860
rect 86212 6804 86268 6860
rect 86660 6804 86716 6860
rect 91812 6804 91868 6860
rect 109508 6804 109564 6860
rect 111300 6804 111356 6860
rect 112084 6804 112140 6860
rect 114324 6804 114380 6860
rect 114660 6804 114716 6860
rect 115332 6804 115388 6860
rect 115668 6804 115724 6860
rect 116564 6804 116620 6860
rect 117460 6804 117516 6860
rect 143220 6804 143276 6860
rect 143780 6804 143836 6860
rect 145124 6804 145180 6860
rect 149156 6804 149212 6860
rect 157108 6804 157164 6860
rect 176148 6804 176204 6860
rect 182644 6804 182700 6860
rect 67060 6692 67116 6748
rect 73668 6692 73724 6748
rect 79268 6692 79324 6748
rect 79492 6692 79548 6748
rect 80388 6692 80444 6748
rect 80612 6692 80668 6748
rect 82516 6692 82572 6748
rect 84644 6692 84700 6748
rect 86884 6692 86940 6748
rect 87108 6692 87164 6748
rect 87556 6692 87612 6748
rect 103236 6692 103292 6748
rect 113988 6692 114044 6748
rect 115556 6692 115612 6748
rect 115780 6692 115836 6748
rect 117124 6692 117180 6748
rect 117348 6692 117404 6748
rect 130788 6692 130844 6748
rect 141316 6692 141372 6748
rect 188244 6692 188300 6748
rect 191716 6692 191772 6748
rect 196420 6692 196476 6748
rect 200004 6692 200060 6748
rect 28756 6580 28812 6636
rect 63700 6580 63756 6636
rect 68628 6580 68684 6636
rect 80836 6580 80892 6636
rect 83076 6580 83132 6636
rect 85876 6580 85932 6636
rect 90580 6580 90636 6636
rect 102340 6580 102396 6636
rect 103124 6580 103180 6636
rect 108276 6580 108332 6636
rect 110292 6580 110348 6636
rect 113652 6580 113708 6636
rect 116564 6580 116620 6636
rect 117460 6580 117516 6636
rect 122276 6580 122332 6636
rect 122500 6580 122556 6636
rect 124964 6580 125020 6636
rect 129556 6580 129612 6636
rect 37716 6468 37772 6524
rect 67060 6468 67116 6524
rect 82516 6468 82572 6524
rect 84308 6468 84364 6524
rect 90692 6468 90748 6524
rect 93268 6468 93324 6524
rect 95844 6468 95900 6524
rect 101108 6468 101164 6524
rect 101332 6468 101388 6524
rect 104692 6468 104748 6524
rect 105700 6468 105756 6524
rect 112196 6468 112252 6524
rect 114100 6468 114156 6524
rect 117236 6468 117292 6524
rect 117796 6468 117852 6524
rect 118020 6468 118076 6524
rect 118580 6468 118636 6524
rect 119140 6468 119196 6524
rect 119364 6468 119420 6524
rect 129220 6468 129276 6524
rect 78708 6356 78764 6412
rect 81956 6356 82012 6412
rect 83860 6356 83916 6412
rect 84084 6356 84140 6412
rect 86548 6356 86604 6412
rect 98196 6356 98252 6412
rect 103572 6356 103628 6412
rect 126644 6356 126700 6412
rect 134260 6580 134316 6636
rect 138628 6580 138684 6636
rect 144116 6580 144172 6636
rect 146020 6580 146076 6636
rect 149380 6580 149436 6636
rect 151732 6580 151788 6636
rect 154420 6580 154476 6636
rect 166852 6580 166908 6636
rect 167636 6580 167692 6636
rect 178276 6580 178332 6636
rect 179620 6580 179676 6636
rect 179844 6580 179900 6636
rect 189812 6580 189868 6636
rect 196532 6580 196588 6636
rect 200900 6580 200956 6636
rect 142660 6468 142716 6524
rect 144228 6468 144284 6524
rect 145460 6468 145516 6524
rect 153524 6468 153580 6524
rect 156324 6468 156380 6524
rect 161028 6468 161084 6524
rect 166292 6468 166348 6524
rect 168644 6468 168700 6524
rect 170996 6468 171052 6524
rect 179732 6468 179788 6524
rect 179956 6468 180012 6524
rect 192836 6468 192892 6524
rect 193732 6468 193788 6524
rect 133028 6356 133084 6412
rect 154756 6356 154812 6412
rect 156772 6356 156828 6412
rect 165172 6356 165228 6412
rect 173796 6356 173852 6412
rect 174132 6356 174188 6412
rect 189364 6356 189420 6412
rect 193172 6356 193228 6412
rect 200900 6356 200956 6412
rect 55540 6244 55596 6300
rect 55644 6244 55700 6300
rect 55748 6244 55804 6300
rect 57428 6244 57484 6300
rect 58436 6244 58492 6300
rect 60004 6244 60060 6300
rect 66836 6244 66892 6300
rect 68180 6244 68236 6300
rect 70868 6244 70924 6300
rect 73108 6244 73164 6300
rect 84980 6244 85036 6300
rect 85652 6244 85708 6300
rect 91476 6244 91532 6300
rect 109620 6244 109676 6300
rect 109868 6244 109924 6300
rect 109972 6244 110028 6300
rect 110076 6244 110132 6300
rect 121828 6244 121884 6300
rect 122948 6244 123004 6300
rect 124964 6244 125020 6300
rect 133476 6244 133532 6300
rect 144004 6244 144060 6300
rect 144452 6244 144508 6300
rect 155988 6244 156044 6300
rect 164196 6244 164252 6300
rect 164300 6244 164356 6300
rect 164404 6244 164460 6300
rect 164612 6244 164668 6300
rect 168644 6244 168700 6300
rect 191828 6244 191884 6300
rect 194292 6244 194348 6300
rect 197764 6244 197820 6300
rect 203252 6244 203308 6300
rect 68628 6132 68684 6188
rect 84420 6132 84476 6188
rect 85204 6132 85260 6188
rect 86436 6132 86492 6188
rect 87556 6132 87612 6188
rect 88900 6132 88956 6188
rect 90692 6132 90748 6188
rect 98532 6132 98588 6188
rect 100100 6132 100156 6188
rect 113876 6132 113932 6188
rect 116004 6132 116060 6188
rect 141764 6132 141820 6188
rect 145348 6132 145404 6188
rect 149268 6132 149324 6188
rect 173908 6132 173964 6188
rect 179620 6132 179676 6188
rect 212548 6132 212604 6188
rect 35588 6020 35644 6076
rect 52052 6020 52108 6076
rect 89796 6020 89852 6076
rect 122164 6020 122220 6076
rect 122612 6020 122668 6076
rect 123508 6020 123564 6076
rect 131460 6020 131516 6076
rect 156772 6020 156828 6076
rect 159236 6020 159292 6076
rect 166516 6020 166572 6076
rect 170996 6020 171052 6076
rect 174692 6020 174748 6076
rect 175140 6020 175196 6076
rect 193284 6020 193340 6076
rect 194852 6020 194908 6076
rect 205716 6020 205772 6076
rect 30100 5908 30156 5964
rect 51828 5908 51884 5964
rect 52164 5908 52220 5964
rect 73780 5908 73836 5964
rect 74004 5908 74060 5964
rect 75460 5908 75516 5964
rect 76468 5908 76524 5964
rect 82404 5908 82460 5964
rect 84644 5908 84700 5964
rect 85764 5908 85820 5964
rect 99428 5908 99484 5964
rect 100660 5908 100716 5964
rect 109620 5908 109676 5964
rect 113764 5908 113820 5964
rect 117012 5908 117068 5964
rect 118804 5908 118860 5964
rect 119028 5908 119084 5964
rect 121268 5908 121324 5964
rect 121828 5908 121884 5964
rect 129556 5908 129612 5964
rect 131236 5908 131292 5964
rect 166404 5908 166460 5964
rect 41748 5796 41804 5852
rect 42420 5796 42476 5852
rect 51604 5796 51660 5852
rect 52052 5796 52108 5852
rect 64596 5796 64652 5852
rect 67284 5796 67340 5852
rect 73556 5796 73612 5852
rect 75908 5796 75964 5852
rect 78596 5796 78652 5852
rect 81508 5796 81564 5852
rect 83300 5796 83356 5852
rect 85204 5796 85260 5852
rect 89236 5796 89292 5852
rect 102116 5796 102172 5852
rect 103236 5796 103292 5852
rect 104468 5796 104524 5852
rect 114212 5796 114268 5852
rect 115444 5796 115500 5852
rect 115892 5796 115948 5852
rect 119364 5796 119420 5852
rect 119924 5796 119980 5852
rect 126644 5796 126700 5852
rect 133140 5796 133196 5852
rect 134260 5796 134316 5852
rect 140980 5796 141036 5852
rect 141204 5796 141260 5852
rect 146244 5796 146300 5852
rect 146916 5796 146972 5852
rect 150276 5796 150332 5852
rect 150948 5796 151004 5852
rect 210308 5796 210364 5852
rect 18116 5684 18172 5740
rect 33908 5684 33964 5740
rect 37716 5684 37772 5740
rect 47012 5684 47068 5740
rect 69412 5684 69468 5740
rect 73108 5684 73164 5740
rect 74788 5684 74844 5740
rect 75012 5684 75068 5740
rect 80052 5684 80108 5740
rect 80724 5684 80780 5740
rect 84644 5684 84700 5740
rect 87108 5684 87164 5740
rect 87332 5684 87388 5740
rect 90468 5684 90524 5740
rect 98196 5684 98252 5740
rect 98420 5684 98476 5740
rect 98980 5684 99036 5740
rect 100772 5684 100828 5740
rect 121156 5684 121212 5740
rect 122276 5684 122332 5740
rect 139412 5684 139468 5740
rect 157220 5684 157276 5740
rect 197764 5684 197820 5740
rect 212548 5684 212604 5740
rect 212772 5684 212828 5740
rect 212996 5684 213052 5740
rect 41748 5572 41804 5628
rect 47460 5572 47516 5628
rect 54180 5572 54236 5628
rect 73668 5572 73724 5628
rect 75796 5572 75852 5628
rect 78708 5572 78764 5628
rect 78932 5572 78988 5628
rect 87892 5572 87948 5628
rect 88340 5572 88396 5628
rect 89796 5572 89852 5628
rect 90020 5572 90076 5628
rect 91700 5572 91756 5628
rect 92260 5572 92316 5628
rect 92596 5572 92652 5628
rect 109508 5572 109564 5628
rect 118580 5572 118636 5628
rect 119028 5572 119084 5628
rect 123508 5572 123564 5628
rect 131012 5572 131068 5628
rect 144788 5572 144844 5628
rect 145348 5572 145404 5628
rect 145684 5572 145740 5628
rect 155988 5572 156044 5628
rect 161476 5572 161532 5628
rect 173796 5572 173852 5628
rect 187908 5572 187964 5628
rect 188692 5572 188748 5628
rect 28376 5460 28432 5516
rect 28480 5460 28536 5516
rect 28584 5460 28640 5516
rect 33908 5460 33964 5516
rect 57428 5460 57484 5516
rect 73220 5460 73276 5516
rect 73444 5460 73500 5516
rect 75012 5460 75068 5516
rect 81396 5460 81452 5516
rect 82704 5460 82760 5516
rect 82808 5460 82864 5516
rect 82912 5460 82968 5516
rect 83524 5460 83580 5516
rect 98196 5460 98252 5516
rect 99428 5460 99484 5516
rect 101444 5460 101500 5516
rect 101668 5460 101724 5516
rect 102340 5460 102396 5516
rect 110292 5460 110348 5516
rect 111972 5460 112028 5516
rect 114212 5460 114268 5516
rect 114660 5460 114716 5516
rect 137032 5460 137088 5516
rect 137136 5460 137192 5516
rect 137240 5460 137296 5516
rect 137508 5460 137564 5516
rect 137844 5460 137900 5516
rect 161140 5460 161196 5516
rect 162260 5460 162316 5516
rect 191360 5460 191416 5516
rect 191464 5460 191520 5516
rect 191568 5460 191624 5516
rect 84308 5348 84364 5404
rect 84532 5348 84588 5404
rect 92372 5348 92428 5404
rect 122724 5348 122780 5404
rect 129332 5348 129388 5404
rect 129556 5348 129612 5404
rect 131236 5348 131292 5404
rect 141092 5348 141148 5404
rect 144004 5348 144060 5404
rect 150276 5348 150332 5404
rect 177940 5348 177996 5404
rect 181300 5348 181356 5404
rect 211316 5348 211372 5404
rect 68404 5236 68460 5292
rect 70868 5236 70924 5292
rect 73780 5236 73836 5292
rect 91476 5236 91532 5292
rect 91700 5236 91756 5292
rect 101220 5236 101276 5292
rect 103012 5236 103068 5292
rect 103236 5236 103292 5292
rect 107380 5236 107436 5292
rect 107604 5236 107660 5292
rect 113204 5236 113260 5292
rect 116676 5236 116732 5292
rect 119028 5236 119084 5292
rect 119252 5236 119308 5292
rect 128548 5236 128604 5292
rect 129668 5236 129724 5292
rect 131348 5236 131404 5292
rect 139188 5236 139244 5292
rect 142548 5236 142604 5292
rect 145684 5236 145740 5292
rect 159572 5236 159628 5292
rect 19236 5124 19292 5180
rect 23044 5124 23100 5180
rect 55972 5124 56028 5180
rect 57428 5124 57484 5180
rect 58660 5124 58716 5180
rect 73332 5124 73388 5180
rect 78708 5124 78764 5180
rect 79044 5124 79100 5180
rect 79716 5124 79772 5180
rect 85092 5124 85148 5180
rect 86212 5124 86268 5180
rect 87444 5124 87500 5180
rect 91924 5124 91980 5180
rect 92260 5124 92316 5180
rect 145124 5124 145180 5180
rect 166740 5124 166796 5180
rect 177716 5124 177772 5180
rect 178052 5124 178108 5180
rect 21140 5012 21196 5068
rect 23380 5012 23436 5068
rect 49812 5012 49868 5068
rect 71428 5012 71484 5068
rect 77140 5012 77196 5068
rect 90020 5012 90076 5068
rect 90244 5012 90300 5068
rect 98868 5012 98924 5068
rect 115668 5012 115724 5068
rect 148596 5012 148652 5068
rect 154532 5012 154588 5068
rect 188916 5012 188972 5068
rect 9604 4900 9660 4956
rect 11620 4900 11676 4956
rect 16436 4900 16492 4956
rect 35700 4900 35756 4956
rect 56196 4900 56252 4956
rect 56644 4900 56700 4956
rect 66836 4900 66892 4956
rect 69748 4900 69804 4956
rect 70084 4900 70140 4956
rect 71204 4900 71260 4956
rect 74788 4900 74844 4956
rect 76804 4900 76860 4956
rect 80388 4900 80444 4956
rect 82180 4900 82236 4956
rect 83972 4900 84028 4956
rect 84532 4900 84588 4956
rect 85764 4900 85820 4956
rect 91700 4900 91756 4956
rect 97300 4900 97356 4956
rect 113204 4900 113260 4956
rect 116452 4900 116508 4956
rect 118804 4900 118860 4956
rect 119028 4900 119084 4956
rect 121156 4900 121212 4956
rect 133588 4900 133644 4956
rect 133812 4900 133868 4956
rect 135940 4900 135996 4956
rect 139412 4900 139468 4956
rect 151060 4900 151116 4956
rect 154644 4900 154700 4956
rect 161364 4900 161420 4956
rect 162484 4900 162540 4956
rect 179396 4900 179452 4956
rect 190036 4900 190092 4956
rect 191940 4900 191996 4956
rect 193172 4900 193228 4956
rect 194852 4900 194908 4956
rect 209972 4900 210028 4956
rect 211764 4900 211820 4956
rect 67284 4788 67340 4844
rect 82404 4788 82460 4844
rect 102788 4788 102844 4844
rect 103012 4788 103068 4844
rect 112084 4788 112140 4844
rect 120036 4788 120092 4844
rect 122836 4788 122892 4844
rect 127204 4788 127260 4844
rect 132356 4788 132412 4844
rect 137396 4788 137452 4844
rect 140980 4788 141036 4844
rect 144228 4788 144284 4844
rect 144676 4788 144732 4844
rect 149492 4788 149548 4844
rect 180180 4788 180236 4844
rect 180404 4788 180460 4844
rect 182196 4788 182252 4844
rect 44772 4676 44828 4732
rect 55540 4676 55596 4732
rect 55644 4676 55700 4732
rect 55748 4676 55804 4732
rect 72212 4676 72268 4732
rect 83076 4676 83132 4732
rect 84980 4676 85036 4732
rect 90804 4676 90860 4732
rect 98644 4676 98700 4732
rect 99204 4676 99260 4732
rect 107492 4676 107548 4732
rect 107716 4676 107772 4732
rect 109868 4676 109924 4732
rect 109972 4676 110028 4732
rect 110076 4676 110132 4732
rect 119588 4676 119644 4732
rect 126980 4676 127036 4732
rect 146692 4676 146748 4732
rect 152292 4676 152348 4732
rect 152628 4676 152684 4732
rect 153524 4676 153580 4732
rect 153748 4676 153804 4732
rect 164196 4676 164252 4732
rect 164300 4676 164356 4732
rect 164404 4676 164460 4732
rect 165172 4676 165228 4732
rect 56196 4564 56252 4620
rect 66836 4564 66892 4620
rect 74340 4564 74396 4620
rect 79716 4564 79772 4620
rect 80500 4564 80556 4620
rect 85876 4564 85932 4620
rect 87444 4564 87500 4620
rect 92708 4564 92764 4620
rect 97188 4564 97244 4620
rect 97412 4564 97468 4620
rect 102116 4564 102172 4620
rect 108724 4564 108780 4620
rect 114772 4564 114828 4620
rect 115556 4564 115612 4620
rect 116340 4564 116396 4620
rect 124292 4564 124348 4620
rect 132132 4564 132188 4620
rect 135828 4564 135884 4620
rect 139188 4564 139244 4620
rect 149604 4564 149660 4620
rect 161364 4564 161420 4620
rect 197876 4676 197932 4732
rect 198436 4676 198492 4732
rect 189252 4564 189308 4620
rect 189588 4564 189644 4620
rect 189924 4564 189980 4620
rect 192164 4564 192220 4620
rect 67956 4452 68012 4508
rect 89572 4452 89628 4508
rect 118132 4452 118188 4508
rect 118356 4452 118412 4508
rect 131012 4452 131068 4508
rect 133476 4452 133532 4508
rect 134372 4452 134428 4508
rect 144340 4452 144396 4508
rect 149492 4452 149548 4508
rect 154868 4452 154924 4508
rect 164724 4452 164780 4508
rect 167860 4452 167916 4508
rect 55300 4340 55356 4396
rect 72548 4340 72604 4396
rect 72772 4340 72828 4396
rect 76692 4340 76748 4396
rect 78484 4340 78540 4396
rect 79828 4340 79884 4396
rect 80052 4340 80108 4396
rect 84308 4340 84364 4396
rect 84644 4340 84700 4396
rect 87668 4340 87724 4396
rect 87892 4340 87948 4396
rect 88900 4340 88956 4396
rect 89124 4340 89180 4396
rect 100548 4340 100604 4396
rect 101220 4340 101276 4396
rect 110740 4340 110796 4396
rect 115668 4340 115724 4396
rect 120372 4340 120428 4396
rect 120596 4340 120652 4396
rect 125412 4340 125468 4396
rect 156548 4340 156604 4396
rect 162820 4340 162876 4396
rect 180404 4340 180460 4396
rect 39396 4228 39452 4284
rect 54964 4228 55020 4284
rect 71428 4228 71484 4284
rect 74228 4228 74284 4284
rect 76132 4228 76188 4284
rect 80724 4228 80780 4284
rect 81620 4228 81676 4284
rect 82964 4228 83020 4284
rect 85540 4228 85596 4284
rect 96740 4228 96796 4284
rect 97188 4228 97244 4284
rect 102340 4228 102396 4284
rect 102564 4228 102620 4284
rect 111524 4228 111580 4284
rect 113092 4228 113148 4284
rect 119364 4228 119420 4284
rect 119588 4228 119644 4284
rect 147700 4228 147756 4284
rect 151060 4228 151116 4284
rect 159460 4228 159516 4284
rect 178276 4228 178332 4284
rect 191492 4228 191548 4284
rect 10052 4116 10108 4172
rect 62580 4116 62636 4172
rect 69188 4116 69244 4172
rect 78036 4116 78092 4172
rect 78260 4116 78316 4172
rect 79716 4116 79772 4172
rect 81508 4116 81564 4172
rect 81844 4116 81900 4172
rect 95732 4116 95788 4172
rect 115444 4116 115500 4172
rect 119924 4116 119980 4172
rect 121268 4116 121324 4172
rect 124180 4116 124236 4172
rect 124404 4116 124460 4172
rect 131012 4116 131068 4172
rect 139412 4116 139468 4172
rect 140644 4116 140700 4172
rect 156548 4116 156604 4172
rect 56980 4004 57036 4060
rect 66276 4004 66332 4060
rect 68292 4004 68348 4060
rect 73108 4004 73164 4060
rect 77364 4004 77420 4060
rect 77812 4004 77868 4060
rect 86660 4004 86716 4060
rect 88900 4004 88956 4060
rect 96964 4004 97020 4060
rect 97412 4004 97468 4060
rect 97636 4004 97692 4060
rect 109172 4004 109228 4060
rect 110292 4004 110348 4060
rect 112756 4004 112812 4060
rect 112980 4004 113036 4060
rect 120148 4004 120204 4060
rect 126980 4004 127036 4060
rect 132244 4004 132300 4060
rect 134596 4004 134652 4060
rect 144228 4004 144284 4060
rect 157444 4004 157500 4060
rect 191492 4004 191548 4060
rect 192052 4004 192108 4060
rect 192276 4004 192332 4060
rect 50372 3892 50428 3948
rect 61684 3892 61740 3948
rect 62580 3892 62636 3948
rect 65268 3892 65324 3948
rect 65492 3892 65548 3948
rect 77140 3892 77196 3948
rect 77700 3892 77756 3948
rect 77924 3892 77980 3948
rect 79156 3892 79212 3948
rect 100660 3892 100716 3948
rect 103460 3892 103516 3948
rect 103796 3892 103852 3948
rect 105028 3892 105084 3948
rect 115780 3892 115836 3948
rect 134260 3892 134316 3948
rect 141204 3892 141260 3948
rect 147364 3892 147420 3948
rect 152852 3892 152908 3948
rect 157556 3892 157612 3948
rect 162820 3892 162876 3948
rect 180180 3892 180236 3948
rect 191716 3892 191772 3948
rect 53844 3780 53900 3836
rect 55300 3780 55356 3836
rect 66724 3780 66780 3836
rect 67060 3780 67116 3836
rect 67284 3780 67340 3836
rect 70532 3780 70588 3836
rect 70756 3780 70812 3836
rect 75348 3780 75404 3836
rect 79044 3780 79100 3836
rect 79380 3780 79436 3836
rect 84420 3780 84476 3836
rect 84644 3780 84700 3836
rect 85428 3780 85484 3836
rect 88340 3780 88396 3836
rect 89348 3780 89404 3836
rect 89572 3780 89628 3836
rect 108948 3780 109004 3836
rect 109172 3780 109228 3836
rect 114996 3780 115052 3836
rect 115220 3780 115276 3836
rect 116116 3780 116172 3836
rect 116340 3780 116396 3836
rect 119252 3780 119308 3836
rect 119700 3780 119756 3836
rect 125860 3780 125916 3836
rect 132020 3780 132076 3836
rect 132692 3780 132748 3836
rect 142772 3780 142828 3836
rect 144452 3780 144508 3836
rect 152964 3780 153020 3836
rect 153188 3780 153244 3836
rect 155092 3780 155148 3836
rect 156212 3780 156268 3836
rect 194964 3780 195020 3836
rect 209636 3780 209692 3836
rect 63700 3668 63756 3724
rect 72996 3668 73052 3724
rect 81172 3668 81228 3724
rect 82740 3668 82796 3724
rect 83412 3668 83468 3724
rect 97748 3668 97804 3724
rect 99764 3668 99820 3724
rect 101444 3668 101500 3724
rect 101668 3668 101724 3724
rect 110628 3668 110684 3724
rect 110852 3668 110908 3724
rect 123284 3668 123340 3724
rect 137396 3668 137452 3724
rect 142212 3668 142268 3724
rect 144228 3668 144284 3724
rect 146132 3668 146188 3724
rect 146692 3668 146748 3724
rect 50372 3556 50428 3612
rect 50596 3556 50652 3612
rect 61684 3556 61740 3612
rect 151060 3668 151116 3724
rect 154308 3668 154364 3724
rect 162820 3668 162876 3724
rect 163044 3668 163100 3724
rect 65380 3556 65436 3612
rect 68628 3556 68684 3612
rect 70084 3556 70140 3612
rect 73220 3556 73276 3612
rect 74788 3556 74844 3612
rect 79156 3556 79212 3612
rect 79380 3556 79436 3612
rect 81956 3556 82012 3612
rect 82852 3556 82908 3612
rect 84084 3556 84140 3612
rect 84308 3556 84364 3612
rect 95620 3556 95676 3612
rect 96068 3556 96124 3612
rect 98084 3556 98140 3612
rect 99092 3556 99148 3612
rect 102116 3556 102172 3612
rect 102676 3556 102732 3612
rect 103460 3556 103516 3612
rect 113652 3556 113708 3612
rect 120708 3556 120764 3612
rect 122388 3556 122444 3612
rect 122948 3556 123004 3612
rect 55300 3444 55356 3500
rect 61908 3444 61964 3500
rect 73108 3444 73164 3500
rect 76692 3444 76748 3500
rect 77252 3444 77308 3500
rect 77812 3444 77868 3500
rect 78932 3444 78988 3500
rect 80612 3444 80668 3500
rect 81732 3444 81788 3500
rect 82068 3444 82124 3500
rect 83524 3444 83580 3500
rect 83748 3444 83804 3500
rect 89012 3444 89068 3500
rect 89236 3444 89292 3500
rect 91588 3444 91644 3500
rect 92484 3444 92540 3500
rect 102564 3444 102620 3500
rect 112980 3444 113036 3500
rect 113204 3444 113260 3500
rect 114772 3444 114828 3500
rect 115220 3444 115276 3500
rect 115668 3444 115724 3500
rect 120148 3444 120204 3500
rect 55300 3220 55356 3276
rect 58772 3220 58828 3276
rect 137844 3556 137900 3612
rect 138628 3556 138684 3612
rect 142772 3556 142828 3612
rect 120596 3444 120652 3500
rect 127428 3444 127484 3500
rect 74900 3332 74956 3388
rect 76804 3332 76860 3388
rect 84420 3332 84476 3388
rect 88900 3332 88956 3388
rect 101332 3332 101388 3388
rect 104468 3332 104524 3388
rect 110404 3332 110460 3388
rect 112756 3332 112812 3388
rect 113540 3332 113596 3388
rect 113764 3332 113820 3388
rect 114324 3332 114380 3388
rect 115108 3332 115164 3388
rect 118020 3332 118076 3388
rect 118244 3332 118300 3388
rect 119140 3332 119196 3388
rect 121604 3332 121660 3388
rect 63700 3220 63756 3276
rect 67172 3220 67228 3276
rect 67396 3220 67452 3276
rect 69972 3220 70028 3276
rect 74340 3220 74396 3276
rect 74564 3220 74620 3276
rect 75572 3220 75628 3276
rect 77476 3220 77532 3276
rect 77700 3220 77756 3276
rect 78260 3220 78316 3276
rect 81508 3220 81564 3276
rect 82964 3220 83020 3276
rect 83972 3220 84028 3276
rect 100212 3220 100268 3276
rect 102676 3220 102732 3276
rect 105700 3220 105756 3276
rect 107380 3220 107436 3276
rect 109284 3220 109340 3276
rect 112868 3220 112924 3276
rect 121156 3220 121212 3276
rect 132580 3220 132636 3276
rect 140980 3444 141036 3500
rect 150948 3444 151004 3500
rect 140868 3332 140924 3388
rect 147700 3332 147756 3388
rect 159684 3332 159740 3388
rect 167076 3332 167132 3388
rect 168644 3332 168700 3388
rect 190148 3332 190204 3388
rect 144228 3220 144284 3276
rect 156212 3220 156268 3276
rect 166404 3220 166460 3276
rect 179620 3220 179676 3276
rect 184660 3220 184716 3276
rect 187348 3220 187404 3276
rect 187796 3220 187852 3276
rect 52724 3108 52780 3164
rect 60004 3108 60060 3164
rect 63924 3108 63980 3164
rect 66276 3108 66332 3164
rect 100660 3108 100716 3164
rect 101220 3108 101276 3164
rect 102452 3108 102508 3164
rect 102900 3108 102956 3164
rect 112308 3108 112364 3164
rect 113652 3108 113708 3164
rect 117348 3108 117404 3164
rect 131460 3108 131516 3164
rect 146244 3108 146300 3164
rect 147700 3108 147756 3164
rect 154756 3108 154812 3164
rect 161140 3108 161196 3164
rect 161364 3108 161420 3164
rect 162260 3108 162316 3164
rect 162484 3108 162540 3164
rect 168756 3108 168812 3164
rect 185220 3108 185276 3164
rect 57092 2996 57148 3052
rect 57428 2996 57484 3052
rect 64148 2996 64204 3052
rect 64708 2996 64764 3052
rect 66948 2996 67004 3052
rect 70756 2996 70812 3052
rect 71652 2996 71708 3052
rect 80164 2996 80220 3052
rect 82516 2996 82572 3052
rect 83188 2996 83244 3052
rect 85428 2996 85484 3052
rect 86212 2996 86268 3052
rect 86436 2996 86492 3052
rect 89684 2996 89740 3052
rect 100996 2996 101052 3052
rect 102340 2996 102396 3052
rect 109620 2996 109676 3052
rect 110404 2996 110460 3052
rect 110740 2996 110796 3052
rect 110964 2996 111020 3052
rect 112196 2996 112252 3052
rect 114324 2996 114380 3052
rect 114772 2996 114828 3052
rect 114996 2996 115052 3052
rect 119028 2996 119084 3052
rect 125636 2996 125692 3052
rect 127092 2996 127148 3052
rect 132468 2996 132524 3052
rect 174132 2996 174188 3052
rect 181860 2996 181916 3052
rect 184436 2996 184492 3052
rect 52948 2884 53004 2940
rect 55300 2884 55356 2940
rect 83860 2884 83916 2940
rect 84084 2884 84140 2940
rect 87668 2884 87724 2940
rect 88788 2884 88844 2940
rect 89012 2884 89068 2940
rect 104132 2884 104188 2940
rect 104356 2884 104412 2940
rect 108724 2884 108780 2940
rect 121044 2884 121100 2940
rect 135828 2884 135884 2940
rect 146020 2884 146076 2940
rect 183092 2884 183148 2940
rect 185892 2884 185948 2940
rect 188916 2884 188972 2940
rect 194068 2884 194124 2940
rect 45892 2772 45948 2828
rect 67060 2772 67116 2828
rect 82852 2772 82908 2828
rect 83188 2772 83244 2828
rect 83636 2772 83692 2828
rect 88900 2772 88956 2828
rect 102228 2772 102284 2828
rect 109620 2772 109676 2828
rect 114436 2772 114492 2828
rect 115332 2772 115388 2828
rect 119476 2772 119532 2828
rect 121828 2772 121884 2828
rect 133028 2772 133084 2828
rect 134260 2772 134316 2828
rect 142548 2772 142604 2828
rect 162484 2772 162540 2828
rect 162708 2772 162764 2828
rect 166292 2772 166348 2828
rect 190596 2772 190652 2828
rect 57316 2660 57372 2716
rect 70084 2660 70140 2716
rect 73332 2660 73388 2716
rect 87668 2660 87724 2716
rect 92372 2660 92428 2716
rect 92596 2660 92652 2716
rect 97524 2660 97580 2716
rect 100436 2660 100492 2716
rect 101444 2660 101500 2716
rect 104356 2660 104412 2716
rect 106596 2660 106652 2716
rect 132692 2660 132748 2716
rect 138516 2660 138572 2716
rect 146020 2660 146076 2716
rect 156211 2660 156267 2716
rect 174132 2660 174188 2716
rect 174356 2660 174412 2716
rect 67172 2548 67228 2604
rect 74340 2548 74396 2604
rect 75684 2548 75740 2604
rect 77924 2548 77980 2604
rect 78820 2548 78876 2604
rect 84644 2548 84700 2604
rect 99316 2548 99372 2604
rect 99988 2548 100044 2604
rect 100772 2548 100828 2604
rect 103348 2548 103404 2604
rect 108388 2548 108444 2604
rect 117908 2548 117964 2604
rect 121156 2548 121212 2604
rect 123060 2548 123116 2604
rect 137732 2548 137788 2604
rect 148260 2548 148316 2604
rect 197540 2548 197596 2604
rect 54964 2436 55020 2492
rect 59892 2436 59948 2492
rect 61572 2436 61628 2492
rect 65380 2436 65436 2492
rect 67620 2436 67676 2492
rect 71316 2436 71372 2492
rect 71540 2436 71596 2492
rect 72660 2436 72716 2492
rect 86884 2436 86940 2492
rect 90580 2436 90636 2492
rect 96292 2436 96348 2492
rect 99764 2436 99820 2492
rect 101668 2436 101724 2492
rect 106596 2436 106652 2492
rect 111972 2436 112028 2492
rect 112196 2436 112252 2492
rect 125636 2436 125692 2492
rect 145684 2436 145740 2492
rect 147588 2436 147644 2492
rect 149492 2436 149548 2492
rect 154420 2436 154476 2492
rect 155876 2436 155932 2492
rect 179060 2436 179116 2492
rect 179284 2436 179340 2492
rect 183092 2436 183148 2492
rect 189252 2436 189308 2492
rect 201572 2436 201628 2492
rect 52948 2324 53004 2380
rect 53172 2324 53228 2380
rect 56980 2324 57036 2380
rect 80836 2324 80892 2380
rect 81396 2324 81452 2380
rect 82068 2324 82124 2380
rect 82292 2324 82348 2380
rect 92596 2324 92652 2380
rect 103348 2324 103404 2380
rect 109171 2324 109227 2380
rect 115556 2324 115612 2380
rect 117236 2324 117292 2380
rect 118580 2324 118636 2380
rect 120596 2324 120652 2380
rect 122052 2324 122108 2380
rect 122612 2324 122668 2380
rect 134260 2324 134316 2380
rect 134596 2324 134652 2380
rect 136388 2324 136444 2380
rect 137732 2324 137788 2380
rect 150612 2324 150668 2380
rect 157780 2324 157836 2380
rect 161251 2324 161307 2380
rect 173124 2324 173180 2380
rect 174916 2324 174972 2380
rect 53508 2212 53564 2268
rect 62131 2212 62187 2268
rect 67620 2212 67676 2268
rect 75572 2212 75628 2268
rect 83636 2212 83692 2268
rect 85764 2212 85820 2268
rect 87220 2212 87276 2268
rect 87444 2212 87500 2268
rect 93940 2212 93996 2268
rect 95620 2212 95676 2268
rect 98196 2212 98252 2268
rect 101556 2212 101612 2268
rect 102900 2212 102956 2268
rect 104244 2212 104300 2268
rect 104468 2212 104524 2268
rect 113204 2212 113260 2268
rect 114100 2212 114156 2268
rect 122500 2212 122556 2268
rect 123844 2212 123900 2268
rect 132804 2212 132860 2268
rect 134148 2212 134204 2268
rect 134484 2212 134540 2268
rect 140084 2212 140140 2268
rect 151172 2212 151228 2268
rect 153860 2212 153916 2268
rect 203588 2212 203644 2268
rect 45892 2100 45948 2156
rect 64708 2100 64764 2156
rect 72100 2100 72156 2156
rect 73220 2100 73276 2156
rect 75236 2100 75292 2156
rect 77700 2100 77756 2156
rect 77924 2100 77980 2156
rect 83076 2100 83132 2156
rect 83412 2100 83468 2156
rect 85204 2100 85260 2156
rect 86324 2100 86380 2156
rect 90244 2100 90300 2156
rect 91140 2100 91196 2156
rect 91924 2100 91980 2156
rect 94388 2100 94444 2156
rect 96292 2100 96348 2156
rect 96516 2100 96572 2156
rect 113316 2100 113372 2156
rect 117572 2100 117628 2156
rect 133252 2100 133308 2156
rect 137732 2100 137788 2156
rect 161028 2100 161084 2156
rect 179284 2100 179340 2156
rect 188692 2100 188748 2156
rect 188916 2100 188972 2156
rect 56980 1988 57036 2044
rect 60788 1988 60844 2044
rect 71652 1988 71708 2044
rect 75460 1988 75516 2044
rect 75684 1988 75740 2044
rect 81396 1988 81452 2044
rect 94276 1988 94332 2044
rect 94500 1988 94556 2044
rect 101332 1988 101388 2044
rect 101556 1988 101612 2044
rect 109732 1988 109788 2044
rect 113652 1988 113708 2044
rect 113876 1988 113932 2044
rect 114772 1988 114828 2044
rect 125860 1988 125916 2044
rect 147924 1988 147980 2044
rect 150052 1988 150108 2044
rect 150724 1988 150780 2044
rect 151060 1988 151116 2044
rect 168084 1988 168140 2044
rect 52724 1876 52780 1932
rect 62468 1876 62524 1932
rect 62804 1876 62860 1932
rect 74564 1876 74620 1932
rect 80724 1876 80780 1932
rect 85540 1876 85596 1932
rect 85764 1876 85820 1932
rect 89684 1876 89740 1932
rect 115444 1876 115500 1932
rect 119364 1876 119420 1932
rect 136164 1876 136220 1932
rect 147364 1876 147420 1932
rect 150836 1876 150892 1932
rect 151508 1876 151564 1932
rect 151732 1876 151788 1932
rect 154420 1876 154476 1932
rect 155988 1876 156044 1932
rect 159572 1876 159628 1932
rect 164724 1876 164780 1932
rect 164948 1876 165004 1932
rect 167972 1876 168028 1932
rect 189924 1876 189980 1932
rect 65380 1764 65436 1820
rect 72996 1764 73052 1820
rect 88676 1764 88732 1820
rect 89236 1764 89292 1820
rect 94052 1764 94108 1820
rect 99652 1764 99708 1820
rect 102788 1764 102844 1820
rect 114772 1764 114828 1820
rect 121268 1764 121324 1820
rect 129332 1764 129388 1820
rect 154644 1764 154700 1820
rect 157780 1764 157836 1820
rect 162820 1764 162876 1820
rect 188692 1764 188748 1820
rect 191716 1764 191772 1820
rect 75236 1652 75292 1708
rect 75460 1652 75516 1708
rect 79716 1652 79772 1708
rect 80052 1652 80108 1708
rect 81396 1652 81452 1708
rect 99764 1652 99820 1708
rect 114996 1652 115052 1708
rect 120932 1652 120988 1708
rect 127204 1652 127260 1708
rect 132020 1652 132076 1708
rect 132804 1652 132860 1708
rect 133028 1652 133084 1708
rect 133700 1652 133756 1708
rect 138516 1652 138572 1708
rect 147924 1652 147980 1708
rect 150276 1652 150332 1708
rect 150724 1652 150780 1708
rect 17780 1540 17836 1596
rect 22708 1540 22764 1596
rect 28756 1540 28812 1596
rect 29988 1540 30044 1596
rect 34244 1540 34300 1596
rect 35476 1540 35532 1596
rect 44772 1540 44828 1596
rect 62131 1540 62187 1596
rect 65940 1540 65996 1596
rect 71540 1540 71596 1596
rect 71764 1540 71820 1596
rect 90356 1540 90412 1596
rect 90580 1540 90636 1596
rect 102452 1540 102508 1596
rect 104020 1540 104076 1596
rect 108836 1540 108892 1596
rect 110292 1540 110348 1596
rect 111524 1540 111580 1596
rect 115892 1540 115948 1596
rect 116116 1540 116172 1596
rect 116564 1540 116620 1596
rect 118020 1540 118076 1596
rect 118468 1540 118524 1596
rect 120484 1540 120540 1596
rect 124628 1540 124684 1596
rect 135716 1540 135772 1596
rect 142436 1540 142492 1596
rect 143444 1540 143500 1596
rect 144004 1540 144060 1596
rect 144452 1540 144508 1596
rect 145012 1540 145068 1596
rect 145236 1540 145292 1596
rect 146132 1540 146188 1596
rect 154308 1540 154364 1596
rect 159684 1540 159740 1596
rect 162708 1540 162764 1596
rect 163156 1540 163212 1596
rect 164836 1540 164892 1596
rect 166516 1540 166572 1596
rect 175140 1540 175196 1596
rect 179396 1540 179452 1596
rect 180404 1540 180460 1596
rect 186116 1540 186172 1596
rect 187908 1540 187964 1596
rect 189140 1540 189196 1596
rect 196420 1540 196476 1596
rect 199444 1540 199500 1596
rect 200116 1540 200172 1596
rect 204372 1540 204428 1596
rect 211652 1540 211708 1596
rect 25172 1428 25228 1484
rect 49700 1428 49756 1484
rect 59780 1428 59836 1484
rect 60340 1428 60396 1484
rect 71988 1428 72044 1484
rect 74900 1428 74956 1484
rect 76244 1428 76300 1484
rect 77252 1428 77308 1484
rect 77476 1428 77532 1484
rect 79492 1428 79548 1484
rect 79716 1428 79772 1484
rect 86996 1428 87052 1484
rect 87220 1428 87276 1484
rect 88004 1428 88060 1484
rect 88676 1428 88732 1484
rect 121044 1428 121100 1484
rect 121604 1428 121660 1484
rect 122500 1428 122556 1484
rect 129332 1428 129388 1484
rect 135604 1428 135660 1484
rect 138628 1428 138684 1484
rect 141652 1428 141708 1484
rect 144340 1428 144396 1484
rect 144676 1428 144732 1484
rect 147924 1428 147980 1484
rect 152180 1428 152236 1484
rect 152852 1428 152908 1484
rect 164500 1428 164556 1484
rect 164724 1428 164780 1484
rect 180628 1428 180684 1484
rect 190596 1428 190652 1484
rect 25620 1316 25676 1372
rect 53620 1316 53676 1372
rect 62580 1316 62636 1372
rect 66836 1316 66892 1372
rect 67060 1316 67116 1372
rect 72100 1316 72156 1372
rect 33684 1204 33740 1260
rect 35588 1204 35644 1260
rect 44436 1204 44492 1260
rect 50596 1204 50652 1260
rect 77028 1316 77084 1372
rect 78932 1316 78988 1372
rect 79940 1316 79996 1372
rect 82852 1316 82908 1372
rect 87556 1316 87612 1372
rect 99204 1316 99260 1372
rect 99428 1316 99484 1372
rect 101220 1316 101276 1372
rect 109060 1316 109116 1372
rect 120260 1316 120316 1372
rect 120708 1316 120764 1372
rect 123284 1316 123340 1372
rect 123508 1316 123564 1372
rect 135044 1316 135100 1372
rect 139412 1316 139468 1372
rect 156100 1316 156156 1372
rect 166180 1316 166236 1372
rect 211092 1316 211148 1372
rect 214452 1316 214508 1372
rect 59220 1204 59276 1260
rect 60452 1204 60508 1260
rect 61908 1204 61964 1260
rect 62132 1204 62188 1260
rect 68068 1204 68124 1260
rect 72548 1204 72604 1260
rect 86996 1204 87052 1260
rect 88564 1204 88620 1260
rect 90356 1204 90412 1260
rect 106036 1204 106092 1260
rect 108836 1204 108892 1260
rect 109396 1204 109452 1260
rect 113988 1204 114044 1260
rect 114212 1204 114268 1260
rect 117012 1204 117068 1260
rect 117572 1204 117628 1260
rect 125972 1204 126028 1260
rect 132692 1204 132748 1260
rect 135828 1204 135884 1260
rect 138068 1204 138124 1260
rect 144004 1204 144060 1260
rect 150164 1204 150220 1260
rect 150388 1204 150444 1260
rect 152740 1204 152796 1260
rect 208292 1204 208348 1260
rect 10164 1092 10220 1148
rect 30660 1092 30716 1148
rect 50148 1092 50204 1148
rect 50372 1092 50428 1148
rect 54068 1092 54124 1148
rect 70532 1092 70588 1148
rect 70756 1092 70812 1148
rect 74116 1092 74172 1148
rect 87220 1092 87276 1148
rect 90580 1092 90636 1148
rect 91028 1092 91084 1148
rect 94052 1092 94108 1148
rect 103236 1092 103292 1148
rect 109620 1092 109676 1148
rect 109844 1092 109900 1148
rect 110964 1092 111020 1148
rect 125860 1092 125916 1148
rect 126196 1092 126252 1148
rect 127428 1092 127484 1148
rect 140308 1092 140364 1148
rect 142884 1092 142940 1148
rect 168644 1092 168700 1148
rect 190596 1092 190652 1148
rect 192836 1092 192892 1148
rect 18452 980 18508 1036
rect 19236 980 19292 1036
rect 39396 980 39452 1036
rect 65380 980 65436 1036
rect 80948 980 81004 1036
rect 84756 980 84812 1036
rect 85764 980 85820 1036
rect 87108 980 87164 1036
rect 87332 980 87388 1036
rect 97524 980 97580 1036
rect 97748 980 97804 1036
rect 100436 980 100492 1036
rect 100772 980 100828 1036
rect 103684 980 103740 1036
rect 106148 980 106204 1036
rect 106372 980 106428 1036
rect 108164 980 108220 1036
rect 110068 980 110124 1036
rect 110292 980 110348 1036
rect 116116 980 116172 1036
rect 119252 980 119308 1036
rect 119924 980 119980 1036
rect 144676 980 144732 1036
rect 147700 980 147756 1036
rect 147924 980 147980 1036
rect 152852 980 152908 1036
rect 153748 980 153804 1036
rect 153972 980 154028 1036
rect 194068 980 194124 1036
rect 195188 980 195244 1036
rect 197092 980 197148 1036
rect 1316 868 1372 924
rect 1988 868 2044 924
rect 2548 868 2604 924
rect 15988 868 16044 924
rect 19684 868 19740 924
rect 40404 868 40460 924
rect 40964 868 41020 924
rect 75236 868 75292 924
rect 75460 868 75516 924
rect 76020 868 76076 924
rect 76244 868 76300 924
rect 80388 868 80444 924
rect 81508 868 81564 924
rect 81844 868 81900 924
rect 82180 868 82236 924
rect 82852 868 82908 924
rect 83076 868 83132 924
rect 123844 868 123900 924
rect 125860 868 125916 924
rect 19348 756 19404 812
rect 44436 756 44492 812
rect 44660 756 44716 812
rect 50372 756 50428 812
rect 50596 756 50652 812
rect 138516 868 138572 924
rect 144452 868 144508 924
rect 151172 868 151228 924
rect 151956 868 152012 924
rect 162820 868 162876 924
rect 171444 868 171500 924
rect 50484 644 50540 700
rect 52052 644 52108 700
rect 57092 644 57148 700
rect 72548 756 72604 812
rect 74116 756 74172 812
rect 81060 756 81116 812
rect 81956 756 82012 812
rect 82292 756 82348 812
rect 107492 756 107548 812
rect 108052 756 108108 812
rect 112308 756 112364 812
rect 197540 1092 197596 1148
rect 216356 1092 216412 1148
rect 197652 980 197708 1036
rect 203028 868 203084 924
rect 205604 868 205660 924
rect 206836 868 206892 924
rect 212884 868 212940 924
rect 217140 868 217196 924
rect 52164 532 52220 588
rect 76244 644 76300 700
rect 76804 644 76860 700
rect 77140 644 77196 700
rect 79268 644 79324 700
rect 80388 644 80444 700
rect 80724 644 80780 700
rect 107940 644 107996 700
rect 117572 644 117628 700
rect 118916 644 118972 700
rect 119140 644 119196 700
rect 134596 644 134652 700
rect 141316 644 141372 700
rect 144452 644 144508 700
rect 144676 644 144732 700
rect 145012 644 145068 700
rect 194068 644 194124 700
rect 56980 532 57036 588
rect 124180 532 124236 588
rect 144900 532 144956 588
rect 150388 532 150444 588
rect 151060 532 151116 588
rect 13972 420 14028 476
rect 49924 420 49980 476
rect 57428 420 57484 476
rect 59780 420 59836 476
rect 72324 420 72380 476
rect 72548 420 72604 476
rect 76580 420 76636 476
rect 77252 420 77308 476
rect 80052 420 80108 476
rect 80276 420 80332 476
rect 81620 420 81676 476
rect 91700 420 91756 476
rect 97300 420 97356 476
rect 97412 420 97468 476
rect 100548 420 100604 476
rect 100772 420 100828 476
rect 102004 420 102060 476
rect 102228 420 102284 476
rect 109844 420 109900 476
rect 110068 420 110124 476
rect 116228 420 116284 476
rect 117572 420 117628 476
rect 117796 420 117852 476
rect 120820 420 120876 476
rect 121940 420 121996 476
rect 130788 420 130844 476
rect 131124 420 131180 476
rect 138516 420 138572 476
rect 57764 308 57820 364
rect 76692 308 76748 364
rect 79604 308 79660 364
rect 81060 308 81116 364
rect 83300 308 83356 364
rect 83524 308 83580 364
rect 85988 308 86044 364
rect 86660 308 86716 364
rect 86884 308 86940 364
rect 99204 308 99260 364
rect 103012 308 103068 364
rect 103236 308 103292 364
rect 110852 308 110908 364
rect 111076 308 111132 364
rect 116676 308 116732 364
rect 121044 308 121100 364
rect 127540 308 127596 364
rect 52052 196 52108 252
rect 52276 196 52332 252
rect 60564 196 60620 252
rect 63588 84 63644 140
rect 65940 84 65996 140
<< metal4 >>
rect 60452 14968 60508 14978
rect 49140 14788 49196 14798
rect 21476 14608 21532 14618
rect 17780 14248 17836 14258
rect 14868 14068 14924 14078
rect 14868 13962 14924 13972
rect 17780 14028 17836 14192
rect 21476 14140 21532 14552
rect 21476 14074 21532 14084
rect 17780 13962 17836 13972
rect 25060 13916 25116 13926
rect 25060 13708 25116 13860
rect 25060 13642 25116 13652
rect 43204 13888 43260 13898
rect 10500 13580 10556 13590
rect 10500 13462 10556 13472
rect 25732 13468 25788 13478
rect 25732 13348 25788 13412
rect 25732 13282 25788 13292
rect 18452 13244 18508 13254
rect 18452 13168 18508 13188
rect 18452 13102 18508 13112
rect 27972 13020 28028 13030
rect 27972 12808 28028 12964
rect 34468 13020 34524 13030
rect 34468 12922 34524 12932
rect 27188 12796 27244 12806
rect 27972 12742 28028 12752
rect 27188 12628 27244 12740
rect 27188 12562 27244 12572
rect 30100 12572 30156 12582
rect 30100 12448 30156 12516
rect 30100 12382 30156 12392
rect 42196 12268 42252 12278
rect 26740 11728 26796 11738
rect 22708 11008 22764 11018
rect 10276 10828 10332 10838
rect 10164 9660 10220 9670
rect 10052 9100 10108 9110
rect 9604 4956 9660 4966
rect 9604 3988 9660 4900
rect 10052 4172 10108 9044
rect 10052 4106 10108 4116
rect 9604 3922 9660 3932
rect 2548 1288 2604 1298
rect 1316 1108 1372 1118
rect 1316 924 1372 1052
rect 1316 858 1372 868
rect 1988 924 2044 934
rect 1988 568 2044 868
rect 2548 924 2604 1232
rect 10164 1148 10220 9604
rect 10276 8316 10332 10772
rect 16212 10288 16268 10298
rect 16212 10108 16268 10232
rect 16212 10042 16268 10052
rect 21700 9928 21756 9938
rect 21700 9324 21756 9872
rect 21700 9258 21756 9268
rect 10276 8250 10332 8260
rect 13972 8092 14028 8102
rect 11620 4956 11676 4966
rect 11620 4348 11676 4900
rect 11620 4282 11676 4292
rect 10164 1082 10220 1092
rect 2548 858 2604 868
rect 1988 502 2044 512
rect 13972 476 14028 8036
rect 19348 8092 19404 8102
rect 18228 7420 18284 7430
rect 18116 5740 18172 5750
rect 16436 4956 16492 4966
rect 16436 4168 16492 4900
rect 16436 4102 16492 4112
rect 17780 2908 17836 2918
rect 17780 1596 17836 2852
rect 17780 1530 17836 1540
rect 13972 410 14028 420
rect 15988 924 16044 934
rect 15988 208 16044 868
rect 18116 748 18172 5684
rect 18228 928 18284 7364
rect 19236 5180 19292 5190
rect 18452 2548 18508 2558
rect 18452 1036 18508 2492
rect 18452 970 18508 980
rect 19236 1036 19292 5124
rect 19236 970 19292 980
rect 18228 862 18284 872
rect 19348 812 19404 8036
rect 21140 5068 21196 5078
rect 21140 1108 21196 5012
rect 22708 1596 22764 10952
rect 26740 10108 26796 11672
rect 29988 10648 30044 10658
rect 28756 10332 28812 10342
rect 26740 10042 26796 10052
rect 28348 10220 28668 10252
rect 28348 10164 28376 10220
rect 28432 10164 28480 10220
rect 28536 10164 28584 10220
rect 28640 10164 28668 10220
rect 28348 9729 28668 10164
rect 28348 9673 28376 9729
rect 28432 9673 28480 9729
rect 28536 9673 28584 9729
rect 28640 9673 28668 9729
rect 28348 9625 28668 9673
rect 28348 9569 28376 9625
rect 28432 9569 28480 9625
rect 28536 9569 28584 9625
rect 28640 9569 28668 9625
rect 28348 9521 28668 9569
rect 28348 9465 28376 9521
rect 28432 9465 28480 9521
rect 28536 9465 28584 9521
rect 28640 9465 28668 9521
rect 26404 8988 26460 8998
rect 25956 7980 26012 7990
rect 25620 7196 25676 7206
rect 22708 1530 22764 1540
rect 23044 5180 23100 5190
rect 23044 1288 23100 5124
rect 23044 1222 23100 1232
rect 23380 5068 23436 5078
rect 21140 1042 21196 1052
rect 19348 746 19404 756
rect 19684 924 19740 934
rect 18116 682 18172 692
rect 19684 388 19740 868
rect 23380 568 23436 5012
rect 25172 2728 25228 2738
rect 25172 1484 25228 2672
rect 25172 1418 25228 1428
rect 25620 1372 25676 7140
rect 25620 1306 25676 1316
rect 23380 502 23436 512
rect 25956 568 26012 7924
rect 26404 1108 26460 8932
rect 28348 8652 28668 9465
rect 28348 8596 28376 8652
rect 28432 8596 28480 8652
rect 28536 8596 28584 8652
rect 28640 8596 28668 8652
rect 28348 8331 28668 8596
rect 28348 8275 28376 8331
rect 28432 8275 28480 8331
rect 28536 8275 28584 8331
rect 28640 8275 28668 8331
rect 28348 8227 28668 8275
rect 28348 8171 28376 8227
rect 28432 8171 28480 8227
rect 28536 8171 28584 8227
rect 28640 8171 28668 8227
rect 28348 8123 28668 8171
rect 28348 8067 28376 8123
rect 28432 8067 28480 8123
rect 28536 8067 28584 8123
rect 28640 8067 28668 8123
rect 28348 7084 28668 8067
rect 28348 7028 28376 7084
rect 28432 7028 28480 7084
rect 28536 7028 28584 7084
rect 28640 7028 28668 7084
rect 28348 6933 28668 7028
rect 28348 6877 28376 6933
rect 28432 6877 28480 6933
rect 28536 6877 28584 6933
rect 28640 6877 28668 6933
rect 28348 6829 28668 6877
rect 28348 6773 28376 6829
rect 28432 6773 28480 6829
rect 28536 6773 28584 6829
rect 28640 6773 28668 6829
rect 28348 6725 28668 6773
rect 28348 6669 28376 6725
rect 28432 6669 28480 6725
rect 28536 6669 28584 6725
rect 28640 6669 28668 6725
rect 28348 5535 28668 6669
rect 28756 6636 28812 10276
rect 28756 6570 28812 6580
rect 28348 5460 28376 5535
rect 28432 5460 28480 5535
rect 28536 5460 28584 5535
rect 28640 5460 28668 5535
rect 28348 5431 28668 5460
rect 28348 5375 28376 5431
rect 28432 5375 28480 5431
rect 28536 5375 28584 5431
rect 28640 5375 28668 5431
rect 28348 5327 28668 5375
rect 28348 5271 28376 5327
rect 28432 5271 28480 5327
rect 28536 5271 28584 5327
rect 28640 5271 28668 5327
rect 28348 4644 28668 5271
rect 28756 3088 28812 3098
rect 28756 1596 28812 3032
rect 28756 1530 28812 1540
rect 29988 1596 30044 10592
rect 36820 10468 36876 10478
rect 36820 10108 36876 10412
rect 36820 10042 36876 10052
rect 30100 8540 30156 8550
rect 30100 5964 30156 8484
rect 42196 7644 42252 12212
rect 43204 9660 43260 13832
rect 44548 11368 44604 11378
rect 44436 10332 44492 10342
rect 44436 10108 44492 10276
rect 44436 10042 44492 10052
rect 43204 9594 43260 9604
rect 44548 9324 44604 11312
rect 46228 11188 46284 11198
rect 46116 10108 46172 10118
rect 46116 9660 46172 10052
rect 46116 9594 46172 9604
rect 44548 9258 44604 9268
rect 42196 7578 42252 7588
rect 46228 7644 46284 11132
rect 49140 10332 49196 14732
rect 53844 14428 53900 14438
rect 53844 13708 53900 14372
rect 57092 13888 57148 13898
rect 57092 13804 57148 13832
rect 57092 13738 57148 13748
rect 53844 13642 53900 13652
rect 56644 13708 56700 13718
rect 53844 13468 53900 13478
rect 53844 13348 53900 13412
rect 53844 13282 53900 13292
rect 54068 13348 54124 13358
rect 53060 13244 53116 13254
rect 53060 12808 53116 13188
rect 53060 12742 53116 12752
rect 53396 12808 53452 12818
rect 51716 11564 51772 11574
rect 51716 11340 51772 11508
rect 51716 11274 51772 11284
rect 51940 11340 51996 11350
rect 49140 10266 49196 10276
rect 51940 10108 51996 11284
rect 53396 10332 53452 12752
rect 53396 10266 53452 10276
rect 51940 10042 51996 10052
rect 47348 9100 47404 9110
rect 47348 8092 47404 9044
rect 52276 8988 52332 8998
rect 47348 8026 47404 8036
rect 48580 8092 48636 8102
rect 46228 7578 46284 7588
rect 30100 5898 30156 5908
rect 30660 7196 30716 7206
rect 29988 1530 30044 1540
rect 30660 1148 30716 7140
rect 34580 7196 34636 7206
rect 33908 5740 33964 5750
rect 33908 5516 33964 5684
rect 33908 3268 33964 5460
rect 33908 3202 33964 3212
rect 34244 3448 34300 3458
rect 33684 2188 33740 2198
rect 33684 1260 33740 2132
rect 34244 1596 34300 3392
rect 34244 1530 34300 1540
rect 34580 1468 34636 7140
rect 44660 7196 44716 7206
rect 37716 6524 37772 6534
rect 35588 6076 35644 6086
rect 35476 3628 35532 3638
rect 35476 1596 35532 3572
rect 35476 1530 35532 1540
rect 34580 1402 34636 1412
rect 33684 1194 33740 1204
rect 35588 1260 35644 6020
rect 37716 5740 37772 6468
rect 37716 5674 37772 5684
rect 41748 5852 41804 5862
rect 41748 5628 41804 5796
rect 41748 5562 41804 5572
rect 42420 5852 42476 5862
rect 35700 4956 35756 4966
rect 35700 4708 35756 4900
rect 35700 4642 35756 4652
rect 35588 1194 35644 1204
rect 39396 4284 39452 4294
rect 30660 1082 30716 1092
rect 26404 1042 26460 1052
rect 39396 1036 39452 4228
rect 42420 1288 42476 5796
rect 42420 1222 42476 1232
rect 44436 1260 44492 1270
rect 39396 970 39452 980
rect 40404 928 40460 962
rect 40404 858 40460 868
rect 40964 924 41020 934
rect 40964 748 41020 868
rect 44436 812 44492 1204
rect 44436 746 44492 756
rect 44660 812 44716 7140
rect 47012 5740 47068 5750
rect 47012 5608 47068 5684
rect 47460 5628 47516 5638
rect 47012 5572 47460 5608
rect 47012 5552 47516 5572
rect 44772 4732 44828 4742
rect 44772 1596 44828 4676
rect 48580 3268 48636 8036
rect 51828 6244 52220 6300
rect 51828 5964 51884 6244
rect 51828 5898 51884 5908
rect 52052 6076 52108 6086
rect 51604 5852 51660 5862
rect 49812 5068 49868 5078
rect 49252 3808 49308 3818
rect 48580 3212 48748 3268
rect 45892 2828 45948 2838
rect 45892 2156 45948 2772
rect 45892 2090 45948 2100
rect 44772 1530 44828 1540
rect 44660 746 44716 756
rect 48692 748 48748 3212
rect 49252 3088 49308 3752
rect 49252 3022 49308 3032
rect 49700 3268 49756 3278
rect 49028 2908 49084 2918
rect 49028 2368 49084 2852
rect 49028 2302 49084 2312
rect 49700 1484 49756 3212
rect 49700 1418 49756 1428
rect 40964 682 41020 692
rect 48692 682 48748 692
rect 25956 502 26012 512
rect 19684 322 19740 332
rect 15988 142 16044 152
rect 49812 208 49868 5012
rect 51604 4888 51660 5796
rect 52052 5852 52108 6020
rect 52164 5964 52220 6244
rect 52164 5898 52220 5908
rect 52052 5786 52108 5796
rect 51604 4822 51660 4832
rect 50372 3948 50428 3958
rect 50372 3612 50428 3892
rect 50372 3546 50428 3556
rect 50596 3612 50652 3622
rect 50596 3387 50652 3556
rect 50484 3331 50652 3387
rect 49924 2728 49980 2738
rect 49924 476 49980 2672
rect 50148 1828 50204 1838
rect 50148 1148 50204 1772
rect 50148 1082 50204 1092
rect 50372 1148 50428 1158
rect 50372 812 50428 1092
rect 50372 746 50428 756
rect 50484 700 50540 3331
rect 50596 1260 50652 1270
rect 50596 812 50652 1204
rect 50596 746 50652 756
rect 50484 634 50540 644
rect 52052 700 52108 710
rect 49924 410 49980 420
rect 52052 252 52108 644
rect 52164 588 52220 598
rect 52164 494 52220 512
rect 52052 186 52108 196
rect 52276 252 52332 8932
rect 53620 7980 53676 7990
rect 53620 6688 53676 7924
rect 54068 7980 54124 13292
rect 56196 12908 56252 12918
rect 55412 12348 55468 12358
rect 55412 12124 55468 12292
rect 55636 12348 55692 12358
rect 55636 12268 55692 12292
rect 55636 12202 55692 12212
rect 55972 12268 56028 12278
rect 55412 12058 55468 12068
rect 55300 11908 55356 11918
rect 55300 11340 55356 11852
rect 55300 11274 55356 11284
rect 55748 11676 55804 11686
rect 55748 10648 55804 11620
rect 55748 10582 55804 10592
rect 54068 7914 54124 7924
rect 55512 9436 55832 10252
rect 55512 9380 55540 9436
rect 55596 9380 55644 9436
rect 55700 9380 55748 9436
rect 55804 9380 55832 9436
rect 55512 9030 55832 9380
rect 55512 8974 55540 9030
rect 55596 8974 55644 9030
rect 55700 8974 55748 9030
rect 55804 8974 55832 9030
rect 55512 8926 55832 8974
rect 55512 8870 55540 8926
rect 55596 8870 55644 8926
rect 55700 8870 55748 8926
rect 55804 8870 55832 8926
rect 55512 8822 55832 8870
rect 55512 8766 55540 8822
rect 55596 8766 55644 8822
rect 55700 8766 55748 8822
rect 55804 8766 55832 8822
rect 55512 7868 55832 8766
rect 55972 8540 56028 12212
rect 56196 12236 56252 12852
rect 56196 12170 56252 12180
rect 56196 11564 56252 11574
rect 56196 11340 56252 11508
rect 56196 11274 56252 11284
rect 56308 11548 56364 11558
rect 56308 10108 56364 11492
rect 56308 10042 56364 10052
rect 55972 8474 56028 8484
rect 55512 7812 55540 7868
rect 55596 7812 55644 7868
rect 55700 7812 55748 7868
rect 55804 7812 55832 7868
rect 55512 7632 55832 7812
rect 55512 7576 55540 7632
rect 55596 7576 55644 7632
rect 55700 7576 55748 7632
rect 55804 7576 55832 7632
rect 55512 7528 55832 7576
rect 55512 7472 55540 7528
rect 55596 7472 55644 7528
rect 55700 7472 55748 7528
rect 55804 7472 55832 7528
rect 55512 7424 55832 7472
rect 55512 7368 55540 7424
rect 55596 7368 55644 7424
rect 55700 7368 55748 7424
rect 55804 7368 55832 7424
rect 53620 6632 53900 6688
rect 53844 3836 53900 6632
rect 55512 6300 55832 7368
rect 55512 6244 55540 6300
rect 55596 6244 55644 6300
rect 55700 6244 55748 6300
rect 55804 6244 55832 6300
rect 55512 6234 55832 6244
rect 55512 6178 55540 6234
rect 55596 6178 55644 6234
rect 55700 6178 55748 6234
rect 55804 6178 55832 6234
rect 55512 6130 55832 6178
rect 55512 6074 55540 6130
rect 55596 6074 55644 6130
rect 55700 6074 55748 6130
rect 55804 6074 55832 6130
rect 55512 6026 55832 6074
rect 55512 5970 55540 6026
rect 55596 5970 55644 6026
rect 55700 5970 55748 6026
rect 55804 5970 55832 6026
rect 54180 5628 54236 5638
rect 54180 4528 54236 5572
rect 55512 4732 55832 5970
rect 55972 5180 56028 5190
rect 56644 5180 56700 13652
rect 60228 12088 60284 12098
rect 57092 11788 57148 11798
rect 57092 11564 57148 11732
rect 57092 11498 57148 11508
rect 57764 11788 57820 11798
rect 56756 10648 56812 10658
rect 56756 10288 56812 10592
rect 56980 10648 57036 10658
rect 56980 10444 57036 10592
rect 56980 10378 57036 10388
rect 56756 10222 56812 10232
rect 57204 10108 57260 10118
rect 57204 8988 57260 10052
rect 57204 8922 57260 8932
rect 57428 7980 57484 7990
rect 57428 6300 57484 7924
rect 57428 6234 57484 6244
rect 56028 5124 56700 5180
rect 55972 5114 56028 5124
rect 55512 4676 55540 4732
rect 55596 4676 55644 4732
rect 55700 4676 55748 4732
rect 55804 4676 55832 4732
rect 55512 4644 55832 4676
rect 56196 4956 56252 4966
rect 56196 4620 56252 4900
rect 56644 4956 56700 5124
rect 57428 5516 57484 5526
rect 57428 5180 57484 5460
rect 57428 5114 57484 5124
rect 56644 4890 56700 4900
rect 56196 4554 56252 4564
rect 54180 4462 54236 4472
rect 55300 4396 55356 4406
rect 53844 3770 53900 3780
rect 54964 4284 55020 4294
rect 52724 3164 52780 3174
rect 52724 1932 52780 3108
rect 52948 2940 53004 2950
rect 52948 2380 53004 2884
rect 54964 2492 55020 4228
rect 55300 4168 55356 4340
rect 55300 4102 55356 4112
rect 55524 4168 55580 4178
rect 55300 3836 55356 3846
rect 55300 3500 55356 3780
rect 55524 3808 55580 4112
rect 55524 3742 55580 3752
rect 56980 4060 57036 4070
rect 55300 3434 55356 3444
rect 55076 3268 55132 3278
rect 55076 3088 55132 3212
rect 55300 3276 55356 3306
rect 55300 3202 55356 3212
rect 55076 3032 55468 3088
rect 54964 2426 55020 2436
rect 55300 2940 55356 2950
rect 52948 2314 53004 2324
rect 53172 2380 53228 2390
rect 53172 2286 53228 2312
rect 52724 1866 52780 1876
rect 53508 2268 53564 2278
rect 53508 1148 53564 2212
rect 55300 2188 55356 2884
rect 55412 2188 55468 3032
rect 56980 2380 57036 4004
rect 56980 2314 57036 2324
rect 57092 3052 57148 3062
rect 55524 2188 55580 2198
rect 55412 2132 55524 2188
rect 55300 2122 55356 2132
rect 55524 2122 55580 2132
rect 56980 2044 57036 2054
rect 53620 2008 53676 2018
rect 53620 1372 53676 1952
rect 53620 1306 53676 1316
rect 54068 1148 54124 1158
rect 53508 1092 54068 1148
rect 54068 1082 54124 1092
rect 56980 588 57036 1988
rect 57092 700 57148 2996
rect 57428 3052 57484 3062
rect 57092 634 57148 644
rect 57316 2716 57372 2726
rect 56980 522 57036 532
rect 57316 568 57372 2660
rect 57316 502 57372 512
rect 57428 476 57484 2996
rect 57428 410 57484 420
rect 57764 364 57820 11732
rect 59556 10668 59612 10678
rect 59556 10108 59612 10612
rect 59556 10042 59612 10052
rect 58660 9772 58716 9782
rect 58436 6508 58492 6518
rect 58436 6300 58492 6452
rect 58436 6234 58492 6244
rect 58660 5180 58716 9716
rect 60228 9100 60284 12032
rect 60452 11908 60508 14912
rect 71428 14968 71484 14978
rect 70196 14812 70252 14822
rect 67844 14788 67900 14798
rect 65604 14588 65660 14598
rect 61460 13916 61516 13926
rect 60452 11842 60508 11852
rect 60788 11908 60844 11918
rect 60228 9034 60284 9044
rect 60340 8988 60396 8998
rect 60396 8932 60508 8988
rect 60340 8922 60396 8932
rect 60004 8204 60060 8214
rect 60004 7420 60060 8148
rect 60452 7868 60508 8932
rect 60676 8540 60732 8550
rect 60676 7980 60732 8484
rect 60676 7914 60732 7924
rect 60452 7802 60508 7812
rect 60788 7756 60844 11852
rect 61460 9884 61516 13860
rect 65604 13692 65660 14532
rect 67620 14428 67676 14438
rect 67620 13888 67676 14372
rect 67844 14428 67900 14732
rect 67844 14362 67900 14372
rect 68516 14788 68572 14798
rect 70252 14756 70364 14812
rect 70196 14746 70252 14756
rect 67620 13822 67676 13832
rect 65604 13626 65660 13636
rect 65940 13692 65996 13702
rect 64036 13580 64092 13590
rect 63252 13528 63308 13538
rect 63252 12460 63308 13472
rect 63252 12394 63308 12404
rect 63700 13528 63756 13538
rect 63476 12124 63532 12134
rect 62132 11788 62188 11798
rect 62132 10444 62188 11732
rect 62132 10378 62188 10388
rect 63364 11008 63420 11018
rect 62916 10108 62972 10118
rect 62916 9928 62972 10052
rect 62916 9862 62972 9872
rect 61460 9818 61516 9828
rect 63252 8428 63308 8438
rect 60788 7690 60844 7700
rect 62580 8092 62636 8102
rect 62580 7644 62636 8036
rect 62580 7578 62636 7588
rect 60004 7354 60060 7364
rect 62804 7420 62860 7430
rect 58660 5114 58716 5124
rect 60004 6300 60060 6310
rect 58772 3276 58828 3286
rect 58772 2548 58828 3220
rect 60004 3164 60060 6244
rect 62804 5068 62860 7364
rect 62804 5002 62860 5012
rect 62580 4172 62636 4182
rect 61684 3948 61740 3958
rect 61684 3612 61740 3892
rect 62580 3948 62636 4116
rect 62580 3882 62636 3892
rect 61684 3546 61740 3556
rect 62132 3808 62188 3818
rect 61908 3500 61964 3510
rect 62132 3448 62188 3752
rect 61964 3444 62188 3448
rect 61908 3392 62188 3444
rect 60004 3098 60060 3108
rect 58772 2482 58828 2492
rect 59220 2908 59276 2918
rect 59220 1260 59276 2852
rect 59892 2492 59948 2502
rect 59892 1648 59948 2436
rect 61572 2492 61628 2502
rect 60340 2368 60396 2378
rect 61572 2368 61628 2436
rect 60396 2312 60508 2368
rect 61572 2312 62187 2368
rect 60340 2302 60396 2312
rect 59892 1582 59948 1592
rect 59220 1194 59276 1204
rect 59780 1484 59836 1494
rect 59780 476 59836 1428
rect 60340 1484 60396 1494
rect 60340 1108 60396 1428
rect 60452 1260 60508 2312
rect 62131 2268 62187 2312
rect 62131 2202 62187 2212
rect 60788 2188 60844 2198
rect 60788 2044 60844 2132
rect 60788 1978 60844 1988
rect 62468 2008 62524 2018
rect 62468 1932 62524 1952
rect 62468 1866 62524 1876
rect 62804 2008 62860 2018
rect 62804 1932 62860 1952
rect 62804 1866 62860 1876
rect 62131 1596 62187 1606
rect 62131 1468 62187 1540
rect 60452 1194 60508 1204
rect 61908 1412 62187 1468
rect 61908 1260 61964 1412
rect 62580 1372 62636 1382
rect 62580 1288 62636 1316
rect 61908 1194 61964 1204
rect 62132 1260 62636 1288
rect 62188 1232 62636 1260
rect 62132 1194 62188 1204
rect 60340 1042 60396 1052
rect 60564 1108 60620 1118
rect 59780 410 59836 420
rect 57764 298 57820 308
rect 52276 186 52332 196
rect 60564 252 60620 1052
rect 60564 186 60620 196
rect 63252 208 63308 8372
rect 63364 7228 63420 10952
rect 63476 8428 63532 12068
rect 63700 12124 63756 13472
rect 63700 12058 63756 12068
rect 63924 13468 63980 13478
rect 63924 11452 63980 13412
rect 64036 13020 64092 13524
rect 65940 13168 65996 13636
rect 67732 13692 68348 13708
rect 67788 13652 68348 13692
rect 67732 13626 67788 13636
rect 68068 13580 68124 13590
rect 68068 13244 68124 13524
rect 68292 13580 68348 13652
rect 68292 13514 68348 13524
rect 68068 13178 68124 13188
rect 65940 13102 65996 13112
rect 66612 13168 66668 13178
rect 64036 12954 64092 12964
rect 65380 11788 65436 11798
rect 65380 11728 65436 11732
rect 65380 11662 65436 11672
rect 65604 11728 65660 11738
rect 63924 11386 63980 11396
rect 65044 11340 65100 11350
rect 63476 8362 63532 8372
rect 63588 9928 63644 9938
rect 63364 7162 63420 7172
rect 63588 6508 63644 9872
rect 63812 7644 63868 7654
rect 63812 6688 63868 7588
rect 63700 6636 63868 6688
rect 63756 6632 63868 6636
rect 64596 7420 64652 7430
rect 63700 6570 63756 6580
rect 63588 6442 63644 6452
rect 64596 5852 64652 7364
rect 63700 5788 63756 5798
rect 64596 5786 64652 5796
rect 63700 4888 63756 5732
rect 63700 4822 63756 4832
rect 63700 3724 63756 3734
rect 63700 3276 63756 3668
rect 63700 3210 63756 3220
rect 63924 3164 63980 3174
rect 63924 1288 63980 3108
rect 64148 3088 64204 3098
rect 64148 2986 64204 2996
rect 64708 3052 64764 3062
rect 64708 2156 64764 2996
rect 65044 2548 65100 11284
rect 65604 4168 65660 11672
rect 66612 11676 66668 13112
rect 68516 12628 68572 14732
rect 69076 14428 69132 14438
rect 68628 13888 68684 13898
rect 68852 13888 68908 13898
rect 68684 13832 68796 13888
rect 68628 13822 68684 13832
rect 68516 12562 68572 12572
rect 67508 12236 67564 12246
rect 66948 11908 67004 11918
rect 66612 11610 66668 11620
rect 66836 11676 66892 11686
rect 66836 11452 66892 11620
rect 66836 11386 66892 11396
rect 66948 10220 67004 11852
rect 67172 11788 67228 11798
rect 67508 11788 67564 12180
rect 67172 11452 67228 11732
rect 67396 11728 67452 11738
rect 67508 11722 67564 11732
rect 68516 11908 68572 11918
rect 67396 11610 67452 11620
rect 68180 11676 68236 11686
rect 67172 11386 67228 11396
rect 68180 10468 68236 11620
rect 68516 11228 68572 11852
rect 68516 11162 68572 11172
rect 68628 11008 68684 11018
rect 68180 10402 68236 10412
rect 68404 10668 68460 10678
rect 68404 10468 68460 10612
rect 68404 10402 68460 10412
rect 68628 10444 68684 10952
rect 68740 10668 68796 13832
rect 68852 12572 68908 13832
rect 68852 12506 68908 12516
rect 68964 12628 69020 12638
rect 68852 12124 68908 12134
rect 68852 11908 68908 12068
rect 68852 11842 68908 11852
rect 68740 10602 68796 10612
rect 68628 10378 68684 10388
rect 66948 10154 67004 10164
rect 67060 10288 67116 10298
rect 66724 8876 66780 8886
rect 66724 8668 66780 8820
rect 67060 8876 67116 10232
rect 67060 8810 67116 8820
rect 68628 10108 68684 10118
rect 66724 8612 67228 8668
rect 66948 8316 67004 8326
rect 65268 4112 65660 4168
rect 66724 6508 66780 6518
rect 65268 3948 65324 4112
rect 66276 4060 66332 4070
rect 65268 3882 65324 3892
rect 65492 3948 65548 3958
rect 65380 3628 65436 3650
rect 65380 3546 65436 3556
rect 65492 3268 65548 3892
rect 65492 3202 65548 3212
rect 66276 3164 66332 4004
rect 66724 3836 66780 6452
rect 66836 6300 66892 6310
rect 66836 4956 66892 6244
rect 66836 4890 66892 4900
rect 66724 3770 66780 3780
rect 66836 4620 66892 4630
rect 66276 3098 66332 3108
rect 65492 2548 65548 2558
rect 65044 2482 65100 2492
rect 65380 2492 65492 2548
rect 65492 2482 65548 2492
rect 65380 2426 65436 2436
rect 64708 2090 64764 2100
rect 63812 1232 63980 1288
rect 65380 1820 65436 1830
rect 63812 748 63868 1232
rect 65380 1036 65436 1764
rect 65380 970 65436 980
rect 65940 1596 65996 1606
rect 49812 142 49868 152
rect 63252 142 63308 152
rect 63588 692 63868 748
rect 63588 140 63644 692
rect 63588 74 63644 84
rect 65940 140 65996 1540
rect 66836 1372 66892 4564
rect 66948 3052 67004 8260
rect 67060 6748 67116 6758
rect 67060 6524 67116 6692
rect 67060 6458 67116 6468
rect 67060 4168 67116 4178
rect 67060 3836 67116 4112
rect 67060 3770 67116 3780
rect 67172 3808 67228 8612
rect 67956 7588 68572 7644
rect 67956 7420 68012 7588
rect 68516 7532 68572 7588
rect 68516 7466 68572 7476
rect 67956 7354 68012 7364
rect 67284 7228 67340 7238
rect 67284 6972 67340 7172
rect 68180 7228 68236 7238
rect 67956 6972 68012 6982
rect 67284 6916 67956 6972
rect 67956 6906 68012 6916
rect 68180 6300 68236 7172
rect 68628 6636 68684 10052
rect 68964 9884 69020 12572
rect 69076 12572 69132 14372
rect 70084 14364 70140 14374
rect 69636 14140 69692 14150
rect 69076 12506 69132 12516
rect 69524 12684 69580 12694
rect 69412 12268 69468 12278
rect 69412 11340 69468 12212
rect 69524 11676 69580 12628
rect 69636 12268 69692 14084
rect 69636 12202 69692 12212
rect 69748 12460 69804 12470
rect 69524 11610 69580 11620
rect 69748 11676 69804 12404
rect 69972 12460 70028 12470
rect 69972 11728 70028 12404
rect 70084 12348 70140 14308
rect 70084 12282 70140 12292
rect 70308 12348 70364 14756
rect 70308 12282 70364 12292
rect 69972 11662 70028 11672
rect 69748 11610 69804 11620
rect 69412 11274 69468 11284
rect 68964 9818 69020 9828
rect 70756 10668 70812 10678
rect 69524 9660 69580 9670
rect 68740 6860 68796 6870
rect 69188 6860 69244 6870
rect 68796 6804 69188 6860
rect 68740 6794 68796 6804
rect 69188 6794 69244 6804
rect 68628 6570 68684 6580
rect 68180 6234 68236 6244
rect 68628 6188 68684 6198
rect 67284 5852 67340 5862
rect 67340 5796 68012 5852
rect 67284 5786 67340 5796
rect 67508 4888 67564 4898
rect 67284 4844 67340 4854
rect 67284 3836 67340 4788
rect 67508 4348 67564 4832
rect 67956 4708 68012 5796
rect 68628 5788 68684 6132
rect 68628 5740 69468 5788
rect 68628 5732 69412 5740
rect 69412 5674 69468 5684
rect 68404 5292 68460 5302
rect 68180 4708 68236 4718
rect 67956 4652 68180 4708
rect 68180 4642 68236 4652
rect 67508 4282 67564 4292
rect 67956 4508 68012 4518
rect 67956 4168 68012 4452
rect 68404 4168 68460 5236
rect 67956 4102 68012 4112
rect 68292 4112 68460 4168
rect 69188 4172 69244 4182
rect 69524 4172 69580 9604
rect 69972 9324 70028 9334
rect 69748 7308 69804 7318
rect 69748 4956 69804 7252
rect 69748 4890 69804 4900
rect 69244 4116 69580 4172
rect 68292 4060 68348 4112
rect 69188 4106 69244 4116
rect 68292 3994 68348 4004
rect 67284 3770 67340 3780
rect 67172 3742 67228 3752
rect 68628 3612 68684 3622
rect 66948 2986 67004 2996
rect 67172 3276 67228 3286
rect 66836 1306 66892 1316
rect 67060 2828 67116 2838
rect 67060 1372 67116 2772
rect 67172 2604 67228 3220
rect 67396 3276 67452 3286
rect 67396 2728 67452 3220
rect 67396 2662 67452 2672
rect 67732 3268 67788 3278
rect 67172 2538 67228 2548
rect 67620 2492 67676 2502
rect 67620 2268 67676 2436
rect 67732 2368 67788 3212
rect 67732 2302 67788 2312
rect 68068 2728 68124 2738
rect 67620 2202 67676 2212
rect 67060 1306 67116 1316
rect 68068 1260 68124 2672
rect 68068 1194 68124 1204
rect 68516 748 68572 758
rect 67732 692 68516 748
rect 67732 208 67788 692
rect 68516 682 68572 692
rect 68628 476 68684 3556
rect 69972 3276 70028 9268
rect 70420 8876 70476 8886
rect 70420 8652 70476 8820
rect 70420 8586 70476 8596
rect 70532 8316 70588 8326
rect 70532 7980 70588 8260
rect 70532 7914 70588 7924
rect 70084 5068 70140 5078
rect 70084 4956 70140 5012
rect 70084 4890 70140 4900
rect 70308 5068 70364 5078
rect 70308 4708 70364 5012
rect 70308 4642 70364 4652
rect 70532 4708 70588 4718
rect 70532 3836 70588 4652
rect 70532 3770 70588 3780
rect 70756 3836 70812 10612
rect 71204 9212 71260 9222
rect 70868 6300 70924 6310
rect 70868 5292 70924 6244
rect 70868 5226 70924 5236
rect 71204 4956 71260 9156
rect 71428 9212 71484 14912
rect 71652 14968 71708 14978
rect 85876 14968 85932 14978
rect 86660 14968 86716 14978
rect 77364 14924 79772 14968
rect 71652 14812 71708 14912
rect 71652 14746 71708 14756
rect 74004 14912 79772 14924
rect 74004 14868 77420 14912
rect 72772 14428 72828 14438
rect 72772 13708 72828 14372
rect 72772 13642 72828 13652
rect 73108 13916 73164 13926
rect 71764 13168 71820 13178
rect 71652 11728 71708 11738
rect 71652 11368 71708 11672
rect 71652 11302 71708 11312
rect 71428 9146 71484 9156
rect 71204 4890 71260 4900
rect 71316 7532 71372 7542
rect 70756 3770 70812 3780
rect 69972 3210 70028 3220
rect 70084 3612 70140 3622
rect 70084 2716 70140 3556
rect 70084 2650 70140 2660
rect 70756 3052 70812 3062
rect 70532 2188 70588 2198
rect 70532 1148 70588 2132
rect 70532 1082 70588 1092
rect 70756 1148 70812 2996
rect 71316 2492 71372 7476
rect 71428 5068 71484 5078
rect 71428 4284 71484 5012
rect 71428 4218 71484 4228
rect 71652 3052 71708 3062
rect 71316 2426 71372 2436
rect 71540 2492 71596 2502
rect 71540 1596 71596 2436
rect 71652 2044 71708 2996
rect 71652 1978 71708 1988
rect 71540 1530 71596 1540
rect 71764 1596 71820 13112
rect 71988 13168 72044 13178
rect 71988 12236 72044 13112
rect 73108 12684 73164 13860
rect 73220 13708 73276 13718
rect 73220 13132 73276 13652
rect 73556 13412 73948 13468
rect 73220 13066 73276 13076
rect 73444 13132 73500 13142
rect 73108 12618 73164 12628
rect 71988 12170 72044 12180
rect 73444 10108 73500 13076
rect 73556 12460 73612 13412
rect 73780 13244 73836 13254
rect 73780 12908 73836 13188
rect 73892 13020 73948 13412
rect 74004 13168 74060 14868
rect 77588 14812 77644 14822
rect 77644 14756 79212 14812
rect 77588 14746 77644 14756
rect 77924 14588 77980 14598
rect 78148 14588 78204 14598
rect 77140 14532 77924 14588
rect 74676 13916 74732 13926
rect 74004 13102 74060 13112
rect 74228 13804 74284 13814
rect 74228 13168 74284 13748
rect 74228 13102 74284 13112
rect 73892 12964 74620 13020
rect 73780 12842 73836 12852
rect 74564 12684 74620 12964
rect 74676 12908 74732 13860
rect 77140 13916 77196 14532
rect 77924 14522 77980 14532
rect 78036 14532 78148 14588
rect 77476 14372 77756 14428
rect 77476 14364 77532 14372
rect 77476 14298 77532 14308
rect 77588 14252 77644 14262
rect 77140 13850 77196 13860
rect 77252 14012 77532 14068
rect 77252 13468 77308 14012
rect 75348 13412 77308 13468
rect 77364 13916 77420 13926
rect 75236 12908 75292 12918
rect 74676 12852 75236 12908
rect 75236 12842 75292 12852
rect 75348 12684 75404 13412
rect 77364 13356 77420 13860
rect 77476 13692 77532 14012
rect 77588 13888 77644 14196
rect 77700 14028 77756 14372
rect 77700 13962 77756 13972
rect 78036 13888 78092 14532
rect 78148 14522 78204 14532
rect 78932 14428 78988 14438
rect 77588 13832 78092 13888
rect 78148 14252 78204 14262
rect 77476 13636 77980 13692
rect 77588 13468 77644 13478
rect 77812 13468 77868 13478
rect 77644 13412 77756 13468
rect 77588 13402 77644 13412
rect 74564 12628 75404 12684
rect 77028 13300 77420 13356
rect 73556 12394 73612 12404
rect 73668 12572 74396 12628
rect 73556 12236 73612 12246
rect 73556 12088 73612 12180
rect 73556 12022 73612 12032
rect 73668 11908 73724 12572
rect 73668 11842 73724 11852
rect 74004 12460 74060 12470
rect 74004 11728 74060 12404
rect 74340 12268 74396 12572
rect 74340 12202 74396 12212
rect 74452 12448 74508 12458
rect 74116 12124 74172 12134
rect 74452 12124 74508 12392
rect 74172 12068 74508 12124
rect 74116 12058 74172 12068
rect 75012 12012 75068 12022
rect 74340 11956 75012 12012
rect 74340 11900 74396 11956
rect 75012 11946 75068 11956
rect 74116 11844 74396 11900
rect 75124 11900 75180 11910
rect 74116 11788 74172 11844
rect 74116 11722 74172 11732
rect 74228 11728 74284 11738
rect 74004 11662 74060 11672
rect 74228 11340 74284 11672
rect 73668 11284 74284 11340
rect 75124 11368 75180 11844
rect 75124 11302 75180 11312
rect 75460 11368 75516 11378
rect 73668 11228 73724 11284
rect 73668 11162 73724 11172
rect 74116 11188 74172 11198
rect 73444 10042 73500 10052
rect 73668 10108 73724 10118
rect 73668 9928 73724 10052
rect 72212 9884 72268 9894
rect 73668 9862 73724 9872
rect 73892 9928 73948 9938
rect 72212 9388 72268 9828
rect 72996 9660 73052 9670
rect 72212 9332 72604 9388
rect 72548 9324 72604 9332
rect 72548 9258 72604 9268
rect 72772 8876 72828 8886
rect 72660 8428 72716 8438
rect 72436 8204 72492 8214
rect 72436 8128 72492 8148
rect 72100 8072 72492 8128
rect 71988 7644 72044 7654
rect 71988 7308 72044 7588
rect 71988 7242 72044 7252
rect 72100 7196 72156 8072
rect 72100 7130 72156 7140
rect 72324 7308 72380 7318
rect 72212 4732 72268 4742
rect 72212 3448 72268 4676
rect 72212 3382 72268 3392
rect 72100 2156 72156 2166
rect 71876 2100 72100 2156
rect 71876 1648 71932 2100
rect 72100 2090 72156 2100
rect 71876 1582 71932 1592
rect 72100 1648 72156 1658
rect 71764 1530 71820 1540
rect 71988 1484 72044 1494
rect 71988 1148 72044 1428
rect 72100 1372 72156 1592
rect 72100 1306 72156 1316
rect 71988 1092 72268 1148
rect 70756 1082 70812 1092
rect 71988 748 72044 758
rect 72212 748 72268 1092
rect 72044 692 72156 748
rect 71988 682 72044 692
rect 72100 568 72156 692
rect 72212 682 72268 692
rect 72100 502 72156 512
rect 67844 420 68684 476
rect 72324 476 72380 7252
rect 72548 4396 72604 4406
rect 72548 1260 72604 4340
rect 72660 2492 72716 8372
rect 72772 4396 72828 8820
rect 72996 8876 73052 9604
rect 72996 8810 73052 8820
rect 72772 4330 72828 4340
rect 72996 8540 73052 8550
rect 72996 3724 73052 8484
rect 73892 7308 73948 9872
rect 73892 7242 73948 7252
rect 73668 6748 73724 6758
rect 73108 6300 73164 6310
rect 73108 5740 73164 6244
rect 73556 5852 73612 5862
rect 73556 5788 73612 5796
rect 73108 5674 73164 5684
rect 73220 5732 73612 5788
rect 73220 5516 73276 5732
rect 73668 5628 73724 6692
rect 73668 5562 73724 5572
rect 73780 5964 73836 5974
rect 73220 5450 73276 5460
rect 73444 5516 73500 5526
rect 73332 5180 73388 5190
rect 73444 5180 73500 5460
rect 73780 5292 73836 5908
rect 73780 5226 73836 5236
rect 74004 5964 74060 5974
rect 73388 5124 73500 5180
rect 73332 5114 73388 5124
rect 74004 4844 74060 5908
rect 73108 4788 74060 4844
rect 73108 4708 73164 4788
rect 73108 4642 73164 4652
rect 73332 4708 73388 4718
rect 72996 3658 73052 3668
rect 73108 4060 73164 4070
rect 73108 3500 73164 4004
rect 72660 2426 72716 2436
rect 72996 3448 73052 3458
rect 73108 3434 73164 3444
rect 73220 3612 73276 3622
rect 72996 1820 73052 3392
rect 73220 2156 73276 3556
rect 73332 2716 73388 4652
rect 74004 4348 74060 4358
rect 74116 4348 74172 11132
rect 75012 10108 75068 10118
rect 75012 9212 75068 10052
rect 75012 9146 75068 9156
rect 74900 8428 74956 8438
rect 74340 8316 74396 8326
rect 74340 7644 74396 8260
rect 74900 8092 74956 8372
rect 74900 8026 74956 8036
rect 75124 8092 75180 8102
rect 74340 7578 74396 7588
rect 74788 7868 74844 7878
rect 74788 5740 74844 7812
rect 75012 7196 75068 7206
rect 74900 7140 75012 7196
rect 74900 6860 74956 7140
rect 75012 7130 75068 7140
rect 74900 6794 74956 6804
rect 74788 5674 74844 5684
rect 75012 5740 75068 5750
rect 75012 5516 75068 5684
rect 75012 5450 75068 5460
rect 74788 4956 74844 4966
rect 74340 4620 74396 4630
rect 74060 4292 74172 4348
rect 74228 4348 74284 4358
rect 74004 4282 74060 4292
rect 74228 4284 74284 4292
rect 74228 4218 74284 4228
rect 74340 3276 74396 4564
rect 74788 3612 74844 4900
rect 75124 3988 75180 8036
rect 75348 7532 75404 7542
rect 75348 6972 75404 7476
rect 75348 6906 75404 6916
rect 75460 5964 75516 11312
rect 76468 10388 76972 10444
rect 76244 10288 76300 10298
rect 76244 9660 76300 10232
rect 76468 10108 76524 10388
rect 76468 10042 76524 10052
rect 76244 9594 76300 9604
rect 76916 8316 76972 10388
rect 77028 9996 77084 13300
rect 77476 13244 77532 13254
rect 77140 13188 77476 13244
rect 77140 13020 77196 13188
rect 77476 13178 77532 13188
rect 77588 13168 77644 13178
rect 77588 13066 77644 13076
rect 77140 12954 77196 12964
rect 77700 12628 77756 13412
rect 77812 12796 77868 13412
rect 77924 13356 77980 13636
rect 78148 13528 78204 14196
rect 78148 13462 78204 13472
rect 78260 14196 78876 14252
rect 78260 13356 78316 14196
rect 78372 14084 78764 14140
rect 78372 13528 78428 14084
rect 78708 14028 78764 14084
rect 78708 13962 78764 13972
rect 78484 13888 78540 13898
rect 78484 13708 78540 13832
rect 78820 13888 78876 14196
rect 78932 13916 78988 14372
rect 79156 14428 79212 14756
rect 79604 14588 79660 14598
rect 79156 14362 79212 14372
rect 79492 14532 79604 14588
rect 79492 14252 79548 14532
rect 79604 14522 79660 14532
rect 79492 14186 79548 14196
rect 79716 14252 79772 14912
rect 80388 14912 81788 14968
rect 80388 14588 80444 14912
rect 80836 14812 80892 14822
rect 80388 14522 80444 14532
rect 80612 14588 80668 14598
rect 79716 14186 79772 14196
rect 79044 14140 79100 14150
rect 79044 14068 79100 14084
rect 79604 14140 79660 14150
rect 79604 14068 79660 14084
rect 80612 14140 80668 14532
rect 80612 14074 80668 14084
rect 80836 14140 80892 14756
rect 81284 14700 81340 14710
rect 81284 14608 81340 14644
rect 81508 14608 81564 14618
rect 81284 14542 81340 14552
rect 81396 14552 81508 14608
rect 81396 14248 81452 14552
rect 81508 14542 81564 14552
rect 80836 14074 80892 14084
rect 81172 14192 81452 14248
rect 81508 14428 81564 14438
rect 81508 14252 81564 14372
rect 81732 14428 81788 14912
rect 82404 14912 84140 14968
rect 82180 14812 82236 14822
rect 81732 14362 81788 14372
rect 82068 14476 82124 14486
rect 82180 14476 82236 14756
rect 82292 14476 82348 14486
rect 82180 14420 82292 14476
rect 81508 14196 82012 14252
rect 79044 14012 79660 14068
rect 81172 13916 81228 14192
rect 81284 14068 81340 14078
rect 81284 13962 81340 13972
rect 81396 14012 81900 14068
rect 78932 13860 81228 13916
rect 78820 13822 78876 13832
rect 81396 13804 81452 14012
rect 78932 13748 81452 13804
rect 81732 13916 81788 13926
rect 78932 13708 78988 13748
rect 78484 13652 78988 13708
rect 78372 13462 78428 13472
rect 77924 13300 78316 13356
rect 81620 13348 81676 13358
rect 79380 13292 81564 13348
rect 77924 13168 77980 13178
rect 79380 13168 79436 13292
rect 77924 13020 77980 13112
rect 77924 12954 77980 12964
rect 78596 13112 79436 13168
rect 80612 13168 80668 13178
rect 81396 13168 81452 13178
rect 78596 12796 78652 13112
rect 78932 13020 78988 13030
rect 78988 12964 80220 13020
rect 78932 12954 78988 12964
rect 79044 12852 80108 12908
rect 77812 12730 77868 12740
rect 78148 12740 78652 12796
rect 78820 12796 78876 12806
rect 77924 12684 77980 12694
rect 77700 12572 77980 12628
rect 78148 12572 78204 12740
rect 78372 12572 78428 12582
rect 78148 12506 78204 12516
rect 78260 12516 78372 12572
rect 77364 12460 77420 12470
rect 77028 9930 77084 9940
rect 77140 12088 77196 12098
rect 77140 9436 77196 12032
rect 77364 12088 77420 12404
rect 77364 12022 77420 12032
rect 78260 12012 78316 12516
rect 78372 12506 78428 12516
rect 78820 12448 78876 12740
rect 78932 12572 78988 12582
rect 79044 12572 79100 12852
rect 80052 12572 80108 12852
rect 78988 12516 79100 12572
rect 79156 12516 79996 12572
rect 78932 12506 78988 12516
rect 79156 12448 79212 12516
rect 78820 12392 79212 12448
rect 79380 12392 79884 12448
rect 77812 11956 78316 12012
rect 78484 12348 78540 12358
rect 77700 11788 77756 11798
rect 77252 11676 77308 11686
rect 77252 9660 77308 11620
rect 77700 11564 77756 11732
rect 77588 11508 77756 11564
rect 77588 10288 77644 11508
rect 77700 11368 77756 11378
rect 77700 10780 77756 11312
rect 77700 10714 77756 10724
rect 77812 10444 77868 11956
rect 78484 11908 78540 12292
rect 79268 12268 79324 12278
rect 78484 11842 78540 11852
rect 78596 12032 78876 12088
rect 77924 11788 77980 11798
rect 77924 11116 77980 11732
rect 78260 11728 78316 11738
rect 78484 11728 78540 11738
rect 78316 11672 78428 11728
rect 78260 11662 78316 11672
rect 77924 11050 77980 11060
rect 78036 11368 78092 11378
rect 77588 10222 77644 10232
rect 77700 10388 77868 10444
rect 77700 9996 77756 10388
rect 77588 9928 77644 9938
rect 77700 9930 77756 9940
rect 77812 10220 77868 10230
rect 77252 9594 77308 9604
rect 77364 9772 77420 9782
rect 77588 9772 77644 9872
rect 77812 9928 77868 10164
rect 77812 9862 77868 9872
rect 77924 9996 77980 10006
rect 77924 9772 77980 9940
rect 77588 9716 77980 9772
rect 77028 9380 77196 9436
rect 77028 8540 77084 9380
rect 77028 8474 77084 8484
rect 77251 8540 77307 8550
rect 77364 8540 77420 9716
rect 78036 9208 78092 11312
rect 78372 11116 78428 11672
rect 78372 11050 78428 11060
rect 78148 10468 78204 10478
rect 78148 9660 78204 10412
rect 78372 10468 78428 10478
rect 78148 9594 78204 9604
rect 78260 10220 78316 10230
rect 77924 9152 78092 9208
rect 77812 8652 77868 8662
rect 77924 8652 77980 9152
rect 78260 9028 78316 10164
rect 78372 9324 78428 10412
rect 78372 9258 78428 9268
rect 77868 8596 77980 8652
rect 78036 8972 78316 9028
rect 77812 8586 77868 8596
rect 77307 8484 77420 8540
rect 77700 8540 77756 8550
rect 77251 8474 77307 8484
rect 77700 8316 77756 8484
rect 76916 8260 77756 8316
rect 78036 8204 78092 8972
rect 78484 8848 78540 11672
rect 77252 8148 78092 8204
rect 78148 8792 78540 8848
rect 77252 7980 77308 8148
rect 77252 7914 77308 7924
rect 77476 7980 77532 7990
rect 77476 7768 77532 7924
rect 77028 7712 77532 7768
rect 75460 5898 75516 5908
rect 75796 7420 75852 7430
rect 75796 5628 75852 7364
rect 75908 7308 75964 7318
rect 75908 5852 75964 7252
rect 76132 7196 76188 7206
rect 76188 7140 76300 7196
rect 76132 7130 76188 7140
rect 76244 6860 76300 7140
rect 76244 6794 76300 6804
rect 75908 5786 75964 5796
rect 76468 5964 76524 5974
rect 75796 5562 75852 5572
rect 76132 4284 76188 4294
rect 75796 4228 76132 4284
rect 75124 3922 75180 3932
rect 75348 3988 75404 3998
rect 75348 3836 75404 3932
rect 75348 3770 75404 3780
rect 74788 3546 74844 3556
rect 74900 3388 74956 3398
rect 74340 3210 74396 3220
rect 74564 3276 74620 3306
rect 74564 3202 74620 3212
rect 74900 3268 74956 3332
rect 74900 3202 74956 3212
rect 75572 3276 75628 3286
rect 75124 3088 75180 3098
rect 73332 2650 73388 2660
rect 73444 3032 74060 3088
rect 73220 2090 73276 2100
rect 73444 2008 73500 3032
rect 73444 1942 73500 1952
rect 73780 2728 73836 2738
rect 73780 2008 73836 2672
rect 74004 2728 74060 3032
rect 74004 2662 74060 2672
rect 73780 1942 73836 1952
rect 74340 2604 74396 2614
rect 72996 1754 73052 1764
rect 74340 1828 74396 2548
rect 74340 1762 74396 1772
rect 74564 1932 74620 1942
rect 74564 1828 74620 1876
rect 74564 1762 74620 1772
rect 72548 1194 72604 1204
rect 74900 1484 74956 1494
rect 74116 1148 74172 1158
rect 67844 388 67900 420
rect 72324 410 72380 420
rect 72548 812 72604 822
rect 72548 476 72604 756
rect 74116 812 74172 1092
rect 74116 746 74172 756
rect 72548 410 72604 420
rect 67844 322 67900 332
rect 74900 252 74956 1428
rect 75124 748 75180 3032
rect 75460 3088 75516 3098
rect 75236 2156 75292 2166
rect 75236 1708 75292 2100
rect 75460 2044 75516 3032
rect 75572 2268 75628 3220
rect 75572 2202 75628 2212
rect 75684 2604 75740 2614
rect 75460 1978 75516 1988
rect 75684 2044 75740 2548
rect 75684 1978 75740 1988
rect 75236 1642 75292 1652
rect 75460 1708 75516 1718
rect 75460 1260 75516 1652
rect 75236 1204 75516 1260
rect 75796 1288 75852 4228
rect 76132 4218 76188 4228
rect 76468 2368 76524 5908
rect 76804 4956 76860 4966
rect 76692 4396 76748 4406
rect 76692 3500 76748 4340
rect 76692 3434 76748 3444
rect 76804 3388 76860 4900
rect 76804 3322 76860 3332
rect 76468 2302 76524 2312
rect 76916 3268 76972 3278
rect 76916 2368 76972 3212
rect 76916 2302 76972 2312
rect 75796 1222 75852 1232
rect 76244 1484 76300 1494
rect 76244 1288 76300 1428
rect 77028 1372 77084 7712
rect 78148 7532 78204 8792
rect 78596 8668 78652 12032
rect 78708 11900 78764 11910
rect 78708 9996 78764 11844
rect 78820 11116 78876 12032
rect 79044 11900 79100 11910
rect 79044 11368 79100 11844
rect 79044 11302 79100 11312
rect 79156 11908 79212 11918
rect 79044 11116 79100 11126
rect 78820 11060 79044 11116
rect 79044 11050 79100 11060
rect 79044 10288 79100 10298
rect 78708 9930 78764 9940
rect 78820 10108 78876 10118
rect 77140 7476 78204 7532
rect 78260 8612 78652 8668
rect 78708 9324 78764 9334
rect 78260 7532 78316 8612
rect 77140 5068 77196 7476
rect 78260 7466 78316 7476
rect 78484 8540 78540 8550
rect 78484 7532 78540 8484
rect 78708 8092 78764 9268
rect 78708 8026 78764 8036
rect 78820 9212 78876 10052
rect 79044 9928 79100 10232
rect 79156 10108 79212 11852
rect 79268 10288 79324 12212
rect 79380 11564 79436 12392
rect 79828 12348 79884 12392
rect 79828 12282 79884 12292
rect 79492 12268 79548 12278
rect 79492 11728 79548 12212
rect 79940 12236 79996 12516
rect 80052 12506 80108 12516
rect 79940 12170 79996 12180
rect 79492 11662 79548 11672
rect 79716 11728 79772 11738
rect 79380 11508 79548 11564
rect 79268 10222 79324 10232
rect 79380 11368 79436 11378
rect 79380 10220 79436 11312
rect 79380 10154 79436 10164
rect 79156 10042 79212 10052
rect 79492 9996 79548 11508
rect 79716 11368 79772 11672
rect 79716 11302 79772 11312
rect 79828 11340 79884 11350
rect 79380 9940 79548 9996
rect 79044 9872 79324 9928
rect 78484 7466 78540 7476
rect 78148 7308 78204 7318
rect 78148 6972 78204 7252
rect 78148 6906 78204 6916
rect 78708 6412 78764 6422
rect 77140 5002 77196 5012
rect 78596 5852 78652 5862
rect 78036 4472 78428 4528
rect 78036 4348 78092 4472
rect 77700 4292 78092 4348
rect 78372 4396 78428 4472
rect 78484 4396 78540 4406
rect 78372 4340 78484 4396
rect 78484 4330 78540 4340
rect 77364 4060 77420 4070
rect 77028 1306 77084 1316
rect 77140 3948 77196 3958
rect 77140 1288 77196 3892
rect 77252 3500 77308 3510
rect 77252 1484 77308 3444
rect 77364 3268 77420 4004
rect 77700 3948 77756 4292
rect 78036 4172 78092 4182
rect 77700 3882 77756 3892
rect 77812 4060 77868 4070
rect 77812 3500 77868 4004
rect 77812 3434 77868 3444
rect 77924 3948 77980 3958
rect 77364 3202 77420 3212
rect 77476 3276 77532 3286
rect 77252 1418 77308 1428
rect 77476 1484 77532 3220
rect 77700 3276 77756 3286
rect 77700 2156 77756 3220
rect 77924 3268 77980 3892
rect 77924 3202 77980 3212
rect 78036 2716 78092 4116
rect 78260 4172 78316 4182
rect 78260 3988 78316 4116
rect 78260 3922 78316 3932
rect 78596 3388 78652 5796
rect 78708 5628 78764 6356
rect 78708 5562 78764 5572
rect 78708 5180 78764 5190
rect 78708 3808 78764 5124
rect 78708 3742 78764 3752
rect 78260 3332 78652 3388
rect 78260 3276 78316 3332
rect 78820 3276 78876 9156
rect 79044 8316 79100 8326
rect 78932 7868 78988 7878
rect 78932 7308 78988 7812
rect 78932 7242 78988 7252
rect 78932 5628 78988 5638
rect 78932 4348 78988 5572
rect 79044 5180 79100 8260
rect 79268 7420 79324 9872
rect 79380 8540 79436 9940
rect 79380 8474 79436 8484
rect 79492 9660 79548 9670
rect 79492 8316 79548 9604
rect 79492 8250 79548 8260
rect 79716 8764 79772 8774
rect 79716 7644 79772 8708
rect 79828 8540 79884 11284
rect 80052 10108 80108 10118
rect 79940 9324 79996 9334
rect 79940 8764 79996 9268
rect 79940 8698 79996 8708
rect 79828 8474 79884 8484
rect 79716 7578 79772 7588
rect 80052 7420 80108 10052
rect 80164 7868 80220 12964
rect 80500 12796 80556 12806
rect 80388 12572 80444 12582
rect 80276 12460 80332 12470
rect 80276 12012 80332 12404
rect 80388 12448 80444 12516
rect 80388 12382 80444 12392
rect 80276 11946 80332 11956
rect 80388 12236 80444 12246
rect 80388 11340 80444 12180
rect 80500 12012 80556 12740
rect 80612 12448 80668 13112
rect 80612 12382 80668 12392
rect 80724 13132 80780 13142
rect 81060 13132 81116 13142
rect 80724 12124 80780 13076
rect 80836 13076 81060 13132
rect 80836 12988 80892 13076
rect 81060 13066 81116 13076
rect 81172 13112 81396 13168
rect 80836 12922 80892 12932
rect 80836 12808 80892 12834
rect 80836 12730 80892 12740
rect 81172 12460 81228 13112
rect 81396 13102 81452 13112
rect 81396 12988 81452 12998
rect 81284 12932 81396 12988
rect 81284 12572 81340 12932
rect 81396 12922 81452 12932
rect 81284 12506 81340 12516
rect 81060 12404 81228 12460
rect 81508 12460 81564 13292
rect 81620 12988 81676 13292
rect 81732 12988 81788 13860
rect 81844 13888 81900 14012
rect 81844 13822 81900 13832
rect 81844 13692 81900 13702
rect 81844 13356 81900 13636
rect 81956 13528 82012 14196
rect 82068 13692 82124 14420
rect 82292 14410 82348 14420
rect 82404 14248 82460 14912
rect 82516 14788 82572 14798
rect 83188 14788 83244 14798
rect 82516 14248 82572 14732
rect 82740 14732 83188 14788
rect 82740 14608 82796 14732
rect 83188 14722 83244 14732
rect 84084 14788 84140 14912
rect 85932 14912 86044 14968
rect 85876 14902 85932 14912
rect 84084 14722 84140 14732
rect 82740 14542 82796 14552
rect 83300 14552 85820 14608
rect 82628 14476 82684 14486
rect 82684 14420 83244 14476
rect 82628 14410 82684 14420
rect 83188 14248 83244 14420
rect 83300 14428 83356 14552
rect 83300 14362 83356 14372
rect 83860 14428 83916 14438
rect 82516 14192 83132 14248
rect 83188 14192 83692 14248
rect 82404 14182 82460 14192
rect 82292 14012 82684 14068
rect 82292 13916 82348 14012
rect 82292 13850 82348 13860
rect 82068 13626 82124 13636
rect 81956 13472 82460 13528
rect 81844 13300 82124 13356
rect 81844 12988 81900 12998
rect 81732 12932 81844 12988
rect 81620 12922 81676 12932
rect 81844 12922 81900 12932
rect 82068 12684 82124 13300
rect 82404 13348 82460 13472
rect 82628 13356 82684 14012
rect 82852 13804 82908 13814
rect 82740 13708 82796 13718
rect 82852 13708 82908 13748
rect 83076 13804 83132 14192
rect 83076 13738 83132 13748
rect 83188 14068 83244 14078
rect 82964 13708 83020 13718
rect 82852 13652 82964 13708
rect 82740 13528 82796 13652
rect 82964 13642 83020 13652
rect 83188 13580 83244 14012
rect 82740 13472 83132 13528
rect 83188 13514 83244 13524
rect 83412 13580 83468 13590
rect 82740 13356 82796 13366
rect 82404 13292 82572 13348
rect 82628 13300 82740 13356
rect 82516 13132 82572 13292
rect 82740 13290 82796 13300
rect 83076 13348 83132 13472
rect 83300 13356 83356 13366
rect 83076 13300 83300 13348
rect 83076 13292 83356 13300
rect 83300 13290 83356 13292
rect 83412 13132 83468 13524
rect 82516 13076 83468 13132
rect 83524 13132 83580 13142
rect 83636 13132 83692 14192
rect 83748 13132 83804 13142
rect 83636 13076 83748 13132
rect 83524 12988 83580 13076
rect 83748 13066 83804 13076
rect 83860 12988 83916 14372
rect 85204 14248 85260 14258
rect 85428 14248 85484 14258
rect 83524 12932 83916 12988
rect 83972 13580 84028 13590
rect 85204 13580 85260 14192
rect 83972 12808 84028 13524
rect 84868 13528 84924 13538
rect 84644 13132 84700 13142
rect 82628 12740 83244 12796
rect 82068 12628 82236 12684
rect 81732 12572 81788 12582
rect 82180 12572 82460 12628
rect 80836 12124 80892 12134
rect 80724 12068 80836 12124
rect 80836 12058 80892 12068
rect 80500 11946 80556 11956
rect 81060 11340 81116 12404
rect 81508 12394 81564 12404
rect 81620 12516 81732 12572
rect 81620 12448 81676 12516
rect 81732 12506 81788 12516
rect 81844 12448 81900 12458
rect 81620 12382 81676 12392
rect 81732 12392 81844 12448
rect 81732 12268 81788 12392
rect 81844 12382 81900 12392
rect 81396 12236 81788 12268
rect 81284 12212 81788 12236
rect 81284 12180 81452 12212
rect 81172 12124 81228 12134
rect 81284 12124 81340 12180
rect 81228 12068 81340 12124
rect 82404 12124 82460 12572
rect 82628 12268 82684 12740
rect 83076 12628 83132 12638
rect 83076 12268 83132 12572
rect 83188 12448 83244 12740
rect 83636 12752 84028 12808
rect 84532 12988 84588 12998
rect 84644 12988 84700 13076
rect 84868 13132 84924 13472
rect 85092 13528 85148 13538
rect 85204 13514 85260 13524
rect 85316 14192 85428 14248
rect 85092 13168 85148 13472
rect 85092 13102 85148 13112
rect 85204 13132 85260 13142
rect 84868 13066 84924 13076
rect 84756 12988 84812 12998
rect 84644 12932 84756 12988
rect 83300 12628 83356 12638
rect 83300 12460 83356 12572
rect 83300 12394 83356 12404
rect 83188 12382 83244 12392
rect 83412 12348 83468 12358
rect 83412 12268 83468 12292
rect 83636 12268 83692 12752
rect 84308 12572 84364 12582
rect 84084 12448 84140 12458
rect 83076 12212 83468 12268
rect 83524 12212 83692 12268
rect 83748 12348 83804 12358
rect 83972 12348 84028 12358
rect 82628 12202 82684 12212
rect 81172 12058 81228 12068
rect 81620 12032 82236 12088
rect 82404 12068 82572 12124
rect 81620 11728 81676 12032
rect 82068 11900 82124 11910
rect 82068 11788 82124 11844
rect 81620 11662 81676 11672
rect 81732 11732 82124 11788
rect 82180 11788 82236 12032
rect 82292 12012 82348 12022
rect 82292 11900 82348 11956
rect 82516 12012 82572 12068
rect 83076 12088 83132 12098
rect 83524 12088 83580 12212
rect 83132 12032 83580 12088
rect 83748 12088 83804 12292
rect 83076 12022 83132 12032
rect 83748 12022 83804 12032
rect 83860 12292 83972 12348
rect 82516 11946 82572 11956
rect 82292 11844 82460 11900
rect 82180 11732 82348 11788
rect 80388 11274 80444 11284
rect 80500 11284 81116 11340
rect 80500 10220 80556 11284
rect 81732 11228 81788 11732
rect 81956 11620 82236 11676
rect 81956 11340 82012 11620
rect 81956 11274 82012 11284
rect 82068 11452 82124 11462
rect 80500 10154 80556 10164
rect 80724 11172 81788 11228
rect 81844 11188 81900 11198
rect 80724 10108 80780 11172
rect 82068 11188 82124 11396
rect 82180 11340 82236 11620
rect 82292 11564 82348 11732
rect 82404 11728 82460 11844
rect 83860 11676 83916 12292
rect 83972 12282 84028 12292
rect 84084 12268 84140 12392
rect 84308 12448 84364 12516
rect 84308 12382 84364 12392
rect 84084 12212 84364 12268
rect 82404 11662 82460 11672
rect 82516 11620 83916 11676
rect 82516 11564 82572 11620
rect 82292 11508 82572 11564
rect 83524 11548 83580 11558
rect 82964 11452 83020 11462
rect 83300 11452 83356 11462
rect 83524 11452 83580 11492
rect 84308 11548 84364 12212
rect 84532 11900 84588 12932
rect 84756 12922 84812 12932
rect 84644 12740 85036 12796
rect 84644 12348 84700 12740
rect 84644 12282 84700 12292
rect 84756 12572 84812 12582
rect 84532 11834 84588 11844
rect 84756 11908 84812 12516
rect 84756 11842 84812 11852
rect 84868 12348 84924 12358
rect 84308 11482 84364 11492
rect 84084 11452 84140 11462
rect 83020 11396 83244 11452
rect 82964 11386 83020 11396
rect 82516 11340 82572 11350
rect 82180 11284 82516 11340
rect 82516 11274 82572 11284
rect 83188 11228 83244 11396
rect 83356 11396 83468 11452
rect 83300 11386 83356 11396
rect 83412 11228 83468 11396
rect 83524 11386 83580 11396
rect 83636 11396 84084 11452
rect 83636 11228 83692 11396
rect 84084 11386 84140 11396
rect 82068 11132 82348 11188
rect 83188 11172 83356 11228
rect 83412 11172 83692 11228
rect 83748 11228 83804 11238
rect 84868 11188 84924 12292
rect 84980 11908 85036 12740
rect 84980 11842 85036 11852
rect 85204 11908 85260 13076
rect 85204 11842 85260 11852
rect 85316 11188 85372 14192
rect 85428 14182 85484 14192
rect 81844 11116 81900 11132
rect 81508 11060 81900 11116
rect 81508 10780 81564 11060
rect 82068 11004 82124 11014
rect 81620 10948 82068 11004
rect 82292 11008 82348 11132
rect 83300 11116 83356 11172
rect 83748 11116 83804 11172
rect 83300 11060 83804 11116
rect 83860 11132 84924 11188
rect 84980 11132 85372 11188
rect 85428 13168 85484 13178
rect 83188 11008 83244 11014
rect 82292 11004 83244 11008
rect 82292 10952 83188 11004
rect 81620 10892 81676 10948
rect 82068 10938 82124 10948
rect 83188 10938 83244 10948
rect 83860 11008 83916 11132
rect 83860 10942 83916 10952
rect 84084 11008 84140 11018
rect 81620 10826 81676 10836
rect 81508 10714 81564 10724
rect 84084 10648 84140 10952
rect 84980 11008 85036 11132
rect 85204 11008 85260 11018
rect 84980 10942 85036 10952
rect 85092 10952 85204 11008
rect 80724 10042 80780 10052
rect 80836 10592 84140 10648
rect 80836 9436 80892 10592
rect 85092 10468 85148 10952
rect 85204 10942 85260 10952
rect 81844 10388 83132 10444
rect 80164 7802 80220 7812
rect 80276 9380 80892 9436
rect 80948 10220 81004 10230
rect 79268 7364 79884 7420
rect 79268 6916 79660 6972
rect 79268 6748 79324 6916
rect 79268 6682 79324 6692
rect 79492 6748 79548 6758
rect 79044 5114 79100 5124
rect 78932 4282 78988 4292
rect 79156 4348 79212 4358
rect 79156 4168 79212 4292
rect 79044 4112 79212 4168
rect 79044 4060 79100 4112
rect 78932 4004 79100 4060
rect 78932 3500 78988 4004
rect 79380 3988 79436 3998
rect 79156 3948 79212 3958
rect 78932 3434 78988 3444
rect 79044 3836 79100 3846
rect 78820 3220 78988 3276
rect 78260 3210 78316 3220
rect 78036 2660 78876 2716
rect 77700 2090 77756 2100
rect 77924 2604 77980 2614
rect 77924 2156 77980 2548
rect 78820 2604 78876 2660
rect 78820 2538 78876 2548
rect 77924 2090 77980 2100
rect 77476 1418 77532 1428
rect 78932 1372 78988 3220
rect 79044 3268 79100 3780
rect 79156 3612 79212 3892
rect 79380 3836 79436 3932
rect 79380 3770 79436 3780
rect 79156 3546 79212 3556
rect 79380 3612 79436 3622
rect 79492 3612 79548 6692
rect 79604 6688 79660 6916
rect 79828 6860 79884 7364
rect 80052 7354 80108 7364
rect 80052 6860 80108 6870
rect 79828 6804 80052 6860
rect 80052 6794 80108 6804
rect 80276 6688 80332 9380
rect 80948 9324 81004 10164
rect 80724 9268 81004 9324
rect 81396 10108 81452 10118
rect 81396 9324 81452 10052
rect 81844 9568 81900 10388
rect 82404 10220 82460 10230
rect 82292 9996 82348 10006
rect 82292 9928 82348 9940
rect 80500 8988 80556 8998
rect 80500 8764 80556 8932
rect 80500 8698 80556 8708
rect 79604 6632 80332 6688
rect 80388 6972 80444 6982
rect 80388 6748 80444 6916
rect 80612 6748 80668 6758
rect 80388 6682 80444 6692
rect 80500 6692 80612 6748
rect 80500 6300 80556 6692
rect 80612 6682 80668 6692
rect 79436 3556 79548 3612
rect 79604 6244 80556 6300
rect 79380 3546 79436 3556
rect 79044 3202 79100 3212
rect 79604 2156 79660 6244
rect 80052 5740 80108 5750
rect 80724 5740 80780 9268
rect 81396 9258 81452 9268
rect 81508 9512 81900 9568
rect 81956 9828 82236 9884
rect 82292 9862 82348 9872
rect 80948 9152 81340 9208
rect 80948 8092 81004 9152
rect 81284 8848 81340 9152
rect 81284 8792 81452 8848
rect 80948 8026 81004 8036
rect 81284 8652 81340 8662
rect 81284 8092 81340 8596
rect 81284 8026 81340 8036
rect 81396 7532 81452 8792
rect 81508 8540 81564 9512
rect 81844 9324 81900 9334
rect 81844 9230 81900 9268
rect 81956 8668 82012 9828
rect 82180 9772 82236 9828
rect 82404 9772 82460 10164
rect 82676 10220 82996 10252
rect 82676 10164 82704 10220
rect 82760 10164 82808 10220
rect 82864 10164 82912 10220
rect 82968 10164 82996 10220
rect 82180 9716 82460 9772
rect 82516 9928 82572 9938
rect 81508 8474 81564 8484
rect 81844 8612 82012 8668
rect 82292 9212 82348 9222
rect 81844 8204 81900 8612
rect 81844 8138 81900 8148
rect 82068 8540 82124 8550
rect 80836 7476 81228 7532
rect 81396 7476 81564 7532
rect 80836 6636 80892 7476
rect 80836 6570 80892 6580
rect 80948 7308 81004 7318
rect 80108 5684 80444 5740
rect 80052 5674 80108 5684
rect 79716 5180 79772 5190
rect 79716 4620 79772 5124
rect 80052 5068 80108 5078
rect 80108 5012 80332 5068
rect 80052 5002 80108 5012
rect 79828 4788 80220 4844
rect 79828 4708 79884 4788
rect 79828 4642 79884 4652
rect 80052 4708 80108 4718
rect 79716 4528 79772 4564
rect 79716 4472 79996 4528
rect 79828 4396 79884 4406
rect 79716 4172 79772 4182
rect 79716 3052 79772 4116
rect 79828 3628 79884 4340
rect 79940 3836 79996 4472
rect 80052 4396 80108 4652
rect 80052 4330 80108 4340
rect 80164 4284 80220 4788
rect 80276 4396 80332 5012
rect 80388 4956 80444 5684
rect 80724 5674 80780 5684
rect 80388 4890 80444 4900
rect 80948 4888 81004 7252
rect 81172 7308 81228 7476
rect 81172 7242 81228 7252
rect 81396 7308 81452 7318
rect 81396 5516 81452 7252
rect 81508 5852 81564 7476
rect 82068 6972 82124 8484
rect 82292 8204 82348 9156
rect 82516 9212 82572 9872
rect 82516 9146 82572 9156
rect 82676 9729 82996 10164
rect 83076 9928 83132 10388
rect 83524 10412 85148 10468
rect 83524 10332 83580 10412
rect 83524 10266 83580 10276
rect 83188 10108 83244 10118
rect 85428 10108 85484 13112
rect 85652 12268 85708 12278
rect 83244 10052 85484 10108
rect 85540 11908 85596 11918
rect 83188 10042 83244 10052
rect 85540 9928 85596 11852
rect 83076 9872 83356 9928
rect 82676 9673 82704 9729
rect 82760 9673 82808 9729
rect 82864 9673 82912 9729
rect 82968 9673 82996 9729
rect 82676 9625 82996 9673
rect 83188 9772 83244 9782
rect 83300 9772 83356 9872
rect 85428 9872 85596 9928
rect 83412 9772 83468 9782
rect 83300 9716 83412 9772
rect 82676 9569 82704 9625
rect 82760 9569 82808 9625
rect 82864 9569 82912 9625
rect 82968 9569 82996 9625
rect 82676 9521 82996 9569
rect 82676 9465 82704 9521
rect 82760 9465 82808 9521
rect 82864 9465 82912 9521
rect 82968 9465 82996 9521
rect 82292 8138 82348 8148
rect 82676 8652 82996 9465
rect 83076 9660 83132 9670
rect 83076 9208 83132 9604
rect 83188 9436 83244 9716
rect 83412 9706 83468 9716
rect 83636 9512 84812 9568
rect 83300 9436 83356 9446
rect 83188 9380 83300 9436
rect 83300 9370 83356 9380
rect 83076 9152 83244 9208
rect 82676 8596 82704 8652
rect 82760 8596 82808 8652
rect 82864 8596 82912 8652
rect 82968 8596 82996 8652
rect 82676 8331 82996 8596
rect 82676 8275 82704 8331
rect 82760 8275 82808 8331
rect 82864 8275 82912 8331
rect 82968 8275 82996 8331
rect 82676 8227 82996 8275
rect 82676 8171 82704 8227
rect 82760 8171 82808 8227
rect 82864 8171 82912 8227
rect 82968 8171 82996 8227
rect 82676 8123 82996 8171
rect 82068 6906 82124 6916
rect 82404 8092 82460 8102
rect 82180 6860 82236 6870
rect 81956 6412 82012 6422
rect 82012 6356 82124 6412
rect 81956 6346 82012 6356
rect 81508 5786 81564 5796
rect 81396 5450 81452 5460
rect 80948 4822 81004 4832
rect 81396 5192 81676 5248
rect 80500 4620 80556 4630
rect 80500 4528 80556 4564
rect 80500 4462 80556 4472
rect 80276 4340 80668 4396
rect 80612 4284 80668 4340
rect 80724 4284 80780 4294
rect 80164 4228 80444 4284
rect 80612 4228 80724 4284
rect 80388 4060 80444 4228
rect 80724 4218 80780 4228
rect 80388 4004 80668 4060
rect 80612 3988 80668 4004
rect 80612 3922 80668 3932
rect 79940 3780 81004 3836
rect 80948 3724 81004 3780
rect 81172 3724 81228 3734
rect 80948 3668 81172 3724
rect 81172 3658 81228 3668
rect 79828 3562 79884 3572
rect 80836 3628 80892 3638
rect 80612 3500 80668 3510
rect 80388 3444 80612 3500
rect 80164 3052 80220 3062
rect 79716 2996 80164 3052
rect 80164 2986 80220 2996
rect 79492 2100 79660 2156
rect 79492 1484 79548 2100
rect 80388 1932 80444 3444
rect 80612 3434 80668 3444
rect 80500 2548 80556 2558
rect 80836 2548 80892 3572
rect 80556 2492 80892 2548
rect 80500 2482 80556 2492
rect 80836 2380 80892 2390
rect 81396 2380 81452 5192
rect 81508 5068 81564 5078
rect 81620 5068 81676 5192
rect 81732 5068 81788 5078
rect 81620 5012 81732 5068
rect 81508 4844 81564 5012
rect 81732 5002 81788 5012
rect 82068 4956 82124 6356
rect 82180 5788 82236 6804
rect 82404 5964 82460 8036
rect 82676 8067 82704 8123
rect 82760 8067 82808 8123
rect 82864 8067 82912 8123
rect 82968 8067 82996 8123
rect 82516 7868 82572 7878
rect 82516 7196 82572 7812
rect 82516 7130 82572 7140
rect 82676 7084 82996 8067
rect 82676 7028 82704 7084
rect 82760 7028 82808 7084
rect 82864 7028 82912 7084
rect 82968 7028 82996 7084
rect 82676 6933 82996 7028
rect 82676 6877 82704 6933
rect 82760 6877 82808 6933
rect 82864 6877 82912 6933
rect 82968 6877 82996 6933
rect 82676 6829 82996 6877
rect 82676 6773 82704 6829
rect 82760 6773 82808 6829
rect 82864 6773 82912 6829
rect 82968 6773 82996 6829
rect 82516 6748 82572 6758
rect 82516 6524 82572 6692
rect 82516 6458 82572 6468
rect 82676 6725 82996 6773
rect 82676 6669 82704 6725
rect 82760 6669 82808 6725
rect 82864 6669 82912 6725
rect 82968 6669 82996 6725
rect 82404 5898 82460 5908
rect 82180 5732 82572 5788
rect 82180 4956 82236 4966
rect 82068 4900 82180 4956
rect 82180 4890 82236 4900
rect 82404 4844 82460 4854
rect 81508 4788 81788 4844
rect 81508 4528 81564 4538
rect 81508 4172 81564 4472
rect 81508 4106 81564 4116
rect 81620 4284 81676 4294
rect 81508 3276 81564 3286
rect 81508 3182 81564 3212
rect 79492 1418 79548 1428
rect 79604 1876 80444 1932
rect 80724 1932 80780 1942
rect 78932 1306 78988 1316
rect 79380 1288 79436 1298
rect 79604 1288 79660 1876
rect 79716 1708 79772 1718
rect 80052 1708 80108 1718
rect 79772 1652 79884 1708
rect 79716 1642 79772 1652
rect 79716 1484 79772 1494
rect 79716 1390 79772 1412
rect 77140 1232 78652 1288
rect 76244 1222 76300 1232
rect 75236 924 75292 1204
rect 78596 1108 78652 1232
rect 79436 1232 79660 1288
rect 79380 1222 79436 1232
rect 79828 1108 79884 1652
rect 79940 1468 79996 1478
rect 79940 1372 79996 1412
rect 79940 1306 79996 1316
rect 76020 1052 78540 1108
rect 78596 1052 79772 1108
rect 75460 924 75516 934
rect 75236 858 75292 868
rect 75348 868 75460 924
rect 75348 748 75404 868
rect 75460 858 75516 868
rect 76020 924 76076 1052
rect 76020 858 76076 868
rect 76244 924 76300 934
rect 75124 692 75404 748
rect 76244 700 76300 868
rect 76356 928 76412 938
rect 76412 872 78428 928
rect 76356 862 76412 872
rect 76244 634 76300 644
rect 76804 748 76860 758
rect 76804 634 76860 644
rect 77140 700 77196 710
rect 76580 476 76636 486
rect 75236 388 75292 398
rect 75124 332 75236 388
rect 75124 252 75180 332
rect 75236 322 75292 332
rect 74900 196 75180 252
rect 76580 208 76636 420
rect 76692 364 76748 374
rect 77140 364 77196 644
rect 76748 308 77196 364
rect 77252 476 77308 486
rect 76692 298 76748 308
rect 77252 208 77308 420
rect 78148 388 78204 398
rect 78148 252 78204 332
rect 78372 388 78428 872
rect 78484 568 78540 1052
rect 79156 868 79660 924
rect 79156 568 79212 868
rect 78484 512 79212 568
rect 79268 700 79324 710
rect 78372 322 78428 332
rect 79268 252 79324 644
rect 79604 364 79660 868
rect 79604 298 79660 308
rect 76580 152 77308 208
rect 77364 208 77420 218
rect 77588 208 77644 218
rect 77420 152 77588 208
rect 78148 196 79324 252
rect 79716 252 79772 1052
rect 79828 1042 79884 1052
rect 80052 476 80108 1652
rect 80388 924 80444 934
rect 80388 700 80444 868
rect 80388 634 80444 644
rect 80724 700 80780 1876
rect 80724 634 80780 644
rect 80276 476 80332 486
rect 80052 410 80108 420
rect 80164 420 80276 476
rect 80164 252 80220 420
rect 80276 410 80332 420
rect 79716 196 80220 252
rect 80836 208 80892 2324
rect 81060 2368 81116 2378
rect 81396 2314 81452 2324
rect 80948 2188 81004 2198
rect 80948 1036 81004 2132
rect 80948 970 81004 980
rect 81060 812 81116 2312
rect 81172 2188 81228 2198
rect 81172 1468 81228 2132
rect 81396 2044 81452 2054
rect 81396 1708 81452 1988
rect 81396 1642 81452 1652
rect 81172 1402 81228 1412
rect 81396 1468 81452 1478
rect 81396 1260 81452 1412
rect 81060 746 81116 756
rect 81172 1204 81452 1260
rect 81060 364 81116 374
rect 81172 364 81228 1204
rect 81116 308 81228 364
rect 81508 924 81564 934
rect 81060 298 81116 308
rect 81508 208 81564 868
rect 81620 476 81676 4228
rect 81732 3500 81788 4788
rect 81732 3434 81788 3444
rect 81844 4172 81900 4182
rect 81844 924 81900 4116
rect 82404 3836 82460 4788
rect 82516 4528 82572 5732
rect 82676 5535 82996 6669
rect 83076 7644 83132 7654
rect 83076 6636 83132 7588
rect 83076 6570 83132 6580
rect 83188 6508 83244 9152
rect 82676 5460 82704 5535
rect 82760 5460 82808 5535
rect 82864 5460 82912 5535
rect 82968 5460 82996 5535
rect 82676 5431 82996 5460
rect 82676 5375 82704 5431
rect 82760 5375 82808 5431
rect 82864 5375 82912 5431
rect 82968 5375 82996 5431
rect 82676 5327 82996 5375
rect 82676 5271 82704 5327
rect 82760 5271 82808 5327
rect 82864 5271 82912 5327
rect 82968 5271 82996 5327
rect 82676 4644 82996 5271
rect 83076 6452 83244 6508
rect 83412 7196 83468 7206
rect 83076 4732 83132 6452
rect 83300 5852 83356 5862
rect 83076 4666 83132 4676
rect 83188 5788 83244 5798
rect 82516 4472 83132 4528
rect 81956 3780 82460 3836
rect 82964 4284 83020 4294
rect 81956 3612 82012 3780
rect 82740 3724 82796 3734
rect 81956 3546 82012 3556
rect 82068 3668 82740 3724
rect 82068 3500 82124 3668
rect 82740 3658 82796 3668
rect 82852 3612 82908 3622
rect 82068 3434 82124 3444
rect 82180 3448 82236 3458
rect 81956 3268 82012 3278
rect 81956 2908 82012 3212
rect 81956 2842 82012 2852
rect 82180 2908 82236 3392
rect 82180 2842 82236 2852
rect 82404 3448 82460 3458
rect 82404 2548 82460 3392
rect 82068 2492 82460 2548
rect 82516 3052 82572 3062
rect 82068 2380 82124 2492
rect 82068 2314 82124 2324
rect 82292 2380 82348 2390
rect 82292 2008 82348 2324
rect 82292 1942 82348 1952
rect 82292 1468 82348 1478
rect 82516 1468 82572 2996
rect 82852 2828 82908 3556
rect 82964 3276 83020 4228
rect 82964 3210 83020 3220
rect 83076 3088 83132 4472
rect 82852 2762 82908 2772
rect 82964 3032 83132 3088
rect 83188 3052 83244 5732
rect 82740 2368 82796 2378
rect 82740 2008 82796 2312
rect 82740 1942 82796 1952
rect 82348 1412 82460 1468
rect 82292 1402 82348 1412
rect 82292 1288 82348 1298
rect 81844 858 81900 868
rect 82180 924 82236 934
rect 81620 410 81676 420
rect 81956 812 82012 822
rect 80836 152 81564 208
rect 81956 208 82012 756
rect 82180 388 82236 868
rect 82292 812 82348 1232
rect 82292 746 82348 756
rect 82404 476 82460 1412
rect 82516 1402 82572 1412
rect 82964 1468 83020 3032
rect 83188 2986 83244 2996
rect 83188 2828 83244 2838
rect 82964 1402 83020 1412
rect 83076 2156 83132 2166
rect 82852 1372 82908 1382
rect 82852 924 82908 1316
rect 82852 858 82908 868
rect 83076 924 83132 2100
rect 83188 1828 83244 2772
rect 83300 2368 83356 5796
rect 83412 5788 83468 7140
rect 83636 7196 83692 9512
rect 84420 9436 84476 9446
rect 83748 8652 83804 8662
rect 83748 7420 83804 8596
rect 83972 8652 84028 8662
rect 83972 8092 84028 8596
rect 83972 8026 84028 8036
rect 84308 7980 84364 7990
rect 83748 7354 83804 7364
rect 83860 7924 84308 7948
rect 83860 7892 84364 7924
rect 83636 7130 83692 7140
rect 83412 5722 83468 5732
rect 83524 6972 83580 6982
rect 83524 5516 83580 6916
rect 83860 6412 83916 7892
rect 83860 6346 83916 6356
rect 83972 7644 84028 7654
rect 83524 5450 83580 5460
rect 83972 4956 84028 7588
rect 84196 7308 84252 7318
rect 83972 4890 84028 4900
rect 84084 6412 84140 6422
rect 83412 3724 83468 3734
rect 83412 3628 83468 3668
rect 83636 3628 83692 3638
rect 83412 3562 83468 3572
rect 83524 3572 83636 3628
rect 83524 3500 83580 3572
rect 83636 3562 83692 3572
rect 84084 3612 84140 6356
rect 84084 3546 84140 3556
rect 83748 3500 83804 3510
rect 83300 2302 83356 2312
rect 83412 3448 83468 3458
rect 83524 3434 83580 3444
rect 83636 3444 83748 3500
rect 83412 2156 83468 3392
rect 83636 2828 83692 3444
rect 83748 3434 83804 3444
rect 83860 3448 83916 3458
rect 83860 2940 83916 3392
rect 83972 3276 84028 3286
rect 84196 3276 84252 7252
rect 84308 6524 84364 6534
rect 84308 5404 84364 6468
rect 84420 6188 84476 9380
rect 84420 6122 84476 6132
rect 84532 8204 84588 8214
rect 84308 5338 84364 5348
rect 84532 5404 84588 8148
rect 84756 8204 84812 9512
rect 84756 8138 84812 8148
rect 84868 8988 84924 8998
rect 84756 7420 84812 7430
rect 84644 7084 84700 7094
rect 84644 6748 84700 7028
rect 84644 6682 84700 6692
rect 84644 5964 84700 5974
rect 84644 5740 84700 5908
rect 84644 5674 84700 5684
rect 84532 5338 84588 5348
rect 84644 5068 84700 5078
rect 84532 4956 84588 4966
rect 84308 4396 84364 4406
rect 84308 3612 84364 4340
rect 84308 3546 84364 3556
rect 84420 3836 84476 3846
rect 84420 3388 84476 3780
rect 84420 3322 84476 3332
rect 84028 3220 84252 3276
rect 83972 3210 84028 3220
rect 84084 2940 84140 2950
rect 83860 2874 83916 2884
rect 83972 2884 84084 2940
rect 83636 2762 83692 2772
rect 83636 2268 83692 2278
rect 83972 2268 84028 2884
rect 84084 2874 84140 2884
rect 83692 2212 84028 2268
rect 83636 2202 83692 2212
rect 83412 2090 83468 2100
rect 83188 1762 83244 1772
rect 84532 1468 84588 4900
rect 84644 4396 84700 5012
rect 84644 4330 84700 4340
rect 84644 3836 84700 3846
rect 84644 2604 84700 3780
rect 84644 2538 84700 2548
rect 84532 1402 84588 1412
rect 84756 1036 84812 7364
rect 84868 6148 84924 8932
rect 85092 8988 85148 8998
rect 85092 7980 85148 8932
rect 85428 8988 85484 9872
rect 85428 8922 85484 8932
rect 85540 9660 85596 9670
rect 85540 8316 85596 9604
rect 85540 8250 85596 8260
rect 85092 7914 85148 7924
rect 85652 7084 85708 12212
rect 85764 9212 85820 14552
rect 85764 9146 85820 9156
rect 85876 10108 85932 10118
rect 85876 7756 85932 10052
rect 85988 8652 86044 14912
rect 86548 12572 86604 12582
rect 86548 12268 86604 12516
rect 86660 12448 86716 14912
rect 102228 14968 102284 14978
rect 102452 14968 102508 14978
rect 102284 14912 102396 14968
rect 102228 14902 102284 14912
rect 98308 14812 98364 14822
rect 92596 14588 92652 14598
rect 87892 14248 87948 14258
rect 86996 13132 87052 13142
rect 86660 12382 86716 12392
rect 86884 12448 86940 12458
rect 86548 12202 86604 12212
rect 86100 11284 86716 11340
rect 86100 10108 86156 11284
rect 86548 11188 86604 11198
rect 86660 11188 86716 11284
rect 86772 11188 86828 11198
rect 86660 11132 86772 11188
rect 86212 10892 86268 10902
rect 86212 10828 86268 10836
rect 86436 10828 86492 10838
rect 86212 10762 86268 10772
rect 86324 10780 86436 10828
rect 86380 10772 86436 10780
rect 86436 10762 86492 10772
rect 86324 10714 86380 10724
rect 86100 10042 86156 10052
rect 85988 8586 86044 8596
rect 86436 8764 86492 8774
rect 85876 7690 85932 7700
rect 86100 7532 86156 7542
rect 85988 7084 86044 7094
rect 85652 7028 85988 7084
rect 85988 7018 86044 7028
rect 85876 6636 85932 6646
rect 85652 6508 85708 6518
rect 84980 6452 85596 6508
rect 84980 6300 85036 6452
rect 84980 6234 85036 6244
rect 85204 6188 85260 6198
rect 84868 6092 85036 6148
rect 84868 5068 84924 5078
rect 84868 2728 84924 5012
rect 84980 4956 85036 6092
rect 85204 5852 85260 6132
rect 85540 6148 85596 6452
rect 85652 6300 85708 6452
rect 85876 6508 85932 6580
rect 85876 6442 85932 6452
rect 85652 6234 85708 6244
rect 85540 6092 85820 6148
rect 85764 5964 85820 6092
rect 85764 5898 85820 5908
rect 85092 5788 85148 5798
rect 85204 5786 85260 5796
rect 85764 5788 85820 5798
rect 85092 5180 85148 5732
rect 85764 5180 85820 5732
rect 85092 5114 85148 5124
rect 85428 5124 85820 5180
rect 84980 4900 85260 4956
rect 84980 4732 85036 4900
rect 84980 4666 85036 4676
rect 84868 2662 84924 2672
rect 85092 3628 85148 3638
rect 85092 1036 85148 3572
rect 85204 2156 85260 4900
rect 85428 3988 85484 5124
rect 85764 4956 85820 4966
rect 86100 4956 86156 7476
rect 86436 6972 86492 8708
rect 86548 7084 86604 11132
rect 86772 11122 86828 11132
rect 86884 9324 86940 12392
rect 86884 9258 86940 9268
rect 86660 8540 86716 8550
rect 86660 7228 86716 8484
rect 86996 8540 87052 13076
rect 87668 12988 87724 12998
rect 87444 10468 87500 10478
rect 87668 10468 87724 12932
rect 87892 12988 87948 14192
rect 89236 14068 89292 14078
rect 89236 13528 89292 14012
rect 92372 14028 92428 14038
rect 89236 13462 89292 13472
rect 91252 13580 91308 13590
rect 87892 12922 87948 12932
rect 89012 13168 89068 13178
rect 89012 12236 89068 13112
rect 89012 12170 89068 12180
rect 89348 13168 89404 13178
rect 89012 12088 89068 12098
rect 89012 12012 89068 12032
rect 89236 12012 89292 12022
rect 89012 11956 89236 12012
rect 89236 11946 89292 11956
rect 89348 11788 89404 13112
rect 91252 13020 91308 13524
rect 92372 13528 92428 13972
rect 92596 14028 92652 14532
rect 92820 14588 92876 14598
rect 92820 14068 92876 14532
rect 98308 14588 98364 14756
rect 102340 14788 102396 14912
rect 138964 14968 139020 14978
rect 151732 14968 151788 14978
rect 102452 14858 102508 14868
rect 103012 14924 103068 14934
rect 115444 14924 115500 14934
rect 120932 14924 120988 14934
rect 102340 14732 102956 14788
rect 100660 14700 100716 14710
rect 98308 14522 98364 14532
rect 98532 14588 98588 14598
rect 92820 14002 92876 14012
rect 93044 14068 93100 14078
rect 92596 13962 92652 13972
rect 92484 13916 92540 13926
rect 92484 13692 92540 13860
rect 92484 13626 92540 13636
rect 92372 13462 92428 13472
rect 91252 12954 91308 12964
rect 92484 13168 92540 13178
rect 92708 13168 92764 13178
rect 91700 12796 91756 12806
rect 90916 12628 90972 12638
rect 89460 12448 89516 12458
rect 89460 12348 89516 12392
rect 89460 12282 89516 12292
rect 89908 12448 89964 12458
rect 88900 11732 89404 11788
rect 88564 11452 88620 11462
rect 88788 11452 88844 11462
rect 88620 11396 88732 11452
rect 88564 11386 88620 11396
rect 87500 10412 87612 10468
rect 87444 10402 87500 10412
rect 87220 8792 87500 8848
rect 86996 8474 87052 8484
rect 87108 8652 87164 8662
rect 86660 7162 86716 7172
rect 86772 8428 86828 8438
rect 86548 7028 86716 7084
rect 86324 6916 86492 6972
rect 86212 6860 86268 6870
rect 86324 6860 86380 6916
rect 86660 6860 86716 7028
rect 86324 6804 86492 6860
rect 86212 6747 86268 6804
rect 86212 6691 86380 6747
rect 85820 4900 86156 4956
rect 86212 5180 86268 5190
rect 85764 4890 85820 4900
rect 85876 4620 85932 4630
rect 85876 4528 85932 4564
rect 85876 4462 85932 4472
rect 86100 4528 86156 4538
rect 85316 3932 85484 3988
rect 85540 4284 85596 4294
rect 85316 3268 85372 3932
rect 85428 3836 85484 3846
rect 85540 3836 85596 4228
rect 85484 3780 85596 3836
rect 85428 3770 85484 3780
rect 86100 3268 86156 4472
rect 86212 3808 86268 5124
rect 86212 3742 86268 3752
rect 86324 3448 86380 6691
rect 86436 6188 86492 6804
rect 86660 6794 86716 6804
rect 86436 6122 86492 6132
rect 86548 6412 86604 6422
rect 86324 3382 86380 3392
rect 86548 3276 86604 6356
rect 86772 5428 86828 8372
rect 86884 7980 86940 7990
rect 86884 7532 86940 7924
rect 87108 7768 87164 8596
rect 87220 7980 87276 8792
rect 87220 7914 87276 7924
rect 87332 8652 87388 8662
rect 87108 7712 87276 7768
rect 86884 7466 86940 7476
rect 86884 6748 86940 6758
rect 87108 6748 87164 6758
rect 86940 6692 87052 6748
rect 86884 6682 86940 6692
rect 86996 5608 87052 6692
rect 87108 5740 87164 6692
rect 87220 5740 87276 7712
rect 87332 7756 87388 8596
rect 87444 8540 87500 8792
rect 87444 8474 87500 8484
rect 87332 7700 87500 7756
rect 87444 7420 87500 7700
rect 87556 7644 87612 10412
rect 87668 10402 87724 10412
rect 87892 11188 87948 11198
rect 87892 9996 87948 11132
rect 88676 10288 88732 11396
rect 88788 11188 88844 11396
rect 88788 11122 88844 11132
rect 88676 10222 88732 10232
rect 87892 9930 87948 9940
rect 88116 10108 88172 10118
rect 88116 9324 88172 10052
rect 88116 9258 88172 9268
rect 88676 8876 88732 8886
rect 88116 8820 88676 8848
rect 88116 8792 88732 8820
rect 88116 8764 88172 8792
rect 88116 8698 88172 8708
rect 88900 8668 88956 11732
rect 89124 9996 89180 10006
rect 89124 9436 89180 9940
rect 89124 9370 89180 9380
rect 89460 9436 89516 9446
rect 89348 9324 89404 9334
rect 88452 8612 88956 8668
rect 89236 9212 89292 9222
rect 88452 8128 88508 8612
rect 88452 8072 88956 8128
rect 87556 7588 87724 7644
rect 87668 7420 87724 7588
rect 87444 7364 87612 7420
rect 87668 7364 88396 7420
rect 87444 6972 87500 6982
rect 87332 5740 87388 5750
rect 87220 5684 87332 5740
rect 87108 5674 87164 5684
rect 87332 5674 87388 5684
rect 86996 5552 87388 5608
rect 86772 5372 87164 5428
rect 85316 3202 85372 3212
rect 85652 3212 86156 3268
rect 86212 3220 86604 3276
rect 86660 4060 86716 4070
rect 85428 3052 85484 3062
rect 85652 3052 85708 3212
rect 85484 2996 85708 3052
rect 86212 3052 86268 3220
rect 85428 2986 85484 2996
rect 86212 2986 86268 2996
rect 86436 3052 86492 3062
rect 85316 2548 85372 2558
rect 85316 2188 85372 2492
rect 85764 2268 85820 2278
rect 85316 2122 85372 2132
rect 85540 2188 85596 2198
rect 85204 2090 85260 2100
rect 85540 1932 85596 2132
rect 85540 1866 85596 1876
rect 85764 1932 85820 2212
rect 86324 2188 86380 2198
rect 86324 2090 86380 2100
rect 85764 1866 85820 1876
rect 86436 1468 86492 2996
rect 86548 2908 86604 2918
rect 86660 2908 86716 4004
rect 86772 2908 86828 2918
rect 86660 2852 86772 2908
rect 86548 2188 86604 2852
rect 86772 2842 86828 2852
rect 86548 2122 86604 2132
rect 86884 2492 86940 2502
rect 86436 1402 86492 1412
rect 85764 1036 85820 1046
rect 85092 980 85764 1036
rect 84756 970 84812 980
rect 85764 970 85820 980
rect 83076 858 83132 868
rect 83188 512 83692 568
rect 83188 476 83244 512
rect 82404 420 83244 476
rect 82180 322 82236 332
rect 83300 388 83356 402
rect 83524 364 83580 374
rect 83300 298 83356 308
rect 83412 308 83524 364
rect 83636 364 83692 512
rect 85988 364 86044 374
rect 83636 308 85988 364
rect 83412 208 83468 308
rect 83524 298 83580 308
rect 85988 298 86044 308
rect 86660 364 86716 374
rect 81956 152 83468 208
rect 86660 208 86716 308
rect 86884 364 86940 2436
rect 86996 1484 87052 1506
rect 86996 1402 87052 1412
rect 87108 1288 87164 5372
rect 87220 2268 87276 2278
rect 87332 2268 87388 5552
rect 87444 5180 87500 6916
rect 87556 6748 87612 7364
rect 88340 7228 88396 7364
rect 88340 7162 88396 7172
rect 88004 7084 88060 7094
rect 88004 6868 88060 7028
rect 87556 6682 87612 6692
rect 87668 6812 88060 6868
rect 88564 6972 88620 6982
rect 87444 5114 87500 5124
rect 87556 6188 87612 6198
rect 87444 4620 87500 4630
rect 87444 4348 87500 4564
rect 87444 4282 87500 4292
rect 87444 2268 87500 2278
rect 87332 2212 87444 2268
rect 87220 1484 87276 2212
rect 87444 2202 87500 2212
rect 87220 1418 87276 1428
rect 87556 1372 87612 6132
rect 87668 4396 87724 6812
rect 87892 5628 87948 5638
rect 88340 5628 88396 5638
rect 87948 5572 88340 5608
rect 87892 5552 88396 5572
rect 88116 4708 88172 4718
rect 87668 4330 87724 4340
rect 87892 4396 87948 4406
rect 87668 2940 87724 2950
rect 87668 2716 87724 2884
rect 87668 2650 87724 2660
rect 87556 1306 87612 1316
rect 86996 1260 87052 1270
rect 87108 1232 87388 1288
rect 86996 1108 87052 1204
rect 86996 1042 87052 1052
rect 87220 1148 87276 1158
rect 87108 1036 87164 1046
rect 87220 1042 87276 1052
rect 87108 388 87164 980
rect 87332 1036 87388 1232
rect 87332 970 87388 980
rect 87892 388 87948 4340
rect 88116 4348 88172 4652
rect 88116 4282 88172 4292
rect 88340 4708 88396 4718
rect 88340 4168 88396 4652
rect 88564 4348 88620 6916
rect 88900 6188 88956 8072
rect 88900 6122 88956 6132
rect 89236 5852 89292 9156
rect 89236 5786 89292 5796
rect 89348 7588 89404 9268
rect 89460 8316 89516 9380
rect 89460 8250 89516 8260
rect 89908 8316 89964 12392
rect 90580 12268 90636 12278
rect 90356 12236 90412 12246
rect 90356 10468 90412 12180
rect 90356 10402 90412 10412
rect 90580 10468 90636 12212
rect 90580 10402 90636 10412
rect 90692 11908 90748 11918
rect 90468 9884 90524 9894
rect 90244 9436 90300 9446
rect 90244 8876 90300 9380
rect 90468 9436 90524 9828
rect 90692 9884 90748 11852
rect 90692 9818 90748 9828
rect 90468 9370 90524 9380
rect 90916 8988 90972 12572
rect 91140 12628 91196 12638
rect 91140 11340 91196 12572
rect 91700 12572 91756 12740
rect 91700 12506 91756 12516
rect 92484 12268 92540 13112
rect 92484 12202 92540 12212
rect 92596 13112 92708 13168
rect 91812 12088 91868 12098
rect 91140 11274 91196 11284
rect 91252 11728 91308 11738
rect 91252 10220 91308 11672
rect 91476 11728 91532 11738
rect 91476 11368 91532 11672
rect 91476 11302 91532 11312
rect 91812 11368 91868 12032
rect 91812 11302 91868 11312
rect 92596 11004 92652 13112
rect 92708 13102 92764 13112
rect 92484 10948 92652 11004
rect 92708 11452 92764 11462
rect 92148 10892 92204 10902
rect 92036 10780 92092 10790
rect 92036 10468 92092 10724
rect 91924 10412 92092 10468
rect 91700 10220 91756 10230
rect 91252 10164 91700 10220
rect 91700 10154 91756 10164
rect 91028 9996 91084 10006
rect 91028 9772 91084 9940
rect 91924 9928 91980 10412
rect 91028 9706 91084 9716
rect 91588 9872 91980 9928
rect 90916 8922 90972 8932
rect 91476 9548 91532 9558
rect 90804 8876 90860 8886
rect 90244 8820 90804 8876
rect 90804 8810 90860 8820
rect 91476 8668 91532 9492
rect 89908 8250 89964 8260
rect 90356 8612 91532 8668
rect 90356 7588 90412 8612
rect 91364 8540 91420 8550
rect 90580 8484 91364 8540
rect 89348 7532 90412 7588
rect 90468 7868 90524 7878
rect 88676 4652 89068 4708
rect 88676 4528 88732 4652
rect 88676 4462 88732 4472
rect 88900 4528 88956 4538
rect 88900 4396 88956 4472
rect 88564 4292 88844 4348
rect 89012 4396 89068 4652
rect 89124 4396 89180 4406
rect 89012 4340 89124 4396
rect 88900 4330 88956 4340
rect 89124 4330 89180 4340
rect 88564 4168 88620 4178
rect 88340 4102 88396 4112
rect 88452 4112 88564 4168
rect 88340 3836 88396 3846
rect 88452 3836 88508 4112
rect 88564 4102 88620 4112
rect 88396 3780 88508 3836
rect 88340 3770 88396 3780
rect 88788 3387 88844 4292
rect 88564 3331 88844 3387
rect 88900 4060 88956 4070
rect 88900 3388 88956 4004
rect 89348 3836 89404 7532
rect 90244 7308 90300 7318
rect 90244 7084 90300 7252
rect 90244 7018 90300 7028
rect 89796 6076 89852 6086
rect 89796 5628 89852 6020
rect 90468 5740 90524 7812
rect 90580 6972 90636 8484
rect 91364 8474 91420 8484
rect 91252 8092 91308 8102
rect 91028 7980 91084 7990
rect 91028 7532 91084 7924
rect 91028 7466 91084 7476
rect 91252 7308 91308 8036
rect 90580 6906 90636 6916
rect 90692 7252 91308 7308
rect 91476 7420 91532 7430
rect 90692 6688 90748 7252
rect 91252 7084 91308 7094
rect 91252 6868 91308 7028
rect 91476 7084 91532 7364
rect 91588 7196 91644 9872
rect 92036 9548 92092 9558
rect 92036 9212 92092 9492
rect 92036 9146 92092 9156
rect 91700 8652 91756 8662
rect 91700 7756 91756 8596
rect 91700 7690 91756 7700
rect 91924 7980 91980 7990
rect 91812 7644 91868 7654
rect 91588 7130 91644 7140
rect 91700 7420 91756 7430
rect 91476 7018 91532 7028
rect 91252 6812 91644 6868
rect 90580 6636 90748 6688
rect 90636 6632 90748 6636
rect 90580 6570 90636 6580
rect 90692 6524 90748 6534
rect 90692 6188 90748 6468
rect 90692 6122 90748 6132
rect 91476 6300 91532 6310
rect 90468 5674 90524 5684
rect 89796 5562 89852 5572
rect 90020 5628 90076 5638
rect 90020 5068 90076 5572
rect 91476 5292 91532 6244
rect 91476 5226 91532 5236
rect 90020 5002 90076 5012
rect 90244 5068 90300 5078
rect 89348 3770 89404 3780
rect 89572 4508 89628 4518
rect 89572 3836 89628 4452
rect 89572 3770 89628 3780
rect 87108 332 87948 388
rect 88004 1484 88060 1494
rect 86884 298 86940 308
rect 88004 252 88060 1428
rect 88564 1260 88620 3331
rect 88900 3322 88956 3332
rect 89012 3500 89068 3510
rect 88788 2940 88844 2950
rect 88788 2380 88844 2884
rect 89012 2940 89068 3444
rect 89012 2874 89068 2884
rect 89236 3500 89292 3510
rect 88900 2828 88956 2838
rect 88900 2548 88956 2772
rect 88900 2482 88956 2492
rect 89124 2548 89180 2558
rect 89124 2380 89180 2492
rect 88788 2324 89180 2380
rect 88676 1820 88732 1830
rect 88676 1484 88732 1764
rect 89236 1820 89292 3444
rect 89684 3052 89740 3062
rect 89684 1932 89740 2996
rect 90244 2156 90300 5012
rect 90804 4732 90860 4742
rect 90804 3628 90860 4676
rect 91476 3628 91532 3638
rect 90804 3572 91476 3628
rect 91476 3562 91532 3572
rect 91588 3500 91644 6812
rect 91700 5628 91756 7364
rect 91812 6860 91868 7588
rect 91924 7196 91980 7924
rect 91924 7130 91980 7140
rect 91812 6794 91868 6804
rect 92148 5968 92204 10836
rect 92260 10828 92316 10838
rect 92260 9212 92316 10772
rect 92260 9146 92316 9156
rect 91700 5562 91756 5572
rect 91812 5912 92204 5968
rect 91700 5292 91756 5302
rect 91700 4956 91756 5236
rect 91700 4890 91756 4900
rect 91588 3434 91644 3444
rect 90580 3268 90636 3278
rect 90580 2492 90636 3212
rect 91252 2908 91308 2918
rect 91308 2852 91644 2908
rect 91252 2842 91308 2852
rect 90580 2426 90636 2436
rect 91028 2548 91084 2558
rect 90244 2090 90300 2100
rect 89684 1866 89740 1876
rect 89236 1754 89292 1764
rect 88676 1418 88732 1428
rect 90356 1596 90412 1606
rect 88564 1194 88620 1204
rect 90356 1260 90412 1540
rect 90356 1194 90412 1204
rect 90580 1596 90636 1606
rect 90580 1148 90636 1540
rect 90580 1082 90636 1092
rect 91028 1148 91084 2492
rect 91140 2188 91196 2198
rect 91140 2090 91196 2100
rect 91476 2188 91532 2198
rect 91476 1828 91532 2132
rect 91588 2008 91644 2852
rect 91812 2368 91868 5912
rect 92484 5788 92540 10948
rect 91924 5732 92540 5788
rect 92596 10828 92652 10838
rect 91924 5180 91980 5732
rect 92260 5628 92316 5638
rect 91924 5114 91980 5124
rect 92148 5572 92260 5628
rect 92148 4348 92204 5572
rect 92260 5562 92316 5572
rect 92596 5628 92652 10772
rect 92596 5562 92652 5572
rect 92372 5404 92428 5414
rect 92148 4282 92204 4292
rect 92260 5180 92316 5190
rect 92260 3988 92316 5124
rect 92372 4348 92428 5348
rect 92708 4620 92764 11396
rect 93044 9660 93100 14012
rect 97300 14028 97356 14038
rect 97076 13580 97132 13590
rect 94948 12684 95004 12694
rect 93044 9594 93100 9604
rect 94052 12088 94108 12098
rect 93268 8204 93324 8214
rect 93268 6524 93324 8148
rect 93268 6458 93324 6468
rect 92708 4554 92764 4564
rect 92372 4282 92428 4292
rect 92260 3922 92316 3932
rect 94052 3628 94108 12032
rect 94724 10468 94780 10478
rect 94500 10108 94556 10118
rect 94500 9928 94556 10052
rect 94500 9862 94556 9872
rect 94724 9928 94780 10412
rect 94948 10468 95004 12628
rect 96068 12684 96124 12694
rect 94948 10402 95004 10412
rect 95284 11900 95340 11910
rect 94724 9862 94780 9872
rect 95284 8540 95340 11844
rect 96068 11788 96124 12628
rect 96068 11722 96124 11732
rect 97076 11788 97132 13524
rect 97300 13580 97356 13972
rect 98532 13888 98588 14532
rect 98532 13822 98588 13832
rect 99876 13916 99932 13926
rect 97300 13514 97356 13524
rect 97636 12628 97692 12638
rect 97636 12460 97692 12572
rect 99876 12460 99932 13860
rect 100660 13888 100716 14644
rect 100660 13822 100716 13832
rect 102116 14608 102172 14618
rect 97636 12394 97692 12404
rect 98756 12448 98812 12458
rect 99876 12394 99932 12404
rect 102004 12684 102060 12694
rect 97076 11722 97132 11732
rect 97636 12236 97692 12246
rect 96740 11368 96796 11378
rect 95284 8474 95340 8484
rect 96068 10220 96124 10230
rect 95844 6524 95900 6534
rect 95732 5068 95788 5078
rect 95844 5068 95900 6468
rect 95956 5068 96012 5078
rect 95844 5012 95956 5068
rect 95732 4172 95788 5012
rect 95956 5002 96012 5012
rect 95732 4106 95788 4116
rect 94052 3562 94108 3572
rect 94276 3628 94332 3638
rect 92484 3500 92540 3510
rect 92372 3444 92484 3500
rect 91812 2302 91868 2312
rect 91924 3088 91980 3098
rect 91924 2156 91980 3032
rect 92372 2716 92428 3444
rect 92484 3434 92540 3444
rect 92372 2650 92428 2660
rect 92596 2716 92652 2726
rect 92596 2380 92652 2660
rect 91924 2090 91980 2100
rect 92036 2368 92092 2378
rect 92596 2314 92652 2324
rect 92036 2008 92092 2312
rect 91588 1952 92092 2008
rect 93940 2268 93996 2278
rect 91476 1762 91532 1772
rect 91700 1828 91756 1838
rect 91028 1082 91084 1092
rect 91700 476 91756 1772
rect 93940 1288 93996 2212
rect 94276 2044 94332 3572
rect 95620 3612 95676 3622
rect 95620 3268 95676 3556
rect 96068 3612 96124 10164
rect 96740 4284 96796 11312
rect 97524 11368 97580 11378
rect 96852 11116 96908 11126
rect 96852 10288 96908 11060
rect 96852 10232 97356 10288
rect 97300 10220 97356 10232
rect 97300 10154 97356 10164
rect 96964 8540 97020 8550
rect 96964 8092 97020 8484
rect 96964 8026 97020 8036
rect 96852 7980 96908 7990
rect 96908 7924 97020 7948
rect 96852 7892 97020 7924
rect 96740 4218 96796 4228
rect 96964 4060 97020 7892
rect 97300 4956 97356 4966
rect 97300 4708 97356 4900
rect 97188 4652 97356 4708
rect 97188 4620 97244 4652
rect 97188 4554 97244 4564
rect 97412 4620 97468 4630
rect 97412 4528 97468 4564
rect 97300 4472 97468 4528
rect 97300 4348 97356 4472
rect 97188 4292 97356 4348
rect 97188 4284 97244 4292
rect 97188 4218 97244 4228
rect 96964 3994 97020 4004
rect 97412 4060 97468 4070
rect 97412 3988 97468 4004
rect 97412 3922 97468 3932
rect 96068 3546 96124 3556
rect 95620 3202 95676 3212
rect 97524 2716 97580 11312
rect 97636 4060 97692 12180
rect 98084 12236 98140 12246
rect 97748 12012 97804 12022
rect 97748 9996 97804 11956
rect 97748 9930 97804 9940
rect 97860 10332 97916 10342
rect 97636 3994 97692 4004
rect 97748 7420 97804 7430
rect 97748 3724 97804 7364
rect 97748 3658 97804 3668
rect 97860 3088 97916 10276
rect 98084 4888 98140 12180
rect 98756 11908 98812 12392
rect 102004 12268 102060 12628
rect 102116 12460 102172 14552
rect 102340 14608 102396 14618
rect 102340 14068 102396 14552
rect 102788 14588 102844 14598
rect 102340 14002 102396 14012
rect 102564 14428 102620 14438
rect 102564 14068 102620 14372
rect 102564 14002 102620 14012
rect 102788 13692 102844 14532
rect 102788 13626 102844 13636
rect 102340 12808 102396 12818
rect 102340 12684 102396 12752
rect 102564 12808 102620 12818
rect 102564 12714 102620 12740
rect 102788 12796 102844 12806
rect 102116 12394 102172 12404
rect 102228 12628 102284 12638
rect 102340 12618 102396 12628
rect 102452 12628 102508 12638
rect 99092 12236 99148 12246
rect 102004 12212 102172 12268
rect 98980 12124 99036 12134
rect 98756 11842 98812 11852
rect 98868 11900 98924 11910
rect 98532 10892 98588 10902
rect 98532 6508 98588 10836
rect 98868 10220 98924 11844
rect 98980 11908 99036 12068
rect 98980 11842 99036 11852
rect 99092 11452 99148 12180
rect 100436 11788 100492 11798
rect 100436 11728 100492 11732
rect 100436 11662 100492 11672
rect 99988 11548 100044 11558
rect 101108 11548 101164 11558
rect 99092 11386 99148 11396
rect 99316 11452 99372 11462
rect 98868 10154 98924 10164
rect 99092 10220 99148 10230
rect 98644 9324 98700 9334
rect 99092 9324 99148 10164
rect 99316 9772 99372 11396
rect 99316 9706 99372 9716
rect 99876 9772 99932 9782
rect 98700 9268 99148 9324
rect 99652 9436 99708 9446
rect 98644 9258 98700 9268
rect 98644 8596 99596 8652
rect 98644 8204 98700 8596
rect 99204 8428 99260 8438
rect 99204 8316 99260 8372
rect 98980 8260 99260 8316
rect 98644 8138 98700 8148
rect 98868 8204 98924 8214
rect 98532 6452 98700 6508
rect 98196 6412 98252 6422
rect 98196 6328 98252 6356
rect 98196 6272 98588 6328
rect 98532 6188 98588 6272
rect 98532 6122 98588 6132
rect 98196 5740 98252 5750
rect 98196 5516 98252 5684
rect 98196 5450 98252 5460
rect 98420 5740 98476 5750
rect 98084 4822 98140 4832
rect 97860 3022 97916 3032
rect 98084 3612 98140 3622
rect 98084 3088 98140 3556
rect 98420 3387 98476 5684
rect 98644 4732 98700 6452
rect 98868 5068 98924 8148
rect 98980 5740 99036 8260
rect 99428 7420 99484 7430
rect 99428 5964 99484 7364
rect 99540 6972 99596 8596
rect 99540 6906 99596 6916
rect 99428 5898 99484 5908
rect 98980 5674 99036 5684
rect 99204 5788 99260 5798
rect 98868 5002 98924 5012
rect 98644 4666 98700 4676
rect 98868 4888 98924 4898
rect 98084 3022 98140 3032
rect 98196 3331 98476 3387
rect 98868 3448 98924 4832
rect 99204 4732 99260 5732
rect 99428 5788 99484 5798
rect 99428 5516 99484 5732
rect 99428 5450 99484 5460
rect 99652 5292 99708 9380
rect 99876 7532 99932 9716
rect 99988 9436 100044 11492
rect 100772 11492 101108 11548
rect 100772 11008 100828 11492
rect 101108 11482 101164 11492
rect 101556 11368 101612 11378
rect 100548 10952 100828 11008
rect 101444 11312 101556 11368
rect 100548 10892 100604 10952
rect 101444 10892 101500 11312
rect 101556 11302 101612 11312
rect 100548 10826 100604 10836
rect 100660 10828 100716 10838
rect 101108 10828 101164 10838
rect 101444 10836 101612 10892
rect 100716 10772 101052 10828
rect 100660 10762 100716 10772
rect 100660 10668 100716 10678
rect 99988 9370 100044 9380
rect 100100 10220 100156 10230
rect 99876 7466 99932 7476
rect 100100 6188 100156 10164
rect 100660 9548 100716 10612
rect 100660 9482 100716 9492
rect 100660 9324 100716 9334
rect 100660 9208 100716 9268
rect 100660 9152 100828 9208
rect 100436 8540 100492 8550
rect 100436 8428 100492 8484
rect 100436 8362 100492 8372
rect 100660 8428 100716 8438
rect 100660 7228 100716 8372
rect 100436 7196 100492 7206
rect 100660 7162 100716 7172
rect 100100 6122 100156 6132
rect 100324 6972 100380 6982
rect 99652 5236 99820 5292
rect 99204 4666 99260 4676
rect 99428 4168 99484 4178
rect 98868 3382 98924 3392
rect 99092 3612 99148 3622
rect 99092 3448 99148 3556
rect 99092 3382 99148 3392
rect 97524 2650 97580 2660
rect 95620 2548 95676 2558
rect 95620 2268 95676 2492
rect 95620 2202 95676 2212
rect 96292 2492 96348 2502
rect 94388 2156 94444 2166
rect 94388 2044 94444 2100
rect 96292 2156 96348 2436
rect 96292 2090 96348 2100
rect 96516 2368 96572 2378
rect 96516 2156 96572 2312
rect 98196 2268 98252 3331
rect 99316 2604 99372 2614
rect 99316 2368 99372 2548
rect 99316 2302 99372 2312
rect 98196 2202 98252 2212
rect 98868 2188 98924 2198
rect 98924 2132 99036 2188
rect 98868 2122 98924 2132
rect 96516 2090 96572 2100
rect 94500 2044 94556 2054
rect 94388 1988 94500 2044
rect 94276 1978 94332 1988
rect 94500 1978 94556 1988
rect 94052 1820 94108 1830
rect 94052 1288 94108 1764
rect 93940 1232 94108 1288
rect 97748 1648 97804 1658
rect 94052 1148 94108 1158
rect 94052 928 94108 1092
rect 94052 862 94108 872
rect 97300 1108 97356 1118
rect 91700 410 91756 420
rect 97300 476 97356 1052
rect 97524 1108 97580 1118
rect 97524 1036 97580 1052
rect 97524 970 97580 980
rect 97748 1036 97804 1592
rect 98980 1648 99036 2132
rect 98980 1582 99036 1592
rect 97748 970 97804 980
rect 99204 1372 99260 1382
rect 97300 410 97356 420
rect 97412 928 97468 938
rect 97412 476 97468 872
rect 97412 410 97468 420
rect 99204 364 99260 1316
rect 99428 1372 99484 4112
rect 99652 4168 99708 4178
rect 99652 3628 99708 4112
rect 99764 3724 99820 5236
rect 99764 3658 99820 3668
rect 99652 3562 99708 3572
rect 100212 3276 100268 3286
rect 99988 2908 100044 2918
rect 99988 2604 100044 2852
rect 100212 2908 100268 3220
rect 100212 2842 100268 2852
rect 99988 2538 100044 2548
rect 99764 2492 99820 2502
rect 99428 1306 99484 1316
rect 99652 1820 99708 1830
rect 99204 298 99260 308
rect 86996 208 88060 252
rect 86660 196 88060 208
rect 99652 252 99708 1764
rect 99764 1708 99820 2436
rect 99764 1642 99820 1652
rect 100324 928 100380 6916
rect 100436 3808 100492 7140
rect 100660 6508 100716 6518
rect 100660 5964 100716 6452
rect 100660 5898 100716 5908
rect 100772 5740 100828 9152
rect 100996 7196 101052 10772
rect 100996 7130 101052 7140
rect 101556 10828 101612 10836
rect 101108 6688 101164 10772
rect 101220 10780 101276 10790
rect 101556 10772 101668 10828
rect 101220 9324 101276 10724
rect 101612 10332 101668 10772
rect 101220 9258 101276 9268
rect 101556 10276 101668 10332
rect 101780 10780 101836 10790
rect 100772 5674 100828 5684
rect 100884 6632 101164 6688
rect 101220 8092 101276 8102
rect 100548 5068 100604 5078
rect 100548 4396 100604 5012
rect 100548 4330 100604 4340
rect 100772 5068 100828 5078
rect 100772 3988 100828 5012
rect 100660 3948 100828 3988
rect 100716 3932 100828 3948
rect 100660 3882 100716 3892
rect 100436 3752 100604 3808
rect 100436 2716 100492 2726
rect 100436 1036 100492 2660
rect 100436 970 100492 980
rect 100324 862 100380 872
rect 100548 928 100604 3752
rect 100884 3387 100940 6632
rect 101108 6524 101164 6546
rect 101108 6442 101164 6452
rect 101220 5292 101276 8036
rect 101444 8092 101500 8102
rect 101220 5226 101276 5236
rect 101332 6524 101388 6534
rect 101220 4396 101276 4406
rect 101332 4396 101388 6468
rect 101444 5516 101500 8036
rect 101444 5450 101500 5460
rect 101276 4340 101388 4396
rect 101220 4330 101276 4340
rect 101444 3724 101500 3734
rect 100660 3331 100940 3387
rect 100996 3628 101052 3638
rect 100660 3164 100716 3331
rect 100660 3098 100716 3108
rect 100996 3052 101052 3572
rect 101332 3388 101388 3398
rect 100996 2986 101052 2996
rect 101220 3164 101276 3174
rect 100772 2604 100828 2614
rect 100772 1036 100828 2548
rect 101220 1372 101276 3108
rect 101332 2044 101388 3332
rect 101444 2716 101500 3668
rect 101444 2650 101500 2660
rect 101556 2268 101612 10276
rect 101780 10220 101836 10724
rect 101668 10164 101836 10220
rect 101892 10468 101948 10478
rect 101668 7228 101724 10164
rect 101892 9548 101948 10412
rect 101892 9482 101948 9492
rect 101668 7162 101724 7172
rect 102004 7196 102060 7206
rect 101668 5788 101724 5798
rect 101668 5516 101724 5732
rect 102004 5788 102060 7140
rect 102116 5852 102172 12212
rect 102228 10892 102284 12572
rect 102788 12572 102844 12740
rect 102452 12088 102508 12572
rect 102564 12516 102844 12572
rect 102564 12236 102620 12516
rect 102564 12170 102620 12180
rect 102788 12448 102844 12458
rect 102452 12032 102620 12088
rect 102564 11728 102620 12032
rect 102228 10826 102284 10836
rect 102340 11676 102396 11686
rect 102340 10648 102396 11620
rect 102228 10592 102396 10648
rect 102452 11672 102620 11728
rect 102228 8092 102284 10592
rect 102228 8026 102284 8036
rect 102340 10468 102396 10478
rect 102340 7420 102396 10412
rect 102452 10108 102508 11672
rect 102564 11548 102620 11558
rect 102564 10108 102620 11492
rect 102676 11340 102732 11350
rect 102676 11116 102732 11284
rect 102676 11050 102732 11060
rect 102676 10108 102732 10118
rect 102564 10052 102676 10108
rect 102452 10042 102508 10052
rect 102676 10042 102732 10052
rect 102788 9928 102844 12392
rect 102900 11548 102956 14732
rect 103012 14428 103068 14868
rect 114324 14868 115444 14924
rect 111412 14812 111468 14822
rect 103012 14362 103068 14372
rect 103908 14700 103964 14710
rect 103348 14252 103404 14262
rect 103404 14196 103852 14252
rect 103348 14186 103404 14196
rect 103796 13580 103852 14196
rect 103796 13514 103852 13524
rect 103236 13356 103292 13366
rect 103908 13348 103964 14644
rect 109172 14608 109228 14618
rect 109228 14552 109452 14608
rect 109172 14542 109228 14552
rect 103012 13132 103068 13142
rect 103012 12236 103068 13076
rect 103236 13020 103292 13300
rect 103684 13292 103964 13348
rect 104692 14428 104748 14438
rect 103236 12954 103292 12964
rect 103572 13020 103628 13030
rect 103012 12170 103068 12180
rect 103236 12448 103292 12458
rect 103236 12088 103292 12392
rect 103460 12088 103516 12098
rect 103236 12022 103292 12032
rect 103348 12032 103460 12088
rect 103348 11788 103404 12032
rect 103460 12022 103516 12032
rect 103012 11732 103404 11788
rect 103012 11676 103068 11732
rect 103012 11610 103068 11620
rect 103460 11728 103516 11738
rect 103460 11564 103516 11672
rect 103460 11498 103516 11508
rect 102900 11482 102956 11492
rect 103572 11340 103628 12964
rect 103684 12908 103740 13292
rect 104132 13020 104188 13030
rect 104188 12964 104412 13020
rect 104132 12954 104188 12964
rect 103684 12842 103740 12852
rect 103908 12908 103964 12918
rect 103908 12808 103964 12852
rect 103908 12742 103964 12752
rect 104244 12808 104300 12818
rect 103572 11274 103628 11284
rect 103908 12348 103964 12358
rect 103908 11188 103964 12292
rect 104244 12088 104300 12752
rect 103012 11132 103964 11188
rect 104020 12032 104300 12088
rect 103012 11004 103068 11132
rect 103012 10938 103068 10948
rect 103236 11004 103292 11014
rect 104020 11004 104076 12032
rect 104244 11900 104300 11910
rect 104132 11228 104188 11238
rect 104132 11122 104188 11132
rect 103236 10828 103292 10948
rect 103012 10772 103292 10828
rect 103348 10948 104076 11004
rect 103012 10220 103068 10772
rect 103124 10444 103180 10454
rect 103124 10220 103180 10388
rect 103236 10220 103292 10230
rect 103124 10164 103236 10220
rect 103012 10154 103068 10164
rect 103236 10154 103292 10164
rect 102676 9872 102844 9928
rect 102452 9548 102508 9558
rect 102452 8652 102508 9492
rect 102452 8586 102508 8596
rect 102676 8652 102732 9872
rect 102788 9772 102844 9782
rect 103348 9772 103404 10948
rect 103684 10780 103740 10790
rect 102844 9716 103404 9772
rect 103572 10332 103628 10342
rect 102788 9706 102844 9716
rect 103012 9100 103068 9110
rect 103068 9044 103404 9100
rect 103012 9034 103068 9044
rect 102676 8586 102732 8596
rect 102340 7354 102396 7364
rect 102900 7868 102956 7878
rect 102116 5786 102172 5796
rect 102228 7196 102284 7206
rect 102004 5722 102060 5732
rect 101668 5450 101724 5460
rect 102228 4888 102284 7140
rect 102340 6636 102396 6646
rect 102340 5516 102396 6580
rect 102340 5450 102396 5460
rect 102228 4822 102284 4832
rect 102788 4844 102844 4854
rect 102116 4620 102172 4630
rect 101668 3724 101724 3734
rect 101668 2492 101724 3668
rect 102116 3612 102172 4564
rect 102340 4472 102732 4528
rect 102340 4284 102396 4472
rect 102564 4284 102620 4294
rect 102340 4218 102396 4228
rect 102452 4228 102564 4284
rect 102452 3612 102508 4228
rect 102564 4218 102620 4228
rect 102116 3546 102172 3556
rect 102228 3556 102508 3612
rect 102676 3612 102732 4472
rect 102228 2828 102284 3556
rect 102676 3546 102732 3556
rect 102564 3500 102620 3510
rect 102620 3444 102732 3448
rect 102564 3392 102732 3444
rect 102340 3268 102396 3278
rect 102340 3052 102396 3212
rect 102564 3268 102620 3278
rect 102340 2986 102396 2996
rect 102452 3164 102508 3174
rect 102228 2762 102284 2772
rect 102452 2604 102508 3108
rect 102564 2908 102620 3212
rect 102676 3276 102732 3392
rect 102676 3210 102732 3220
rect 102564 2842 102620 2852
rect 102788 2908 102844 4788
rect 102900 3164 102956 7812
rect 103012 7228 103068 7238
rect 103012 6412 103068 7172
rect 103236 7228 103292 7238
rect 103236 6748 103292 7172
rect 103348 7196 103404 9044
rect 103460 8876 103516 8886
rect 103460 7532 103516 8820
rect 103460 7466 103516 7476
rect 103348 7130 103404 7140
rect 103236 6682 103292 6692
rect 103124 6636 103180 6646
rect 103572 6636 103628 10276
rect 103684 9996 103740 10724
rect 104244 10332 104300 11844
rect 104356 11728 104412 12964
rect 104692 12908 104748 14372
rect 109284 14428 109340 14438
rect 109396 14428 109452 14552
rect 109620 14428 109676 14438
rect 109396 14372 109620 14428
rect 104692 12842 104748 12852
rect 108612 13168 108668 13178
rect 104356 11662 104412 11672
rect 104468 12348 104524 12358
rect 104244 10266 104300 10276
rect 103684 9930 103740 9940
rect 104244 9772 104300 9782
rect 103124 6524 103180 6580
rect 103348 6580 103628 6636
rect 103684 8540 103740 8550
rect 103348 6524 103404 6580
rect 103124 6468 103404 6524
rect 103572 6412 103628 6422
rect 103012 6356 103572 6412
rect 103572 6346 103628 6356
rect 103236 5852 103292 5862
rect 103012 5292 103068 5302
rect 103012 4844 103068 5236
rect 103236 5292 103292 5796
rect 103236 5226 103292 5236
rect 103012 4778 103068 4788
rect 103684 4168 103740 8484
rect 104132 8316 104188 8326
rect 104132 7868 104188 8260
rect 104132 7802 104188 7812
rect 103796 7420 103852 7430
rect 103796 7084 103852 7364
rect 103908 7196 103964 7206
rect 103964 7140 104188 7196
rect 103908 7130 103964 7140
rect 103796 7018 103852 7028
rect 102900 3098 102956 3108
rect 103348 4112 103740 4168
rect 103908 4708 103964 4718
rect 102788 2842 102844 2852
rect 103348 2604 103404 4112
rect 103684 3988 103740 3998
rect 103460 3948 103516 3958
rect 103460 3612 103516 3892
rect 103460 3546 103516 3556
rect 102452 2548 103180 2604
rect 101668 2426 101724 2436
rect 103124 2380 103180 2548
rect 103460 2728 103516 2738
rect 103460 2604 103516 2672
rect 103684 2728 103740 3932
rect 103684 2662 103740 2672
rect 103796 3948 103852 3958
rect 103796 2604 103852 3892
rect 103460 2548 103852 2604
rect 103348 2538 103404 2548
rect 103348 2380 103404 2390
rect 103124 2324 103348 2380
rect 103348 2314 103404 2324
rect 103908 2368 103964 4652
rect 104132 4168 104188 7140
rect 104132 4102 104188 4112
rect 104132 2940 104188 2950
rect 103908 2302 103964 2312
rect 104020 2548 104076 2558
rect 101556 2202 101612 2212
rect 102900 2268 102956 2278
rect 101332 1978 101388 1988
rect 101556 2044 101612 2054
rect 101220 1306 101276 1316
rect 101556 1108 101612 1988
rect 102228 1828 102284 1838
rect 101556 1042 101612 1052
rect 101780 1108 101836 1118
rect 100772 970 100828 980
rect 100548 476 100604 872
rect 101780 748 101836 1052
rect 101780 682 101836 692
rect 102004 748 102060 758
rect 100772 476 100828 486
rect 100548 410 100604 420
rect 100660 420 100772 476
rect 100660 252 100716 420
rect 100772 410 100828 420
rect 102004 476 102060 692
rect 102004 410 102060 420
rect 102228 476 102284 1772
rect 102452 1828 102508 1838
rect 102452 1596 102508 1772
rect 102788 1820 102844 1830
rect 102900 1820 102956 2212
rect 102844 1764 102956 1820
rect 102788 1754 102844 1764
rect 102452 1530 102508 1540
rect 104020 1596 104076 2492
rect 104132 2368 104188 2884
rect 104132 2302 104188 2312
rect 104244 2268 104300 9716
rect 104468 5852 104524 12292
rect 106148 12124 106204 12134
rect 105924 11908 105980 11918
rect 105476 11852 105924 11908
rect 105476 11728 105532 11852
rect 105924 11842 105980 11852
rect 106148 11788 106204 12068
rect 106148 11722 106204 11732
rect 106708 12088 106764 12098
rect 105476 11662 105532 11672
rect 106260 11548 106316 11558
rect 104580 11368 104636 11378
rect 104580 10108 104636 11312
rect 104804 11340 104860 11350
rect 104580 10042 104636 10052
rect 104692 10780 104748 10790
rect 104580 9436 104636 9446
rect 104580 8540 104636 9380
rect 104580 8474 104636 8484
rect 104692 6524 104748 10724
rect 104804 8092 104860 11284
rect 104804 8026 104860 8036
rect 105028 11340 105084 11350
rect 104692 6458 104748 6468
rect 104468 5786 104524 5796
rect 105028 3948 105084 11284
rect 106036 10828 106092 10838
rect 105924 10556 105980 10566
rect 105812 10108 105868 10118
rect 105812 10014 105868 10052
rect 105924 9772 105980 10500
rect 106036 10108 106092 10772
rect 106260 10828 106316 11492
rect 106708 11368 106764 12032
rect 106708 11302 106764 11312
rect 106932 12088 106988 12098
rect 106260 10762 106316 10772
rect 106036 10042 106092 10052
rect 106708 10556 106764 10566
rect 106484 9996 106540 10006
rect 106148 9940 106484 9996
rect 106036 9884 106092 9894
rect 106148 9884 106204 9940
rect 106484 9930 106540 9940
rect 106092 9828 106204 9884
rect 106036 9818 106092 9828
rect 105924 9706 105980 9716
rect 106596 8876 106652 8886
rect 106372 8652 106428 8662
rect 106148 7644 106204 7654
rect 105140 7532 105196 7542
rect 105140 6972 105196 7476
rect 105140 6906 105196 6916
rect 105700 7308 105756 7318
rect 105700 6524 105756 7252
rect 106148 7308 106204 7588
rect 106372 7644 106428 8596
rect 106596 8652 106652 8820
rect 106596 8586 106652 8596
rect 106372 7578 106428 7588
rect 106148 7242 106204 7252
rect 105700 6458 105756 6468
rect 105028 3882 105084 3892
rect 105700 4528 105756 4538
rect 104468 3388 104524 3398
rect 104356 2940 104412 2950
rect 104356 2716 104412 2884
rect 104356 2650 104412 2660
rect 104244 2202 104300 2212
rect 104468 2268 104524 3332
rect 105700 3276 105756 4472
rect 105924 4528 105980 4538
rect 105924 4168 105980 4472
rect 105924 4102 105980 4112
rect 106148 4168 106204 4178
rect 105700 3210 105756 3220
rect 106148 3088 106204 4112
rect 106148 3022 106204 3032
rect 106596 2716 106652 2726
rect 104468 2202 104524 2212
rect 106148 2548 106204 2558
rect 104020 1530 104076 1540
rect 106036 1260 106092 1270
rect 102228 410 102284 420
rect 103236 1148 103292 1158
rect 99652 196 100716 252
rect 103012 364 103068 374
rect 103012 208 103068 308
rect 103236 364 103292 1092
rect 103684 1036 103740 1046
rect 103236 298 103292 308
rect 103348 980 103684 1036
rect 103348 208 103404 980
rect 103684 970 103740 980
rect 106036 748 106092 1204
rect 106148 1036 106204 2492
rect 106596 2492 106652 2660
rect 106596 2426 106652 2436
rect 106708 2188 106764 10500
rect 106932 6972 106988 12032
rect 107492 11900 107548 11910
rect 107492 9660 107548 11844
rect 108612 11788 108668 13112
rect 108836 13168 108892 13178
rect 108836 12808 108892 13112
rect 108836 12742 108892 12752
rect 109171 12808 109227 12818
rect 109171 12684 109227 12752
rect 108724 12628 109227 12684
rect 108724 12012 108780 12628
rect 109284 12448 109340 14372
rect 109620 14362 109676 14372
rect 109620 13020 109676 13030
rect 109171 12348 109228 12448
rect 109284 12382 109340 12392
rect 109396 12964 109620 13020
rect 108724 11946 108780 11956
rect 108836 12292 109228 12348
rect 108836 11788 108892 12292
rect 108948 12012 109004 12022
rect 108948 11908 109004 11956
rect 108948 11842 109004 11852
rect 108612 11732 108892 11788
rect 107940 11564 107996 11574
rect 107492 9594 107548 9604
rect 107716 10892 107772 10902
rect 107492 8876 107548 8886
rect 107492 7980 107548 8820
rect 107492 7914 107548 7924
rect 107716 7980 107772 10836
rect 107940 10892 107996 11508
rect 107940 10826 107996 10836
rect 109060 11564 109116 11574
rect 107716 7914 107772 7924
rect 108388 10668 108444 10678
rect 106932 6906 106988 6916
rect 108276 7868 108332 7878
rect 108276 6636 108332 7812
rect 108276 6570 108332 6580
rect 107380 5372 107772 5428
rect 107380 5292 107436 5372
rect 107380 5226 107436 5236
rect 107604 5292 107660 5302
rect 107492 4732 107548 4742
rect 107380 3276 107436 3286
rect 107380 3088 107436 3220
rect 107380 3022 107436 3032
rect 106708 2122 106764 2132
rect 107492 2008 107548 4676
rect 107604 3988 107660 5236
rect 107716 4732 107772 5372
rect 107716 4666 107772 4676
rect 107604 3922 107660 3932
rect 107716 3448 107772 3458
rect 107716 3276 107772 3392
rect 107940 3448 107996 3458
rect 107940 3276 107996 3392
rect 107716 3220 107996 3276
rect 108388 2604 108444 10612
rect 109060 9436 109116 11508
rect 109060 9370 109116 9380
rect 109172 8652 109228 12292
rect 109396 12236 109452 12964
rect 109620 12954 109676 12964
rect 110740 12628 110796 12638
rect 109396 12170 109452 12180
rect 109620 12448 109676 12458
rect 109172 8586 109228 8596
rect 109284 12012 109340 12022
rect 108612 8540 108668 8550
rect 108612 8204 108668 8484
rect 108612 8138 108668 8148
rect 109284 7532 109340 11956
rect 109396 11908 109452 11918
rect 109396 9436 109452 11852
rect 109396 9370 109452 9380
rect 109508 11340 109564 11350
rect 109060 7476 109340 7532
rect 109060 4732 109116 7476
rect 109396 6972 109452 6982
rect 109396 5788 109452 6916
rect 109508 6860 109564 11284
rect 109508 6794 109564 6804
rect 109620 6300 109676 12392
rect 110404 11728 110460 11738
rect 110740 11728 110796 12572
rect 110964 12628 111020 12638
rect 110740 11672 110908 11728
rect 109620 6234 109676 6244
rect 109840 9436 110160 10252
rect 110404 9996 110460 11672
rect 110404 9930 110460 9940
rect 109840 9380 109868 9436
rect 109924 9380 109972 9436
rect 110028 9380 110076 9436
rect 110132 9380 110160 9436
rect 109840 9030 110160 9380
rect 110852 9436 110908 11672
rect 110964 11564 111020 12572
rect 110964 11498 111020 11508
rect 111076 11340 111132 11350
rect 110852 9370 110908 9380
rect 110964 10332 111020 10342
rect 110740 9212 110796 9222
rect 109840 8974 109868 9030
rect 109924 8974 109972 9030
rect 110028 8974 110076 9030
rect 110132 8974 110160 9030
rect 109840 8926 110160 8974
rect 110404 9100 110460 9110
rect 110404 9028 110460 9044
rect 110404 8972 110572 9028
rect 109840 8870 109868 8926
rect 109924 8870 109972 8926
rect 110028 8870 110076 8926
rect 110132 8870 110160 8926
rect 109840 8822 110160 8870
rect 109840 8766 109868 8822
rect 109924 8766 109972 8822
rect 110028 8766 110076 8822
rect 110132 8766 110160 8822
rect 109840 7868 110160 8766
rect 109840 7812 109868 7868
rect 109924 7812 109972 7868
rect 110028 7812 110076 7868
rect 110132 7812 110160 7868
rect 109840 7632 110160 7812
rect 109840 7576 109868 7632
rect 109924 7576 109972 7632
rect 110028 7576 110076 7632
rect 110132 7576 110160 7632
rect 109840 7528 110160 7576
rect 109840 7472 109868 7528
rect 109924 7472 109972 7528
rect 110028 7472 110076 7528
rect 110132 7472 110160 7528
rect 109840 7424 110160 7472
rect 109840 7368 109868 7424
rect 109924 7368 109972 7424
rect 110028 7368 110076 7424
rect 110132 7368 110160 7424
rect 109840 6300 110160 7368
rect 110404 8316 110460 8326
rect 109840 6244 109868 6300
rect 109924 6244 109972 6300
rect 110028 6244 110076 6300
rect 110132 6244 110160 6300
rect 109840 6234 110160 6244
rect 109840 6178 109868 6234
rect 109924 6178 109972 6234
rect 110028 6178 110076 6234
rect 110132 6178 110160 6234
rect 109840 6130 110160 6178
rect 109840 6074 109868 6130
rect 109924 6074 109972 6130
rect 110028 6074 110076 6130
rect 110132 6074 110160 6130
rect 109840 6026 110160 6074
rect 109620 5964 109676 5974
rect 109396 5722 109452 5732
rect 109508 5908 109620 5964
rect 109508 5628 109564 5908
rect 109620 5898 109676 5908
rect 109840 5970 109868 6026
rect 109924 5970 109972 6026
rect 110028 5970 110076 6026
rect 110132 5970 110160 6026
rect 109508 5562 109564 5572
rect 109620 5788 109676 5798
rect 109060 4676 109228 4732
rect 108724 4620 108780 4630
rect 108780 4564 109116 4620
rect 108724 4554 108780 4564
rect 108948 3836 109004 3846
rect 109060 3836 109116 4564
rect 109172 4060 109228 4676
rect 109620 4708 109676 5732
rect 109620 4642 109676 4652
rect 109840 4732 110160 5970
rect 110292 6636 110348 6646
rect 110292 5516 110348 6580
rect 110292 5450 110348 5460
rect 109840 4676 109868 4732
rect 109924 4676 109972 4732
rect 110028 4676 110076 4732
rect 110132 4676 110160 4732
rect 109840 4644 110160 4676
rect 109732 4528 109788 4538
rect 109284 4348 109340 4358
rect 109340 4292 109452 4348
rect 109284 4282 109340 4292
rect 109172 3994 109228 4004
rect 109396 3988 109452 4292
rect 109396 3922 109452 3932
rect 109172 3836 109228 3846
rect 109060 3780 109172 3836
rect 108948 3276 109004 3780
rect 109172 3770 109228 3780
rect 109284 3276 109340 3286
rect 108948 3220 109284 3276
rect 109284 3210 109340 3220
rect 109620 3052 109676 3062
rect 108724 2940 108780 2950
rect 108388 2538 108444 2548
rect 108500 2548 108556 2558
rect 108500 2044 108556 2492
rect 108724 2368 108780 2884
rect 109620 2828 109676 2996
rect 109620 2762 109676 2772
rect 109171 2380 109227 2390
rect 108724 2324 109171 2368
rect 108724 2312 109227 2324
rect 108836 2188 108892 2198
rect 108724 2132 108836 2188
rect 108724 2044 108780 2132
rect 108836 2122 108892 2132
rect 107492 1952 107996 2008
rect 108500 1988 108780 2044
rect 109732 2044 109788 4472
rect 110292 4060 110348 4070
rect 110292 3808 110348 4004
rect 110292 3742 110348 3752
rect 110404 3388 110460 8260
rect 110516 4396 110572 8972
rect 110740 8316 110796 9156
rect 110740 8250 110796 8260
rect 110852 9100 110908 9110
rect 110852 7084 110908 9044
rect 110852 7018 110908 7028
rect 110740 4396 110796 4406
rect 110516 4340 110740 4396
rect 110740 4330 110796 4340
rect 110628 3808 110684 3818
rect 110628 3724 110684 3752
rect 110628 3658 110684 3668
rect 110852 3724 110908 3734
rect 110404 3322 110460 3332
rect 110852 3268 110908 3668
rect 110628 3212 110908 3268
rect 110404 3052 110460 3062
rect 110404 2548 110460 2996
rect 110628 2728 110684 3212
rect 110740 3052 110796 3062
rect 110740 2908 110796 2996
rect 110964 3052 111020 10276
rect 111076 8092 111132 11284
rect 111188 9884 111244 9894
rect 111188 9548 111244 9828
rect 111188 9482 111244 9492
rect 111076 8026 111132 8036
rect 111300 8092 111356 8102
rect 111300 6860 111356 8036
rect 111300 6794 111356 6804
rect 110964 2986 111020 2996
rect 110740 2852 111244 2908
rect 110628 2672 110908 2728
rect 110404 2482 110460 2492
rect 109732 1978 109788 1988
rect 107604 1288 107660 1298
rect 106148 970 106204 980
rect 106372 1036 106428 1046
rect 106372 928 106428 980
rect 106372 862 106428 872
rect 107492 928 107548 938
rect 107492 812 107548 872
rect 107492 746 107548 756
rect 107604 748 107660 1232
rect 106036 682 106092 692
rect 107604 682 107660 692
rect 107940 700 107996 1952
rect 108836 1596 108892 1606
rect 108836 1260 108892 1540
rect 110292 1596 110348 1606
rect 109060 1372 109116 1382
rect 109060 1288 109116 1316
rect 109060 1222 109116 1232
rect 109396 1288 109452 1298
rect 109620 1288 109676 1298
rect 108836 1194 108892 1204
rect 109396 1194 109452 1204
rect 109508 1232 109620 1288
rect 108164 1036 108220 1046
rect 108052 980 108164 1036
rect 108052 812 108108 980
rect 108164 970 108220 980
rect 108052 746 108108 756
rect 107940 634 107996 644
rect 109396 568 109452 578
rect 109508 568 109564 1232
rect 109620 1222 109676 1232
rect 109452 512 109564 568
rect 109620 1148 109676 1158
rect 109620 568 109676 1092
rect 109396 502 109452 512
rect 109620 502 109676 512
rect 109844 1148 109900 1158
rect 109844 476 109900 1092
rect 109844 410 109900 420
rect 110068 1036 110124 1046
rect 110068 476 110124 980
rect 110292 1036 110348 1540
rect 110292 970 110348 980
rect 110068 410 110124 420
rect 110852 364 110908 2672
rect 110964 2188 111020 2198
rect 111188 2188 111244 2852
rect 111300 2188 111356 2198
rect 111188 2132 111300 2188
rect 110964 1148 111020 2132
rect 111300 2122 111356 2132
rect 110964 1082 111020 1092
rect 110852 298 110908 308
rect 111076 568 111132 578
rect 111076 364 111132 512
rect 111412 568 111468 14756
rect 113540 14732 113932 14788
rect 112644 12740 113036 12796
rect 112644 12628 112700 12740
rect 111748 12572 111804 12582
rect 112644 12562 112700 12572
rect 112980 12572 113036 12740
rect 112980 12516 113260 12572
rect 111748 11728 111804 12516
rect 113092 12448 113148 12458
rect 113204 12448 113260 12516
rect 113204 12392 113372 12448
rect 111748 11662 111804 11672
rect 112196 12268 112252 12278
rect 112420 12268 112476 12278
rect 112084 6860 112140 6870
rect 111972 5516 112028 5526
rect 111524 4284 111580 4294
rect 111524 1596 111580 4228
rect 111972 2492 112028 5460
rect 112084 4844 112140 6804
rect 112196 6524 112252 12212
rect 112308 12212 112420 12268
rect 112308 11908 112364 12212
rect 112420 12202 112476 12212
rect 112308 11842 112364 11852
rect 112532 11908 112588 11918
rect 112532 11564 112588 11852
rect 112532 11498 112588 11508
rect 112756 11676 112812 11686
rect 112756 10108 112812 11620
rect 113092 11008 113148 12392
rect 113316 11788 113372 12392
rect 113092 10942 113148 10952
rect 113204 11728 113260 11738
rect 113316 11722 113372 11732
rect 112756 10042 112812 10052
rect 112980 9884 113036 9894
rect 112980 8204 113036 9828
rect 113204 8540 113260 11672
rect 113540 11452 113596 14732
rect 113876 14588 113932 14732
rect 113988 14588 114044 14598
rect 113876 14532 113988 14588
rect 113988 14522 114044 14532
rect 114324 14428 114380 14868
rect 115444 14858 115500 14868
rect 120596 14868 120932 14924
rect 114436 14608 114492 14618
rect 119588 14608 119644 14618
rect 120596 14608 120652 14868
rect 120932 14858 120988 14868
rect 114492 14552 115164 14608
rect 114436 14542 114492 14552
rect 114996 14476 115052 14486
rect 114212 14364 114268 14374
rect 114324 14362 114380 14372
rect 114660 14428 114716 14438
rect 114212 14140 114268 14308
rect 114212 14084 114604 14140
rect 114324 12908 114380 12918
rect 113540 11386 113596 11396
rect 113652 12348 113708 12358
rect 113204 8474 113260 8484
rect 113316 11008 113372 11018
rect 112980 8138 113036 8148
rect 112196 6458 112252 6468
rect 112308 8092 112364 8102
rect 112084 4778 112140 4788
rect 112308 3387 112364 8036
rect 113092 6508 113148 6518
rect 112868 5788 112924 5798
rect 112868 4732 112924 5732
rect 113092 5788 113148 6452
rect 113092 5722 113148 5732
rect 113204 5292 113260 5302
rect 113204 4956 113260 5236
rect 113204 4890 113260 4900
rect 112868 4676 113260 4732
rect 112532 4528 112588 4538
rect 112532 3628 112588 4472
rect 113092 4284 113148 4294
rect 112756 4228 113092 4284
rect 112756 4060 112812 4228
rect 113092 4218 113148 4228
rect 112756 3994 112812 4004
rect 112980 4060 113036 4070
rect 113204 4060 113260 4676
rect 112532 3562 112588 3572
rect 112756 3628 112812 3638
rect 112756 3388 112812 3572
rect 112980 3500 113036 4004
rect 112980 3434 113036 3444
rect 113092 4004 113260 4060
rect 112308 3331 112476 3387
rect 112308 3164 112364 3174
rect 111972 2426 112028 2436
rect 112196 3052 112252 3062
rect 112196 2492 112252 2996
rect 112196 2426 112252 2436
rect 111524 1530 111580 1540
rect 112308 812 112364 3108
rect 112420 3088 112476 3331
rect 112756 3322 112812 3332
rect 112868 3276 112924 3286
rect 112868 3088 112924 3220
rect 112420 3032 112924 3088
rect 113092 2008 113148 4004
rect 113204 3500 113260 3510
rect 113204 2268 113260 3444
rect 113204 2202 113260 2212
rect 113316 2156 113372 10952
rect 113652 11004 113708 12292
rect 114212 12348 114268 12358
rect 114100 12124 114156 12134
rect 113988 11564 114044 11574
rect 113988 11228 114044 11508
rect 114100 11548 114156 12068
rect 114100 11482 114156 11492
rect 114212 11368 114268 12292
rect 114324 12124 114380 12852
rect 114548 12908 114604 14084
rect 114548 12842 114604 12852
rect 114324 12058 114380 12068
rect 114436 12572 114492 12582
rect 114436 12088 114492 12516
rect 114436 12022 114492 12032
rect 114548 12460 114604 12470
rect 114212 11302 114268 11312
rect 114324 11564 114380 11574
rect 114324 11228 114380 11508
rect 113988 11172 114380 11228
rect 114436 11368 114492 11378
rect 113652 10938 113708 10948
rect 114436 11008 114492 11312
rect 114436 10942 114492 10952
rect 113764 10828 113820 10838
rect 113540 10468 113596 10478
rect 113540 6508 113596 10412
rect 113764 10468 113820 10772
rect 113764 10402 113820 10412
rect 114324 10828 114380 10838
rect 114324 8204 114380 10772
rect 113652 8148 114380 8204
rect 114436 10108 114492 10118
rect 113652 6636 113708 8148
rect 113876 7980 113932 7990
rect 113876 7756 113932 7924
rect 114324 7868 114380 7878
rect 114100 7756 114156 7766
rect 113876 7700 114100 7756
rect 114100 7690 114156 7700
rect 114324 7308 114380 7812
rect 114324 7242 114380 7252
rect 113652 6570 113708 6580
rect 113764 6916 114156 6972
rect 113540 6442 113596 6452
rect 113764 6300 113820 6916
rect 114100 6860 114156 6916
rect 114324 6860 114380 6870
rect 114100 6804 114324 6860
rect 114324 6794 114380 6804
rect 113988 6748 114044 6758
rect 113988 6688 114044 6692
rect 113988 6632 114268 6688
rect 114100 6524 114156 6546
rect 114212 6508 114268 6632
rect 114324 6508 114380 6518
rect 114212 6452 114324 6508
rect 114100 6442 114156 6452
rect 114324 6442 114380 6452
rect 113540 6244 113820 6300
rect 113540 3388 113596 6244
rect 113876 6188 113932 6198
rect 113764 6132 113876 6188
rect 113764 5964 113820 6132
rect 113876 6122 113932 6132
rect 113764 5898 113820 5908
rect 114212 5852 114268 5862
rect 114212 5516 114268 5796
rect 114212 5450 114268 5460
rect 113764 3988 113820 3998
rect 113540 3322 113596 3332
rect 113652 3612 113708 3622
rect 113652 3164 113708 3556
rect 113764 3388 113820 3932
rect 113764 3322 113820 3332
rect 113988 3988 114044 3998
rect 113652 3098 113708 3108
rect 113876 2188 113932 2198
rect 113316 2090 113372 2100
rect 113428 2132 113820 2188
rect 113428 2008 113484 2132
rect 113092 1952 113484 2008
rect 113652 2044 113708 2054
rect 112308 746 112364 756
rect 111412 502 111468 512
rect 111076 298 111132 308
rect 86660 152 87052 196
rect 103012 152 103404 208
rect 113652 208 113708 1988
rect 113764 1108 113820 2132
rect 113876 2044 113932 2132
rect 113876 1978 113932 1988
rect 113988 1260 114044 3932
rect 114324 3388 114380 3398
rect 114212 3268 114268 3278
rect 114100 2268 114156 2278
rect 114100 1260 114156 2212
rect 114212 2188 114268 3212
rect 114324 3052 114380 3332
rect 114324 2986 114380 2996
rect 114436 2828 114492 10052
rect 114548 4348 114604 12404
rect 114660 6860 114716 14372
rect 114996 14252 115052 14420
rect 115108 14428 115164 14552
rect 115108 14362 115164 14372
rect 115220 14532 117404 14588
rect 115220 14252 115276 14532
rect 116564 14428 116620 14438
rect 114996 14196 115276 14252
rect 116340 14252 116396 14262
rect 116340 14068 116396 14196
rect 116564 14252 116620 14372
rect 116564 14186 116620 14196
rect 116788 14428 116844 14438
rect 115444 14028 115500 14038
rect 115332 13972 115444 14028
rect 114772 13916 114828 13926
rect 114828 13860 115052 13916
rect 114772 13850 114828 13860
rect 114772 12684 114828 12694
rect 114996 12684 115052 13860
rect 114828 12628 114940 12684
rect 114772 12618 114828 12628
rect 114772 12460 114828 12470
rect 114884 12460 114940 12628
rect 114996 12618 115052 12628
rect 114884 12404 115164 12460
rect 114772 11728 114828 12404
rect 114772 11662 114828 11672
rect 114996 11728 115052 11738
rect 114772 11228 114828 11238
rect 114772 9660 114828 11172
rect 114996 10288 115052 11672
rect 115108 10288 115164 12404
rect 115220 12012 115276 12022
rect 115220 11188 115276 11956
rect 115220 11122 115276 11132
rect 115220 10288 115276 10298
rect 115108 10232 115220 10288
rect 114772 9594 114828 9604
rect 114884 10220 114940 10230
rect 114996 10222 115052 10232
rect 115220 10222 115276 10232
rect 114884 7868 114940 10164
rect 115332 9028 115388 13972
rect 115444 13962 115500 13972
rect 116004 14028 116060 14038
rect 116340 14012 116508 14068
rect 116004 13888 116060 13972
rect 115444 13832 116060 13888
rect 115444 13168 115500 13832
rect 116452 13692 116508 14012
rect 116452 13626 116508 13636
rect 115668 13168 115724 13178
rect 115444 13102 115500 13112
rect 115556 13112 115668 13168
rect 114884 7802 114940 7812
rect 115108 8972 115388 9028
rect 115444 10220 115500 10230
rect 115108 7756 115164 8972
rect 115444 8652 115500 10164
rect 115444 8586 115500 8596
rect 115556 7948 115612 13112
rect 115668 13102 115724 13112
rect 116788 13020 116844 14372
rect 115668 12964 116844 13020
rect 116900 14372 117180 14428
rect 115668 12124 115724 12964
rect 116900 12796 116956 14372
rect 117012 14248 117068 14258
rect 117012 13916 117068 14192
rect 117124 14068 117180 14372
rect 117236 14252 117292 14286
rect 117348 14252 117404 14532
rect 117572 14532 117964 14588
rect 117572 14428 117628 14532
rect 117796 14428 117852 14438
rect 117572 14362 117628 14372
rect 117684 14372 117796 14428
rect 117684 14252 117740 14372
rect 117796 14362 117852 14372
rect 117348 14196 117740 14252
rect 117796 14252 117852 14262
rect 117908 14252 117964 14532
rect 118132 14552 119588 14608
rect 118132 14252 118188 14552
rect 119588 14542 119644 14552
rect 119700 14552 120092 14608
rect 118804 14476 118860 14486
rect 119364 14476 119420 14486
rect 118356 14252 118412 14262
rect 117908 14196 118188 14252
rect 118244 14196 118356 14252
rect 117236 14182 117292 14192
rect 117796 14068 117852 14196
rect 117124 14012 117852 14068
rect 117908 13916 117964 13926
rect 117012 13860 117908 13916
rect 117908 13850 117964 13860
rect 118132 13916 118188 13926
rect 118132 13822 118188 13832
rect 118244 13692 118300 14196
rect 118356 14186 118412 14196
rect 118804 13916 118860 14420
rect 119140 14428 119196 14438
rect 119140 14252 119196 14372
rect 119364 14362 119420 14372
rect 119700 14252 119756 14552
rect 119924 14476 119980 14486
rect 119140 14196 119756 14252
rect 119812 14248 119868 14258
rect 117796 13636 118300 13692
rect 118356 13888 118412 13898
rect 118804 13850 118860 13860
rect 119700 13916 119756 13926
rect 117796 13468 117852 13636
rect 117796 13402 117852 13412
rect 118356 12908 118412 13832
rect 119476 13580 119532 13590
rect 118580 13524 119476 13580
rect 118580 13168 118636 13524
rect 119476 13514 119532 13524
rect 118804 13168 118860 13178
rect 118580 13102 118636 13112
rect 118692 13112 118804 13168
rect 115668 12058 115724 12068
rect 115780 12740 116956 12796
rect 117012 12852 118412 12908
rect 115780 11728 115836 12740
rect 117012 12572 117068 12852
rect 116452 12516 117068 12572
rect 116004 12268 116060 12278
rect 115108 7690 115164 7700
rect 115220 7892 115612 7948
rect 115668 11672 115836 11728
rect 115892 12124 115948 12134
rect 115220 7644 115276 7892
rect 115220 7578 115276 7588
rect 115332 7756 115388 7766
rect 115220 7420 115276 7430
rect 115220 7196 115276 7364
rect 115220 7130 115276 7140
rect 115332 7048 115388 7700
rect 114660 6794 114716 6804
rect 114772 6992 115388 7048
rect 115444 7196 115500 7206
rect 114660 6508 114716 6518
rect 114660 5516 114716 6452
rect 114660 5450 114716 5460
rect 114772 4620 114828 6992
rect 115332 6860 115388 6870
rect 115332 6508 115388 6804
rect 115332 6442 115388 6452
rect 115444 5852 115500 7140
rect 115668 7048 115724 11672
rect 115780 11564 115836 11574
rect 115780 9996 115836 11508
rect 115892 10648 115948 12068
rect 116004 11676 116060 12212
rect 116340 11900 116396 11910
rect 116228 11676 116284 11686
rect 116004 11610 116060 11620
rect 116116 11620 116228 11676
rect 115892 10582 115948 10592
rect 115780 9930 115836 9940
rect 115556 6992 115724 7048
rect 115780 9324 115836 9334
rect 115556 6748 115612 6992
rect 115556 6682 115612 6692
rect 115668 6860 115724 6870
rect 115444 5786 115500 5796
rect 114772 4554 114828 4564
rect 115556 5068 115612 5078
rect 115556 4620 115612 5012
rect 115668 5068 115724 6804
rect 115780 6748 115836 9268
rect 116004 9212 116060 9222
rect 116116 9212 116172 11620
rect 116228 11610 116284 11620
rect 116340 11564 116396 11844
rect 116340 11498 116396 11508
rect 116228 11340 116284 11350
rect 116228 10444 116284 11284
rect 116228 10378 116284 10388
rect 116340 10648 116396 10658
rect 116060 9156 116172 9212
rect 116004 9146 116060 9156
rect 116340 7868 116396 10592
rect 116452 8204 116508 12516
rect 116788 12348 116844 12358
rect 117908 12348 117964 12358
rect 116844 12292 117852 12348
rect 116788 12282 116844 12292
rect 117348 12124 117404 12134
rect 117012 12068 117348 12124
rect 116788 11676 116844 11686
rect 116676 11620 116788 11676
rect 116452 8138 116508 8148
rect 116564 11564 116620 11574
rect 115780 6682 115836 6692
rect 116004 7812 116396 7868
rect 116004 6188 116060 7812
rect 116564 7756 116620 11508
rect 116676 7868 116732 11620
rect 116788 11610 116844 11620
rect 116788 9884 116844 9894
rect 117012 9884 117068 12068
rect 117348 12058 117404 12068
rect 117124 11788 117180 11798
rect 117796 11788 117852 12292
rect 117908 11908 117964 12292
rect 118244 12124 118300 12134
rect 118692 12124 118748 13112
rect 118804 13102 118860 13112
rect 118916 13076 119308 13132
rect 118916 12268 118972 13076
rect 119140 12908 119196 12918
rect 119252 12908 119308 13076
rect 119364 12908 119420 12918
rect 119252 12852 119364 12908
rect 118916 12202 118972 12212
rect 119028 12460 119084 12470
rect 118300 12068 118748 12124
rect 118244 12058 118300 12068
rect 117908 11852 118972 11908
rect 117796 11732 118300 11788
rect 117124 11728 117180 11732
rect 117124 11672 117740 11728
rect 117684 11564 117740 11672
rect 117684 11498 117740 11508
rect 117572 11004 117628 11014
rect 116844 9828 117068 9884
rect 117236 10948 117572 11004
rect 116788 9818 116844 9828
rect 117236 9748 117292 10948
rect 117572 10938 117628 10948
rect 117348 10780 117404 10790
rect 117348 10444 117404 10724
rect 117348 10378 117404 10388
rect 117460 10724 118076 10780
rect 116676 7802 116732 7812
rect 116788 9692 117292 9748
rect 116004 6122 116060 6132
rect 116116 7700 116620 7756
rect 115668 5002 115724 5012
rect 115892 5852 115948 5862
rect 115556 4554 115612 4564
rect 115780 4888 115836 4898
rect 115668 4528 115724 4538
rect 115668 4396 115724 4472
rect 114548 4292 115612 4348
rect 115668 4330 115724 4340
rect 115444 4172 115500 4182
rect 114996 3836 115052 3846
rect 115220 3836 115276 3846
rect 114772 3500 114828 3510
rect 114772 3382 114828 3392
rect 114772 3052 114828 3062
rect 114772 2908 114828 2996
rect 114996 3052 115052 3780
rect 115108 3780 115220 3836
rect 115108 3388 115164 3780
rect 115220 3770 115276 3780
rect 115108 3322 115164 3332
rect 115220 3500 115276 3510
rect 114996 2986 115052 2996
rect 115220 2908 115276 3444
rect 114772 2852 115276 2908
rect 115444 2940 115500 4116
rect 115556 3808 115612 4292
rect 115780 3948 115836 4832
rect 115780 3882 115836 3892
rect 115556 3752 115836 3808
rect 115668 3500 115724 3510
rect 115668 3088 115724 3444
rect 115780 3088 115836 3752
rect 115892 3612 115948 5796
rect 116004 4528 116060 4538
rect 116004 4168 116060 4472
rect 116004 4102 116060 4112
rect 116116 3836 116172 7700
rect 116788 7308 116844 9692
rect 117460 9388 117516 10724
rect 118020 10668 118076 10724
rect 117684 10592 117964 10648
rect 118020 10602 118076 10612
rect 117684 10444 117740 10592
rect 117684 10378 117740 10388
rect 117796 10468 117852 10478
rect 117908 10468 117964 10592
rect 118020 10468 118076 10478
rect 117908 10412 118020 10468
rect 116900 9332 117516 9388
rect 117572 9772 117628 9782
rect 116900 9212 116956 9332
rect 117124 9212 117180 9222
rect 116900 9146 116956 9156
rect 117012 9156 117124 9212
rect 116564 7252 116844 7308
rect 116564 6860 116620 7252
rect 116564 6794 116620 6804
rect 116564 6636 116620 6646
rect 116452 5068 116508 5078
rect 116452 4956 116508 5012
rect 116116 3770 116172 3780
rect 116228 4888 116284 4898
rect 116452 4890 116508 4900
rect 115892 3556 116172 3612
rect 115892 3088 115948 3098
rect 115780 3032 115892 3088
rect 115668 3022 115724 3032
rect 115892 3022 115948 3032
rect 115444 2884 115724 2940
rect 114436 2762 114492 2772
rect 115332 2828 115388 2838
rect 115332 2716 115388 2772
rect 114772 2660 115388 2716
rect 114772 2548 114828 2660
rect 114772 2482 114828 2492
rect 114996 2548 115052 2558
rect 114212 2122 114268 2132
rect 114772 2044 114828 2054
rect 114772 1820 114828 1988
rect 114772 1754 114828 1764
rect 114996 1708 115052 2492
rect 115556 2380 115612 2390
rect 115220 2008 115276 2018
rect 115276 1952 115500 2008
rect 115220 1942 115276 1952
rect 115444 1932 115500 1952
rect 115444 1866 115500 1876
rect 114996 1642 115052 1652
rect 115444 1288 115500 1298
rect 115556 1288 115612 2324
rect 114212 1260 114268 1270
rect 114100 1204 114212 1260
rect 115500 1232 115612 1288
rect 115668 1288 115724 2884
rect 116116 2368 116172 3556
rect 115892 2312 116172 2368
rect 115444 1222 115500 1232
rect 115668 1222 115724 1232
rect 115780 2188 115836 2198
rect 113988 1194 114044 1204
rect 114212 1194 114268 1204
rect 115780 1108 115836 2132
rect 115892 1596 115948 2312
rect 115892 1530 115948 1540
rect 116116 1596 116172 1606
rect 113764 1052 115836 1108
rect 116116 1036 116172 1540
rect 116116 970 116172 980
rect 116228 476 116284 4832
rect 116340 4620 116396 4630
rect 116340 3988 116396 4564
rect 116452 3988 116508 3998
rect 116340 3932 116452 3988
rect 116452 3922 116508 3932
rect 116340 3836 116396 3846
rect 116340 3628 116396 3780
rect 116340 3562 116396 3572
rect 116564 1596 116620 6580
rect 117012 5964 117068 9156
rect 117124 9146 117180 9156
rect 117124 8316 117180 8326
rect 117124 7868 117180 8260
rect 117124 7802 117180 7812
rect 117348 7532 117404 7542
rect 117012 5898 117068 5908
rect 117124 6748 117180 6758
rect 117012 5788 117068 5798
rect 116564 1530 116620 1540
rect 116676 5292 116732 5302
rect 116228 410 116284 420
rect 116676 364 116732 5236
rect 116788 2188 116844 2198
rect 116788 1484 116844 2132
rect 117012 2188 117068 5732
rect 117012 2122 117068 2132
rect 117124 1648 117180 6692
rect 117348 6748 117404 7476
rect 117460 7228 117516 7238
rect 117460 6860 117516 7172
rect 117460 6794 117516 6804
rect 117348 6682 117404 6692
rect 117460 6636 117516 6646
rect 117572 6636 117628 9716
rect 117684 9324 117740 9334
rect 117684 8316 117740 9268
rect 117684 8250 117740 8260
rect 117684 7868 117740 7878
rect 117684 7408 117740 7812
rect 117796 7644 117852 10412
rect 118020 10402 118076 10412
rect 118244 10444 118300 11732
rect 118244 10378 118300 10388
rect 118580 11452 118636 11462
rect 118244 10288 118300 10298
rect 118244 9748 118300 10232
rect 118468 10288 118524 10298
rect 118020 9692 118300 9748
rect 118356 10108 118412 10118
rect 117796 7578 117852 7588
rect 117908 8204 117964 8214
rect 117684 7352 117852 7408
rect 117516 6580 117628 6636
rect 117684 7196 117740 7206
rect 117460 6570 117516 6580
rect 117236 6524 117292 6534
rect 117236 5788 117292 6468
rect 117236 5722 117292 5732
rect 117684 4888 117740 7140
rect 117796 6524 117852 7352
rect 117796 6458 117852 6468
rect 117684 4822 117740 4832
rect 117348 4348 117404 4358
rect 117236 3628 117292 3638
rect 117236 2380 117292 3572
rect 117348 3164 117404 4292
rect 117348 3098 117404 3108
rect 117460 3808 117516 3818
rect 117236 2314 117292 2324
rect 117124 1582 117180 1592
rect 117348 2008 117404 2018
rect 117348 1484 117404 1952
rect 117460 1648 117516 3752
rect 117684 2908 117740 2918
rect 117572 2368 117628 2378
rect 117572 2156 117628 2312
rect 117572 2090 117628 2100
rect 117684 2008 117740 2852
rect 117908 2604 117964 8148
rect 118020 7228 118076 9692
rect 118244 9436 118300 9446
rect 118132 8988 118188 8998
rect 118132 8652 118188 8932
rect 118132 8586 118188 8596
rect 118244 8428 118300 9380
rect 118244 8362 118300 8372
rect 118244 8092 118300 8102
rect 118244 7532 118300 8036
rect 118244 7466 118300 7476
rect 118020 7162 118076 7172
rect 118020 6524 118076 6534
rect 118020 4168 118076 6468
rect 118244 5068 118300 5078
rect 118132 4888 118188 4898
rect 118132 4508 118188 4832
rect 118132 4442 118188 4452
rect 118020 4112 118188 4168
rect 117908 2538 117964 2548
rect 118020 3388 118076 3398
rect 117684 1942 117740 1952
rect 117460 1582 117516 1592
rect 118020 1596 118076 3332
rect 118132 2908 118188 4112
rect 118244 3388 118300 5012
rect 118356 4508 118412 10052
rect 118468 8764 118524 10232
rect 118468 8698 118524 8708
rect 118356 4442 118412 4452
rect 118468 7420 118524 7430
rect 118244 3322 118300 3332
rect 118132 2842 118188 2852
rect 118020 1530 118076 1540
rect 118468 1596 118524 7364
rect 118580 6524 118636 11396
rect 118804 11340 118860 11350
rect 118692 11284 118804 11340
rect 118692 11188 118748 11284
rect 118804 11274 118860 11284
rect 118692 11122 118748 11132
rect 118916 11188 118972 11852
rect 118916 11122 118972 11132
rect 119028 9436 119084 12404
rect 119140 12268 119196 12852
rect 119364 12842 119420 12852
rect 119364 12628 119420 12638
rect 119364 12460 119420 12572
rect 119364 12394 119420 12404
rect 119588 12628 119644 12638
rect 119140 12202 119196 12212
rect 119140 11908 119196 11918
rect 119140 11452 119196 11852
rect 119140 11386 119196 11396
rect 119252 11900 119308 11910
rect 119028 9370 119084 9380
rect 118692 8988 118748 8998
rect 118692 8540 118748 8932
rect 118692 8474 118748 8484
rect 118804 8428 118860 8438
rect 118580 6458 118636 6468
rect 118692 7644 118748 7654
rect 118580 5628 118636 5638
rect 118580 3988 118636 5572
rect 118692 4732 118748 7588
rect 118804 5964 118860 8372
rect 119252 6688 119308 11844
rect 119364 11908 119420 11918
rect 119364 11788 119420 11852
rect 119364 11722 119420 11732
rect 119588 10108 119644 12572
rect 119588 10042 119644 10052
rect 119364 9324 119420 9334
rect 119364 8764 119420 9268
rect 119364 8698 119420 8708
rect 119588 9324 119644 9334
rect 119588 8092 119644 9268
rect 119364 8036 119644 8092
rect 119364 7644 119420 8036
rect 119364 7578 119420 7588
rect 119476 7868 119532 7878
rect 118804 5898 118860 5908
rect 119028 6632 119308 6688
rect 119028 5964 119084 6632
rect 119140 6524 119196 6534
rect 119364 6524 119420 6534
rect 119196 6468 119308 6524
rect 119140 6458 119196 6468
rect 119028 5898 119084 5908
rect 119028 5628 119084 5638
rect 119028 5292 119084 5572
rect 119028 5226 119084 5236
rect 119252 5292 119308 6468
rect 119364 5852 119420 6468
rect 119364 5786 119420 5796
rect 119252 5226 119308 5236
rect 118804 5068 118860 5078
rect 118804 4956 118860 5012
rect 118804 4890 118860 4900
rect 119028 4956 119084 4966
rect 119028 4888 119084 4900
rect 119028 4822 119084 4832
rect 119364 4888 119420 4898
rect 118692 4676 119084 4732
rect 118580 3932 118860 3988
rect 118580 3088 118636 3098
rect 118580 2380 118636 3032
rect 118580 2314 118636 2324
rect 118468 1530 118524 1540
rect 116788 1428 117180 1484
rect 117348 1428 117628 1484
rect 116676 298 116732 308
rect 117012 1260 117068 1270
rect 117012 208 117068 1204
rect 117124 1108 117180 1428
rect 117572 1260 117628 1428
rect 117572 1194 117628 1204
rect 117124 1052 117964 1108
rect 117572 700 117628 710
rect 117572 476 117628 644
rect 117572 410 117628 420
rect 117796 568 117852 578
rect 117796 476 117852 512
rect 117796 410 117852 420
rect 117908 388 117964 1052
rect 118804 568 118860 3932
rect 118916 3808 118972 3818
rect 118916 700 118972 3752
rect 119028 3052 119084 4676
rect 119252 4348 119308 4358
rect 119252 3836 119308 4292
rect 119364 4284 119420 4832
rect 119364 4218 119420 4228
rect 119252 3770 119308 3780
rect 119364 3448 119420 3458
rect 119028 2986 119084 2996
rect 119140 3388 119196 3398
rect 119140 2368 119196 3332
rect 119140 2302 119196 2312
rect 119252 3088 119308 3098
rect 119252 1036 119308 3032
rect 119364 1932 119420 3392
rect 119476 2828 119532 7812
rect 119588 4732 119644 4742
rect 119588 4284 119644 4676
rect 119588 4218 119644 4228
rect 119700 3836 119756 13860
rect 119812 8092 119868 14192
rect 119924 13692 119980 14420
rect 120036 14248 120092 14552
rect 120372 14588 120652 14608
rect 120428 14552 120652 14588
rect 121044 14700 121100 14710
rect 120372 14522 120428 14532
rect 120484 14476 120540 14486
rect 120036 14182 120092 14192
rect 120148 14428 120204 14438
rect 119924 13636 120092 13692
rect 119924 13132 119980 13142
rect 119924 11676 119980 13076
rect 120036 11676 120092 13636
rect 120148 12088 120204 14372
rect 120372 13580 120428 13590
rect 120484 13580 120540 14420
rect 120708 14364 120764 14374
rect 120428 13524 120540 13580
rect 120596 13804 120652 13814
rect 120596 13580 120652 13748
rect 120372 13514 120428 13524
rect 120596 13514 120652 13524
rect 120708 12572 120764 14308
rect 121044 14364 121100 14644
rect 121044 14298 121100 14308
rect 121268 14700 121324 14710
rect 120820 14248 120876 14258
rect 120820 13804 120876 14192
rect 120820 13738 120876 13748
rect 120708 12506 120764 12516
rect 120932 12796 120988 12806
rect 120372 12448 120428 12458
rect 120148 12022 120204 12032
rect 120260 12236 120316 12246
rect 120148 11676 120204 11686
rect 120036 11620 120148 11676
rect 119924 11610 119980 11620
rect 120148 11610 120204 11620
rect 120260 10648 120316 12180
rect 120148 10592 120316 10648
rect 120036 10220 120092 10230
rect 120036 9928 120092 10164
rect 120036 9862 120092 9872
rect 119812 8026 119868 8036
rect 119924 9772 119980 9782
rect 119924 5852 119980 9716
rect 120036 9548 120092 9558
rect 120036 9324 120092 9492
rect 120036 9258 120092 9268
rect 119924 5786 119980 5796
rect 120036 7756 120092 7766
rect 120036 4844 120092 7700
rect 120036 4778 120092 4788
rect 120036 4708 120092 4718
rect 119700 3770 119756 3780
rect 119924 4172 119980 4182
rect 119476 2762 119532 2772
rect 119364 1866 119420 1876
rect 119252 970 119308 980
rect 119924 1036 119980 4116
rect 120036 3448 120092 4652
rect 120148 4060 120204 10592
rect 120260 10468 120316 10478
rect 120260 8204 120316 10412
rect 120260 8138 120316 8148
rect 120372 6972 120428 12392
rect 120596 12236 120652 12246
rect 120596 11908 120652 12180
rect 120596 11842 120652 11852
rect 120932 11788 120988 12740
rect 121044 12448 121100 12458
rect 121044 12348 121100 12392
rect 121044 12282 121100 12292
rect 120932 11722 120988 11732
rect 121156 12268 121212 12278
rect 120484 11368 120540 11378
rect 120540 11312 120764 11368
rect 120484 11302 120540 11312
rect 120596 11008 120652 11018
rect 120708 11008 120764 11312
rect 120820 11008 120876 11018
rect 120708 10952 120820 11008
rect 120596 10828 120652 10952
rect 120820 10942 120876 10952
rect 121156 11004 121212 12212
rect 121156 10938 121212 10948
rect 120596 10772 120988 10828
rect 120932 10332 120988 10772
rect 121268 10648 121324 14644
rect 124628 14700 124684 14710
rect 124404 14608 124460 14618
rect 124404 14476 124460 14552
rect 124628 14608 124684 14644
rect 124628 14542 124684 14552
rect 132804 14608 132860 14618
rect 124628 14476 124684 14486
rect 124404 14410 124460 14420
rect 124516 14420 124628 14476
rect 124516 14140 124572 14420
rect 124628 14410 124684 14420
rect 124516 14074 124572 14084
rect 124740 14140 124796 14150
rect 123284 13888 123340 13898
rect 123060 13168 123116 13178
rect 122724 13020 122780 13030
rect 122164 12808 122220 12818
rect 121380 12268 121436 12278
rect 121380 11900 121436 12212
rect 121380 11834 121436 11844
rect 121716 11908 121772 11918
rect 121268 10582 121324 10592
rect 120820 10276 120988 10332
rect 120708 9324 120764 9334
rect 120596 7980 120652 7990
rect 120596 7644 120652 7924
rect 120708 7768 120764 9268
rect 120820 8204 120876 10276
rect 121044 10220 121100 10230
rect 120820 8138 120876 8148
rect 120932 10108 120988 10118
rect 120932 7980 120988 10052
rect 121044 9928 121100 10164
rect 121268 10220 121324 10230
rect 121156 9928 121212 9938
rect 121044 9872 121156 9928
rect 121156 9862 121212 9872
rect 121268 9212 121324 10164
rect 121268 9146 121324 9156
rect 121380 10108 121436 10118
rect 120932 7914 120988 7924
rect 120708 7712 121100 7768
rect 120596 7588 120988 7644
rect 120708 7228 120764 7238
rect 120372 6916 120652 6972
rect 120484 4888 120540 4898
rect 120372 4832 120484 4888
rect 120372 4396 120428 4832
rect 120484 4822 120540 4832
rect 120372 4330 120428 4340
rect 120596 4396 120652 6916
rect 120596 4330 120652 4340
rect 120148 3994 120204 4004
rect 120596 3988 120652 3998
rect 120708 3988 120764 7172
rect 120932 7228 120988 7588
rect 121044 7408 121100 7712
rect 121044 7352 121212 7408
rect 121156 7308 121212 7352
rect 121268 7308 121324 7318
rect 121156 7252 121268 7308
rect 121268 7242 121324 7252
rect 120932 7162 120988 7172
rect 121156 7084 121212 7094
rect 121156 5740 121212 7028
rect 121156 5674 121212 5684
rect 121268 5964 121324 5974
rect 121156 4956 121212 4966
rect 121156 4348 121212 4900
rect 121268 4888 121324 5908
rect 121268 4822 121324 4832
rect 121380 4528 121436 10052
rect 121604 9996 121660 10006
rect 121604 9212 121660 9940
rect 121604 9146 121660 9156
rect 121492 8092 121548 8102
rect 121492 4888 121548 8036
rect 121492 4822 121548 4832
rect 121604 7420 121660 7430
rect 121380 4462 121436 4472
rect 121156 4292 121324 4348
rect 121268 4172 121324 4292
rect 121268 4106 121324 4116
rect 120820 3988 120876 3998
rect 120708 3932 120820 3988
rect 120148 3500 120204 3510
rect 120596 3500 120652 3932
rect 120820 3922 120876 3932
rect 121604 3836 121660 7364
rect 120820 3780 121660 3836
rect 120204 3444 120540 3500
rect 120148 3434 120204 3444
rect 120036 3382 120092 3392
rect 120484 3276 120540 3444
rect 120596 3434 120652 3444
rect 120708 3612 120764 3622
rect 120708 3448 120764 3556
rect 120708 3382 120764 3392
rect 120820 3276 120876 3780
rect 120484 3220 120876 3276
rect 120932 3448 120988 3458
rect 121716 3448 121772 11852
rect 122052 10648 122108 10658
rect 121828 10288 121884 10298
rect 121828 9996 121884 10232
rect 122052 10107 122108 10592
rect 121828 9930 121884 9940
rect 121940 10051 122108 10107
rect 121828 8316 121884 8326
rect 121828 7196 121884 8260
rect 121940 7228 121996 10051
rect 121940 7172 122108 7228
rect 121828 7130 121884 7140
rect 121940 7084 121996 7094
rect 121828 6300 121884 6310
rect 121828 5964 121884 6244
rect 121828 5898 121884 5908
rect 120932 2548 120988 3392
rect 121604 3392 121772 3448
rect 121604 3388 121660 3392
rect 121604 3322 121660 3332
rect 121156 3276 121212 3286
rect 121044 3220 121156 3276
rect 121940 3268 121996 7028
rect 121044 2940 121100 3220
rect 121156 3210 121212 3220
rect 121716 3212 121996 3268
rect 121716 3088 121772 3212
rect 121940 3088 121996 3098
rect 121716 3022 121772 3032
rect 121828 3032 121940 3088
rect 121044 2874 121100 2884
rect 121828 2828 121884 3032
rect 121940 3022 121996 3032
rect 121828 2762 121884 2772
rect 121940 2728 121996 2738
rect 120260 2492 120764 2548
rect 120260 1372 120316 2492
rect 120596 2380 120652 2390
rect 120484 2324 120596 2380
rect 120484 1596 120540 2324
rect 120596 2314 120652 2324
rect 120708 2268 120764 2492
rect 120932 2482 120988 2492
rect 121156 2604 121212 2614
rect 121156 2482 121212 2492
rect 120708 2212 121660 2268
rect 121268 1820 121324 1830
rect 120932 1764 121268 1820
rect 120932 1708 120988 1764
rect 121268 1754 121324 1764
rect 120932 1642 120988 1652
rect 120484 1530 120540 1540
rect 121044 1484 121100 1494
rect 120260 1306 120316 1316
rect 120708 1372 120764 1382
rect 120372 1108 120428 1118
rect 120708 1108 120764 1316
rect 120428 1052 120764 1108
rect 120820 1288 120876 1298
rect 120372 1042 120428 1052
rect 119924 970 119980 980
rect 118916 634 118972 644
rect 119140 700 119196 710
rect 118804 502 118860 512
rect 119140 388 119196 644
rect 120820 476 120876 1232
rect 120820 410 120876 420
rect 117908 332 119196 388
rect 121044 364 121100 1428
rect 121604 1484 121660 2212
rect 121604 1418 121660 1428
rect 121940 476 121996 2672
rect 122052 2380 122108 7172
rect 122164 6076 122220 12752
rect 122724 12460 122780 12964
rect 122724 12394 122780 12404
rect 122276 11788 122332 11798
rect 122276 7644 122332 11732
rect 122500 11788 122556 11798
rect 122500 11008 122556 11732
rect 122500 10942 122556 10952
rect 122724 11008 122780 11018
rect 122724 9884 122780 10952
rect 122724 9818 122780 9828
rect 122276 7588 122556 7644
rect 122500 7532 122556 7588
rect 122500 7476 122668 7532
rect 122500 7196 122556 7206
rect 122500 6972 122556 7140
rect 122500 6906 122556 6916
rect 122164 6010 122220 6020
rect 122276 6636 122332 6646
rect 122276 5740 122332 6580
rect 122276 5674 122332 5684
rect 122500 6636 122556 6646
rect 122388 3612 122444 3622
rect 122388 2728 122444 3556
rect 122388 2662 122444 2672
rect 122500 2604 122556 6580
rect 122612 6076 122668 7476
rect 122612 6010 122668 6020
rect 122724 6972 122780 6982
rect 122724 5404 122780 6916
rect 122724 5338 122780 5348
rect 122948 6300 123004 6310
rect 122836 4844 122892 4854
rect 122052 2314 122108 2324
rect 122276 2548 122556 2604
rect 122612 3628 122668 3638
rect 122276 1108 122332 2548
rect 122612 2380 122668 3572
rect 122612 2314 122668 2324
rect 122500 2268 122556 2278
rect 122388 2188 122444 2198
rect 122500 2188 122556 2212
rect 122612 2188 122668 2198
rect 122500 2132 122612 2188
rect 122388 2044 122444 2132
rect 122612 2122 122668 2132
rect 122388 1988 122780 2044
rect 122500 1828 122556 1838
rect 122500 1484 122556 1772
rect 122724 1828 122780 1988
rect 122724 1762 122780 1772
rect 122500 1418 122556 1428
rect 122276 1042 122332 1052
rect 122836 1108 122892 4788
rect 122948 3612 123004 6244
rect 122948 3546 123004 3556
rect 123060 2604 123116 13112
rect 123284 13168 123340 13832
rect 124292 13804 124348 13814
rect 124348 13748 124572 13804
rect 124292 13738 124348 13748
rect 123284 13102 123340 13112
rect 123508 12448 123564 12458
rect 123396 11728 123452 11738
rect 123396 8092 123452 11672
rect 123508 8652 123564 12392
rect 124516 10892 124572 13748
rect 124740 13468 124796 14084
rect 126756 14068 126812 14078
rect 124740 13402 124796 13412
rect 126196 13888 126252 13898
rect 126196 12808 126252 13832
rect 126196 12742 126252 12752
rect 126756 12808 126812 14012
rect 126980 13916 127036 13926
rect 126980 13528 127036 13860
rect 126756 12742 126812 12752
rect 126868 13472 127036 13528
rect 126868 12628 126924 13472
rect 132692 13132 132748 13142
rect 127540 12988 127596 12998
rect 127764 12988 127820 12998
rect 127596 12932 127708 12988
rect 127540 12922 127596 12932
rect 126532 12572 126924 12628
rect 125524 12460 125580 12470
rect 125524 12236 125580 12404
rect 126532 12460 126588 12572
rect 126532 12394 126588 12404
rect 125524 12170 125580 12180
rect 125748 12236 125804 12246
rect 124516 10826 124572 10836
rect 125748 10220 125804 12180
rect 127652 12088 127708 12932
rect 127652 12022 127708 12032
rect 126308 11900 126364 11910
rect 126308 11340 126364 11844
rect 126308 11274 126364 11284
rect 126532 11564 126588 11574
rect 126532 11340 126588 11508
rect 126532 11274 126588 11284
rect 126308 10780 126364 10790
rect 125748 10154 125804 10164
rect 126084 10332 126140 10342
rect 126084 10108 126140 10276
rect 126084 10042 126140 10052
rect 126308 10108 126364 10724
rect 126308 10042 126364 10052
rect 124628 9660 124684 9670
rect 124628 9100 124684 9604
rect 124628 9034 124684 9044
rect 124852 9660 124908 9670
rect 123508 8586 123564 8596
rect 124852 8428 124908 9604
rect 126980 8988 127036 8998
rect 126980 8540 127036 8932
rect 126980 8474 127036 8484
rect 127204 8988 127260 8998
rect 124852 8362 124908 8372
rect 123396 8026 123452 8036
rect 127092 8092 127148 8102
rect 126868 7756 126924 7766
rect 126868 7308 126924 7700
rect 127092 7756 127148 8036
rect 127204 7868 127260 8932
rect 127204 7802 127260 7812
rect 127092 7690 127148 7700
rect 127092 7532 127148 7542
rect 126980 7308 127036 7318
rect 126868 7252 126980 7308
rect 126980 7242 127036 7252
rect 126084 7196 126140 7206
rect 124964 6636 125020 6646
rect 124964 6300 125020 6580
rect 124964 6234 125020 6244
rect 123508 6076 123564 6086
rect 123508 5628 123564 6020
rect 123508 5562 123564 5572
rect 124292 4620 124348 4630
rect 124292 4528 124348 4564
rect 124292 4462 124348 4472
rect 125412 4396 125468 4406
rect 124180 4172 124236 4182
rect 124180 4078 124236 4112
rect 124404 4172 124460 4182
rect 123060 2538 123116 2548
rect 123284 3724 123340 3734
rect 123284 1372 123340 3668
rect 124292 3628 124348 3638
rect 123844 2268 123900 2278
rect 123284 1306 123340 1316
rect 123508 1372 123564 1382
rect 123508 1288 123564 1316
rect 123508 1222 123564 1232
rect 122836 1042 122892 1052
rect 123844 924 123900 2212
rect 124292 1648 124348 3572
rect 124404 3268 124460 4116
rect 125412 3836 125468 4340
rect 126084 3988 126140 7140
rect 127092 7084 127148 7476
rect 127764 7228 127820 12932
rect 130788 12348 130844 12358
rect 130788 12268 130844 12292
rect 130788 12212 131068 12268
rect 128324 12088 128380 12098
rect 127988 8876 128044 8886
rect 127988 8428 128044 8820
rect 127988 8362 128044 8372
rect 127764 7162 127820 7172
rect 127092 7018 127148 7028
rect 126644 6412 126700 6422
rect 126644 5852 126700 6356
rect 126644 5786 126700 5796
rect 127204 4844 127260 4854
rect 126980 4732 127036 4742
rect 126308 4348 126364 4358
rect 126308 4168 126364 4292
rect 126868 4168 126924 4178
rect 126308 4112 126868 4168
rect 126868 4102 126924 4112
rect 126980 4060 127036 4676
rect 126980 3994 127036 4004
rect 126084 3922 126140 3932
rect 125860 3836 125916 3846
rect 125412 3780 125860 3836
rect 125860 3770 125916 3780
rect 127092 3448 127148 3458
rect 124404 3202 124460 3212
rect 124628 3268 124684 3278
rect 124292 1582 124348 1592
rect 124628 1596 124684 3212
rect 125636 3052 125692 3062
rect 125636 2492 125692 2996
rect 127092 3052 127148 3392
rect 127092 2986 127148 2996
rect 125636 2426 125692 2436
rect 125972 2188 126028 2198
rect 124628 1530 124684 1540
rect 125860 2044 125916 2054
rect 123844 858 123900 868
rect 123956 1288 124012 1298
rect 123956 568 124012 1232
rect 125860 1148 125916 1988
rect 125972 1260 126028 2132
rect 125972 1194 126028 1204
rect 126196 1828 126252 1838
rect 125860 1082 125916 1092
rect 126196 1148 126252 1772
rect 127204 1708 127260 4788
rect 127204 1642 127260 1652
rect 127428 3500 127484 3510
rect 126196 1082 126252 1092
rect 127428 1148 127484 3444
rect 128324 3387 128380 12032
rect 131012 11728 131068 12212
rect 131460 12236 131516 12246
rect 131460 11900 131516 12180
rect 131460 11834 131516 11844
rect 132468 12236 132524 12246
rect 131012 11672 131516 11728
rect 130900 11548 130956 11558
rect 129444 11228 129500 11238
rect 128436 8316 128492 8326
rect 128436 7756 128492 8260
rect 129444 8204 129500 11172
rect 130900 10668 130956 11492
rect 130900 10602 130956 10612
rect 131012 11116 131068 11126
rect 129444 8138 129500 8148
rect 129780 10444 129836 10454
rect 128436 7690 128492 7700
rect 129220 7868 129276 7878
rect 129220 6524 129276 7812
rect 129220 6458 129276 6468
rect 129332 7084 129388 7094
rect 129332 5404 129388 7028
rect 129556 6636 129612 6646
rect 129780 6636 129836 10388
rect 130900 10332 130956 10342
rect 131012 10332 131068 11060
rect 130956 10276 131068 10332
rect 131124 11004 131180 11014
rect 130900 10266 130956 10276
rect 131012 9212 131068 9222
rect 129612 6580 129836 6636
rect 130788 6748 130844 6758
rect 129556 6570 129612 6580
rect 129332 5338 129388 5348
rect 129556 5964 129612 5974
rect 129556 5404 129612 5908
rect 129556 5338 129612 5348
rect 128548 5292 128604 5302
rect 129668 5292 129724 5302
rect 128604 5236 129668 5248
rect 128548 5192 129724 5236
rect 128324 3331 128492 3387
rect 127428 1082 127484 1092
rect 127540 1468 127596 1478
rect 125860 928 125916 962
rect 125860 858 125916 868
rect 123956 502 124012 512
rect 124180 588 124236 606
rect 124180 502 124236 512
rect 121940 410 121996 420
rect 121044 298 121100 308
rect 127540 364 127596 1412
rect 128436 1468 128492 3331
rect 129668 3268 129724 3278
rect 129668 2728 129724 3212
rect 129668 2662 129724 2672
rect 129332 1820 129388 1830
rect 129332 1484 129388 1764
rect 129332 1418 129388 1428
rect 128436 1402 128492 1412
rect 130788 476 130844 6692
rect 131012 5628 131068 9156
rect 131124 8652 131180 10948
rect 131124 8586 131180 8596
rect 131348 10648 131404 10658
rect 131012 5562 131068 5572
rect 131236 5964 131292 5974
rect 131236 5404 131292 5908
rect 131236 5338 131292 5348
rect 131348 5292 131404 10592
rect 131460 6076 131516 11672
rect 132244 11548 132300 11558
rect 131460 6010 131516 6020
rect 132132 11004 132188 11014
rect 131348 5226 131404 5236
rect 131012 5068 131068 5078
rect 131012 4508 131068 5012
rect 131012 4442 131068 4452
rect 131124 4888 131180 4898
rect 131012 4172 131068 4182
rect 131012 3808 131068 4116
rect 131012 3742 131068 3752
rect 130788 410 130844 420
rect 131124 476 131180 4832
rect 131460 4888 131516 4898
rect 131460 3988 131516 4832
rect 132132 4620 132188 10948
rect 132132 4554 132188 4564
rect 131460 3922 131516 3932
rect 131684 4348 131740 4358
rect 131684 3988 131740 4292
rect 132244 4060 132300 11492
rect 132468 9100 132524 12180
rect 132692 11788 132748 13076
rect 132692 11722 132748 11732
rect 132804 11548 132860 14552
rect 133140 14068 133196 14078
rect 132692 11492 132860 11548
rect 132916 11728 132972 11738
rect 132692 11188 132748 11492
rect 132692 11132 132860 11188
rect 132468 9034 132524 9044
rect 132244 3994 132300 4004
rect 132356 4844 132412 4854
rect 131684 3922 131740 3932
rect 132020 3836 132076 3846
rect 132020 3628 132076 3780
rect 132020 3562 132076 3572
rect 131460 3164 131516 3174
rect 131460 1708 131516 3108
rect 132356 2188 132412 4788
rect 132692 3836 132748 3846
rect 132580 3276 132636 3286
rect 132580 3088 132636 3220
rect 132692 3268 132748 3780
rect 132804 3808 132860 11132
rect 132916 8092 132972 11672
rect 133028 11548 133084 11558
rect 133028 11340 133084 11492
rect 133028 11274 133084 11284
rect 132916 8026 132972 8036
rect 133028 10892 133084 10902
rect 133028 6412 133084 10836
rect 133028 6346 133084 6356
rect 133140 5852 133196 14012
rect 134036 14028 134092 14038
rect 133476 13244 133532 13254
rect 133364 9436 133420 9446
rect 133364 8764 133420 9380
rect 133364 8698 133420 8708
rect 133364 7756 133420 7766
rect 133364 7420 133420 7700
rect 133364 7354 133420 7364
rect 133476 6300 133532 13188
rect 133924 11548 133980 11558
rect 133476 6234 133532 6244
rect 133588 11116 133644 11126
rect 133140 5786 133196 5796
rect 133476 5068 133532 5078
rect 133476 4508 133532 5012
rect 133588 4956 133644 11060
rect 133700 10892 133756 10902
rect 133700 8316 133756 10836
rect 133924 10556 133980 11492
rect 133924 10490 133980 10500
rect 134036 8876 134092 13972
rect 134260 14028 134316 14038
rect 134260 13244 134316 13972
rect 138068 13916 138124 13926
rect 137172 13888 137228 13898
rect 136500 13468 136556 13478
rect 134260 13178 134316 13188
rect 135604 13244 135660 13254
rect 134260 12268 134316 12278
rect 134148 11908 134204 11918
rect 134148 9884 134204 11852
rect 134260 11676 134316 12212
rect 135492 11900 135548 11910
rect 135492 11787 135548 11844
rect 134260 11610 134316 11620
rect 135044 11731 135548 11787
rect 134260 11188 134316 11198
rect 134260 10444 134316 11132
rect 134260 10378 134316 10388
rect 134820 10828 134876 10838
rect 134260 10288 134316 10298
rect 134260 10108 134316 10232
rect 134260 10042 134316 10052
rect 134148 9818 134204 9828
rect 134036 8810 134092 8820
rect 133700 8250 133756 8260
rect 134820 7980 134876 10772
rect 134932 9928 134988 9938
rect 134932 8204 134988 9872
rect 134932 8138 134988 8148
rect 134820 7914 134876 7924
rect 134260 7644 134316 7654
rect 134260 7228 134316 7588
rect 134260 7162 134316 7172
rect 134260 6972 134316 6982
rect 134260 6636 134316 6916
rect 134260 6570 134316 6580
rect 134260 5852 134316 5862
rect 134260 5788 134316 5796
rect 134260 5722 134316 5732
rect 133588 4890 133644 4900
rect 133812 4956 133868 4966
rect 133476 4442 133532 4452
rect 132804 3742 132860 3752
rect 133812 3387 133868 4900
rect 134372 4528 134428 4538
rect 134372 4434 134428 4452
rect 134596 4060 134652 4070
rect 132692 3202 132748 3212
rect 133700 3331 133868 3387
rect 134260 3948 134316 3958
rect 132468 3052 132636 3088
rect 132524 3032 132636 3052
rect 132468 2986 132524 2996
rect 133028 2828 133084 2838
rect 133028 2728 133084 2772
rect 132692 2716 133084 2728
rect 132748 2672 133084 2716
rect 132692 2650 132748 2660
rect 132804 2268 132860 2278
rect 132804 2188 132860 2212
rect 132356 2132 132748 2188
rect 132804 2156 133308 2188
rect 132804 2132 133252 2156
rect 132020 1708 132076 1718
rect 131460 1652 132020 1708
rect 132020 1642 132076 1652
rect 132692 1260 132748 2132
rect 133252 2090 133308 2100
rect 132804 1772 133084 1828
rect 132804 1708 132860 1772
rect 132804 1642 132860 1652
rect 133028 1708 133084 1772
rect 133028 1642 133084 1652
rect 133700 1708 133756 3331
rect 134260 2828 134316 3892
rect 134596 2908 134652 4004
rect 134596 2842 134652 2852
rect 134260 2762 134316 2772
rect 134260 2380 134316 2406
rect 134260 2302 134316 2312
rect 134596 2380 134652 2390
rect 133700 1642 133756 1652
rect 134148 2268 134204 2278
rect 134148 1648 134204 2212
rect 134148 1582 134204 1592
rect 134484 2268 134540 2278
rect 134484 1288 134540 2212
rect 134484 1222 134540 1232
rect 132692 1194 132748 1204
rect 134596 700 134652 2324
rect 135044 1372 135100 11731
rect 135268 9772 135324 9782
rect 135268 9436 135324 9716
rect 135268 9370 135324 9380
rect 135604 8764 135660 13188
rect 135940 11340 136108 11368
rect 135996 11312 136108 11340
rect 135940 11274 135996 11284
rect 136052 10828 136108 11312
rect 136052 10762 136108 10772
rect 135940 10468 135996 10478
rect 135940 9212 135996 10412
rect 135940 9146 135996 9156
rect 135604 8698 135660 8708
rect 135828 8092 135884 8102
rect 135828 4620 135884 8036
rect 136500 8092 136556 13412
rect 137172 11728 137228 13832
rect 137956 13468 138012 13478
rect 137620 12908 137676 12918
rect 137620 12684 137676 12852
rect 137620 12618 137676 12628
rect 137844 12684 137900 12694
rect 137172 11662 137228 11672
rect 137732 11788 137788 11798
rect 136500 8026 136556 8036
rect 136724 11340 136780 11350
rect 135940 6972 135996 6982
rect 135940 6508 135996 6916
rect 135940 6442 135996 6452
rect 135940 4956 135996 4966
rect 135940 4888 135996 4900
rect 135940 4822 135996 4832
rect 136276 4888 136332 4898
rect 135828 4554 135884 4564
rect 136164 4708 136220 4718
rect 136052 4348 136108 4358
rect 136052 3088 136108 4292
rect 136052 3022 136108 3032
rect 135828 2940 135884 2950
rect 135716 2548 135772 2558
rect 135716 1596 135772 2492
rect 135716 1530 135772 1540
rect 135604 1484 135660 1494
rect 135604 1390 135660 1412
rect 135044 1306 135100 1316
rect 135828 1260 135884 2884
rect 135940 2908 135996 2918
rect 135940 2548 135996 2852
rect 136164 2908 136220 4652
rect 136164 2842 136220 2852
rect 135940 2482 135996 2492
rect 136276 2188 136332 4832
rect 136388 4708 136444 4718
rect 136388 2380 136444 4652
rect 136724 3387 136780 11284
rect 137732 10780 137788 11732
rect 137844 11548 137900 12628
rect 137844 11482 137900 11492
rect 137732 10714 137788 10724
rect 137956 10648 138012 13412
rect 138068 11728 138124 13860
rect 138964 12628 139020 14912
rect 150836 14924 151676 14968
rect 150836 14912 151620 14924
rect 149044 14732 149772 14788
rect 138964 12562 139020 12572
rect 139412 14364 139468 14374
rect 138292 12348 138348 12358
rect 138068 11662 138124 11672
rect 138180 12012 138236 12022
rect 138180 11188 138236 11956
rect 138180 11122 138236 11132
rect 138292 11116 138348 12292
rect 138628 11452 138684 11462
rect 138292 11050 138348 11060
rect 138404 11188 138460 11198
rect 138180 10648 138236 10658
rect 137956 10582 138012 10592
rect 138068 10592 138180 10648
rect 138068 10468 138124 10592
rect 138180 10582 138236 10592
rect 137620 10412 138124 10468
rect 137004 10220 137324 10252
rect 137004 10164 137032 10220
rect 137088 10164 137136 10220
rect 137192 10164 137240 10220
rect 137296 10164 137324 10220
rect 137004 9729 137324 10164
rect 137004 9673 137032 9729
rect 137088 9673 137136 9729
rect 137192 9673 137240 9729
rect 137296 9673 137324 9729
rect 137004 9625 137324 9673
rect 137004 9569 137032 9625
rect 137088 9569 137136 9625
rect 137192 9569 137240 9625
rect 137296 9569 137324 9625
rect 137004 9521 137324 9569
rect 137004 9465 137032 9521
rect 137088 9465 137136 9521
rect 137192 9465 137240 9521
rect 137296 9465 137324 9521
rect 137004 8652 137324 9465
rect 137004 8596 137032 8652
rect 137088 8596 137136 8652
rect 137192 8596 137240 8652
rect 137296 8596 137324 8652
rect 137004 8331 137324 8596
rect 137004 8275 137032 8331
rect 137088 8275 137136 8331
rect 137192 8275 137240 8331
rect 137296 8275 137324 8331
rect 137004 8227 137324 8275
rect 137004 8171 137032 8227
rect 137088 8171 137136 8227
rect 137192 8171 137240 8227
rect 137296 8171 137324 8227
rect 137004 8123 137324 8171
rect 137004 8067 137032 8123
rect 137088 8067 137136 8123
rect 137192 8067 137240 8123
rect 137296 8067 137324 8123
rect 136836 7756 136892 7766
rect 136836 7084 136892 7700
rect 136836 7018 136892 7028
rect 137004 7084 137324 8067
rect 137004 7028 137032 7084
rect 137088 7028 137136 7084
rect 137192 7028 137240 7084
rect 137296 7028 137324 7084
rect 137004 6933 137324 7028
rect 137004 6877 137032 6933
rect 137088 6877 137136 6933
rect 137192 6877 137240 6933
rect 137296 6877 137324 6933
rect 137004 6829 137324 6877
rect 137004 6773 137032 6829
rect 137088 6773 137136 6829
rect 137192 6773 137240 6829
rect 137296 6773 137324 6829
rect 137004 6725 137324 6773
rect 137004 6669 137032 6725
rect 137088 6669 137136 6725
rect 137192 6669 137240 6725
rect 137296 6669 137324 6725
rect 137004 5535 137324 6669
rect 137004 5460 137032 5535
rect 137088 5460 137136 5535
rect 137192 5460 137240 5535
rect 137296 5460 137324 5535
rect 137004 5431 137324 5460
rect 137508 8092 137564 8102
rect 137508 5516 137564 8036
rect 137620 6972 137676 10412
rect 138068 10288 138124 10298
rect 137956 8092 138012 8102
rect 137956 7868 138012 8036
rect 137956 7802 138012 7812
rect 137620 6906 137676 6916
rect 137508 5450 137564 5460
rect 137844 5516 137900 5526
rect 137004 5375 137032 5431
rect 137088 5375 137136 5431
rect 137192 5375 137240 5431
rect 137296 5375 137324 5431
rect 137004 5327 137324 5375
rect 137004 5271 137032 5327
rect 137088 5271 137136 5327
rect 137192 5271 137240 5327
rect 137296 5271 137324 5327
rect 137004 4644 137324 5271
rect 137396 4844 137452 4854
rect 137396 3724 137452 4788
rect 137844 3808 137900 5460
rect 137396 3658 137452 3668
rect 137732 3752 137900 3808
rect 137620 3628 137676 3638
rect 137732 3628 137788 3752
rect 137676 3572 137788 3628
rect 137844 3612 137900 3622
rect 137620 3562 137676 3572
rect 136724 3331 136892 3387
rect 136836 2728 136892 3331
rect 136836 2662 136892 2672
rect 136388 2314 136444 2324
rect 137732 2604 137788 2614
rect 137732 2380 137788 2548
rect 137732 2314 137788 2324
rect 135828 1194 135884 1204
rect 135940 2132 136332 2188
rect 137844 2188 137900 3556
rect 137732 2156 137788 2166
rect 135940 1108 135996 2132
rect 137844 2122 137900 2132
rect 136164 1932 136220 1942
rect 136164 1468 136220 1876
rect 136164 1402 136220 1412
rect 135940 1042 135996 1052
rect 137732 928 137788 2100
rect 138068 1260 138124 10232
rect 138180 7420 138236 7430
rect 138180 6972 138236 7364
rect 138180 6906 138236 6916
rect 138404 5068 138460 11132
rect 138516 9100 138572 9110
rect 138516 8540 138572 9044
rect 138516 8474 138572 8484
rect 138628 6636 138684 11396
rect 138628 6570 138684 6580
rect 138740 10108 138796 10118
rect 138404 5002 138460 5012
rect 138740 4888 138796 10052
rect 139412 9884 139468 14308
rect 142660 14252 142716 14262
rect 139524 14068 139580 14078
rect 139524 13916 139580 14012
rect 142660 14068 142716 14196
rect 142660 14002 142716 14012
rect 145684 14248 145740 14258
rect 139524 13850 139580 13860
rect 141092 13348 141148 13358
rect 141092 12988 141148 13292
rect 141092 12922 141148 12932
rect 142996 13348 143052 13358
rect 142436 12908 142492 12918
rect 141092 12808 141148 12818
rect 139748 12268 139804 12278
rect 139412 9818 139468 9828
rect 139524 12088 139580 12098
rect 139524 7768 139580 12032
rect 139636 10892 139692 10902
rect 139636 10668 139692 10836
rect 139636 10602 139692 10612
rect 139748 10444 139804 12212
rect 139748 10378 139804 10388
rect 140420 11728 140476 11738
rect 140308 9212 140364 9222
rect 139412 7712 139580 7768
rect 139748 8540 139804 8550
rect 139412 7228 139468 7712
rect 139412 7162 139468 7172
rect 139524 7644 139580 7654
rect 139412 5740 139468 5750
rect 138740 4822 138796 4832
rect 139188 5292 139244 5302
rect 139188 4620 139244 5236
rect 139412 4956 139468 5684
rect 139412 4890 139468 4900
rect 139524 4888 139580 7588
rect 139748 7644 139804 8484
rect 139748 7578 139804 7588
rect 140308 5788 140364 9156
rect 140308 5722 140364 5732
rect 139524 4822 139580 4832
rect 139188 4554 139244 4564
rect 139412 4172 139468 4182
rect 138628 3612 138684 3622
rect 138516 2716 138572 2726
rect 138516 1708 138572 2660
rect 138516 1642 138572 1652
rect 138628 1484 138684 3556
rect 138740 3268 138796 3278
rect 138740 2008 138796 3212
rect 138740 1942 138796 1952
rect 138628 1418 138684 1428
rect 139412 1372 139468 4116
rect 140084 4168 140140 4178
rect 140084 2268 140140 4112
rect 140084 2202 140140 2212
rect 140308 4168 140364 4178
rect 139412 1306 139468 1316
rect 138068 1194 138124 1204
rect 140308 1148 140364 4112
rect 140420 1648 140476 11672
rect 140756 11564 140812 11586
rect 140756 11482 140812 11492
rect 141092 11004 141148 12752
rect 141204 12236 141260 12246
rect 141204 11728 141260 12180
rect 141204 11662 141260 11672
rect 141316 11900 141372 11910
rect 141316 11452 141372 11844
rect 141316 11386 141372 11396
rect 141540 11900 141596 11910
rect 141092 10938 141148 10948
rect 141428 10892 141484 10902
rect 140980 10444 141036 10454
rect 140980 10108 141036 10388
rect 141428 10332 141484 10836
rect 141428 10266 141484 10276
rect 140980 10042 141036 10052
rect 141428 10108 141484 10118
rect 140980 9772 141036 9782
rect 140532 7196 140588 7206
rect 140532 3988 140588 7140
rect 140980 6076 141036 9716
rect 141204 7980 141260 7990
rect 141204 7756 141260 7924
rect 141204 7690 141260 7700
rect 141316 6748 141372 6758
rect 140980 6020 141260 6076
rect 140980 5852 141036 5862
rect 140980 4844 141036 5796
rect 141204 5852 141260 6020
rect 141204 5786 141260 5796
rect 140980 4778 141036 4788
rect 141092 5404 141148 5414
rect 141092 4348 141148 5348
rect 141092 4282 141148 4292
rect 140532 3922 140588 3932
rect 140644 4172 140700 4182
rect 140644 3448 140700 4116
rect 141316 3988 141372 6692
rect 141204 3948 141260 3958
rect 141316 3922 141372 3932
rect 140980 3500 141036 3510
rect 140644 3392 140924 3448
rect 140868 3388 140924 3392
rect 140980 3382 141036 3392
rect 141204 3448 141260 3892
rect 141204 3382 141260 3392
rect 141428 3387 141484 10052
rect 141540 4168 141596 11844
rect 141540 4102 141596 4112
rect 141652 10108 141708 10118
rect 140868 3322 140924 3332
rect 141316 3331 141484 3387
rect 140420 1582 140476 1592
rect 140308 1082 140364 1092
rect 137732 862 137788 872
rect 138516 924 138572 934
rect 134596 634 134652 644
rect 131124 410 131180 420
rect 138516 476 138572 868
rect 141316 700 141372 3331
rect 141652 1484 141708 10052
rect 142436 9884 142492 12852
rect 142772 12908 142828 12918
rect 142772 12808 142828 12852
rect 142772 12742 142828 12752
rect 142884 12628 142940 12638
rect 142436 9818 142492 9828
rect 142660 11908 142716 11918
rect 141764 8764 141820 8774
rect 141764 6188 141820 8708
rect 142548 7756 142604 7766
rect 142436 7420 142492 7430
rect 142436 7196 142492 7364
rect 142436 7130 142492 7140
rect 141764 6122 141820 6132
rect 142548 5292 142604 7700
rect 142660 7408 142716 11852
rect 142772 10468 142828 10478
rect 142772 9996 142828 10412
rect 142884 10108 142940 12572
rect 142884 10042 142940 10052
rect 142772 9772 142828 9940
rect 142772 9706 142828 9716
rect 142772 9436 142828 9446
rect 142772 7756 142828 9380
rect 142996 7980 143052 13292
rect 145124 13168 145180 13178
rect 144116 12448 144172 12458
rect 142996 7914 143052 7924
rect 143892 11728 143948 11738
rect 142772 7690 142828 7700
rect 143556 7644 143612 7654
rect 142660 7352 142828 7408
rect 142660 7196 142716 7206
rect 142660 6524 142716 7140
rect 142660 6458 142716 6468
rect 142772 6508 142828 7352
rect 143556 7228 143612 7588
rect 143556 7172 143836 7228
rect 142772 6442 142828 6452
rect 143220 6860 143276 6870
rect 142548 5226 142604 5236
rect 142436 5068 142492 5078
rect 141652 1418 141708 1428
rect 142212 3724 142268 3734
rect 142212 1288 142268 3668
rect 142436 1596 142492 5012
rect 143220 4708 143276 6804
rect 143780 6860 143836 7172
rect 143780 6794 143836 6804
rect 143892 5608 143948 11672
rect 144004 7228 144060 7238
rect 144004 6300 144060 7172
rect 144116 6636 144172 12392
rect 144228 11728 144284 11738
rect 144228 11340 144284 11672
rect 144228 11274 144284 11284
rect 144340 11228 144396 11238
rect 144340 10108 144396 11172
rect 144340 10042 144396 10052
rect 144900 10288 144956 10298
rect 144228 9660 144284 9670
rect 144228 7980 144284 9604
rect 144228 7914 144284 7924
rect 144452 9436 144508 9446
rect 144452 7084 144508 9380
rect 144676 8540 144732 8550
rect 144452 7018 144508 7028
rect 144564 8316 144620 8326
rect 144116 6570 144172 6580
rect 144004 6234 144060 6244
rect 144228 6524 144284 6534
rect 143892 5552 144172 5608
rect 144004 5404 144060 5414
rect 143220 4642 143276 4652
rect 143444 4708 143500 4718
rect 142660 3988 142716 3998
rect 142548 3808 142604 3818
rect 142548 2828 142604 3752
rect 142660 3387 142716 3932
rect 142772 3836 142828 3846
rect 142772 3612 142828 3780
rect 142772 3546 142828 3556
rect 142660 3331 142828 3387
rect 142548 2762 142604 2772
rect 142772 2548 142828 3331
rect 142772 2482 142828 2492
rect 142884 2728 142940 2738
rect 142436 1530 142492 1540
rect 142212 1222 142268 1232
rect 142884 1148 142940 2672
rect 143444 1596 143500 4652
rect 144004 4528 144060 5348
rect 143892 4472 144060 4528
rect 143892 3628 143948 4472
rect 143892 3562 143948 3572
rect 144004 3988 144060 3998
rect 143444 1530 143500 1540
rect 144004 1596 144060 3932
rect 144116 3387 144172 5552
rect 144228 4844 144284 6468
rect 144452 6300 144508 6310
rect 144228 4778 144284 4788
rect 144340 4888 144396 4898
rect 144340 4508 144396 4832
rect 144340 4442 144396 4452
rect 144340 4348 144396 4358
rect 144452 4348 144508 6244
rect 144396 4292 144508 4348
rect 144340 4282 144396 4292
rect 144228 4060 144284 4070
rect 144228 3724 144284 4004
rect 144228 3658 144284 3668
rect 144452 3836 144508 3846
rect 144452 3628 144508 3780
rect 144340 3572 144508 3628
rect 144116 3331 144284 3387
rect 144228 3276 144284 3331
rect 144228 3210 144284 3220
rect 144004 1530 144060 1540
rect 144340 1484 144396 3572
rect 144564 3387 144620 8260
rect 144676 7308 144732 8484
rect 144676 7242 144732 7252
rect 144788 8092 144844 8102
rect 144788 5628 144844 8036
rect 144788 5562 144844 5572
rect 144900 5068 144956 10232
rect 144900 5002 144956 5012
rect 145012 8204 145068 8214
rect 144676 4888 144732 4898
rect 144676 4778 144732 4788
rect 144564 3331 144732 3387
rect 144340 1418 144396 1428
rect 144452 1596 144508 1606
rect 144004 1288 144060 1298
rect 144004 1194 144060 1204
rect 142884 1082 142940 1092
rect 144452 924 144508 1540
rect 144676 1484 144732 3331
rect 145012 1596 145068 8148
rect 145124 6860 145180 13112
rect 145684 9772 145740 14192
rect 146132 14248 146188 14258
rect 146132 13708 146188 14192
rect 149044 14068 149100 14732
rect 149268 14608 149324 14618
rect 149268 14252 149324 14552
rect 149380 14588 149548 14608
rect 149436 14552 149548 14588
rect 149380 14522 149436 14532
rect 149268 14186 149324 14196
rect 149044 14002 149100 14012
rect 149268 14068 149324 14078
rect 146020 13692 146188 13708
rect 148708 13708 148764 13718
rect 146076 13652 146188 13692
rect 147924 13692 147980 13702
rect 146020 13626 146076 13636
rect 147924 13528 147980 13636
rect 147924 13462 147980 13472
rect 148148 13692 148204 13702
rect 148148 13468 148204 13636
rect 148148 13402 148204 13412
rect 148372 13468 148428 13478
rect 148372 13348 148428 13412
rect 148372 13282 148428 13292
rect 146916 13244 146972 13254
rect 146916 13020 146972 13188
rect 146916 12954 146972 12964
rect 147588 12808 147644 12818
rect 147476 12012 147532 12022
rect 145796 11908 145852 11918
rect 145796 10444 145852 11852
rect 146132 11900 146188 11910
rect 146132 11676 146188 11844
rect 145908 11620 146188 11676
rect 145908 11368 145964 11620
rect 146020 11548 146076 11558
rect 146020 11452 146076 11492
rect 146020 11386 146076 11396
rect 145908 11302 145964 11312
rect 146132 11368 146188 11378
rect 146132 10648 146188 11312
rect 146020 10592 146188 10648
rect 146244 11228 146300 11238
rect 146020 10556 146076 10592
rect 146020 10490 146076 10500
rect 145796 10378 145852 10388
rect 145684 9706 145740 9716
rect 146132 9660 146188 9670
rect 146020 9604 146132 9660
rect 145124 6794 145180 6804
rect 145460 8428 145516 8438
rect 145460 6524 145516 8372
rect 146020 8204 146076 9604
rect 146132 9594 146188 9604
rect 146020 8138 146076 8148
rect 146020 7532 146076 7542
rect 146020 6636 146076 7476
rect 146020 6570 146076 6580
rect 145460 6458 145516 6468
rect 145348 6188 145404 6198
rect 145124 5788 145180 5798
rect 145124 5180 145180 5732
rect 145348 5628 145404 6132
rect 146244 5852 146300 11172
rect 146244 5786 146300 5796
rect 146916 7644 146972 7654
rect 146916 5852 146972 7588
rect 146916 5786 146972 5796
rect 145348 5562 145404 5572
rect 145684 5628 145740 5638
rect 145684 5292 145740 5572
rect 145684 5226 145740 5236
rect 145124 5114 145180 5124
rect 146692 4732 146748 4742
rect 146132 3724 146188 3734
rect 145572 3268 145628 3278
rect 145572 2728 145628 3212
rect 146020 3088 146076 3098
rect 146020 2940 146076 3032
rect 146020 2874 146076 2884
rect 145572 2662 145628 2672
rect 146020 2716 146076 2726
rect 146020 2548 146076 2660
rect 145684 2492 145740 2502
rect 146020 2482 146076 2492
rect 145012 1530 145068 1540
rect 145236 2008 145292 2018
rect 145236 1596 145292 1952
rect 145236 1530 145292 1540
rect 144676 1418 144732 1428
rect 145012 1288 145068 1298
rect 144452 858 144508 868
rect 144676 1036 144732 1046
rect 141316 634 141372 644
rect 144452 700 144508 710
rect 144452 568 144508 644
rect 144676 700 144732 980
rect 144676 634 144732 644
rect 145012 700 145068 1232
rect 145684 1108 145740 2436
rect 146132 1596 146188 3668
rect 146692 3724 146748 4676
rect 147364 3948 147420 3958
rect 147364 3808 147420 3892
rect 147364 3742 147420 3752
rect 146692 3658 146748 3668
rect 147476 3387 147532 11956
rect 147588 7532 147644 12752
rect 148708 12572 148764 13652
rect 149156 13132 149212 13142
rect 148708 12506 148764 12516
rect 148932 13020 148988 13030
rect 149156 12988 149212 13076
rect 148036 11900 148092 11910
rect 147700 10780 147756 10790
rect 147700 10468 147756 10724
rect 147700 10402 147756 10412
rect 147812 10648 147868 10658
rect 147812 10108 147868 10592
rect 147812 10042 147868 10052
rect 147700 9928 147756 9938
rect 147700 7980 147756 9872
rect 147700 7914 147756 7924
rect 147924 7980 147980 7990
rect 147588 7466 147644 7476
rect 147924 4348 147980 7924
rect 148036 7228 148092 11844
rect 148036 7162 148092 7172
rect 148260 11548 148316 11558
rect 147700 4292 147980 4348
rect 148036 4888 148092 4898
rect 147700 4284 147756 4292
rect 147700 4218 147756 4228
rect 147924 4168 147980 4178
rect 147812 3988 147868 3998
rect 147364 3331 147532 3387
rect 147700 3388 147756 3398
rect 147812 3387 147868 3932
rect 147756 3332 147868 3387
rect 147700 3331 147868 3332
rect 146244 3164 146300 3174
rect 146244 2548 146300 3108
rect 146244 2482 146300 2492
rect 147364 1932 147420 3331
rect 147700 3322 147756 3331
rect 147700 3164 147756 3174
rect 147588 2492 147644 2502
rect 147588 2008 147644 2436
rect 147588 1942 147644 1952
rect 147364 1866 147420 1876
rect 147700 1828 147756 3108
rect 147924 2044 147980 4112
rect 148036 3088 148092 4832
rect 148036 3022 148092 3032
rect 148260 2604 148316 11492
rect 148932 10892 148988 12964
rect 149044 12932 149212 12988
rect 149044 12012 149100 12932
rect 149044 11946 149100 11956
rect 149156 12796 149212 12806
rect 149156 11900 149212 12740
rect 149268 12684 149324 14012
rect 149492 13528 149548 14552
rect 149492 13462 149548 13472
rect 149492 13132 149548 13142
rect 149492 12796 149548 13076
rect 149492 12730 149548 12740
rect 149268 12618 149324 12628
rect 149380 12572 149660 12628
rect 149268 12448 149324 12458
rect 149380 12448 149436 12572
rect 149324 12392 149436 12448
rect 149492 12448 149548 12458
rect 149268 12382 149324 12392
rect 149156 11834 149212 11844
rect 149380 12012 149436 12022
rect 149380 11908 149436 11956
rect 149380 11842 149436 11852
rect 148932 10826 148988 10836
rect 149156 10220 149212 10230
rect 149044 9660 149100 9670
rect 148820 9604 149044 9660
rect 148484 8540 148540 8550
rect 148484 8316 148540 8484
rect 148484 8250 148540 8260
rect 148820 7644 148876 9604
rect 149044 9594 149100 9604
rect 148820 7578 148876 7588
rect 149044 7644 149100 7654
rect 149044 7084 149100 7588
rect 149044 7018 149100 7028
rect 149156 6860 149212 10164
rect 149492 9436 149548 12392
rect 149604 11908 149660 12572
rect 149604 11842 149660 11852
rect 149716 11728 149772 14732
rect 150276 14608 150332 14618
rect 150164 13708 150220 13718
rect 149492 9370 149548 9380
rect 149604 11672 149772 11728
rect 149828 13356 149884 13366
rect 149380 8428 149436 8438
rect 149380 7868 149436 8372
rect 149380 7802 149436 7812
rect 149156 6794 149212 6804
rect 149268 7420 149324 7430
rect 149268 6188 149324 7364
rect 149604 7420 149660 11672
rect 149604 7354 149660 7364
rect 149716 10780 149772 10790
rect 149492 7084 149548 7094
rect 149380 6636 149436 6646
rect 149492 6636 149548 7028
rect 149436 6580 149548 6636
rect 149380 6570 149436 6580
rect 149268 6122 149324 6132
rect 148596 5068 148652 5078
rect 148596 4974 148652 5012
rect 149492 4844 149548 4854
rect 149380 4788 149492 4844
rect 149380 4708 149436 4788
rect 149492 4778 149548 4788
rect 149380 4642 149436 4652
rect 149716 4708 149772 10724
rect 149828 4888 149884 13300
rect 149940 12684 149996 12694
rect 149940 6972 149996 12628
rect 150052 11008 150108 11018
rect 150052 10648 150108 10952
rect 150052 10582 150108 10592
rect 149940 6906 149996 6916
rect 150052 7308 150108 7318
rect 149828 4822 149884 4832
rect 149716 4642 149772 4652
rect 149604 4620 149660 4630
rect 149604 4528 149660 4564
rect 149492 4508 149548 4518
rect 149380 4452 149492 4508
rect 149604 4462 149660 4472
rect 149380 3808 149436 4452
rect 149492 4442 149548 4452
rect 149380 3742 149436 3752
rect 148260 2538 148316 2548
rect 149492 2492 149548 2502
rect 149492 2368 149548 2436
rect 149492 2302 149548 2312
rect 147700 1762 147756 1772
rect 147812 2008 147868 2018
rect 147924 1978 147980 1988
rect 150052 2044 150108 7252
rect 150052 1978 150108 1988
rect 147812 1648 147868 1952
rect 146132 1530 146188 1540
rect 147700 1592 147868 1648
rect 147924 1828 147980 1838
rect 147924 1708 147980 1772
rect 147924 1642 147980 1652
rect 145684 1042 145740 1052
rect 147700 1036 147756 1592
rect 147700 970 147756 980
rect 147924 1484 147980 1494
rect 147924 1036 147980 1428
rect 150164 1260 150220 13652
rect 150276 13168 150332 14552
rect 150276 13102 150332 13112
rect 150500 13168 150556 13178
rect 150500 12808 150556 13112
rect 150500 12742 150556 12752
rect 150276 10468 150332 10478
rect 150276 10108 150332 10412
rect 150276 10042 150332 10052
rect 150388 9436 150444 9446
rect 150388 7980 150444 9380
rect 150388 7914 150444 7924
rect 150276 5852 150332 5862
rect 150276 5404 150332 5796
rect 150276 5338 150332 5348
rect 150836 5068 150892 14912
rect 151620 14858 151676 14868
rect 151060 14700 151116 14710
rect 151060 12808 151116 14644
rect 151284 14252 151340 14262
rect 151172 14028 151228 14038
rect 151172 13888 151228 13972
rect 151172 13822 151228 13832
rect 150948 12796 151116 12808
rect 151004 12752 151116 12796
rect 150948 12730 151004 12740
rect 151284 12684 151340 14196
rect 151284 12618 151340 12628
rect 151396 13888 151452 13898
rect 151396 12268 151452 13832
rect 151396 12202 151452 12212
rect 151172 11900 151228 11910
rect 151060 11188 151116 11198
rect 151060 10668 151116 11132
rect 151172 11008 151228 11844
rect 151172 10942 151228 10952
rect 151508 11368 151564 11378
rect 151060 10602 151116 10612
rect 151284 10892 151340 10902
rect 151284 9660 151340 10836
rect 151508 10780 151564 11312
rect 151508 10714 151564 10724
rect 151284 9594 151340 9604
rect 151732 6636 151788 14912
rect 152740 14788 152796 14798
rect 152740 14252 152796 14732
rect 154420 14788 154476 14798
rect 152740 14186 152796 14196
rect 153076 14700 153132 14710
rect 153076 14252 153132 14644
rect 153076 14186 153132 14196
rect 153524 14700 153580 14710
rect 152292 13468 152348 13478
rect 151732 6570 151788 6580
rect 152180 10108 152236 10118
rect 150836 5002 150892 5012
rect 150948 5852 151004 5862
rect 150948 4888 151004 5796
rect 150948 4822 151004 4832
rect 151060 4956 151116 4966
rect 151060 4528 151116 4900
rect 151060 4462 151116 4472
rect 151060 4284 151116 4294
rect 151060 3988 151116 4228
rect 151060 3922 151116 3932
rect 150948 3808 151004 3818
rect 150612 3628 150668 3638
rect 150276 3088 150332 3098
rect 150276 1708 150332 3032
rect 150612 2380 150668 3572
rect 150948 3500 151004 3752
rect 150948 3434 151004 3444
rect 151060 3724 151116 3734
rect 151060 3268 151116 3668
rect 151060 3202 151116 3212
rect 151284 3268 151340 3278
rect 151284 2728 151340 3212
rect 151284 2662 151340 2672
rect 151508 2728 151564 2738
rect 150612 2314 150668 2324
rect 150836 2368 150892 2378
rect 150276 1642 150332 1652
rect 150724 2044 150780 2054
rect 150724 1708 150780 1988
rect 150836 1932 150892 2312
rect 151172 2268 151228 2278
rect 151060 2044 151116 2054
rect 151060 1942 151116 1952
rect 150836 1866 150892 1876
rect 150724 1642 150780 1652
rect 150164 1194 150220 1204
rect 150388 1260 150444 1270
rect 147924 970 147980 980
rect 145012 634 145068 644
rect 144900 588 144956 598
rect 144452 532 144900 568
rect 144452 512 144956 532
rect 150388 588 150444 1204
rect 151172 924 151228 2212
rect 151508 1932 151564 2672
rect 151956 2008 152012 2018
rect 151508 1866 151564 1876
rect 151732 1932 151788 1942
rect 151732 1828 151788 1876
rect 151732 1762 151788 1772
rect 151172 858 151228 868
rect 151956 924 152012 1952
rect 152180 1484 152236 10052
rect 152292 4732 152348 13412
rect 152852 12908 152908 12918
rect 152740 11564 152796 11574
rect 152740 11470 152796 11492
rect 152852 9996 152908 12852
rect 153188 11908 153244 11918
rect 153412 11908 153468 11918
rect 153244 11852 153356 11908
rect 153188 11842 153244 11852
rect 152964 11548 153020 11558
rect 152964 10288 153020 11492
rect 152964 10222 153020 10232
rect 153188 10444 153244 10454
rect 153188 10288 153244 10388
rect 153188 10222 153244 10232
rect 152852 9930 152908 9940
rect 152852 9660 152908 9670
rect 153300 9660 153356 11852
rect 153412 10108 153468 11852
rect 153524 11900 153580 14644
rect 154084 14140 154140 14150
rect 154084 12460 154140 14084
rect 154084 12394 154140 12404
rect 154308 13132 154364 13142
rect 154308 12460 154364 13076
rect 154308 12394 154364 12404
rect 153524 11834 153580 11844
rect 153412 10042 153468 10052
rect 153300 9604 154028 9660
rect 152740 8428 152796 8438
rect 152740 7532 152796 8372
rect 152852 8316 152908 9604
rect 152852 8250 152908 8260
rect 152740 7466 152796 7476
rect 153524 6524 153580 6534
rect 152740 4788 153132 4844
rect 152292 4666 152348 4676
rect 152628 4732 152684 4742
rect 152628 3448 152684 4676
rect 152740 4708 152796 4788
rect 152740 4642 152796 4652
rect 152964 4708 153020 4718
rect 152852 4348 152908 4358
rect 152852 3948 152908 4292
rect 152852 3882 152908 3892
rect 152964 3836 153020 4652
rect 153076 4528 153132 4788
rect 153524 4732 153580 6468
rect 153524 4666 153580 4676
rect 153748 4732 153804 4742
rect 153748 4528 153804 4676
rect 153076 4472 153804 4528
rect 153860 3988 153916 3998
rect 153188 3836 153244 3846
rect 152964 3770 153020 3780
rect 153076 3780 153188 3836
rect 153076 3628 153132 3780
rect 153188 3770 153244 3780
rect 152628 3382 152684 3392
rect 152740 3572 153132 3628
rect 152180 1418 152236 1428
rect 152740 1260 152796 3572
rect 153860 2268 153916 3932
rect 153860 2202 153916 2212
rect 153748 1828 153804 1838
rect 152740 1194 152796 1204
rect 152852 1484 152908 1494
rect 152852 1036 152908 1428
rect 152852 970 152908 980
rect 153748 1036 153804 1772
rect 153748 970 153804 980
rect 153972 1036 154028 9604
rect 154196 7756 154252 7766
rect 154084 7420 154140 7430
rect 154084 4888 154140 7364
rect 154196 7084 154252 7700
rect 154196 7018 154252 7028
rect 154420 6636 154476 14732
rect 156436 14788 156492 14798
rect 156100 14700 156156 14710
rect 156100 14428 156156 14644
rect 156100 14362 156156 14372
rect 156212 14476 156268 14486
rect 156212 14248 156268 14420
rect 156436 14476 156492 14732
rect 162708 14608 162764 14618
rect 156436 14410 156492 14420
rect 162036 14428 162092 14438
rect 156772 14364 156828 14374
rect 156212 14192 156492 14248
rect 156436 14028 156492 14192
rect 156436 13962 156492 13972
rect 155876 13804 155932 13814
rect 154420 6570 154476 6580
rect 154532 12808 154588 12818
rect 154532 5068 154588 12752
rect 155764 12460 155820 12470
rect 154532 5002 154588 5012
rect 154756 12268 154812 12278
rect 154756 6412 154812 12212
rect 155764 11908 155820 12404
rect 155876 12088 155932 13748
rect 156212 12460 156268 12470
rect 155876 12022 155932 12032
rect 156100 12448 156156 12458
rect 156100 12088 156156 12392
rect 156212 12236 156268 12404
rect 156212 12170 156268 12180
rect 156100 12022 156156 12032
rect 156324 12088 156380 12098
rect 155764 11842 155820 11852
rect 154644 4956 154700 4966
rect 154644 4888 154700 4900
rect 154084 4832 154700 4888
rect 154756 4888 154812 6356
rect 154756 4822 154812 4832
rect 154868 11788 154924 11798
rect 154868 4508 154924 11732
rect 155092 11788 155148 11798
rect 154980 11116 155036 11126
rect 154980 10892 155036 11060
rect 154980 10826 155036 10836
rect 154868 4442 154924 4452
rect 155092 3836 155148 11732
rect 156100 11728 156156 11738
rect 156100 11116 156156 11672
rect 156100 11050 156156 11060
rect 156212 11676 156268 11686
rect 156212 10220 156268 11620
rect 156212 10154 156268 10164
rect 156100 10108 156156 10118
rect 155988 9928 156044 9938
rect 155988 7756 156044 9872
rect 156100 8428 156156 10052
rect 156212 9928 156268 9938
rect 156324 9928 156380 12032
rect 156268 9872 156380 9928
rect 156548 9928 156604 9938
rect 156212 9862 156268 9872
rect 156100 8362 156156 8372
rect 155988 7690 156044 7700
rect 156548 7756 156604 9872
rect 156548 7690 156604 7700
rect 156324 6524 156380 6534
rect 155988 6300 156044 6310
rect 155988 5628 156044 6244
rect 156324 5788 156380 6468
rect 156772 6412 156828 14308
rect 158676 14252 158732 14262
rect 158340 13916 158396 13926
rect 158340 13822 158396 13832
rect 158564 13888 158620 13898
rect 157780 11728 157836 11738
rect 157556 10220 157612 10230
rect 157444 8540 157500 8550
rect 157108 7644 157164 7654
rect 157108 6860 157164 7588
rect 157108 6794 157164 6804
rect 156772 6076 156828 6356
rect 156772 6010 156828 6020
rect 156324 5740 157276 5788
rect 156324 5732 157220 5740
rect 157220 5674 157276 5684
rect 155988 5562 156044 5572
rect 156548 4396 156604 4406
rect 156548 4172 156604 4340
rect 156548 4106 156604 4116
rect 157444 4060 157500 8484
rect 157444 3994 157500 4004
rect 157556 3948 157612 10164
rect 157780 9772 157836 11672
rect 158564 11676 158620 13832
rect 158676 12460 158732 14196
rect 159460 14248 159516 14258
rect 159460 14028 159516 14192
rect 159460 13962 159516 13972
rect 161924 13708 161980 13718
rect 158676 12394 158732 12404
rect 161028 13244 161084 13254
rect 160580 12348 160636 12358
rect 160580 11908 160636 12292
rect 160580 11842 160636 11852
rect 158564 11610 158620 11620
rect 158788 11676 158844 11686
rect 158788 11228 158844 11620
rect 158788 11162 158844 11172
rect 159012 11228 159068 11238
rect 159012 10668 159068 11172
rect 159012 10602 159068 10612
rect 160916 11116 160972 11126
rect 157780 9706 157836 9716
rect 157892 10108 157948 10118
rect 157892 8488 157948 10052
rect 158004 10108 158060 10118
rect 158004 9884 158060 10052
rect 158004 9818 158060 9828
rect 157780 8432 157948 8488
rect 158340 9100 158396 9110
rect 157780 7868 157836 8432
rect 158340 8316 158396 9044
rect 158340 8250 158396 8260
rect 157780 7802 157836 7812
rect 159236 6076 159292 6086
rect 159236 5248 159292 6020
rect 159572 5292 159628 5302
rect 159236 5236 159572 5248
rect 159236 5192 159628 5236
rect 159460 5068 159516 5078
rect 159460 4284 159516 5012
rect 159460 4218 159516 4228
rect 160916 4168 160972 11060
rect 161028 6524 161084 13188
rect 161924 12448 161980 13652
rect 162036 13528 162092 14372
rect 162372 14248 162428 14258
rect 162036 13462 162092 13472
rect 162260 13580 162316 13590
rect 161924 12382 161980 12392
rect 162148 12908 162204 12918
rect 162036 12124 162092 12134
rect 162036 11548 162092 12068
rect 162148 12012 162204 12852
rect 162148 11946 162204 11956
rect 162260 11676 162316 13524
rect 162260 11610 162316 11620
rect 162036 11482 162092 11492
rect 162148 11340 162204 11350
rect 162148 10556 162204 11284
rect 162148 10490 162204 10500
rect 161140 10444 161196 10454
rect 161140 10108 161196 10388
rect 161140 10042 161196 10052
rect 161028 6458 161084 6468
rect 161476 5628 161532 5638
rect 161140 5516 161196 5526
rect 161140 4888 161196 5460
rect 161140 4822 161196 4832
rect 161364 4956 161420 4966
rect 161364 4620 161420 4900
rect 161364 4554 161420 4564
rect 161476 4528 161532 5572
rect 161476 4462 161532 4472
rect 162260 5516 162316 5526
rect 160916 4102 160972 4112
rect 162260 3988 162316 5460
rect 162260 3922 162316 3932
rect 157556 3882 157612 3892
rect 155092 3770 155148 3780
rect 156212 3836 156268 3846
rect 154308 3724 154364 3734
rect 154308 1596 154364 3668
rect 154644 3628 154700 3638
rect 154532 3268 154588 3278
rect 154420 2908 154476 2918
rect 154420 2492 154476 2852
rect 154420 2426 154476 2436
rect 154532 2008 154588 3212
rect 154420 1952 154588 2008
rect 154420 1932 154476 1952
rect 154420 1866 154476 1876
rect 154644 1820 154700 3572
rect 154756 3448 154812 3458
rect 154756 3164 154812 3392
rect 156212 3276 156268 3780
rect 156212 3210 156268 3220
rect 159572 3628 159628 3638
rect 154756 3098 154812 3108
rect 155876 2716 156267 2728
rect 155876 2672 156211 2716
rect 155876 2492 155932 2672
rect 156211 2650 156267 2660
rect 155876 2426 155932 2436
rect 155988 2548 156044 2558
rect 155988 1932 156044 2492
rect 156211 2548 156267 2558
rect 156211 2188 156267 2492
rect 155988 1866 156044 1876
rect 156100 2132 156267 2188
rect 157780 2380 157836 2390
rect 157780 2188 157836 2324
rect 158004 2188 158060 2198
rect 154644 1754 154700 1764
rect 154308 1530 154364 1540
rect 156100 1372 156156 2132
rect 157780 2122 157836 2132
rect 157892 2132 158004 2188
rect 157780 1828 157836 1830
rect 157892 1828 157948 2132
rect 158004 2122 158060 2132
rect 159572 1932 159628 3572
rect 159572 1866 159628 1876
rect 159684 3388 159740 3398
rect 162372 3387 162428 14192
rect 162708 14028 162764 14552
rect 178276 14428 178332 14438
rect 174132 14248 174188 14258
rect 162708 13962 162764 13972
rect 166180 14068 166236 14078
rect 172564 14068 172620 14078
rect 162596 13888 162652 13898
rect 162596 13244 162652 13832
rect 162596 13178 162652 13188
rect 163044 13528 163100 13538
rect 162708 12348 162764 12358
rect 162484 12012 162540 12022
rect 162484 4956 162540 11956
rect 162484 4890 162540 4900
rect 157780 1820 157948 1828
rect 157836 1772 157948 1820
rect 157780 1754 157836 1764
rect 159684 1596 159740 3332
rect 162260 3331 162428 3387
rect 161140 3212 161420 3268
rect 161140 3164 161196 3212
rect 161140 3098 161196 3108
rect 161364 3164 161420 3212
rect 161364 3098 161420 3108
rect 162260 3164 162316 3331
rect 162260 3098 162316 3108
rect 162484 3164 162540 3174
rect 162484 2828 162540 3108
rect 162484 2762 162540 2772
rect 162708 2828 162764 12292
rect 162932 11728 162988 11738
rect 162820 10648 162876 10658
rect 162820 10220 162876 10592
rect 162932 10288 162988 11672
rect 162932 10222 162988 10232
rect 162820 10154 162876 10164
rect 163044 8540 163100 13472
rect 165396 13356 165452 13366
rect 164948 13244 165004 13254
rect 164948 13168 165004 13188
rect 164948 13102 165004 13112
rect 165396 13020 165452 13300
rect 165396 12954 165452 12964
rect 165732 13020 165788 13030
rect 165732 12808 165788 12964
rect 165732 12742 165788 12752
rect 165956 12808 166012 12818
rect 164276 12460 164332 12470
rect 164276 12124 164332 12404
rect 164276 12058 164332 12068
rect 164500 12124 164556 12134
rect 164500 12022 164556 12032
rect 165172 12088 165228 12098
rect 163716 12012 163772 12022
rect 163380 11908 163436 11918
rect 163380 10892 163436 11852
rect 163380 10826 163436 10836
rect 162820 8484 163100 8540
rect 162820 6508 162876 8484
rect 162932 7980 162988 7990
rect 162932 7308 162988 7924
rect 162932 7242 162988 7252
rect 162820 6442 162876 6452
rect 162820 4396 162876 4406
rect 162820 3948 162876 4340
rect 162820 3882 162876 3892
rect 163156 4168 163212 4178
rect 162820 3724 162876 3734
rect 162820 3448 162876 3668
rect 162820 3382 162876 3392
rect 163044 3724 163100 3734
rect 163044 3268 163100 3668
rect 162708 2762 162764 2772
rect 162820 3212 163100 3268
rect 161251 2380 161307 2390
rect 161028 2324 161251 2368
rect 161028 2312 161307 2324
rect 161028 2156 161084 2312
rect 161028 2090 161084 2100
rect 162820 2008 162876 3212
rect 159684 1530 159740 1540
rect 162708 1952 162876 2008
rect 162708 1596 162764 1952
rect 162708 1530 162764 1540
rect 162820 1820 162876 1830
rect 156100 1306 156156 1316
rect 153972 970 154028 980
rect 151956 858 152012 868
rect 162820 924 162876 1764
rect 163156 1596 163212 4112
rect 163716 2728 163772 11956
rect 164836 11452 164892 11462
rect 164612 11004 164668 11014
rect 164612 10648 164668 10948
rect 164612 10582 164668 10592
rect 164836 10332 164892 11396
rect 164836 10266 164892 10276
rect 164948 10556 165004 10566
rect 164168 9436 164488 10252
rect 164948 10220 165004 10500
rect 164948 10154 165004 10164
rect 164168 9380 164196 9436
rect 164252 9380 164300 9436
rect 164356 9380 164404 9436
rect 164460 9380 164488 9436
rect 164168 9030 164488 9380
rect 164168 8974 164196 9030
rect 164252 8974 164300 9030
rect 164356 8974 164404 9030
rect 164460 8974 164488 9030
rect 164168 8926 164488 8974
rect 164168 8870 164196 8926
rect 164252 8870 164300 8926
rect 164356 8870 164404 8926
rect 164460 8870 164488 8926
rect 164168 8822 164488 8870
rect 164168 8766 164196 8822
rect 164252 8766 164300 8822
rect 164356 8766 164404 8822
rect 164460 8766 164488 8822
rect 164168 7868 164488 8766
rect 164168 7812 164196 7868
rect 164252 7812 164300 7868
rect 164356 7812 164404 7868
rect 164460 7812 164488 7868
rect 164168 7632 164488 7812
rect 164168 7576 164196 7632
rect 164252 7576 164300 7632
rect 164356 7576 164404 7632
rect 164460 7576 164488 7632
rect 164168 7528 164488 7576
rect 164168 7472 164196 7528
rect 164252 7472 164300 7528
rect 164356 7472 164404 7528
rect 164460 7472 164488 7528
rect 164168 7424 164488 7472
rect 164168 7368 164196 7424
rect 164252 7368 164300 7424
rect 164356 7368 164404 7424
rect 164460 7368 164488 7424
rect 164168 6300 164488 7368
rect 164724 10108 164780 10118
rect 164168 6244 164196 6300
rect 164252 6244 164300 6300
rect 164356 6244 164404 6300
rect 164460 6244 164488 6300
rect 164168 6234 164488 6244
rect 164168 6178 164196 6234
rect 164252 6178 164300 6234
rect 164356 6178 164404 6234
rect 164460 6178 164488 6234
rect 164168 6130 164488 6178
rect 164168 6074 164196 6130
rect 164252 6074 164300 6130
rect 164356 6074 164404 6130
rect 164460 6074 164488 6130
rect 164168 6026 164488 6074
rect 164168 5970 164196 6026
rect 164252 5970 164300 6026
rect 164356 5970 164404 6026
rect 164460 5970 164488 6026
rect 164168 4732 164488 5970
rect 164612 6300 164668 6310
rect 164612 4888 164668 6244
rect 164612 4822 164668 4832
rect 164168 4676 164196 4732
rect 164252 4676 164300 4732
rect 164356 4676 164404 4732
rect 164460 4676 164488 4732
rect 164168 4644 164488 4676
rect 164724 4508 164780 10052
rect 165172 6412 165228 12032
rect 165956 10468 166012 12752
rect 166180 11548 166236 14012
rect 166852 14028 166908 14038
rect 166292 13168 166348 13178
rect 166292 12012 166348 13112
rect 166292 11946 166348 11956
rect 166516 12460 166572 12470
rect 166516 12012 166572 12404
rect 166516 11946 166572 11956
rect 166628 11908 166684 11918
rect 166180 11492 166460 11548
rect 165956 10402 166012 10412
rect 166292 9996 166348 10006
rect 166292 7868 166348 9940
rect 166404 7980 166460 11492
rect 166628 11004 166684 11852
rect 166740 11340 166796 11350
rect 166740 11116 166796 11284
rect 166740 11050 166796 11060
rect 166628 10938 166684 10948
rect 166404 7914 166460 7924
rect 166628 10332 166684 10342
rect 166292 7802 166348 7812
rect 165172 4732 165228 6356
rect 166292 6524 166348 6534
rect 166292 4888 166348 6468
rect 166516 6076 166572 6086
rect 165172 4666 165228 4676
rect 166180 4832 166348 4888
rect 166404 5964 166460 5974
rect 164724 4442 164780 4452
rect 164836 4528 164892 4538
rect 163716 2662 163772 2672
rect 163156 1530 163212 1540
rect 164724 1932 164780 1942
rect 164500 1484 164556 1494
rect 164724 1484 164780 1876
rect 164836 1596 164892 4472
rect 165620 3808 165676 3818
rect 165620 2728 165676 3752
rect 165620 2662 165676 2672
rect 164836 1530 164892 1540
rect 164948 1932 165004 1942
rect 164556 1428 164668 1468
rect 164500 1412 164668 1428
rect 164724 1418 164780 1428
rect 164612 1288 164668 1412
rect 164948 1288 165004 1876
rect 166180 1372 166236 4832
rect 166292 3448 166348 3458
rect 166292 2828 166348 3392
rect 166404 3276 166460 5908
rect 166404 3210 166460 3220
rect 166292 2762 166348 2772
rect 166516 1596 166572 6020
rect 166628 2908 166684 10276
rect 166852 6636 166908 13972
rect 172452 13916 172508 13926
rect 167972 13468 168028 13478
rect 167748 13348 167804 13358
rect 167972 13348 168028 13412
rect 167804 13292 168028 13348
rect 172452 13356 172508 13860
rect 167748 13282 167804 13292
rect 166852 6570 166908 6580
rect 167636 11908 167692 11918
rect 167636 6636 167692 11852
rect 167860 10332 167916 13292
rect 172452 13290 172508 13300
rect 168532 12448 168588 12458
rect 168532 11564 168588 12392
rect 171220 12448 171276 12458
rect 171220 12348 171276 12392
rect 171220 12282 171276 12292
rect 172228 12348 172284 12358
rect 172228 12268 172284 12292
rect 172228 12202 172284 12212
rect 168532 11498 168588 11508
rect 168868 11900 168924 11910
rect 167860 10266 167916 10276
rect 167860 8316 167916 8326
rect 167860 7756 167916 8260
rect 167860 7690 167916 7700
rect 167636 6570 167692 6580
rect 168644 6524 168700 6534
rect 168644 6300 168700 6468
rect 168644 6234 168700 6244
rect 166740 5180 166796 5190
rect 166740 5068 166796 5124
rect 166740 5002 166796 5012
rect 167860 4508 167916 4518
rect 166628 2842 166684 2852
rect 167076 3388 167132 3398
rect 167076 2908 167132 3332
rect 167860 3088 167916 4452
rect 167860 3022 167916 3032
rect 168084 3988 168140 3998
rect 167076 2842 167132 2852
rect 168084 2044 168140 3932
rect 168084 1978 168140 1988
rect 168644 3388 168700 3398
rect 168868 3387 168924 11844
rect 172564 11900 172620 14012
rect 174020 13692 174076 13702
rect 173572 13580 173628 13590
rect 173572 13168 173628 13524
rect 173572 13112 173740 13168
rect 173684 12796 173740 13112
rect 173684 12730 173740 12740
rect 173796 12908 173852 12918
rect 172564 11834 172620 11844
rect 173796 11900 173852 12852
rect 174020 12684 174076 13636
rect 174020 12618 174076 12628
rect 174132 13168 174188 14192
rect 174468 13916 174524 13926
rect 174468 13822 174524 13832
rect 175028 13888 175084 13898
rect 173796 11834 173852 11844
rect 170996 11564 171052 11574
rect 168980 9212 169036 9222
rect 168980 8988 169036 9156
rect 168980 8922 169036 8932
rect 170996 9100 171052 11508
rect 173348 10648 173404 10658
rect 166516 1530 166572 1540
rect 167972 1932 168028 1942
rect 167972 1468 168028 1876
rect 167972 1402 168028 1412
rect 166180 1306 166236 1316
rect 164612 1232 165004 1288
rect 168644 1148 168700 3332
rect 168756 3331 168924 3387
rect 170436 8540 170492 8550
rect 168756 3164 168812 3331
rect 170436 3268 170492 8484
rect 170996 6688 171052 9044
rect 173124 10332 173180 10342
rect 172900 8764 172956 8774
rect 172900 7308 172956 8708
rect 172900 7242 172956 7252
rect 170884 6632 171052 6688
rect 170884 4708 170940 6632
rect 170996 6524 171052 6534
rect 170996 6076 171052 6468
rect 170996 6010 171052 6020
rect 170884 4642 170940 4652
rect 171444 4708 171500 4718
rect 170436 3202 170492 3212
rect 168756 3098 168812 3108
rect 168644 1082 168700 1092
rect 162820 858 162876 868
rect 171444 924 171500 4652
rect 173124 2380 173180 10276
rect 173348 10108 173404 10592
rect 173348 9100 173404 10052
rect 173348 9034 173404 9044
rect 173908 7084 173964 7094
rect 173796 6412 173852 6422
rect 173796 5628 173852 6356
rect 173908 6188 173964 7028
rect 174132 6412 174188 13112
rect 174244 12684 174300 12694
rect 174244 12460 174300 12628
rect 174244 12394 174300 12404
rect 174468 12460 174524 12470
rect 174132 6346 174188 6356
rect 174356 12268 174412 12278
rect 173908 6122 173964 6132
rect 173796 5562 173852 5572
rect 174132 3052 174188 3062
rect 174132 2716 174188 2996
rect 174132 2650 174188 2660
rect 174356 2716 174412 12212
rect 174468 11788 174524 12404
rect 174468 11722 174524 11732
rect 174692 9884 174748 9894
rect 174692 6076 174748 9828
rect 175028 8092 175084 13832
rect 178052 13528 178108 13538
rect 175028 8026 175084 8036
rect 175140 12988 175196 12998
rect 174692 6010 174748 6020
rect 175140 6076 175196 12932
rect 177716 12988 177772 12998
rect 177716 7756 177772 12932
rect 178052 9996 178108 13472
rect 178052 9930 178108 9940
rect 178164 10468 178220 10478
rect 177716 7690 177772 7700
rect 178164 9212 178220 10412
rect 176148 7644 176204 7654
rect 176148 6860 176204 7588
rect 176148 6794 176204 6804
rect 177940 7308 177996 7318
rect 175140 6010 175196 6020
rect 177940 5404 177996 7252
rect 177940 5338 177996 5348
rect 177716 5180 177772 5190
rect 177716 4888 177772 5124
rect 177716 4822 177772 4832
rect 178052 5180 178108 5190
rect 174356 2650 174412 2660
rect 174916 4348 174972 4358
rect 173124 2314 173180 2324
rect 174916 2380 174972 4292
rect 178052 3988 178108 5124
rect 178052 3922 178108 3932
rect 174916 2314 174972 2324
rect 175140 3808 175196 3818
rect 175140 1596 175196 3752
rect 178164 2368 178220 9156
rect 178276 6636 178332 14372
rect 182756 14364 182812 14374
rect 179620 13528 179676 13538
rect 178836 12236 178892 12246
rect 178836 12088 178892 12180
rect 178836 12022 178892 12032
rect 179620 11116 179676 13472
rect 180852 12684 180908 12694
rect 180852 12348 180908 12628
rect 180852 12282 180908 12292
rect 178836 9928 178892 9938
rect 178836 6972 178892 9872
rect 178836 6906 178892 6916
rect 179060 9928 179116 9938
rect 178276 6570 178332 6580
rect 178276 4284 178332 4294
rect 178276 4168 178332 4228
rect 178276 4102 178332 4112
rect 179060 2492 179116 9872
rect 179620 6636 179676 11060
rect 180404 11908 180460 11918
rect 179620 6570 179676 6580
rect 179844 6636 179900 6646
rect 179732 6524 179788 6534
rect 179844 6508 179900 6580
rect 179788 6468 179900 6508
rect 179732 6452 179900 6468
rect 179956 6524 180012 6534
rect 179620 6188 179676 6198
rect 179956 6148 180012 6468
rect 179676 6132 180012 6148
rect 179620 6092 180012 6132
rect 179396 4956 179452 4966
rect 179396 4348 179452 4900
rect 179060 2426 179116 2436
rect 179284 2492 179340 2502
rect 178164 2302 178220 2312
rect 179284 2156 179340 2436
rect 179284 2090 179340 2100
rect 175140 1530 175196 1540
rect 179396 1596 179452 4292
rect 180180 4844 180236 4854
rect 180180 3948 180236 4788
rect 180404 4844 180460 11852
rect 182644 11908 182700 11918
rect 180852 11368 180908 11378
rect 180852 9212 180908 11312
rect 180964 10892 181020 10902
rect 180964 10332 181020 10836
rect 180964 10266 181020 10276
rect 180852 9146 180908 9156
rect 181300 8540 181356 8550
rect 181076 8092 181132 8102
rect 181076 7868 181132 8036
rect 181300 8092 181356 8484
rect 181300 8026 181356 8036
rect 181860 8540 181916 8550
rect 181076 7802 181132 7812
rect 181300 5404 181356 5414
rect 180404 4778 180460 4788
rect 180628 4888 180684 4898
rect 180180 3882 180236 3892
rect 180404 4396 180460 4406
rect 180404 4168 180460 4340
rect 179620 3276 179676 3286
rect 179620 2368 179676 3220
rect 179620 2302 179676 2312
rect 179396 1530 179452 1540
rect 180404 1596 180460 4112
rect 180404 1530 180460 1540
rect 180628 1484 180684 4832
rect 181300 3448 181356 5348
rect 181524 3988 181580 3998
rect 181300 3382 181356 3392
rect 181412 3628 181468 3638
rect 181412 3088 181468 3572
rect 181412 3022 181468 3032
rect 181524 2548 181580 3932
rect 181860 3052 181916 8484
rect 182644 6860 182700 11852
rect 182756 10648 182812 14308
rect 191156 14068 191212 14078
rect 191156 13962 191212 13972
rect 193396 13916 193452 13926
rect 193396 13822 193452 13832
rect 183204 13804 183260 13814
rect 183204 13708 183260 13748
rect 183204 13642 183260 13652
rect 191828 13528 191884 13538
rect 187572 13468 187628 13478
rect 185332 13020 185388 13030
rect 185332 12448 185388 12964
rect 185332 12382 185388 12392
rect 187012 12348 187068 12358
rect 187012 11900 187068 12292
rect 187012 11834 187068 11844
rect 185108 11728 185164 11738
rect 182980 11676 183036 11686
rect 182756 9884 182812 10592
rect 182756 9818 182812 9828
rect 182868 11228 182924 11238
rect 182868 9548 182924 11172
rect 182868 9482 182924 9492
rect 182980 9436 183036 11620
rect 183428 11452 183484 11462
rect 183428 10444 183484 11396
rect 183428 10378 183484 10388
rect 183988 11368 184044 11378
rect 183988 10288 184044 11312
rect 184996 11188 185052 11198
rect 182980 9370 183036 9380
rect 183764 10220 183820 10230
rect 183988 10222 184044 10232
rect 184324 10892 184380 10902
rect 183764 9436 183820 10164
rect 184324 10108 184380 10836
rect 184324 10042 184380 10052
rect 184996 10288 185052 11132
rect 184996 9884 185052 10232
rect 184996 9818 185052 9828
rect 183764 9370 183820 9380
rect 185108 8316 185164 11672
rect 187572 11548 187628 13412
rect 190036 12448 190092 12458
rect 187460 11116 187516 11126
rect 186452 10108 186508 10118
rect 186452 9884 186508 10052
rect 186452 9818 186508 9828
rect 185108 8250 185164 8260
rect 182644 6794 182700 6804
rect 182980 7756 183036 7766
rect 182196 4844 182252 4854
rect 182196 4528 182252 4788
rect 182196 4462 182252 4472
rect 182980 3988 183036 7700
rect 186340 7172 186620 7228
rect 182980 3922 183036 3932
rect 183092 4528 183148 4538
rect 181860 2986 181916 2996
rect 183092 2940 183148 4472
rect 186340 4168 186396 7172
rect 186564 7084 186620 7172
rect 186788 7084 186844 7094
rect 186564 7028 186788 7084
rect 186788 7018 186844 7028
rect 186340 4102 186396 4112
rect 186452 6972 186508 6982
rect 184660 3392 184828 3448
rect 184660 3276 184716 3392
rect 184772 3387 184828 3392
rect 184772 3331 185276 3387
rect 184660 3210 184716 3220
rect 185220 3164 185276 3331
rect 185220 3098 185276 3108
rect 186116 3268 186172 3278
rect 183092 2874 183148 2884
rect 184436 3052 184492 3062
rect 181524 2482 181580 2492
rect 183092 2548 183148 2558
rect 184436 2548 184492 2996
rect 184436 2482 184492 2492
rect 185892 2940 185948 2950
rect 183092 2426 183148 2436
rect 185892 2008 185948 2884
rect 185892 1942 185948 1952
rect 186116 1596 186172 3212
rect 186452 2008 186508 6916
rect 187460 3387 187516 11060
rect 187572 8316 187628 11492
rect 187908 12088 187964 12098
rect 187572 8250 187628 8260
rect 187796 11004 187852 11014
rect 187460 3331 187740 3387
rect 186452 1942 186508 1952
rect 187348 3276 187404 3306
rect 187348 1828 187404 3212
rect 187348 1762 187404 1772
rect 187684 1828 187740 3331
rect 187796 3276 187852 10948
rect 187908 5628 187964 12032
rect 189812 11452 189868 11462
rect 188356 11368 188412 11378
rect 188020 10668 188076 10678
rect 188020 8764 188076 10612
rect 188020 8698 188076 8708
rect 188244 9660 188300 9670
rect 188244 6748 188300 9604
rect 188244 6682 188300 6692
rect 187908 5562 187964 5572
rect 187796 3210 187852 3220
rect 187684 1762 187740 1772
rect 187908 2908 187964 2918
rect 186116 1530 186172 1540
rect 187908 1596 187964 2852
rect 188356 2908 188412 11312
rect 189812 11188 189868 11396
rect 189812 11122 189868 11132
rect 189924 9660 189980 9670
rect 188916 7756 188972 7766
rect 188356 2842 188412 2852
rect 188692 5628 188748 5638
rect 188692 2156 188748 5572
rect 188916 5068 188972 7700
rect 189812 6636 189868 6646
rect 189812 6508 189868 6580
rect 189364 6452 189868 6508
rect 189364 6412 189420 6452
rect 189364 6346 189420 6356
rect 188916 4528 188972 5012
rect 188916 4462 188972 4472
rect 189252 4620 189308 4630
rect 189252 4528 189308 4564
rect 189252 4462 189308 4472
rect 189588 4620 189644 4630
rect 189588 3448 189644 4564
rect 189924 4620 189980 9604
rect 190036 4956 190092 12392
rect 190036 4890 190092 4900
rect 190148 11728 190204 11738
rect 189924 4554 189980 4564
rect 189588 3382 189644 3392
rect 190148 3388 190204 11672
rect 191716 11564 191772 11574
rect 190820 11188 190876 11198
rect 190148 3322 190204 3332
rect 190596 10108 190652 10118
rect 188468 2008 188524 2018
rect 188468 1828 188524 1952
rect 188692 2008 188748 2100
rect 188916 2940 188972 2950
rect 188916 2156 188972 2884
rect 190596 2828 190652 10052
rect 190820 7644 190876 11132
rect 190932 10220 190988 10230
rect 190932 10108 190988 10164
rect 190932 9212 190988 10052
rect 191332 10220 191652 10252
rect 191332 10164 191360 10220
rect 191416 10164 191464 10220
rect 191520 10164 191568 10220
rect 191624 10164 191652 10220
rect 191332 9729 191652 10164
rect 191332 9673 191360 9729
rect 191416 9673 191464 9729
rect 191520 9673 191568 9729
rect 191624 9673 191652 9729
rect 191332 9625 191652 9673
rect 191332 9569 191360 9625
rect 191416 9569 191464 9625
rect 191520 9569 191568 9625
rect 191624 9569 191652 9625
rect 191332 9521 191652 9569
rect 191332 9465 191360 9521
rect 191416 9465 191464 9521
rect 191520 9465 191568 9521
rect 191624 9465 191652 9521
rect 190932 9146 190988 9156
rect 191044 9324 191100 9334
rect 191044 8428 191100 9268
rect 191044 8362 191100 8372
rect 191332 8652 191652 9465
rect 191332 8596 191360 8652
rect 191416 8596 191464 8652
rect 191520 8596 191568 8652
rect 191624 8596 191652 8652
rect 190820 7578 190876 7588
rect 191332 8331 191652 8596
rect 191332 8275 191360 8331
rect 191416 8275 191464 8331
rect 191520 8275 191568 8331
rect 191624 8275 191652 8331
rect 191332 8227 191652 8275
rect 191332 8171 191360 8227
rect 191416 8171 191464 8227
rect 191520 8171 191568 8227
rect 191624 8171 191652 8227
rect 191332 8123 191652 8171
rect 191332 8067 191360 8123
rect 191416 8067 191464 8123
rect 191520 8067 191568 8123
rect 191624 8067 191652 8123
rect 191332 7084 191652 8067
rect 191332 7028 191360 7084
rect 191416 7028 191464 7084
rect 191520 7028 191568 7084
rect 191624 7028 191652 7084
rect 191332 6933 191652 7028
rect 191332 6877 191360 6933
rect 191416 6877 191464 6933
rect 191520 6877 191568 6933
rect 191624 6877 191652 6933
rect 191332 6829 191652 6877
rect 191332 6773 191360 6829
rect 191416 6773 191464 6829
rect 191520 6773 191568 6829
rect 191624 6773 191652 6829
rect 191332 6725 191652 6773
rect 191332 6669 191360 6725
rect 191416 6669 191464 6725
rect 191520 6669 191568 6725
rect 191624 6669 191652 6725
rect 191716 7756 191772 11508
rect 191716 6748 191772 7700
rect 191716 6682 191772 6692
rect 191332 5535 191652 6669
rect 191828 6300 191884 13472
rect 197540 13348 197596 13358
rect 193284 13168 193340 13178
rect 192164 10288 192220 10298
rect 192164 9772 192220 10232
rect 192164 9706 192220 9716
rect 193060 9928 193116 9938
rect 193060 8092 193116 9872
rect 193060 8026 193116 8036
rect 193172 8764 193228 8774
rect 192836 7532 192892 7542
rect 192836 6524 192892 7476
rect 192836 6458 192892 6468
rect 193172 6412 193228 8708
rect 193172 6346 193228 6356
rect 191828 6234 191884 6244
rect 193284 6076 193340 13112
rect 195524 13020 195580 13030
rect 195524 12922 195580 12932
rect 196532 12908 196588 12918
rect 193844 12684 193900 12694
rect 193844 12460 193900 12628
rect 193844 12394 193900 12404
rect 195412 12572 195468 12582
rect 194852 12124 194908 12134
rect 194740 11548 194796 11558
rect 193844 10828 193900 10838
rect 193844 9212 193900 10772
rect 193844 9146 193900 9156
rect 194292 10444 194348 10454
rect 193732 8540 193788 8550
rect 193732 6524 193788 8484
rect 193732 6458 193788 6468
rect 194292 6300 194348 10388
rect 194740 9772 194796 11492
rect 194740 9706 194796 9716
rect 194292 6234 194348 6244
rect 193284 6010 193340 6020
rect 194852 6076 194908 12068
rect 195412 9212 195468 12516
rect 195412 9146 195468 9156
rect 194852 6010 194908 6020
rect 196420 7756 196476 7766
rect 196420 6748 196476 7700
rect 191332 5460 191360 5535
rect 191416 5460 191464 5535
rect 191520 5460 191568 5535
rect 191624 5460 191652 5535
rect 191332 5431 191652 5460
rect 191332 5375 191360 5431
rect 191416 5375 191464 5431
rect 191520 5375 191568 5431
rect 191624 5375 191652 5431
rect 191332 5327 191652 5375
rect 191332 5271 191360 5327
rect 191416 5271 191464 5327
rect 191520 5271 191568 5327
rect 191624 5271 191652 5327
rect 191332 4644 191652 5271
rect 191940 4956 191996 4966
rect 191940 4888 191996 4900
rect 191940 4822 191996 4832
rect 193172 4956 193228 4966
rect 192164 4620 192220 4630
rect 192164 4528 192220 4564
rect 192052 4472 192220 4528
rect 191492 4292 191772 4348
rect 191492 4284 191548 4292
rect 191492 4218 191548 4228
rect 191492 4060 191548 4070
rect 190596 2762 190652 2772
rect 190708 2908 190764 2918
rect 188916 2090 188972 2100
rect 189140 2728 189196 2738
rect 188692 1942 188748 1952
rect 188692 1828 188748 1830
rect 188468 1820 188748 1828
rect 188468 1772 188692 1820
rect 188692 1754 188748 1764
rect 187908 1530 187964 1540
rect 189140 1596 189196 2672
rect 190708 2548 190764 2852
rect 189252 2492 189308 2502
rect 190708 2482 190764 2492
rect 189252 2008 189308 2436
rect 191492 2188 191548 4004
rect 191716 3948 191772 4292
rect 192052 4060 192108 4472
rect 193172 4348 193228 4900
rect 193172 4282 193228 4292
rect 194852 4956 194908 4966
rect 192052 3994 192108 4004
rect 192276 4060 192332 4070
rect 191716 3882 191772 3892
rect 192276 3387 192332 4004
rect 194852 3988 194908 4900
rect 194852 3922 194908 3932
rect 194964 3836 195020 3846
rect 194964 3628 195020 3780
rect 194964 3562 195020 3572
rect 191604 3331 192332 3387
rect 191604 2368 191660 3331
rect 191604 2302 191660 2312
rect 194068 2940 194124 2950
rect 191492 2122 191548 2132
rect 191716 2188 191772 2198
rect 189252 1952 189980 2008
rect 189924 1932 189980 1952
rect 189924 1866 189980 1876
rect 191716 1820 191772 2132
rect 191716 1754 191772 1764
rect 189140 1530 189196 1540
rect 180628 1418 180684 1428
rect 190596 1484 190652 1494
rect 190596 1148 190652 1428
rect 194068 1288 194124 2884
rect 196420 1596 196476 6692
rect 196532 6636 196588 12852
rect 197316 11228 197372 11238
rect 196644 10648 196700 10658
rect 196644 7644 196700 10592
rect 197316 10108 197372 11172
rect 197316 10042 197372 10052
rect 197540 8316 197596 13292
rect 211652 13356 211708 13366
rect 203252 12808 203308 12818
rect 200900 12684 200956 12694
rect 197764 12124 197820 12134
rect 197764 11908 197820 12068
rect 197764 11842 197820 11852
rect 198436 11900 198492 11910
rect 198212 10468 198268 10478
rect 197988 10108 198044 10118
rect 197540 8250 197596 8260
rect 197764 9660 197820 9670
rect 196644 7578 196700 7588
rect 196532 6570 196588 6580
rect 197764 6300 197820 9604
rect 197988 9660 198044 10052
rect 198212 9884 198268 10412
rect 198212 9818 198268 9828
rect 197988 9212 198044 9604
rect 197988 9146 198044 9156
rect 197764 5740 197820 6244
rect 197764 5674 197820 5684
rect 198212 7420 198268 7430
rect 197876 4732 197932 4742
rect 197876 4638 197932 4652
rect 198212 2908 198268 7364
rect 198436 4732 198492 11844
rect 200340 10288 200396 10298
rect 200340 9884 200396 10232
rect 200340 9818 200396 9828
rect 199892 9436 199948 9446
rect 198436 4666 198492 4676
rect 199444 8652 199500 8662
rect 198212 2842 198268 2852
rect 197652 2728 197708 2738
rect 197540 2604 197596 2614
rect 196420 1530 196476 1540
rect 197316 2188 197372 2198
rect 194068 1222 194124 1232
rect 190596 1082 190652 1092
rect 192836 1148 192892 1158
rect 171444 858 171500 868
rect 192836 928 192892 1092
rect 195188 1108 195244 1118
rect 192836 862 192892 872
rect 194068 1036 194124 1046
rect 150388 522 150444 532
rect 151060 748 151116 758
rect 151060 588 151116 692
rect 194068 700 194124 980
rect 195188 1036 195244 1052
rect 195188 970 195244 980
rect 197092 1036 197148 1046
rect 194068 634 194124 644
rect 151060 522 151116 532
rect 138516 410 138572 420
rect 197092 388 197148 980
rect 197092 322 197148 332
rect 197316 388 197372 2132
rect 197540 1148 197596 2548
rect 197540 1082 197596 1092
rect 197652 1036 197708 2672
rect 197652 970 197708 980
rect 198212 1828 198268 1838
rect 198212 928 198268 1772
rect 199444 1596 199500 8596
rect 199892 8316 199948 9380
rect 199892 8250 199948 8260
rect 200116 8540 200172 8550
rect 200004 7308 200060 7318
rect 200004 6748 200060 7252
rect 200004 6682 200060 6692
rect 199444 1530 199500 1540
rect 200116 1596 200172 8484
rect 200900 6636 200956 12628
rect 201908 8988 201964 8998
rect 201908 8652 201964 8932
rect 201908 8586 201964 8596
rect 200900 6412 200956 6580
rect 200900 6346 200956 6356
rect 201572 7420 201628 7430
rect 201572 3268 201628 7364
rect 203252 6300 203308 12752
rect 208292 12628 208348 12638
rect 206948 12088 207004 12098
rect 206948 11900 207004 12032
rect 206948 11834 207004 11844
rect 204484 11008 204540 11018
rect 204484 9772 204540 10952
rect 204484 9706 204540 9716
rect 205716 9548 205772 9558
rect 203252 6234 203308 6244
rect 203700 7980 203756 7990
rect 203700 4888 203756 7924
rect 203924 7980 203980 7990
rect 203924 7532 203980 7924
rect 203924 7466 203980 7476
rect 205716 6076 205772 9492
rect 206388 9548 206444 9558
rect 206388 8988 206444 9492
rect 206388 8922 206444 8932
rect 205716 6010 205772 6020
rect 203700 4822 203756 4832
rect 201572 3202 201628 3212
rect 200116 1530 200172 1540
rect 201572 2492 201628 2502
rect 201572 1468 201628 2436
rect 203588 2268 203644 2278
rect 203588 2188 203644 2212
rect 203588 2122 203644 2132
rect 204372 1648 204428 1658
rect 204372 1530 204428 1540
rect 201572 1402 201628 1412
rect 198212 862 198268 872
rect 203028 1288 203084 1298
rect 203028 924 203084 1232
rect 208292 1260 208348 12572
rect 210308 12268 210364 12278
rect 208404 8988 208460 8998
rect 208404 7868 208460 8932
rect 208404 7802 208460 7812
rect 210308 5852 210364 12212
rect 211204 10288 211260 10298
rect 211204 7420 211260 10232
rect 211204 7354 211260 7364
rect 210308 5786 210364 5796
rect 211316 5404 211372 5414
rect 209972 4956 210028 4966
rect 209972 4528 210028 4900
rect 209972 4462 210028 4472
rect 209636 3836 209692 3846
rect 209636 3742 209692 3752
rect 211316 3088 211372 5348
rect 211316 3022 211372 3032
rect 211652 1596 211708 13300
rect 212996 12236 213052 12246
rect 212548 9212 212604 9222
rect 212548 8764 212604 9156
rect 212548 8698 212604 8708
rect 212548 6188 212604 6198
rect 212548 5740 212604 6132
rect 212548 5674 212604 5684
rect 212772 5740 212828 5750
rect 211764 4956 211820 4966
rect 211764 4888 211820 4900
rect 211764 4822 211820 4832
rect 212772 3448 212828 5684
rect 212996 5740 213052 12180
rect 216356 8092 216412 8102
rect 212996 5674 213052 5684
rect 214452 7420 214508 7430
rect 212772 3382 212828 3392
rect 211652 1530 211708 1540
rect 211092 1468 211148 1478
rect 211092 1372 211148 1412
rect 211092 1306 211148 1316
rect 214452 1372 214508 7364
rect 214452 1306 214508 1316
rect 208292 1194 208348 1204
rect 216356 1148 216412 8036
rect 216356 1082 216412 1092
rect 203028 858 203084 868
rect 205604 924 205660 934
rect 205604 568 205660 868
rect 205604 502 205660 512
rect 206836 924 206892 934
rect 197316 322 197372 332
rect 127540 298 127596 308
rect 113652 152 117068 208
rect 206836 208 206892 868
rect 212884 928 212940 962
rect 212884 858 212940 868
rect 217140 924 217196 934
rect 217140 388 217196 868
rect 217140 322 217196 332
rect 67732 142 67788 152
rect 77364 142 77420 152
rect 77588 142 77644 152
rect 206836 142 206892 152
rect 65940 74 65996 84
<< via4 >>
rect 60452 14912 60508 14968
rect 49140 14732 49196 14788
rect 21476 14552 21532 14608
rect 17780 14192 17836 14248
rect 14868 14028 14924 14068
rect 14868 14012 14924 14028
rect 25060 13652 25116 13708
rect 43204 13832 43260 13888
rect 10500 13524 10556 13528
rect 10500 13472 10556 13524
rect 25732 13292 25788 13348
rect 18452 13112 18508 13168
rect 34468 12964 34524 12988
rect 34468 12932 34524 12964
rect 27972 12752 28028 12808
rect 27188 12572 27244 12628
rect 30100 12392 30156 12448
rect 42196 12212 42252 12268
rect 26740 11672 26796 11728
rect 22708 10952 22764 11008
rect 10276 10772 10332 10828
rect 9604 3932 9660 3988
rect 2548 1232 2604 1288
rect 1316 1052 1372 1108
rect 16212 10232 16268 10288
rect 21700 9872 21756 9928
rect 11620 4292 11676 4348
rect 1988 512 2044 568
rect 16436 4112 16492 4168
rect 17780 2852 17836 2908
rect 18452 2492 18508 2548
rect 18228 872 18284 928
rect 18116 692 18172 748
rect 29988 10592 30044 10648
rect 28376 9673 28432 9729
rect 28480 9673 28536 9729
rect 28584 9673 28640 9729
rect 28376 9569 28432 9625
rect 28480 9569 28536 9625
rect 28584 9569 28640 9625
rect 28376 9465 28432 9521
rect 28480 9465 28536 9521
rect 28584 9465 28640 9521
rect 23044 1232 23100 1288
rect 21140 1052 21196 1108
rect 25172 2672 25228 2728
rect 23380 512 23436 568
rect 28376 8275 28432 8331
rect 28480 8275 28536 8331
rect 28584 8275 28640 8331
rect 28376 8171 28432 8227
rect 28480 8171 28536 8227
rect 28584 8171 28640 8227
rect 28376 8067 28432 8123
rect 28480 8067 28536 8123
rect 28584 8067 28640 8123
rect 28376 6877 28432 6933
rect 28480 6877 28536 6933
rect 28584 6877 28640 6933
rect 28376 6773 28432 6829
rect 28480 6773 28536 6829
rect 28584 6773 28640 6829
rect 28376 6669 28432 6725
rect 28480 6669 28536 6725
rect 28584 6669 28640 6725
rect 28376 5516 28432 5535
rect 28376 5479 28432 5516
rect 28480 5516 28536 5535
rect 28480 5479 28536 5516
rect 28584 5516 28640 5535
rect 28584 5479 28640 5516
rect 28376 5375 28432 5431
rect 28480 5375 28536 5431
rect 28584 5375 28640 5431
rect 28376 5271 28432 5327
rect 28480 5271 28536 5327
rect 28584 5271 28640 5327
rect 28756 3032 28812 3088
rect 36820 10412 36876 10468
rect 44548 11312 44604 11368
rect 46228 11132 46284 11188
rect 46116 10052 46172 10108
rect 53844 14372 53900 14428
rect 57092 13832 57148 13888
rect 53844 13652 53900 13708
rect 56644 13652 56700 13708
rect 53844 13292 53900 13348
rect 54068 13292 54124 13348
rect 53060 12752 53116 12808
rect 53396 12752 53452 12808
rect 26404 1052 26460 1108
rect 33908 3212 33964 3268
rect 34244 3392 34300 3448
rect 33684 2132 33740 2188
rect 35476 3572 35532 3628
rect 34580 1412 34636 1468
rect 35700 4652 35756 4708
rect 42420 1232 42476 1288
rect 40404 924 40460 928
rect 40404 872 40460 924
rect 40964 692 41020 748
rect 49252 3752 49308 3808
rect 49252 3032 49308 3088
rect 49700 3212 49756 3268
rect 49028 2852 49084 2908
rect 49028 2312 49084 2368
rect 48692 692 48748 748
rect 25956 512 26012 568
rect 19684 332 19740 388
rect 15988 152 16044 208
rect 51604 4832 51660 4888
rect 49924 2672 49980 2728
rect 50148 1772 50204 1828
rect 49812 152 49868 208
rect 52164 532 52220 568
rect 52164 512 52220 532
rect 55636 12212 55692 12268
rect 55972 12212 56028 12268
rect 55300 11852 55356 11908
rect 55748 10592 55804 10648
rect 55540 8974 55596 9030
rect 55644 8974 55700 9030
rect 55748 8974 55804 9030
rect 55540 8870 55596 8926
rect 55644 8870 55700 8926
rect 55748 8870 55804 8926
rect 55540 8766 55596 8822
rect 55644 8766 55700 8822
rect 55748 8766 55804 8822
rect 56308 11492 56364 11548
rect 56308 10052 56364 10108
rect 55540 7576 55596 7632
rect 55644 7576 55700 7632
rect 55748 7576 55804 7632
rect 55540 7472 55596 7528
rect 55644 7472 55700 7528
rect 55748 7472 55804 7528
rect 55540 7368 55596 7424
rect 55644 7368 55700 7424
rect 55748 7368 55804 7424
rect 55540 6178 55596 6234
rect 55644 6178 55700 6234
rect 55748 6178 55804 6234
rect 55540 6074 55596 6130
rect 55644 6074 55700 6130
rect 55748 6074 55804 6130
rect 55540 5970 55596 6026
rect 55644 5970 55700 6026
rect 55748 5970 55804 6026
rect 60228 12032 60284 12088
rect 56756 10592 56812 10648
rect 56980 10592 57036 10648
rect 56756 10232 56812 10288
rect 54180 4472 54236 4528
rect 55300 4112 55356 4168
rect 55524 4112 55580 4168
rect 55524 3752 55580 3808
rect 55076 3212 55132 3268
rect 55300 3220 55356 3268
rect 55300 3212 55356 3220
rect 53172 2324 53228 2368
rect 53172 2312 53228 2324
rect 55300 2132 55356 2188
rect 55524 2132 55580 2188
rect 53620 1952 53676 2008
rect 57316 512 57372 568
rect 59556 10052 59612 10108
rect 58436 6452 58492 6508
rect 71428 14912 71484 14968
rect 67844 14732 67900 14788
rect 60452 11852 60508 11908
rect 60788 11852 60844 11908
rect 67620 14372 67676 14428
rect 67844 14372 67900 14428
rect 68516 14732 68572 14788
rect 67620 13832 67676 13888
rect 63252 13472 63308 13528
rect 63700 13472 63756 13528
rect 63364 10952 63420 11008
rect 62916 9872 62972 9928
rect 62804 5012 62860 5068
rect 62132 3752 62188 3808
rect 58772 2492 58828 2548
rect 59220 2852 59276 2908
rect 60340 2312 60396 2368
rect 59892 1592 59948 1648
rect 60788 2132 60844 2188
rect 62468 1952 62524 2008
rect 62804 1952 62860 2008
rect 60340 1052 60396 1108
rect 60564 1052 60620 1108
rect 65940 13112 65996 13168
rect 66612 13112 66668 13168
rect 65380 11672 65436 11728
rect 65604 11672 65660 11728
rect 63588 9872 63644 9928
rect 63364 7172 63420 7228
rect 63588 6452 63644 6508
rect 63700 5732 63756 5788
rect 63700 4832 63756 4888
rect 64148 3052 64204 3088
rect 64148 3032 64204 3052
rect 69076 14372 69132 14428
rect 68628 13832 68684 13888
rect 68516 12572 68572 12628
rect 66948 11852 67004 11908
rect 67396 11676 67452 11728
rect 68516 11852 68572 11908
rect 67396 11672 67452 11676
rect 68628 10952 68684 11008
rect 68180 10412 68236 10468
rect 68404 10412 68460 10468
rect 68852 13832 68908 13888
rect 68964 12572 69020 12628
rect 68852 11852 68908 11908
rect 67060 10232 67116 10288
rect 68628 10052 68684 10108
rect 66724 6452 66780 6508
rect 65380 3612 65436 3628
rect 65380 3572 65436 3612
rect 65492 3212 65548 3268
rect 65044 2492 65100 2548
rect 65492 2492 65548 2548
rect 63252 152 63308 208
rect 67060 4112 67116 4168
rect 67284 7172 67340 7228
rect 68180 7172 68236 7228
rect 69412 12212 69468 12268
rect 69636 12212 69692 12268
rect 69972 11672 70028 11728
rect 67172 3752 67228 3808
rect 67508 4832 67564 4888
rect 68180 4652 68236 4708
rect 67508 4292 67564 4348
rect 67956 4112 68012 4168
rect 67396 2672 67452 2728
rect 67732 3212 67788 3268
rect 67732 2312 67788 2368
rect 68068 2672 68124 2728
rect 68516 692 68572 748
rect 70084 5012 70140 5068
rect 70308 5012 70364 5068
rect 70308 4652 70364 4708
rect 70532 4652 70588 4708
rect 71652 14912 71708 14968
rect 72772 14372 72828 14428
rect 72772 13652 72828 13708
rect 71764 13112 71820 13168
rect 71652 11672 71708 11728
rect 71652 11312 71708 11368
rect 70532 2132 70588 2188
rect 71988 13112 72044 13168
rect 73220 13652 73276 13708
rect 74004 13112 74060 13168
rect 74228 13112 74284 13168
rect 78932 14372 78988 14428
rect 73556 12032 73612 12088
rect 73668 11852 73724 11908
rect 74340 12212 74396 12268
rect 74452 12392 74508 12448
rect 74004 11672 74060 11728
rect 74228 11672 74284 11728
rect 75124 11312 75180 11368
rect 75460 11312 75516 11368
rect 74116 11132 74172 11188
rect 73668 9872 73724 9928
rect 73892 9872 73948 9928
rect 72212 3392 72268 3448
rect 71876 1592 71932 1648
rect 72100 1592 72156 1648
rect 71988 692 72044 748
rect 72212 692 72268 748
rect 72100 512 72156 568
rect 73108 4652 73164 4708
rect 73332 4652 73388 4708
rect 72996 3392 73052 3448
rect 74788 7812 74844 7868
rect 74004 4292 74060 4348
rect 74228 4292 74284 4348
rect 76244 10232 76300 10288
rect 77588 13132 77644 13168
rect 77588 13112 77644 13132
rect 78148 13472 78204 13528
rect 78484 13832 78540 13888
rect 78820 13832 78876 13888
rect 79156 14372 79212 14428
rect 81284 14552 81340 14608
rect 81508 14552 81564 14608
rect 81508 14372 81564 14428
rect 81732 14372 81788 14428
rect 81284 14028 81340 14068
rect 81284 14012 81340 14028
rect 78372 13472 78428 13528
rect 77924 13112 77980 13168
rect 80612 13112 80668 13168
rect 77140 12032 77196 12088
rect 77364 12032 77420 12088
rect 77700 11312 77756 11368
rect 79268 12212 79324 12268
rect 78484 11852 78540 11908
rect 78260 11672 78316 11728
rect 78036 11312 78092 11368
rect 77588 10232 77644 10288
rect 77588 9872 77644 9928
rect 77812 9872 77868 9928
rect 77028 8484 77084 8540
rect 78484 11672 78540 11728
rect 78148 10412 78204 10468
rect 78372 10412 78428 10468
rect 77251 8484 77307 8540
rect 77700 8484 77756 8540
rect 75124 3932 75180 3988
rect 75348 3932 75404 3988
rect 74564 3220 74620 3268
rect 74564 3212 74620 3220
rect 74900 3212 74956 3268
rect 73444 1952 73500 2008
rect 73780 2672 73836 2728
rect 74004 2672 74060 2728
rect 75124 3032 75180 3088
rect 73780 1952 73836 2008
rect 74340 1772 74396 1828
rect 74564 1772 74620 1828
rect 67844 332 67900 388
rect 67732 152 67788 208
rect 75460 3032 75516 3088
rect 76468 2312 76524 2368
rect 76916 3212 76972 3268
rect 76916 2312 76972 2368
rect 75796 1232 75852 1288
rect 79044 11312 79100 11368
rect 79156 11852 79212 11908
rect 79044 10232 79100 10288
rect 78708 9268 78764 9324
rect 79492 12212 79548 12268
rect 79492 11672 79548 11728
rect 79716 11672 79772 11728
rect 79268 10232 79324 10288
rect 79380 11312 79436 11368
rect 79156 10052 79212 10108
rect 79716 11312 79772 11368
rect 76244 1232 76300 1288
rect 77364 3212 77420 3268
rect 77924 3212 77980 3268
rect 78260 3932 78316 3988
rect 78708 3752 78764 3808
rect 78932 7812 78988 7868
rect 79380 8484 79436 8540
rect 80052 10052 80108 10108
rect 79828 8484 79884 8540
rect 80388 12392 80444 12448
rect 80612 12392 80668 12448
rect 81396 13112 81452 13168
rect 80836 12932 80892 12988
rect 80836 12796 80892 12808
rect 80836 12752 80892 12796
rect 81396 12932 81452 12988
rect 81620 13292 81676 13348
rect 81620 12932 81676 12988
rect 81844 13832 81900 13888
rect 82404 14192 82460 14248
rect 82516 14732 82572 14788
rect 83188 14732 83244 14788
rect 85876 14912 85932 14968
rect 84084 14732 84140 14788
rect 82740 14552 82796 14608
rect 83300 14372 83356 14428
rect 83860 14372 83916 14428
rect 81844 12932 81900 12988
rect 82740 13652 82796 13708
rect 83188 14012 83244 14068
rect 82964 13652 83020 13708
rect 85204 14192 85260 14248
rect 84868 13472 84924 13528
rect 81620 12392 81676 12448
rect 81844 12392 81900 12448
rect 82628 12212 82684 12268
rect 83076 12572 83132 12628
rect 84532 12932 84588 12988
rect 85092 13472 85148 13528
rect 85428 14192 85484 14248
rect 85092 13112 85148 13168
rect 84756 12932 84812 12988
rect 83188 12392 83244 12448
rect 83300 12572 83356 12628
rect 84084 12392 84140 12448
rect 81620 11672 81676 11728
rect 83076 12032 83132 12088
rect 83748 12032 83804 12088
rect 81844 11132 81900 11188
rect 82404 11672 82460 11728
rect 84308 12392 84364 12448
rect 83524 11492 83580 11548
rect 84756 11852 84812 11908
rect 84308 11492 84364 11548
rect 84980 11852 85036 11908
rect 85204 11852 85260 11908
rect 85428 13112 85484 13168
rect 83860 10952 83916 11008
rect 84084 10952 84140 11008
rect 84980 10952 85036 11008
rect 85204 10952 85260 11008
rect 80164 7812 80220 7868
rect 78932 4292 78988 4348
rect 79156 4292 79212 4348
rect 79380 3932 79436 3988
rect 81396 9268 81452 9324
rect 79044 3212 79100 3268
rect 82292 9872 82348 9928
rect 81844 9268 81900 9324
rect 82516 9872 82572 9928
rect 81508 8484 81564 8540
rect 82068 8484 82124 8540
rect 80052 5012 80108 5068
rect 79828 4652 79884 4708
rect 80052 4652 80108 4708
rect 85652 12212 85708 12268
rect 85540 11852 85596 11908
rect 82704 9673 82760 9729
rect 82808 9673 82864 9729
rect 82912 9673 82968 9729
rect 82704 9569 82760 9625
rect 82808 9569 82864 9625
rect 82912 9569 82968 9625
rect 82704 9465 82760 9521
rect 82808 9465 82864 9521
rect 82912 9465 82968 9521
rect 82704 8275 82760 8331
rect 82808 8275 82864 8331
rect 82912 8275 82968 8331
rect 82704 8171 82760 8227
rect 82808 8171 82864 8227
rect 82912 8171 82968 8227
rect 80948 4832 81004 4888
rect 80500 4472 80556 4528
rect 80612 3932 80668 3988
rect 79828 3572 79884 3628
rect 80836 3572 80892 3628
rect 80500 2492 80556 2548
rect 81508 5012 81564 5068
rect 81732 5012 81788 5068
rect 82704 8067 82760 8123
rect 82808 8067 82864 8123
rect 82912 8067 82968 8123
rect 82516 7812 82572 7868
rect 82704 6877 82760 6933
rect 82808 6877 82864 6933
rect 82912 6877 82968 6933
rect 82704 6773 82760 6829
rect 82808 6773 82864 6829
rect 82912 6773 82968 6829
rect 82704 6669 82760 6725
rect 82808 6669 82864 6725
rect 82912 6669 82968 6725
rect 81508 4472 81564 4528
rect 81508 3220 81564 3268
rect 81508 3212 81564 3220
rect 79716 1428 79772 1468
rect 79716 1412 79772 1428
rect 79380 1232 79436 1288
rect 79940 1412 79996 1468
rect 76356 872 76412 928
rect 76804 700 76860 748
rect 76804 692 76860 700
rect 75236 332 75292 388
rect 78148 332 78204 388
rect 78372 332 78428 388
rect 77364 152 77420 208
rect 77588 152 77644 208
rect 79828 1052 79884 1108
rect 81060 2312 81116 2368
rect 80948 2132 81004 2188
rect 81172 2132 81228 2188
rect 81172 1412 81228 1468
rect 81396 1412 81452 1468
rect 82704 5516 82760 5535
rect 82704 5479 82760 5516
rect 82808 5516 82864 5535
rect 82808 5479 82864 5516
rect 82912 5516 82968 5535
rect 82912 5479 82968 5516
rect 82704 5375 82760 5431
rect 82808 5375 82864 5431
rect 82912 5375 82968 5431
rect 82704 5271 82760 5327
rect 82808 5271 82864 5327
rect 82912 5271 82968 5327
rect 83188 5732 83244 5788
rect 82180 3392 82236 3448
rect 81956 3212 82012 3268
rect 81956 2852 82012 2908
rect 82180 2852 82236 2908
rect 82404 3392 82460 3448
rect 82292 1952 82348 2008
rect 82740 2312 82796 2368
rect 82740 1952 82796 2008
rect 82292 1412 82348 1468
rect 82292 1232 82348 1288
rect 82516 1412 82572 1468
rect 82964 1412 83020 1468
rect 83412 5732 83468 5788
rect 83412 3572 83468 3628
rect 83636 3572 83692 3628
rect 83300 2312 83356 2368
rect 83412 3392 83468 3448
rect 83860 3392 83916 3448
rect 84644 5012 84700 5068
rect 83188 1772 83244 1828
rect 84532 1412 84588 1468
rect 86660 14912 86716 14968
rect 102228 14912 102284 14968
rect 87892 14192 87948 14248
rect 86660 12392 86716 12448
rect 86884 12392 86940 12448
rect 86548 12212 86604 12268
rect 86548 11132 86604 11188
rect 86772 11132 86828 11188
rect 86212 10772 86268 10828
rect 86436 10772 86492 10828
rect 84868 5012 84924 5068
rect 85652 6452 85708 6508
rect 85876 6452 85932 6508
rect 85092 5732 85148 5788
rect 85764 5732 85820 5788
rect 84868 2672 84924 2728
rect 85092 3572 85148 3628
rect 86884 9268 86940 9324
rect 87668 12932 87724 12988
rect 89236 14012 89292 14068
rect 89236 13472 89292 13528
rect 87892 12932 87948 12988
rect 89012 13112 89068 13168
rect 89348 13112 89404 13168
rect 89012 12032 89068 12088
rect 102452 14924 102508 14968
rect 102452 14912 102508 14924
rect 92820 14012 92876 14068
rect 93044 14012 93100 14068
rect 92372 13472 92428 13528
rect 92484 13112 92540 13168
rect 90916 12572 90972 12628
rect 89460 12392 89516 12448
rect 89908 12392 89964 12448
rect 87444 10412 87500 10468
rect 86996 8484 87052 8540
rect 86660 7172 86716 7228
rect 85876 4472 85932 4528
rect 86100 4472 86156 4528
rect 86212 3752 86268 3808
rect 86324 3392 86380 3448
rect 87668 10412 87724 10468
rect 87892 11132 87948 11188
rect 88788 11132 88844 11188
rect 88676 10232 88732 10288
rect 88116 10052 88172 10108
rect 88116 9268 88172 9324
rect 89348 9268 89404 9324
rect 85316 3212 85372 3268
rect 85316 2492 85372 2548
rect 85316 2132 85372 2188
rect 85540 2132 85596 2188
rect 86324 2156 86380 2188
rect 86324 2132 86380 2156
rect 86548 2852 86604 2908
rect 86772 2852 86828 2908
rect 86548 2132 86604 2188
rect 86436 1412 86492 1468
rect 82180 332 82236 388
rect 83300 364 83356 388
rect 83300 332 83356 364
rect 86996 1428 87052 1468
rect 86996 1412 87052 1428
rect 88340 7172 88396 7228
rect 87444 4292 87500 4348
rect 88116 4652 88172 4708
rect 86996 1052 87052 1108
rect 87220 1092 87276 1108
rect 87220 1052 87276 1092
rect 88116 4292 88172 4348
rect 88340 4652 88396 4708
rect 90356 10412 90412 10468
rect 90580 12212 90636 12268
rect 90580 10412 90636 10468
rect 90692 11852 90748 11908
rect 91140 12572 91196 12628
rect 92484 12212 92540 12268
rect 92708 13112 92764 13168
rect 91812 12032 91868 12088
rect 91252 11672 91308 11728
rect 91476 11672 91532 11728
rect 91476 11312 91532 11368
rect 91812 11312 91868 11368
rect 88676 4472 88732 4528
rect 88900 4472 88956 4528
rect 88340 4112 88396 4168
rect 88564 4112 88620 4168
rect 88900 2492 88956 2548
rect 89124 2492 89180 2548
rect 91476 3572 91532 3628
rect 92260 10772 92316 10828
rect 90580 3212 90636 3268
rect 91252 2852 91308 2908
rect 91028 2492 91084 2548
rect 91140 2156 91196 2188
rect 91140 2132 91196 2156
rect 91476 2132 91532 2188
rect 92596 10772 92652 10828
rect 92148 4292 92204 4348
rect 94052 12032 94108 12088
rect 92372 4292 92428 4348
rect 92260 3932 92316 3988
rect 94724 10412 94780 10468
rect 94500 9872 94556 9928
rect 94948 10412 95004 10468
rect 94724 9872 94780 9928
rect 98532 13832 98588 13888
rect 97636 12572 97692 12628
rect 100660 13832 100716 13888
rect 102116 14552 102172 14608
rect 98756 12392 98812 12448
rect 96740 11312 96796 11368
rect 95732 5012 95788 5068
rect 95956 5012 96012 5068
rect 94052 3572 94108 3628
rect 94276 3572 94332 3628
rect 91812 2312 91868 2368
rect 91924 3032 91980 3088
rect 92036 2312 92092 2368
rect 91476 1772 91532 1828
rect 91700 1772 91756 1828
rect 97524 11312 97580 11368
rect 97412 3932 97468 3988
rect 95620 3212 95676 3268
rect 102340 14552 102396 14608
rect 102340 14012 102396 14068
rect 102564 14372 102620 14428
rect 102564 14012 102620 14068
rect 102340 12752 102396 12808
rect 102564 12796 102620 12808
rect 102564 12752 102620 12796
rect 102228 12572 102284 12628
rect 98756 11852 98812 11908
rect 98980 11852 99036 11908
rect 100436 11672 100492 11728
rect 99988 11492 100044 11548
rect 98084 4832 98140 4888
rect 97860 3032 97916 3088
rect 99204 5732 99260 5788
rect 98868 4832 98924 4888
rect 98084 3032 98140 3088
rect 99428 5732 99484 5788
rect 101108 11492 101164 11548
rect 101556 11312 101612 11368
rect 100660 10772 100716 10828
rect 100436 8484 100492 8540
rect 100660 7172 100716 7228
rect 99428 4112 99484 4168
rect 98868 3392 98924 3448
rect 99092 3392 99148 3448
rect 95620 2492 95676 2548
rect 96516 2312 96572 2368
rect 99316 2312 99372 2368
rect 98868 2132 98924 2188
rect 97748 1592 97804 1648
rect 94052 872 94108 928
rect 97300 1052 97356 1108
rect 97524 1052 97580 1108
rect 98980 1592 99036 1648
rect 97412 872 97468 928
rect 99652 4112 99708 4168
rect 99652 3572 99708 3628
rect 99988 2852 100044 2908
rect 100212 2852 100268 2908
rect 100660 6452 100716 6508
rect 101108 10772 101164 10828
rect 100548 5012 100604 5068
rect 100772 5012 100828 5068
rect 100324 872 100380 928
rect 101108 6468 101164 6508
rect 101108 6452 101164 6468
rect 100996 3572 101052 3628
rect 101892 10412 101948 10468
rect 101668 7172 101724 7228
rect 101668 5732 101724 5788
rect 102004 5732 102060 5788
rect 102452 12572 102508 12628
rect 102788 12392 102844 12448
rect 102340 10412 102396 10468
rect 102452 10052 102508 10108
rect 102564 11492 102620 11548
rect 102676 10052 102732 10108
rect 103012 14372 103068 14428
rect 109172 14552 109228 14608
rect 104692 14372 104748 14428
rect 103236 12392 103292 12448
rect 103236 12032 103292 12088
rect 103460 12032 103516 12088
rect 103460 11672 103516 11728
rect 102900 11492 102956 11548
rect 103908 12752 103964 12808
rect 104244 12752 104300 12808
rect 104132 11172 104188 11188
rect 104132 11132 104188 11172
rect 102228 4832 102284 4888
rect 102340 3212 102396 3268
rect 102564 3212 102620 3268
rect 102564 2852 102620 2908
rect 103012 7172 103068 7228
rect 103236 7172 103292 7228
rect 109284 14372 109340 14428
rect 109620 14372 109676 14428
rect 108612 13112 108668 13168
rect 104356 11672 104412 11728
rect 103908 4652 103964 4708
rect 102788 2852 102844 2908
rect 103684 3932 103740 3988
rect 103460 2672 103516 2728
rect 103684 2672 103740 2728
rect 104132 4112 104188 4168
rect 103908 2312 103964 2368
rect 104020 2492 104076 2548
rect 102228 1772 102284 1828
rect 101556 1052 101612 1108
rect 101780 1052 101836 1108
rect 100548 872 100604 928
rect 101780 692 101836 748
rect 102004 692 102060 748
rect 102452 1772 102508 1828
rect 104132 2312 104188 2368
rect 105924 11852 105980 11908
rect 105476 11672 105532 11728
rect 106708 12032 106764 12088
rect 106260 11492 106316 11548
rect 104580 11312 104636 11368
rect 104580 10052 104636 10108
rect 104580 8484 104636 8540
rect 106036 10772 106092 10828
rect 105812 10052 105868 10108
rect 106708 11312 106764 11368
rect 106932 12032 106988 12088
rect 106260 10772 106316 10828
rect 105700 4472 105756 4528
rect 105924 4472 105980 4528
rect 105924 4112 105980 4168
rect 106148 4112 106204 4168
rect 106148 3032 106204 3088
rect 106148 2492 106204 2548
rect 108836 13112 108892 13168
rect 108836 12752 108892 12808
rect 109171 12752 109227 12808
rect 109284 12392 109340 12448
rect 108948 11852 109004 11908
rect 107380 3032 107436 3088
rect 106708 2132 106764 2188
rect 107604 3932 107660 3988
rect 107716 3392 107772 3448
rect 107940 3392 107996 3448
rect 110740 12572 110796 12628
rect 109620 12392 109676 12448
rect 109396 11852 109452 11908
rect 110404 11672 110460 11728
rect 110964 12572 111020 12628
rect 109868 8974 109924 9030
rect 109972 8974 110028 9030
rect 110076 8974 110132 9030
rect 109868 8870 109924 8926
rect 109972 8870 110028 8926
rect 110076 8870 110132 8926
rect 109868 8766 109924 8822
rect 109972 8766 110028 8822
rect 110076 8766 110132 8822
rect 109868 7576 109924 7632
rect 109972 7576 110028 7632
rect 110076 7576 110132 7632
rect 109868 7472 109924 7528
rect 109972 7472 110028 7528
rect 110076 7472 110132 7528
rect 109868 7368 109924 7424
rect 109972 7368 110028 7424
rect 110076 7368 110132 7424
rect 109868 6178 109924 6234
rect 109972 6178 110028 6234
rect 110076 6178 110132 6234
rect 109868 6074 109924 6130
rect 109972 6074 110028 6130
rect 110076 6074 110132 6130
rect 109396 5732 109452 5788
rect 109868 5970 109924 6026
rect 109972 5970 110028 6026
rect 110076 5970 110132 6026
rect 109620 5732 109676 5788
rect 109620 4652 109676 4708
rect 109732 4472 109788 4528
rect 109284 4292 109340 4348
rect 109396 3932 109452 3988
rect 108500 2492 108556 2548
rect 108836 2132 108892 2188
rect 110292 3752 110348 3808
rect 110628 3752 110684 3808
rect 110404 2492 110460 2548
rect 107604 1232 107660 1288
rect 106372 872 106428 928
rect 107492 872 107548 928
rect 106036 692 106092 748
rect 107604 692 107660 748
rect 109060 1232 109116 1288
rect 109396 1260 109452 1288
rect 109396 1232 109452 1260
rect 109620 1232 109676 1288
rect 109396 512 109452 568
rect 109620 512 109676 568
rect 110964 2132 111020 2188
rect 111300 2132 111356 2188
rect 111076 512 111132 568
rect 112644 12572 112700 12628
rect 113092 12392 113148 12448
rect 111748 11672 111804 11728
rect 112196 12212 112252 12268
rect 112420 12212 112476 12268
rect 112308 11852 112364 11908
rect 112532 11852 112588 11908
rect 113092 10952 113148 11008
rect 113204 11672 113260 11728
rect 138964 14912 139020 14968
rect 114436 14552 114492 14608
rect 114324 14372 114380 14428
rect 114660 14372 114716 14428
rect 113204 8484 113260 8540
rect 113316 10952 113372 11008
rect 113092 6452 113148 6508
rect 112868 5732 112924 5788
rect 113092 5732 113148 5788
rect 112532 4472 112588 4528
rect 112532 3572 112588 3628
rect 112756 3572 112812 3628
rect 114100 11492 114156 11548
rect 114436 12032 114492 12088
rect 114212 11312 114268 11368
rect 114436 11312 114492 11368
rect 114436 10952 114492 11008
rect 113764 10772 113820 10828
rect 113540 10412 113596 10468
rect 113764 10412 113820 10468
rect 114324 10772 114380 10828
rect 113540 6452 113596 6508
rect 114100 6468 114156 6508
rect 114100 6452 114156 6468
rect 114324 6452 114380 6508
rect 113764 3932 113820 3988
rect 113988 3932 114044 3988
rect 111412 512 111468 568
rect 113876 2132 113932 2188
rect 114212 3212 114268 3268
rect 115108 14372 115164 14428
rect 116564 14372 116620 14428
rect 116788 14372 116844 14428
rect 114772 11672 114828 11728
rect 114996 11672 115052 11728
rect 114996 10232 115052 10288
rect 115220 11132 115276 11188
rect 115220 10232 115276 10288
rect 115444 13112 115500 13168
rect 115668 13112 115724 13168
rect 114884 7812 114940 7868
rect 117012 14192 117068 14248
rect 117236 14196 117292 14248
rect 117572 14372 117628 14428
rect 117796 14372 117852 14428
rect 119588 14552 119644 14608
rect 117236 14192 117292 14196
rect 118132 13860 118188 13888
rect 118132 13832 118188 13860
rect 119140 14372 119196 14428
rect 119364 14420 119420 14428
rect 119364 14372 119420 14420
rect 119812 14192 119868 14248
rect 118356 13832 118412 13888
rect 118580 13112 118636 13168
rect 118804 13112 118860 13168
rect 116004 12212 116060 12268
rect 114660 6452 114716 6508
rect 115332 6452 115388 6508
rect 115892 10592 115948 10648
rect 115556 5012 115612 5068
rect 116340 10592 116396 10648
rect 118916 12212 118972 12268
rect 115780 4832 115836 4888
rect 115668 4472 115724 4528
rect 114772 3444 114828 3448
rect 114772 3392 114828 3444
rect 115668 3032 115724 3088
rect 116004 4472 116060 4528
rect 116004 4112 116060 4168
rect 117796 10412 117852 10468
rect 118020 10412 118076 10468
rect 116452 5012 116508 5068
rect 116228 4832 116284 4888
rect 115892 3032 115948 3088
rect 114772 2492 114828 2548
rect 114996 2492 115052 2548
rect 114212 2132 114268 2188
rect 115220 1952 115276 2008
rect 115444 1232 115500 1288
rect 115668 1232 115724 1288
rect 115780 2132 115836 2188
rect 116452 3932 116508 3988
rect 116340 3572 116396 3628
rect 117012 5732 117068 5788
rect 116788 2132 116844 2188
rect 117012 2132 117068 2188
rect 117460 7172 117516 7228
rect 117684 7812 117740 7868
rect 118244 10232 118300 10288
rect 118468 10232 118524 10288
rect 117236 5732 117292 5788
rect 117684 4832 117740 4888
rect 117348 4292 117404 4348
rect 117236 3572 117292 3628
rect 117460 3752 117516 3808
rect 117124 1592 117180 1648
rect 117348 1952 117404 2008
rect 117684 2852 117740 2908
rect 117572 2312 117628 2368
rect 118020 7172 118076 7228
rect 118244 5012 118300 5068
rect 118132 4832 118188 4888
rect 117684 1952 117740 2008
rect 117460 1592 117516 1648
rect 118132 2852 118188 2908
rect 118692 11132 118748 11188
rect 118916 11132 118972 11188
rect 119364 12572 119420 12628
rect 119588 12572 119644 12628
rect 119140 12212 119196 12268
rect 119140 11852 119196 11908
rect 118692 8484 118748 8540
rect 119364 11852 119420 11908
rect 119588 10052 119644 10108
rect 118804 5012 118860 5068
rect 119028 4832 119084 4888
rect 119364 4832 119420 4888
rect 118580 3032 118636 3088
rect 117796 512 117852 568
rect 118916 3752 118972 3808
rect 119252 4292 119308 4348
rect 119364 3392 119420 3448
rect 119140 2312 119196 2368
rect 119252 3032 119308 3088
rect 120036 14192 120092 14248
rect 120148 14372 120204 14428
rect 120820 14192 120876 14248
rect 120372 12392 120428 12448
rect 120148 12032 120204 12088
rect 120036 9872 120092 9928
rect 120036 4652 120092 4708
rect 120260 10412 120316 10468
rect 120596 11852 120652 11908
rect 121044 12392 121100 12448
rect 121156 12212 121212 12268
rect 120484 11312 120540 11368
rect 120596 10952 120652 11008
rect 120820 10952 120876 11008
rect 124404 14552 124460 14608
rect 124628 14552 124684 14608
rect 132804 14552 132860 14608
rect 123284 13832 123340 13888
rect 123060 13112 123116 13168
rect 122164 12752 122220 12808
rect 121380 12212 121436 12268
rect 121716 11852 121772 11908
rect 121268 10592 121324 10648
rect 120932 10052 120988 10108
rect 121156 9872 121212 9928
rect 121380 10052 121436 10108
rect 120708 7172 120764 7228
rect 120484 4832 120540 4888
rect 120596 3932 120652 3988
rect 120932 7172 120988 7228
rect 121268 4832 121324 4888
rect 121492 4832 121548 4888
rect 121380 4472 121436 4528
rect 120820 3932 120876 3988
rect 120036 3392 120092 3448
rect 120708 3392 120764 3448
rect 122052 10592 122108 10648
rect 121828 10232 121884 10288
rect 120932 3392 120988 3448
rect 121716 3032 121772 3088
rect 121940 3032 121996 3088
rect 121940 2672 121996 2728
rect 120932 2492 120988 2548
rect 121156 2492 121212 2548
rect 120372 1052 120428 1108
rect 120820 1232 120876 1288
rect 118804 512 118860 568
rect 122500 10952 122556 11008
rect 122724 10952 122780 11008
rect 122388 2672 122444 2728
rect 122612 3572 122668 3628
rect 122388 2132 122444 2188
rect 122612 2132 122668 2188
rect 122500 1772 122556 1828
rect 122724 1772 122780 1828
rect 122276 1052 122332 1108
rect 123284 13112 123340 13168
rect 123508 12392 123564 12448
rect 123396 11672 123452 11728
rect 126756 14012 126812 14068
rect 126196 13832 126252 13888
rect 126196 12752 126252 12808
rect 126756 12752 126812 12808
rect 127540 12932 127596 12988
rect 127652 12032 127708 12088
rect 127764 12932 127820 12988
rect 126084 10052 126140 10108
rect 126308 10052 126364 10108
rect 124292 4472 124348 4528
rect 124180 4116 124236 4168
rect 124180 4112 124236 4116
rect 124292 3572 124348 3628
rect 123508 1232 123564 1288
rect 122836 1052 122892 1108
rect 128324 12032 128380 12088
rect 127764 7172 127820 7228
rect 126308 4292 126364 4348
rect 126868 4112 126924 4168
rect 126084 3932 126140 3988
rect 127092 3392 127148 3448
rect 124404 3212 124460 3268
rect 124628 3212 124684 3268
rect 124292 1592 124348 1648
rect 125972 2132 126028 2188
rect 123956 1232 124012 1288
rect 126196 1772 126252 1828
rect 130900 11492 130956 11548
rect 127540 1412 127596 1468
rect 125860 924 125916 928
rect 125860 872 125916 924
rect 123956 512 124012 568
rect 124180 532 124236 568
rect 124180 512 124236 532
rect 129668 3212 129724 3268
rect 129668 2672 129724 2728
rect 128436 1412 128492 1468
rect 131348 10592 131404 10648
rect 132244 11492 132300 11548
rect 131012 5012 131068 5068
rect 131124 4832 131180 4888
rect 131012 3752 131068 3808
rect 131460 4832 131516 4888
rect 131460 3932 131516 3988
rect 131684 4292 131740 4348
rect 133140 14012 133196 14068
rect 132916 11672 132972 11728
rect 131684 3932 131740 3988
rect 132020 3572 132076 3628
rect 133028 11492 133084 11548
rect 133924 11492 133980 11548
rect 133476 5012 133532 5068
rect 137172 13832 137228 13888
rect 134260 12212 134316 12268
rect 134148 11852 134204 11908
rect 134260 11132 134316 11188
rect 134820 10772 134876 10828
rect 134260 10232 134316 10288
rect 134932 9872 134988 9928
rect 134260 7172 134316 7228
rect 134260 5732 134316 5788
rect 132804 3752 132860 3808
rect 134372 4508 134428 4528
rect 134372 4472 134428 4508
rect 132692 3212 132748 3268
rect 134596 2852 134652 2908
rect 134260 2324 134316 2368
rect 134260 2312 134316 2324
rect 134148 1592 134204 1648
rect 134484 1232 134540 1288
rect 136052 10772 136108 10828
rect 135940 10412 135996 10468
rect 137172 11672 137228 11728
rect 135940 6452 135996 6508
rect 135940 4832 135996 4888
rect 136276 4832 136332 4888
rect 136164 4652 136220 4708
rect 136052 4292 136108 4348
rect 136052 3032 136108 3088
rect 135716 2492 135772 2548
rect 135604 1428 135660 1468
rect 135604 1412 135660 1428
rect 135940 2852 135996 2908
rect 136164 2852 136220 2908
rect 135940 2492 135996 2548
rect 136388 4652 136444 4708
rect 137844 11492 137900 11548
rect 138964 12572 139020 12628
rect 138068 11672 138124 11728
rect 138180 11132 138236 11188
rect 138404 11132 138460 11188
rect 137956 10592 138012 10648
rect 138180 10592 138236 10648
rect 137032 9673 137088 9729
rect 137136 9673 137192 9729
rect 137240 9673 137296 9729
rect 137032 9569 137088 9625
rect 137136 9569 137192 9625
rect 137240 9569 137296 9625
rect 137032 9465 137088 9521
rect 137136 9465 137192 9521
rect 137240 9465 137296 9521
rect 137032 8275 137088 8331
rect 137136 8275 137192 8331
rect 137240 8275 137296 8331
rect 137032 8171 137088 8227
rect 137136 8171 137192 8227
rect 137240 8171 137296 8227
rect 137032 8067 137088 8123
rect 137136 8067 137192 8123
rect 137240 8067 137296 8123
rect 137032 6877 137088 6933
rect 137136 6877 137192 6933
rect 137240 6877 137296 6933
rect 137032 6773 137088 6829
rect 137136 6773 137192 6829
rect 137240 6773 137296 6829
rect 137032 6669 137088 6725
rect 137136 6669 137192 6725
rect 137240 6669 137296 6725
rect 137032 5516 137088 5535
rect 137032 5479 137088 5516
rect 137136 5516 137192 5535
rect 137136 5479 137192 5516
rect 137240 5516 137296 5535
rect 137240 5479 137296 5516
rect 138068 10232 138124 10288
rect 137032 5375 137088 5431
rect 137136 5375 137192 5431
rect 137240 5375 137296 5431
rect 137032 5271 137088 5327
rect 137136 5271 137192 5327
rect 137240 5271 137296 5327
rect 137620 3572 137676 3628
rect 136836 2672 136892 2728
rect 137844 2132 137900 2188
rect 136164 1412 136220 1468
rect 135940 1052 135996 1108
rect 138740 10052 138796 10108
rect 138404 5012 138460 5068
rect 139524 14012 139580 14068
rect 142660 14012 142716 14068
rect 145684 14192 145740 14248
rect 141092 13292 141148 13348
rect 141092 12932 141148 12988
rect 142996 13292 143052 13348
rect 141092 12752 141148 12808
rect 139748 12212 139804 12268
rect 139524 12032 139580 12088
rect 140420 11672 140476 11728
rect 139412 7172 139468 7228
rect 138740 4832 138796 4888
rect 140308 5732 140364 5788
rect 139524 4832 139580 4888
rect 138740 3212 138796 3268
rect 138740 1952 138796 2008
rect 140084 4112 140140 4168
rect 140308 4112 140364 4168
rect 140756 11508 140812 11548
rect 140756 11492 140812 11508
rect 141204 11672 141260 11728
rect 140980 10052 141036 10108
rect 141092 4292 141148 4348
rect 140532 3932 140588 3988
rect 141316 3932 141372 3988
rect 140980 3444 141036 3448
rect 140980 3392 141036 3444
rect 141204 3392 141260 3448
rect 141540 4112 141596 4168
rect 141652 10052 141708 10108
rect 140420 1592 140476 1648
rect 137732 872 137788 928
rect 142772 12752 142828 12808
rect 142884 12572 142940 12628
rect 142660 11852 142716 11908
rect 142772 10412 142828 10468
rect 142884 10052 142940 10108
rect 145124 13112 145180 13168
rect 144116 12392 144172 12448
rect 143892 11672 143948 11728
rect 142772 6452 142828 6508
rect 142436 5012 142492 5068
rect 144004 7172 144060 7228
rect 144228 11672 144284 11728
rect 144340 10052 144396 10108
rect 144900 10232 144956 10288
rect 143220 4652 143276 4708
rect 143444 4652 143500 4708
rect 142660 3932 142716 3988
rect 142548 3752 142604 3808
rect 142772 2492 142828 2548
rect 142884 2672 142940 2728
rect 142212 1232 142268 1288
rect 143892 3572 143948 3628
rect 144004 3932 144060 3988
rect 144340 4832 144396 4888
rect 144340 4292 144396 4348
rect 144900 5012 144956 5068
rect 144676 4844 144732 4888
rect 144676 4832 144732 4844
rect 144004 1260 144060 1288
rect 144004 1232 144060 1260
rect 146132 14192 146188 14248
rect 149268 14552 149324 14608
rect 149044 14012 149100 14068
rect 149268 14012 149324 14068
rect 147924 13472 147980 13528
rect 148708 13652 148764 13708
rect 148372 13292 148428 13348
rect 147588 12752 147644 12808
rect 145796 11852 145852 11908
rect 146020 11492 146076 11548
rect 145908 11312 145964 11368
rect 146132 11312 146188 11368
rect 145124 5732 145180 5788
rect 145572 3212 145628 3268
rect 146020 3032 146076 3088
rect 145572 2672 145628 2728
rect 146020 2492 146076 2548
rect 145236 1952 145292 2008
rect 145012 1232 145068 1288
rect 147364 3752 147420 3808
rect 147700 10412 147756 10468
rect 147812 10592 147868 10648
rect 147700 9872 147756 9928
rect 148036 7172 148092 7228
rect 148260 11492 148316 11548
rect 148036 4832 148092 4888
rect 147924 4112 147980 4168
rect 147812 3932 147868 3988
rect 146244 2492 146300 2548
rect 147588 1952 147644 2008
rect 148036 3032 148092 3088
rect 149492 13472 149548 13528
rect 149268 12392 149324 12448
rect 149492 12392 149548 12448
rect 149380 11852 149436 11908
rect 149604 11852 149660 11908
rect 150276 14552 150332 14608
rect 150164 13652 150220 13708
rect 148596 5012 148652 5068
rect 149380 4652 149436 4708
rect 150052 10952 150108 11008
rect 150052 10592 150108 10648
rect 149828 4832 149884 4888
rect 149716 4652 149772 4708
rect 149604 4472 149660 4528
rect 149380 3752 149436 3808
rect 149492 2312 149548 2368
rect 147700 1772 147756 1828
rect 147812 1952 147868 2008
rect 147924 1772 147980 1828
rect 145684 1052 145740 1108
rect 150276 13112 150332 13168
rect 150500 13112 150556 13168
rect 150500 12752 150556 12808
rect 150276 10412 150332 10468
rect 150276 10052 150332 10108
rect 151732 14912 151788 14968
rect 151172 13832 151228 13888
rect 151396 13832 151452 13888
rect 151396 12212 151452 12268
rect 151060 11132 151116 11188
rect 151172 10952 151228 11008
rect 151508 11312 151564 11368
rect 152740 14732 152796 14788
rect 154420 14732 154476 14788
rect 150836 5012 150892 5068
rect 150948 4832 151004 4888
rect 151060 4472 151116 4528
rect 151060 3932 151116 3988
rect 150948 3752 151004 3808
rect 150612 3572 150668 3628
rect 150276 3032 150332 3088
rect 151060 3212 151116 3268
rect 151284 3212 151340 3268
rect 151284 2672 151340 2728
rect 151508 2672 151564 2728
rect 150836 2312 150892 2368
rect 151060 1988 151116 2008
rect 151060 1952 151116 1988
rect 151956 1952 152012 2008
rect 151732 1772 151788 1828
rect 152740 11508 152796 11548
rect 152740 11492 152796 11508
rect 153188 11852 153244 11908
rect 152964 11492 153020 11548
rect 152964 10232 153020 10288
rect 153188 10232 153244 10288
rect 153412 11852 153468 11908
rect 152740 4652 152796 4708
rect 152964 4652 153020 4708
rect 152852 4292 152908 4348
rect 153860 3932 153916 3988
rect 152628 3392 152684 3448
rect 153748 1772 153804 1828
rect 156436 14732 156492 14788
rect 156100 14372 156156 14428
rect 162708 14552 162764 14608
rect 154532 12752 154588 12808
rect 154756 12212 154812 12268
rect 155876 12032 155932 12088
rect 156100 12392 156156 12448
rect 156100 12032 156156 12088
rect 156324 12032 156380 12088
rect 155764 11852 155820 11908
rect 154756 4832 154812 4888
rect 156100 11672 156156 11728
rect 156100 10052 156156 10108
rect 155988 9872 156044 9928
rect 156212 9872 156268 9928
rect 156548 9872 156604 9928
rect 162036 14372 162092 14428
rect 158340 13860 158396 13888
rect 158340 13832 158396 13860
rect 158564 13832 158620 13888
rect 157780 11672 157836 11728
rect 159460 14192 159516 14248
rect 161924 13652 161980 13708
rect 160580 11852 160636 11908
rect 158004 10052 158060 10108
rect 159460 5012 159516 5068
rect 162372 14192 162428 14248
rect 162036 13472 162092 13528
rect 161924 12392 161980 12448
rect 162036 11492 162092 11548
rect 161140 10052 161196 10108
rect 161140 4832 161196 4888
rect 161476 4472 161532 4528
rect 160916 4112 160972 4168
rect 162260 3932 162316 3988
rect 154644 3572 154700 3628
rect 154532 3212 154588 3268
rect 154420 2852 154476 2908
rect 154756 3392 154812 3448
rect 159572 3572 159628 3628
rect 155988 2492 156044 2548
rect 156211 2492 156267 2548
rect 157780 2132 157836 2188
rect 158004 2132 158060 2188
rect 178276 14372 178332 14428
rect 174132 14192 174188 14248
rect 166180 14012 166236 14068
rect 162596 13832 162652 13888
rect 163044 13472 163100 13528
rect 162932 11672 162988 11728
rect 162820 10592 162876 10648
rect 162932 10232 162988 10288
rect 164948 13112 165004 13168
rect 165732 12752 165788 12808
rect 165956 12752 166012 12808
rect 164500 12068 164556 12088
rect 164500 12032 164556 12068
rect 165172 12032 165228 12088
rect 163380 11852 163436 11908
rect 162820 6452 162876 6508
rect 163156 4112 163212 4168
rect 162820 3392 162876 3448
rect 164612 10592 164668 10648
rect 164196 8974 164252 9030
rect 164300 8974 164356 9030
rect 164404 8974 164460 9030
rect 164196 8870 164252 8926
rect 164300 8870 164356 8926
rect 164404 8870 164460 8926
rect 164196 8766 164252 8822
rect 164300 8766 164356 8822
rect 164404 8766 164460 8822
rect 164196 7576 164252 7632
rect 164300 7576 164356 7632
rect 164404 7576 164460 7632
rect 164196 7472 164252 7528
rect 164300 7472 164356 7528
rect 164404 7472 164460 7528
rect 164196 7368 164252 7424
rect 164300 7368 164356 7424
rect 164404 7368 164460 7424
rect 164724 10052 164780 10108
rect 164196 6178 164252 6234
rect 164300 6178 164356 6234
rect 164404 6178 164460 6234
rect 164196 6074 164252 6130
rect 164300 6074 164356 6130
rect 164404 6074 164460 6130
rect 164196 5970 164252 6026
rect 164300 5970 164356 6026
rect 164404 5970 164460 6026
rect 164612 4832 164668 4888
rect 166292 13112 166348 13168
rect 166628 11852 166684 11908
rect 165956 10412 166012 10468
rect 164836 4472 164892 4528
rect 163716 2672 163772 2728
rect 165620 3752 165676 3808
rect 165620 2672 165676 2728
rect 166292 3392 166348 3448
rect 172564 14012 172620 14068
rect 167748 13292 167804 13348
rect 167636 11852 167692 11908
rect 168532 12392 168588 12448
rect 171220 12392 171276 12448
rect 172228 12212 172284 12268
rect 166740 5012 166796 5068
rect 166628 2852 166684 2908
rect 167860 3032 167916 3088
rect 168084 3932 168140 3988
rect 167076 2852 167132 2908
rect 174468 13860 174524 13888
rect 174468 13832 174524 13860
rect 175028 13832 175084 13888
rect 174132 13112 174188 13168
rect 173348 10592 173404 10648
rect 167972 1412 168028 1468
rect 170884 4652 170940 4708
rect 171444 4652 171500 4708
rect 170436 3212 170492 3268
rect 173348 10052 173404 10108
rect 174356 12212 174412 12268
rect 178052 13472 178108 13528
rect 175140 12932 175196 12988
rect 177716 12932 177772 12988
rect 178164 10412 178220 10468
rect 177716 4832 177772 4888
rect 174916 4292 174972 4348
rect 178052 3932 178108 3988
rect 175140 3752 175196 3808
rect 179620 13472 179676 13528
rect 178836 12032 178892 12088
rect 178836 9872 178892 9928
rect 179060 9872 179116 9928
rect 178276 4112 178332 4168
rect 180404 11852 180460 11908
rect 179396 4292 179452 4348
rect 178164 2312 178220 2368
rect 182644 11852 182700 11908
rect 180852 11312 180908 11368
rect 180628 4832 180684 4888
rect 180404 4112 180460 4168
rect 179620 2312 179676 2368
rect 181524 3932 181580 3988
rect 181300 3392 181356 3448
rect 181412 3572 181468 3628
rect 181412 3032 181468 3088
rect 191156 14028 191212 14068
rect 191156 14012 191212 14028
rect 193396 13860 193452 13888
rect 193396 13832 193452 13860
rect 183204 13652 183260 13708
rect 185332 12392 185388 12448
rect 182756 10592 182812 10648
rect 185108 11672 185164 11728
rect 183988 11312 184044 11368
rect 184996 11132 185052 11188
rect 183988 10232 184044 10288
rect 184996 10232 185052 10288
rect 191828 13472 191884 13528
rect 190036 12392 190092 12448
rect 187572 11492 187628 11548
rect 186452 10052 186508 10108
rect 182196 4472 182252 4528
rect 182980 3932 183036 3988
rect 183092 4472 183148 4528
rect 186340 4112 186396 4168
rect 186116 3212 186172 3268
rect 181524 2492 181580 2548
rect 183092 2492 183148 2548
rect 184436 2492 184492 2548
rect 185892 1952 185948 2008
rect 187908 12032 187964 12088
rect 186452 1952 186508 2008
rect 187348 3220 187404 3268
rect 187348 3212 187404 3220
rect 187348 1772 187404 1828
rect 188356 11312 188412 11368
rect 187684 1772 187740 1828
rect 187908 2852 187964 2908
rect 189812 11132 189868 11188
rect 188356 2852 188412 2908
rect 188916 5012 188972 5068
rect 188916 4472 188972 4528
rect 189252 4472 189308 4528
rect 190148 11672 190204 11728
rect 189588 3392 189644 3448
rect 190820 11132 190876 11188
rect 188468 1952 188524 2008
rect 190932 10052 190988 10108
rect 191360 9673 191416 9729
rect 191464 9673 191520 9729
rect 191568 9673 191624 9729
rect 191360 9569 191416 9625
rect 191464 9569 191520 9625
rect 191568 9569 191624 9625
rect 191360 9465 191416 9521
rect 191464 9465 191520 9521
rect 191568 9465 191624 9521
rect 191360 8275 191416 8331
rect 191464 8275 191520 8331
rect 191568 8275 191624 8331
rect 191360 8171 191416 8227
rect 191464 8171 191520 8227
rect 191568 8171 191624 8227
rect 191360 8067 191416 8123
rect 191464 8067 191520 8123
rect 191568 8067 191624 8123
rect 191360 6877 191416 6933
rect 191464 6877 191520 6933
rect 191568 6877 191624 6933
rect 191360 6773 191416 6829
rect 191464 6773 191520 6829
rect 191568 6773 191624 6829
rect 191360 6669 191416 6725
rect 191464 6669 191520 6725
rect 191568 6669 191624 6725
rect 197540 13292 197596 13348
rect 193284 13112 193340 13168
rect 192164 10232 192220 10288
rect 193060 9872 193116 9928
rect 195524 12964 195580 12988
rect 195524 12932 195580 12964
rect 194740 11492 194796 11548
rect 193844 10772 193900 10828
rect 191360 5516 191416 5535
rect 191360 5479 191416 5516
rect 191464 5516 191520 5535
rect 191464 5479 191520 5516
rect 191568 5516 191624 5535
rect 191568 5479 191624 5516
rect 191360 5375 191416 5431
rect 191464 5375 191520 5431
rect 191568 5375 191624 5431
rect 191360 5271 191416 5327
rect 191464 5271 191520 5327
rect 191568 5271 191624 5327
rect 191940 4832 191996 4888
rect 190708 2852 190764 2908
rect 189140 2672 189196 2728
rect 188692 1952 188748 2008
rect 190708 2492 190764 2548
rect 193172 4292 193228 4348
rect 194852 3932 194908 3988
rect 194964 3572 195020 3628
rect 191604 2312 191660 2368
rect 191492 2132 191548 2188
rect 191716 2132 191772 2188
rect 196644 10592 196700 10648
rect 203252 12752 203308 12808
rect 197764 11852 197820 11908
rect 198212 10412 198268 10468
rect 197988 10052 198044 10108
rect 197876 4676 197932 4708
rect 197876 4652 197932 4676
rect 200340 10232 200396 10288
rect 198212 2852 198268 2908
rect 197652 2672 197708 2728
rect 197316 2132 197372 2188
rect 194068 1232 194124 1288
rect 195188 1052 195244 1108
rect 192836 872 192892 928
rect 151060 692 151116 748
rect 197092 332 197148 388
rect 198212 1772 198268 1828
rect 208292 12572 208348 12628
rect 206948 12032 207004 12088
rect 204484 10952 204540 11008
rect 203700 4832 203756 4888
rect 201572 3212 201628 3268
rect 203588 2132 203644 2188
rect 204372 1596 204428 1648
rect 204372 1592 204428 1596
rect 201572 1412 201628 1468
rect 198212 872 198268 928
rect 203028 1232 203084 1288
rect 210308 12212 210364 12268
rect 211204 10232 211260 10288
rect 209972 4472 210028 4528
rect 209636 3780 209692 3808
rect 209636 3752 209692 3780
rect 211316 3032 211372 3088
rect 211764 4832 211820 4888
rect 212772 3392 212828 3448
rect 211092 1412 211148 1468
rect 205604 512 205660 568
rect 197316 332 197372 388
rect 212884 924 212940 928
rect 212884 872 212940 924
rect 217140 332 217196 388
rect 206836 152 206892 208
<< metal5 >>
rect 60436 14968 71500 14984
rect 60436 14912 60452 14968
rect 60508 14912 71428 14968
rect 71484 14912 71500 14968
rect 60436 14896 71500 14912
rect 71636 14968 83036 14984
rect 71636 14912 71652 14968
rect 71708 14912 83036 14968
rect 71636 14896 83036 14912
rect 49124 14788 67916 14804
rect 49124 14732 49140 14788
rect 49196 14732 67844 14788
rect 67900 14732 67916 14788
rect 49124 14716 67916 14732
rect 68500 14788 82588 14804
rect 68500 14732 68516 14788
rect 68572 14732 82516 14788
rect 82572 14732 82588 14788
rect 68500 14716 82588 14732
rect 82948 14624 83036 14896
rect 83172 14968 85948 14984
rect 83172 14912 85876 14968
rect 85932 14912 85948 14968
rect 83172 14896 85948 14912
rect 86644 14968 102300 14984
rect 86644 14912 86660 14968
rect 86716 14912 102228 14968
rect 102284 14912 102300 14968
rect 86644 14896 102300 14912
rect 102436 14968 138812 14984
rect 102436 14912 102452 14968
rect 102508 14912 138812 14968
rect 102436 14896 138812 14912
rect 138948 14968 151804 14984
rect 138948 14912 138964 14968
rect 139020 14912 151732 14968
rect 151788 14912 151804 14968
rect 138948 14896 151804 14912
rect 83172 14788 83260 14896
rect 138724 14804 138812 14896
rect 83172 14732 83188 14788
rect 83244 14732 83260 14788
rect 83172 14716 83260 14732
rect 84068 14788 138588 14804
rect 84068 14732 84084 14788
rect 84140 14732 138588 14788
rect 84068 14716 138588 14732
rect 138724 14788 152812 14804
rect 138724 14732 152740 14788
rect 152796 14732 152812 14788
rect 138724 14716 152812 14732
rect 154404 14788 156508 14804
rect 154404 14732 154420 14788
rect 154476 14732 156436 14788
rect 156492 14732 156508 14788
rect 154404 14716 156508 14732
rect 138500 14624 138588 14716
rect 21460 14608 81356 14624
rect 21460 14552 21476 14608
rect 21532 14552 81284 14608
rect 81340 14552 81356 14608
rect 21460 14536 81356 14552
rect 81492 14608 82812 14624
rect 81492 14552 81508 14608
rect 81564 14552 82740 14608
rect 82796 14552 82812 14608
rect 81492 14536 82812 14552
rect 82948 14608 102188 14624
rect 82948 14552 102116 14608
rect 102172 14552 102188 14608
rect 82948 14536 102188 14552
rect 102324 14608 109244 14624
rect 102324 14552 102340 14608
rect 102396 14552 109172 14608
rect 109228 14552 109244 14608
rect 102324 14536 109244 14552
rect 109380 14608 114508 14624
rect 109380 14552 114436 14608
rect 114492 14552 114508 14608
rect 109380 14536 114508 14552
rect 114644 14536 119436 14624
rect 119572 14608 124476 14624
rect 119572 14552 119588 14608
rect 119644 14552 124404 14608
rect 124460 14552 124476 14608
rect 119572 14536 124476 14552
rect 124612 14608 132876 14624
rect 124612 14552 124628 14608
rect 124684 14552 132804 14608
rect 132860 14552 132876 14608
rect 124612 14536 132876 14552
rect 138500 14608 149340 14624
rect 138500 14552 149268 14608
rect 149324 14552 149340 14608
rect 138500 14536 149340 14552
rect 150260 14608 162780 14624
rect 150260 14552 150276 14608
rect 150332 14552 162708 14608
rect 162764 14552 162780 14608
rect 150260 14536 162780 14552
rect 109380 14444 109468 14536
rect 53828 14428 67692 14444
rect 53828 14372 53844 14428
rect 53900 14372 67620 14428
rect 67676 14372 67692 14428
rect 53828 14356 67692 14372
rect 67828 14428 69148 14444
rect 67828 14372 67844 14428
rect 67900 14372 69076 14428
rect 69132 14372 69148 14428
rect 67828 14356 69148 14372
rect 72756 14428 79004 14444
rect 72756 14372 72772 14428
rect 72828 14372 78932 14428
rect 78988 14372 79004 14428
rect 72756 14356 79004 14372
rect 79140 14428 81580 14444
rect 79140 14372 79156 14428
rect 79212 14372 81508 14428
rect 81564 14372 81580 14428
rect 79140 14356 81580 14372
rect 81716 14428 83372 14444
rect 81716 14372 81732 14428
rect 81788 14372 83300 14428
rect 83356 14372 83372 14428
rect 81716 14356 83372 14372
rect 83844 14428 102636 14444
rect 83844 14372 83860 14428
rect 83916 14372 102564 14428
rect 102620 14372 102636 14428
rect 83844 14356 102636 14372
rect 102996 14428 104764 14444
rect 102996 14372 103012 14428
rect 103068 14372 104692 14428
rect 104748 14372 104764 14428
rect 102996 14356 104764 14372
rect 109268 14428 109468 14444
rect 109268 14372 109284 14428
rect 109340 14372 109468 14428
rect 109268 14356 109468 14372
rect 109604 14428 114396 14444
rect 109604 14372 109620 14428
rect 109676 14372 114324 14428
rect 114380 14372 114396 14428
rect 109604 14356 114396 14372
rect 114644 14428 114732 14536
rect 114644 14372 114660 14428
rect 114716 14372 114732 14428
rect 114644 14356 114732 14372
rect 115092 14428 116636 14444
rect 115092 14372 115108 14428
rect 115164 14372 116564 14428
rect 116620 14372 116636 14428
rect 115092 14356 116636 14372
rect 116772 14428 117644 14444
rect 116772 14372 116788 14428
rect 116844 14372 117572 14428
rect 117628 14372 117644 14428
rect 116772 14356 117644 14372
rect 117780 14428 119212 14444
rect 117780 14372 117796 14428
rect 117852 14372 119140 14428
rect 119196 14372 119212 14428
rect 117780 14356 119212 14372
rect 119348 14428 119436 14536
rect 119348 14372 119364 14428
rect 119420 14372 119436 14428
rect 119348 14356 119436 14372
rect 120132 14428 156172 14444
rect 120132 14372 120148 14428
rect 120204 14372 156100 14428
rect 156156 14372 156172 14428
rect 120132 14356 156172 14372
rect 162020 14428 178348 14444
rect 162020 14372 162036 14428
rect 162092 14372 178276 14428
rect 178332 14372 178348 14428
rect 162020 14356 178348 14372
rect 17764 14248 82476 14264
rect 17764 14192 17780 14248
rect 17836 14192 82404 14248
rect 82460 14192 82476 14248
rect 17764 14176 82476 14192
rect 82612 14248 85276 14264
rect 82612 14192 85204 14248
rect 85260 14192 85276 14248
rect 82612 14176 85276 14192
rect 85412 14248 87964 14264
rect 85412 14192 85428 14248
rect 85484 14192 87892 14248
rect 87948 14192 87964 14248
rect 85412 14176 87964 14192
rect 88996 14248 117084 14264
rect 88996 14192 117012 14248
rect 117068 14192 117084 14248
rect 88996 14176 117084 14192
rect 117220 14248 119884 14264
rect 117220 14192 117236 14248
rect 117292 14192 119812 14248
rect 119868 14192 119884 14248
rect 117220 14176 119884 14192
rect 120020 14248 120892 14264
rect 120020 14192 120036 14248
rect 120092 14192 120820 14248
rect 120876 14192 120892 14248
rect 120020 14176 120892 14192
rect 132675 14248 145756 14264
rect 132675 14192 145684 14248
rect 145740 14192 145756 14248
rect 132675 14176 145756 14192
rect 146116 14248 159532 14264
rect 146116 14192 146132 14248
rect 146188 14192 159460 14248
rect 159516 14192 159532 14248
rect 146116 14176 159532 14192
rect 162356 14248 174204 14264
rect 162356 14192 162372 14248
rect 162428 14192 174132 14248
rect 174188 14192 174204 14248
rect 162356 14176 174204 14192
rect 82612 14084 82700 14176
rect 88996 14084 89084 14176
rect 14852 14068 81356 14084
rect 14852 14012 14868 14068
rect 14924 14012 81284 14068
rect 81340 14012 81356 14068
rect 14852 13996 81356 14012
rect 81492 13996 82700 14084
rect 83172 14068 89084 14084
rect 83172 14012 83188 14068
rect 83244 14012 89084 14068
rect 83172 13996 89084 14012
rect 89220 14068 92892 14084
rect 89220 14012 89236 14068
rect 89292 14012 92820 14068
rect 92876 14012 92892 14068
rect 89220 13996 92892 14012
rect 93028 14068 102412 14084
rect 93028 14012 93044 14068
rect 93100 14012 102340 14068
rect 102396 14012 102412 14068
rect 93028 13996 102412 14012
rect 102548 14068 126828 14084
rect 102548 14012 102564 14068
rect 102620 14012 126756 14068
rect 126812 14012 126828 14068
rect 102548 13996 126828 14012
rect 81492 13904 81580 13996
rect 132675 13904 132763 14176
rect 133124 14068 139596 14084
rect 133124 14012 133140 14068
rect 133196 14012 139524 14068
rect 139580 14012 139596 14068
rect 133124 13996 139596 14012
rect 142644 14068 149116 14084
rect 142644 14012 142660 14068
rect 142716 14012 149044 14068
rect 149100 14012 149116 14068
rect 142644 13996 149116 14012
rect 149252 14068 166252 14084
rect 149252 14012 149268 14068
rect 149324 14012 166180 14068
rect 166236 14012 166252 14068
rect 149252 13996 166252 14012
rect 172548 14068 191228 14084
rect 172548 14012 172564 14068
rect 172620 14012 191156 14068
rect 191212 14012 191228 14068
rect 172548 13996 191228 14012
rect 43188 13888 57164 13904
rect 43188 13832 43204 13888
rect 43260 13832 57092 13888
rect 57148 13832 57164 13888
rect 43188 13816 57164 13832
rect 67604 13888 68700 13904
rect 67604 13832 67620 13888
rect 67676 13832 68628 13888
rect 68684 13832 68700 13888
rect 67604 13816 68700 13832
rect 68836 13888 78556 13904
rect 68836 13832 68852 13888
rect 68908 13832 78484 13888
rect 78540 13832 78556 13888
rect 68836 13816 78556 13832
rect 78804 13888 81580 13904
rect 78804 13832 78820 13888
rect 78876 13832 81580 13888
rect 78804 13816 81580 13832
rect 81828 13888 98604 13904
rect 81828 13832 81844 13888
rect 81900 13832 98532 13888
rect 98588 13832 98604 13888
rect 81828 13816 98604 13832
rect 100644 13888 118204 13904
rect 100644 13832 100660 13888
rect 100716 13832 118132 13888
rect 118188 13832 118204 13888
rect 100644 13816 118204 13832
rect 118340 13888 123356 13904
rect 118340 13832 118356 13888
rect 118412 13832 123284 13888
rect 123340 13832 123356 13888
rect 118340 13816 123356 13832
rect 126180 13888 132763 13904
rect 126180 13832 126196 13888
rect 126252 13832 132763 13888
rect 126180 13816 132763 13832
rect 137156 13888 151244 13904
rect 137156 13832 137172 13888
rect 137228 13832 151172 13888
rect 151228 13832 151244 13888
rect 137156 13816 151244 13832
rect 151380 13888 158412 13904
rect 151380 13832 151396 13888
rect 151452 13832 158340 13888
rect 158396 13832 158412 13888
rect 151380 13816 158412 13832
rect 158548 13888 162444 13904
rect 158548 13832 158564 13888
rect 158620 13832 162444 13888
rect 158548 13816 162444 13832
rect 162580 13888 174540 13904
rect 162580 13832 162596 13888
rect 162652 13832 174468 13888
rect 174524 13832 174540 13888
rect 162580 13816 174540 13832
rect 175012 13888 193468 13904
rect 175012 13832 175028 13888
rect 175084 13832 193396 13888
rect 193452 13832 193468 13888
rect 175012 13816 193468 13832
rect 162356 13724 162444 13816
rect 25044 13708 53916 13724
rect 25044 13652 25060 13708
rect 25116 13652 53844 13708
rect 53900 13652 53916 13708
rect 25044 13636 53916 13652
rect 56628 13708 72844 13724
rect 56628 13652 56644 13708
rect 56700 13652 72772 13708
rect 72828 13652 72844 13708
rect 56628 13636 72844 13652
rect 73204 13708 82812 13724
rect 73204 13652 73220 13708
rect 73276 13652 82740 13708
rect 82796 13652 82812 13708
rect 73204 13636 82812 13652
rect 82948 13708 148780 13724
rect 82948 13652 82964 13708
rect 83020 13652 148708 13708
rect 148764 13652 148780 13708
rect 82948 13636 148780 13652
rect 150148 13708 161996 13724
rect 150148 13652 150164 13708
rect 150220 13652 161924 13708
rect 161980 13652 161996 13708
rect 150148 13636 161996 13652
rect 162356 13708 183276 13724
rect 162356 13652 183204 13708
rect 183260 13652 183276 13708
rect 162356 13636 183276 13652
rect 10484 13528 63324 13544
rect 10484 13472 10500 13528
rect 10556 13472 63252 13528
rect 63308 13472 63324 13528
rect 10484 13456 63324 13472
rect 63684 13528 78220 13544
rect 63684 13472 63700 13528
rect 63756 13472 78148 13528
rect 78204 13472 78220 13528
rect 63684 13456 78220 13472
rect 78356 13528 84940 13544
rect 78356 13472 78372 13528
rect 78428 13472 84868 13528
rect 84924 13472 84940 13528
rect 78356 13456 84940 13472
rect 85076 13528 89308 13544
rect 85076 13472 85092 13528
rect 85148 13472 89236 13528
rect 89292 13472 89308 13528
rect 85076 13456 89308 13472
rect 92356 13528 147996 13544
rect 92356 13472 92372 13528
rect 92428 13472 147924 13528
rect 147980 13472 147996 13528
rect 92356 13456 147996 13472
rect 149476 13528 162108 13544
rect 149476 13472 149492 13528
rect 149548 13472 162036 13528
rect 162092 13472 162108 13528
rect 149476 13456 162108 13472
rect 163028 13528 178124 13544
rect 163028 13472 163044 13528
rect 163100 13472 178052 13528
rect 178108 13472 178124 13528
rect 163028 13456 178124 13472
rect 179604 13528 191900 13544
rect 179604 13472 179620 13528
rect 179676 13472 191828 13528
rect 191884 13472 191900 13528
rect 179604 13456 191900 13472
rect 25716 13348 53916 13364
rect 25716 13292 25732 13348
rect 25788 13292 53844 13348
rect 53900 13292 53916 13348
rect 25716 13276 53916 13292
rect 54052 13348 81244 13364
rect 54052 13292 54068 13348
rect 54124 13292 81244 13348
rect 54052 13276 81244 13292
rect 81604 13348 141164 13364
rect 81604 13292 81620 13348
rect 81676 13292 141092 13348
rect 141148 13292 141164 13348
rect 81604 13276 141164 13292
rect 142980 13348 148220 13364
rect 142980 13292 142996 13348
rect 143052 13292 148220 13348
rect 142980 13276 148220 13292
rect 148356 13348 167820 13364
rect 148356 13292 148372 13348
rect 148428 13292 167748 13348
rect 167804 13292 167820 13348
rect 148356 13276 167820 13292
rect 167955 13348 197612 13364
rect 167955 13292 197540 13348
rect 197596 13292 197612 13348
rect 167955 13276 197612 13292
rect 18436 13168 66012 13184
rect 18436 13112 18452 13168
rect 18508 13112 65940 13168
rect 65996 13112 66012 13168
rect 18436 13096 66012 13112
rect 66596 13168 71836 13184
rect 66596 13112 66612 13168
rect 66668 13112 71764 13168
rect 71820 13112 71836 13168
rect 66596 13096 71836 13112
rect 71972 13168 74076 13184
rect 71972 13112 71988 13168
rect 72044 13112 74004 13168
rect 74060 13112 74076 13168
rect 71972 13096 74076 13112
rect 74212 13168 77660 13184
rect 74212 13112 74228 13168
rect 74284 13112 77588 13168
rect 77644 13112 77660 13168
rect 74212 13096 77660 13112
rect 77908 13168 80684 13184
rect 77908 13112 77924 13168
rect 77980 13112 80612 13168
rect 80668 13112 80684 13168
rect 77908 13096 80684 13112
rect 34452 12988 80908 13004
rect 34452 12932 34468 12988
rect 34524 12932 80836 12988
rect 80892 12932 80908 12988
rect 34452 12916 80908 12932
rect 81156 12824 81244 13276
rect 148132 13184 148220 13276
rect 167955 13184 168043 13276
rect 81380 13168 85164 13184
rect 81380 13112 81396 13168
rect 81452 13112 85092 13168
rect 85148 13112 85164 13168
rect 81380 13096 85164 13112
rect 85412 13168 89084 13184
rect 85412 13112 85428 13168
rect 85484 13112 89012 13168
rect 89068 13112 89084 13168
rect 85412 13096 89084 13112
rect 89332 13168 92556 13184
rect 89332 13112 89348 13168
rect 89404 13112 92484 13168
rect 92540 13112 92556 13168
rect 89332 13096 92556 13112
rect 92692 13168 108684 13184
rect 92692 13112 92708 13168
rect 92764 13112 108612 13168
rect 108668 13112 108684 13168
rect 92692 13096 108684 13112
rect 108820 13168 115516 13184
rect 108820 13112 108836 13168
rect 108892 13112 115444 13168
rect 115500 13112 115516 13168
rect 108820 13096 115516 13112
rect 115652 13168 118652 13184
rect 115652 13112 115668 13168
rect 115724 13112 118580 13168
rect 118636 13112 118652 13168
rect 115652 13096 118652 13112
rect 118788 13168 123132 13184
rect 118788 13112 118804 13168
rect 118860 13112 123060 13168
rect 123116 13112 123132 13168
rect 118788 13096 123132 13112
rect 123268 13168 145196 13184
rect 123268 13112 123284 13168
rect 123340 13112 145124 13168
rect 145180 13112 145196 13168
rect 123268 13096 145196 13112
rect 148132 13168 150348 13184
rect 148132 13112 150276 13168
rect 150332 13112 150348 13168
rect 148132 13096 150348 13112
rect 150484 13168 165020 13184
rect 150484 13112 150500 13168
rect 150556 13112 164948 13168
rect 165004 13112 165020 13168
rect 150484 13096 165020 13112
rect 166276 13168 168043 13184
rect 166276 13112 166292 13168
rect 166348 13112 168043 13168
rect 166276 13096 168043 13112
rect 174116 13168 193356 13184
rect 174116 13112 174132 13168
rect 174188 13112 193284 13168
rect 193340 13112 193356 13168
rect 174116 13096 193356 13112
rect 81380 12988 81692 13004
rect 81380 12932 81396 12988
rect 81452 12932 81620 12988
rect 81676 12932 81692 12988
rect 81380 12916 81692 12932
rect 81828 12988 84604 13004
rect 81828 12932 81844 12988
rect 81900 12932 84532 12988
rect 84588 12932 84604 12988
rect 81828 12916 84604 12932
rect 84740 12988 87740 13004
rect 84740 12932 84756 12988
rect 84812 12932 87668 12988
rect 87724 12932 87740 12988
rect 84740 12916 87740 12932
rect 87876 12988 127612 13004
rect 87876 12932 87892 12988
rect 87948 12932 127540 12988
rect 127596 12932 127612 12988
rect 87876 12916 127612 12932
rect 127748 12988 138588 13004
rect 127748 12932 127764 12988
rect 127820 12932 138588 12988
rect 127748 12916 138588 12932
rect 141076 12988 175212 13004
rect 141076 12932 141092 12988
rect 141148 12932 175140 12988
rect 175196 12932 175212 12988
rect 141076 12916 175212 12932
rect 177700 12988 195596 13004
rect 177700 12932 177716 12988
rect 177772 12932 195524 12988
rect 195580 12932 195596 12988
rect 177700 12916 195596 12932
rect 138500 12824 138588 12916
rect 27956 12808 53132 12824
rect 27956 12752 27972 12808
rect 28028 12752 53060 12808
rect 53116 12752 53132 12808
rect 27956 12736 53132 12752
rect 53380 12808 80908 12824
rect 53380 12752 53396 12808
rect 53452 12752 80836 12808
rect 80892 12752 80908 12808
rect 53380 12736 80908 12752
rect 81156 12808 102412 12824
rect 81156 12752 102340 12808
rect 102396 12752 102412 12808
rect 81156 12736 102412 12752
rect 102548 12808 103980 12824
rect 102548 12752 102564 12808
rect 102620 12752 103908 12808
rect 103964 12752 103980 12808
rect 102548 12736 103980 12752
rect 104228 12808 108908 12824
rect 104228 12752 104244 12808
rect 104300 12752 108836 12808
rect 108892 12752 108908 12808
rect 104228 12736 108908 12752
rect 109155 12808 121003 12824
rect 109155 12752 109171 12808
rect 109227 12752 121003 12808
rect 109155 12736 121003 12752
rect 122148 12808 126268 12824
rect 122148 12752 122164 12808
rect 122220 12752 126196 12808
rect 126252 12752 126268 12808
rect 122148 12736 126268 12752
rect 126740 12808 138364 12824
rect 126740 12752 126756 12808
rect 126812 12752 138364 12808
rect 126740 12736 138364 12752
rect 138500 12808 141164 12824
rect 138500 12752 141092 12808
rect 141148 12752 141164 12808
rect 138500 12736 141164 12752
rect 142756 12808 147324 12824
rect 142756 12752 142772 12808
rect 142828 12752 147324 12808
rect 142756 12736 147324 12752
rect 147572 12808 150572 12824
rect 147572 12752 147588 12808
rect 147644 12752 150500 12808
rect 150556 12752 150572 12808
rect 147572 12736 150572 12752
rect 154516 12808 165804 12824
rect 154516 12752 154532 12808
rect 154588 12752 165732 12808
rect 165788 12752 165804 12808
rect 154516 12736 165804 12752
rect 165940 12808 203324 12824
rect 165940 12752 165956 12808
rect 166012 12752 203252 12808
rect 203308 12752 203324 12808
rect 165940 12736 203324 12752
rect 120915 12644 121003 12736
rect 138276 12644 138364 12736
rect 147236 12644 147324 12736
rect 27172 12628 68588 12644
rect 27172 12572 27188 12628
rect 27244 12572 68516 12628
rect 68572 12572 68588 12628
rect 27172 12556 68588 12572
rect 68948 12628 83148 12644
rect 68948 12572 68964 12628
rect 69020 12572 83076 12628
rect 83132 12572 83148 12628
rect 68948 12556 83148 12572
rect 83284 12628 90988 12644
rect 83284 12572 83300 12628
rect 83356 12572 90916 12628
rect 90972 12572 90988 12628
rect 83284 12556 90988 12572
rect 91124 12628 97708 12644
rect 91124 12572 91140 12628
rect 91196 12572 97636 12628
rect 97692 12572 97708 12628
rect 91124 12556 97708 12572
rect 98516 12628 102300 12644
rect 98516 12572 102228 12628
rect 102284 12572 102300 12628
rect 98516 12556 102300 12572
rect 102436 12628 110812 12644
rect 102436 12572 102452 12628
rect 102508 12572 110740 12628
rect 110796 12572 110812 12628
rect 102436 12556 110812 12572
rect 110948 12628 112716 12644
rect 110948 12572 110964 12628
rect 111020 12572 112644 12628
rect 112700 12572 112716 12628
rect 110948 12556 112716 12572
rect 112852 12628 119436 12644
rect 112852 12572 119364 12628
rect 119420 12572 119436 12628
rect 112852 12556 119436 12572
rect 119572 12628 120668 12644
rect 119572 12572 119588 12628
rect 119644 12572 120668 12628
rect 119572 12556 120668 12572
rect 120915 12556 138140 12644
rect 138276 12628 139036 12644
rect 138276 12572 138964 12628
rect 139020 12572 139036 12628
rect 138276 12556 139036 12572
rect 142868 12628 144523 12644
rect 142868 12572 142884 12628
rect 142940 12572 144523 12628
rect 142868 12556 144523 12572
rect 147236 12628 208364 12644
rect 147236 12572 208292 12628
rect 208348 12572 208364 12628
rect 147236 12556 208364 12572
rect 98516 12464 98604 12556
rect 112852 12464 112940 12556
rect 120580 12464 120668 12556
rect 138052 12464 138140 12556
rect 144435 12464 144523 12556
rect 30084 12448 74188 12464
rect 30084 12392 30100 12448
rect 30156 12392 74188 12448
rect 30084 12376 74188 12392
rect 74436 12448 80460 12464
rect 74436 12392 74452 12448
rect 74508 12392 80388 12448
rect 80444 12392 80460 12448
rect 74436 12376 80460 12392
rect 80596 12448 81692 12464
rect 80596 12392 80612 12448
rect 80668 12392 81620 12448
rect 81676 12392 81692 12448
rect 80596 12376 81692 12392
rect 81828 12448 82924 12464
rect 81828 12392 81844 12448
rect 81900 12392 82924 12448
rect 81828 12376 82924 12392
rect 83172 12448 84156 12464
rect 83172 12392 83188 12448
rect 83244 12392 84084 12448
rect 84140 12392 84156 12448
rect 83172 12376 84156 12392
rect 84292 12448 86732 12464
rect 84292 12392 84308 12448
rect 84364 12392 86660 12448
rect 86716 12392 86732 12448
rect 84292 12376 86732 12392
rect 86868 12448 89532 12464
rect 86868 12392 86884 12448
rect 86940 12392 89460 12448
rect 89516 12392 89532 12448
rect 86868 12376 89532 12392
rect 89892 12448 98604 12464
rect 89892 12392 89908 12448
rect 89964 12392 98604 12448
rect 89892 12376 98604 12392
rect 98740 12448 102860 12464
rect 98740 12392 98756 12448
rect 98812 12392 102788 12448
rect 102844 12392 102860 12448
rect 98740 12376 102860 12392
rect 103220 12448 109356 12464
rect 103220 12392 103236 12448
rect 103292 12392 109284 12448
rect 109340 12392 109356 12448
rect 103220 12376 109356 12392
rect 109604 12448 112940 12464
rect 109604 12392 109620 12448
rect 109676 12392 112940 12448
rect 109604 12376 112940 12392
rect 113076 12448 120444 12464
rect 113076 12392 113092 12448
rect 113148 12392 120372 12448
rect 120428 12392 120444 12448
rect 113076 12376 120444 12392
rect 120580 12448 121116 12464
rect 120580 12392 121044 12448
rect 121100 12392 121116 12448
rect 120580 12376 121116 12392
rect 123492 12448 137916 12464
rect 123492 12392 123508 12448
rect 123564 12392 137916 12448
rect 123492 12376 137916 12392
rect 138052 12448 144188 12464
rect 138052 12392 144116 12448
rect 144172 12392 144188 12448
rect 138052 12376 144188 12392
rect 144435 12448 149340 12464
rect 144435 12392 149268 12448
rect 149324 12392 149340 12448
rect 144435 12376 149340 12392
rect 149476 12448 156172 12464
rect 149476 12392 149492 12448
rect 149548 12392 156100 12448
rect 156156 12392 156172 12448
rect 149476 12376 156172 12392
rect 161908 12448 168604 12464
rect 161908 12392 161924 12448
rect 161980 12392 168532 12448
rect 168588 12392 168604 12448
rect 161908 12376 168604 12392
rect 171204 12448 190108 12464
rect 171204 12392 171220 12448
rect 171276 12392 185332 12448
rect 185388 12392 190036 12448
rect 190092 12392 190108 12448
rect 171204 12376 190108 12392
rect 42180 12268 55708 12284
rect 42180 12212 42196 12268
rect 42252 12212 55636 12268
rect 55692 12212 55708 12268
rect 42180 12196 55708 12212
rect 55956 12268 69484 12284
rect 55956 12212 55972 12268
rect 56028 12212 69412 12268
rect 69468 12212 69484 12268
rect 55956 12196 69484 12212
rect 69620 12268 73963 12284
rect 69620 12212 69636 12268
rect 69692 12212 73963 12268
rect 69620 12196 73963 12212
rect 60212 12088 73628 12104
rect 60212 12032 60228 12088
rect 60284 12032 73556 12088
rect 73612 12032 73628 12088
rect 60212 12016 73628 12032
rect 73875 11924 73963 12196
rect 74100 12104 74188 12376
rect 82836 12284 82924 12376
rect 74324 12268 79340 12284
rect 74324 12212 74340 12268
rect 74396 12212 79268 12268
rect 79324 12212 79340 12268
rect 74324 12196 79340 12212
rect 79476 12268 82700 12284
rect 79476 12212 79492 12268
rect 79548 12212 82628 12268
rect 82684 12212 82700 12268
rect 79476 12196 82700 12212
rect 82836 12268 85724 12284
rect 82836 12212 85652 12268
rect 85708 12212 85724 12268
rect 82836 12196 85724 12212
rect 86532 12268 90652 12284
rect 86532 12212 86548 12268
rect 86604 12212 90580 12268
rect 90636 12212 90652 12268
rect 86532 12196 90652 12212
rect 92468 12268 112268 12284
rect 92468 12212 92484 12268
rect 92540 12212 112196 12268
rect 112252 12212 112268 12268
rect 92468 12196 112268 12212
rect 112404 12268 115516 12284
rect 112404 12212 112420 12268
rect 112476 12212 115516 12268
rect 112404 12196 115516 12212
rect 115988 12268 118988 12284
rect 115988 12212 116004 12268
rect 116060 12212 118916 12268
rect 118972 12212 118988 12268
rect 115988 12196 118988 12212
rect 119124 12268 121228 12284
rect 119124 12212 119140 12268
rect 119196 12212 121156 12268
rect 121212 12212 121228 12268
rect 119124 12196 121228 12212
rect 121364 12268 134332 12284
rect 121364 12212 121380 12268
rect 121436 12212 134260 12268
rect 134316 12212 134332 12268
rect 121364 12196 134332 12212
rect 115428 12104 115516 12196
rect 74100 12088 77212 12104
rect 74100 12032 77140 12088
rect 77196 12032 77212 12088
rect 74100 12016 77212 12032
rect 77348 12088 83148 12104
rect 77348 12032 77364 12088
rect 77420 12032 83076 12088
rect 83132 12032 83148 12088
rect 77348 12016 83148 12032
rect 83732 12088 89084 12104
rect 83732 12032 83748 12088
rect 83804 12032 89012 12088
rect 89068 12032 89084 12088
rect 83732 12016 89084 12032
rect 89220 12088 91884 12104
rect 89220 12032 91812 12088
rect 91868 12032 91884 12088
rect 89220 12016 91884 12032
rect 94036 12088 103308 12104
rect 94036 12032 94052 12088
rect 94108 12032 103236 12088
rect 103292 12032 103308 12088
rect 94036 12016 103308 12032
rect 103444 12088 106780 12104
rect 103444 12032 103460 12088
rect 103516 12032 106708 12088
rect 106764 12032 106780 12088
rect 103444 12016 106780 12032
rect 106916 12088 114508 12104
rect 106916 12032 106932 12088
rect 106988 12032 114436 12088
rect 114492 12032 114508 12088
rect 106916 12016 114508 12032
rect 114644 12016 115292 12104
rect 115428 12088 120220 12104
rect 115428 12032 120148 12088
rect 120204 12032 120220 12088
rect 115428 12016 120220 12032
rect 127636 12088 128396 12104
rect 127636 12032 127652 12088
rect 127708 12032 128324 12088
rect 128380 12032 128396 12088
rect 127636 12016 128396 12032
rect 89220 11924 89308 12016
rect 114644 11924 114732 12016
rect 55284 11908 60524 11924
rect 55284 11852 55300 11908
rect 55356 11852 60452 11908
rect 60508 11852 60524 11908
rect 55284 11836 60524 11852
rect 60772 11908 67020 11924
rect 60772 11852 60788 11908
rect 60844 11852 66948 11908
rect 67004 11852 67020 11908
rect 60772 11836 67020 11852
rect 67156 11908 68588 11924
rect 67156 11852 68516 11908
rect 68572 11852 68588 11908
rect 67156 11836 68588 11852
rect 68836 11908 73740 11924
rect 68836 11852 68852 11908
rect 68908 11852 73668 11908
rect 73724 11852 73740 11908
rect 68836 11836 73740 11852
rect 73875 11908 78556 11924
rect 73875 11852 78484 11908
rect 78540 11852 78556 11908
rect 73875 11836 78556 11852
rect 79140 11908 84828 11924
rect 79140 11852 79156 11908
rect 79212 11852 84756 11908
rect 84812 11852 84828 11908
rect 79140 11836 84828 11852
rect 84964 11908 85276 11924
rect 84964 11852 84980 11908
rect 85036 11852 85204 11908
rect 85260 11852 85276 11908
rect 84964 11836 85276 11852
rect 85524 11908 89308 11924
rect 85524 11852 85540 11908
rect 85596 11852 89308 11908
rect 85524 11836 89308 11852
rect 90676 11908 98828 11924
rect 90676 11852 90692 11908
rect 90748 11852 98756 11908
rect 98812 11852 98828 11908
rect 90676 11836 98828 11852
rect 98964 11908 105772 11924
rect 98964 11852 98980 11908
rect 99036 11852 105772 11908
rect 98964 11836 105772 11852
rect 105908 11908 109020 11924
rect 105908 11852 105924 11908
rect 105980 11852 108948 11908
rect 109004 11852 109020 11908
rect 105908 11836 109020 11852
rect 109380 11908 112380 11924
rect 109380 11852 109396 11908
rect 109452 11852 112308 11908
rect 112364 11852 112380 11908
rect 109380 11836 112380 11852
rect 112516 11908 114732 11924
rect 112516 11852 112532 11908
rect 112588 11852 114732 11908
rect 112516 11836 114732 11852
rect 115204 11924 115292 12016
rect 137828 11924 137916 12376
rect 139732 12268 151468 12284
rect 139732 12212 139748 12268
rect 139804 12212 151396 12268
rect 151452 12212 151468 12268
rect 139732 12196 151468 12212
rect 154740 12268 172300 12284
rect 154740 12212 154756 12268
rect 154812 12212 172228 12268
rect 172284 12212 172300 12268
rect 154740 12196 172300 12212
rect 174340 12268 210380 12284
rect 174340 12212 174356 12268
rect 174412 12212 210308 12268
rect 210364 12212 210380 12268
rect 174340 12196 210380 12212
rect 139508 12088 155948 12104
rect 139508 12032 139524 12088
rect 139580 12032 155876 12088
rect 155932 12032 155948 12088
rect 139508 12016 155948 12032
rect 156084 12088 156172 12104
rect 156084 12032 156100 12088
rect 156156 12032 156172 12088
rect 156084 11924 156172 12032
rect 156308 12088 164572 12104
rect 156308 12032 156324 12088
rect 156380 12032 164500 12088
rect 164556 12032 164572 12088
rect 156308 12016 164572 12032
rect 165156 12088 178908 12104
rect 165156 12032 165172 12088
rect 165228 12032 178836 12088
rect 178892 12032 178908 12088
rect 165156 12016 178908 12032
rect 187892 12088 207020 12104
rect 187892 12032 187908 12088
rect 187964 12032 206948 12088
rect 207004 12032 207020 12088
rect 187892 12016 207020 12032
rect 115204 11908 119212 11924
rect 115204 11852 119140 11908
rect 119196 11852 119212 11908
rect 115204 11836 119212 11852
rect 119348 11908 120668 11924
rect 119348 11852 119364 11908
rect 119420 11852 120596 11908
rect 120652 11852 120668 11908
rect 119348 11836 120668 11852
rect 121700 11908 134220 11924
rect 121700 11852 121716 11908
rect 121772 11852 134148 11908
rect 134204 11852 134220 11908
rect 121700 11836 134220 11852
rect 137828 11908 142732 11924
rect 137828 11852 142660 11908
rect 142716 11852 142732 11908
rect 137828 11836 142732 11852
rect 145780 11908 149452 11924
rect 145780 11852 145796 11908
rect 145852 11852 149380 11908
rect 149436 11852 149452 11908
rect 145780 11836 149452 11852
rect 149588 11908 153260 11924
rect 149588 11852 149604 11908
rect 149660 11852 153188 11908
rect 153244 11852 153260 11908
rect 149588 11836 153260 11852
rect 153396 11908 155836 11924
rect 153396 11852 153412 11908
rect 153468 11852 155764 11908
rect 155820 11852 155836 11908
rect 153396 11836 155836 11852
rect 156084 11908 160652 11924
rect 156084 11852 160580 11908
rect 160636 11852 160652 11908
rect 156084 11836 160652 11852
rect 161572 11836 163228 11924
rect 163364 11908 166700 11924
rect 163364 11852 163380 11908
rect 163436 11852 166628 11908
rect 166684 11852 166700 11908
rect 163364 11836 166700 11852
rect 167620 11908 180476 11924
rect 167620 11852 167636 11908
rect 167692 11852 180404 11908
rect 180460 11852 180476 11908
rect 167620 11836 180476 11852
rect 182628 11908 197836 11924
rect 182628 11852 182644 11908
rect 182700 11852 197764 11908
rect 197820 11852 197836 11908
rect 182628 11836 197836 11852
rect 67156 11744 67244 11836
rect 105684 11744 105772 11836
rect 161572 11744 161660 11836
rect 163140 11744 163228 11836
rect 26724 11728 65452 11744
rect 26724 11672 26740 11728
rect 26796 11672 65380 11728
rect 65436 11672 65452 11728
rect 26724 11656 65452 11672
rect 65588 11728 67244 11744
rect 65588 11672 65604 11728
rect 65660 11672 67244 11728
rect 65588 11656 67244 11672
rect 67380 11728 70044 11744
rect 67380 11672 67396 11728
rect 67452 11672 69972 11728
rect 70028 11672 70044 11728
rect 67380 11656 70044 11672
rect 71636 11728 74076 11744
rect 71636 11672 71652 11728
rect 71708 11672 74004 11728
rect 74060 11672 74076 11728
rect 71636 11656 74076 11672
rect 74212 11728 78332 11744
rect 74212 11672 74228 11728
rect 74284 11672 78260 11728
rect 78316 11672 78332 11728
rect 74212 11656 78332 11672
rect 78468 11728 79564 11744
rect 78468 11672 78484 11728
rect 78540 11672 79492 11728
rect 79548 11672 79564 11728
rect 78468 11656 79564 11672
rect 79700 11728 81692 11744
rect 79700 11672 79716 11728
rect 79772 11672 81620 11728
rect 81676 11672 81692 11728
rect 79700 11656 81692 11672
rect 82388 11728 91324 11744
rect 82388 11672 82404 11728
rect 82460 11672 91252 11728
rect 91308 11672 91324 11728
rect 82388 11656 91324 11672
rect 91460 11728 100508 11744
rect 91460 11672 91476 11728
rect 91532 11672 100436 11728
rect 100492 11672 100508 11728
rect 91460 11656 100508 11672
rect 100644 11728 103532 11744
rect 100644 11672 103460 11728
rect 103516 11672 103532 11728
rect 100644 11656 103532 11672
rect 104340 11728 105548 11744
rect 104340 11672 104356 11728
rect 104412 11672 105476 11728
rect 105532 11672 105548 11728
rect 104340 11656 105548 11672
rect 105684 11728 110476 11744
rect 105684 11672 110404 11728
rect 110460 11672 110476 11728
rect 105684 11656 110476 11672
rect 111732 11728 113276 11744
rect 111732 11672 111748 11728
rect 111804 11672 113204 11728
rect 113260 11672 113276 11728
rect 111732 11656 113276 11672
rect 113860 11728 114844 11744
rect 113860 11672 114772 11728
rect 114828 11672 114844 11728
rect 113860 11656 114844 11672
rect 114980 11728 123468 11744
rect 114980 11672 114996 11728
rect 115052 11672 123396 11728
rect 123452 11672 123468 11728
rect 114980 11656 123468 11672
rect 132900 11728 137244 11744
rect 132900 11672 132916 11728
rect 132972 11672 137172 11728
rect 137228 11672 137244 11728
rect 132900 11656 137244 11672
rect 138052 11728 140492 11744
rect 138052 11672 138068 11728
rect 138124 11672 140420 11728
rect 140476 11672 140492 11728
rect 138052 11656 140492 11672
rect 141188 11728 143964 11744
rect 141188 11672 141204 11728
rect 141260 11672 143892 11728
rect 143948 11672 143964 11728
rect 141188 11656 143964 11672
rect 144212 11728 156172 11744
rect 144212 11672 144228 11728
rect 144284 11672 156100 11728
rect 156156 11672 156172 11728
rect 144212 11656 156172 11672
rect 157764 11728 161660 11744
rect 157764 11672 157780 11728
rect 157836 11672 161660 11728
rect 157764 11656 161660 11672
rect 161796 11728 163004 11744
rect 161796 11672 162932 11728
rect 162988 11672 163004 11728
rect 161796 11656 163004 11672
rect 163140 11728 185180 11744
rect 163140 11672 185108 11728
rect 185164 11672 185180 11728
rect 163140 11656 185180 11672
rect 185540 11728 190220 11744
rect 185540 11672 190148 11728
rect 190204 11672 190220 11728
rect 185540 11656 190220 11672
rect 56292 11548 83596 11564
rect 56292 11492 56308 11548
rect 56364 11492 83524 11548
rect 83580 11492 83596 11548
rect 56292 11476 83596 11492
rect 84292 11548 100060 11564
rect 84292 11492 84308 11548
rect 84364 11492 99988 11548
rect 100044 11492 100060 11548
rect 84292 11476 100060 11492
rect 100644 11384 100732 11656
rect 113860 11564 113948 11656
rect 161796 11564 161884 11656
rect 185540 11564 185628 11656
rect 101092 11548 102636 11564
rect 101092 11492 101108 11548
rect 101164 11492 102564 11548
rect 102620 11492 102636 11548
rect 101092 11476 102636 11492
rect 102884 11548 106332 11564
rect 102884 11492 102900 11548
rect 102956 11492 106260 11548
rect 106316 11492 106332 11548
rect 102884 11476 106332 11492
rect 106468 11476 113948 11564
rect 114084 11548 130972 11564
rect 114084 11492 114100 11548
rect 114156 11492 130900 11548
rect 130956 11492 130972 11548
rect 114084 11476 130972 11492
rect 132228 11548 133100 11564
rect 132228 11492 132244 11548
rect 132300 11492 133028 11548
rect 133084 11492 133100 11548
rect 132228 11476 133100 11492
rect 133908 11548 137916 11564
rect 133908 11492 133924 11548
rect 133980 11492 137844 11548
rect 137900 11492 137916 11548
rect 133908 11476 137916 11492
rect 140740 11548 146092 11564
rect 140740 11492 140756 11548
rect 140812 11492 146020 11548
rect 146076 11492 146092 11548
rect 140740 11476 146092 11492
rect 148244 11548 152812 11564
rect 148244 11492 148260 11548
rect 148316 11492 152740 11548
rect 152796 11492 152812 11548
rect 148244 11476 152812 11492
rect 152948 11548 161884 11564
rect 152948 11492 152964 11548
rect 153020 11492 161884 11548
rect 152948 11476 161884 11492
rect 162020 11548 185628 11564
rect 162020 11492 162036 11548
rect 162092 11492 185628 11548
rect 162020 11476 185628 11492
rect 187556 11548 194812 11564
rect 187556 11492 187572 11548
rect 187628 11492 194740 11548
rect 194796 11492 194812 11548
rect 187556 11476 194812 11492
rect 106468 11384 106556 11476
rect 44532 11368 71724 11384
rect 44532 11312 44548 11368
rect 44604 11312 71652 11368
rect 71708 11312 71724 11368
rect 44532 11296 71724 11312
rect 71860 11368 75196 11384
rect 71860 11312 75124 11368
rect 75180 11312 75196 11368
rect 71860 11296 75196 11312
rect 75444 11368 77772 11384
rect 75444 11312 75460 11368
rect 75516 11312 77700 11368
rect 77756 11312 77772 11368
rect 75444 11296 77772 11312
rect 78020 11368 79116 11384
rect 78020 11312 78036 11368
rect 78092 11312 79044 11368
rect 79100 11312 79116 11368
rect 78020 11296 79116 11312
rect 79364 11368 79788 11384
rect 79364 11312 79380 11368
rect 79436 11312 79716 11368
rect 79772 11312 79788 11368
rect 79364 11296 79788 11312
rect 80148 11368 91548 11384
rect 80148 11312 91476 11368
rect 91532 11312 91548 11368
rect 80148 11296 91548 11312
rect 91796 11368 96812 11384
rect 91796 11312 91812 11368
rect 91868 11312 96740 11368
rect 96796 11312 96812 11368
rect 91796 11296 96812 11312
rect 97508 11368 100732 11384
rect 97508 11312 97524 11368
rect 97580 11312 100732 11368
rect 97508 11296 100732 11312
rect 101540 11368 104428 11384
rect 101540 11312 101556 11368
rect 101612 11312 104428 11368
rect 101540 11296 104428 11312
rect 104564 11368 106556 11384
rect 104564 11312 104580 11368
rect 104636 11312 106556 11368
rect 104564 11296 106556 11312
rect 106692 11368 114284 11384
rect 106692 11312 106708 11368
rect 106764 11312 114212 11368
rect 114268 11312 114284 11368
rect 106692 11296 114284 11312
rect 114420 11368 120556 11384
rect 114420 11312 114436 11368
rect 114492 11312 120484 11368
rect 120540 11312 120556 11368
rect 114420 11296 120556 11312
rect 130995 11368 145980 11384
rect 130995 11312 145908 11368
rect 145964 11312 145980 11368
rect 130995 11296 145980 11312
rect 146116 11368 151356 11384
rect 146116 11312 146132 11368
rect 146188 11312 151356 11368
rect 146116 11296 151356 11312
rect 151492 11368 180924 11384
rect 151492 11312 151508 11368
rect 151564 11312 180852 11368
rect 180908 11312 180924 11368
rect 151492 11296 180924 11312
rect 183972 11368 188428 11384
rect 183972 11312 183988 11368
rect 184044 11312 188356 11368
rect 188412 11312 188428 11368
rect 183972 11296 188428 11312
rect 71860 11204 71948 11296
rect 80148 11204 80236 11296
rect 104340 11204 104428 11296
rect 130995 11204 131083 11296
rect 151268 11204 151356 11296
rect 46212 11188 71948 11204
rect 46212 11132 46228 11188
rect 46284 11132 71948 11188
rect 46212 11116 71948 11132
rect 74100 11188 80236 11204
rect 74100 11132 74116 11188
rect 74172 11132 80236 11188
rect 74100 11116 80236 11132
rect 81828 11188 86620 11204
rect 81828 11132 81844 11188
rect 81900 11132 86548 11188
rect 86604 11132 86620 11188
rect 81828 11116 86620 11132
rect 86756 11188 87964 11204
rect 86756 11132 86772 11188
rect 86828 11132 87892 11188
rect 87948 11132 87964 11188
rect 86756 11116 87964 11132
rect 88772 11188 104204 11204
rect 88772 11132 88788 11188
rect 88844 11132 104132 11188
rect 104188 11132 104204 11188
rect 88772 11116 104204 11132
rect 104340 11116 115068 11204
rect 115204 11188 118764 11204
rect 115204 11132 115220 11188
rect 115276 11132 118692 11188
rect 118748 11132 118764 11188
rect 115204 11116 118764 11132
rect 118900 11188 131083 11204
rect 118900 11132 118916 11188
rect 118972 11132 131083 11188
rect 118900 11116 131083 11132
rect 134244 11188 138252 11204
rect 134244 11132 134260 11188
rect 134316 11132 138180 11188
rect 138236 11132 138252 11188
rect 134244 11116 138252 11132
rect 138388 11188 151132 11204
rect 138388 11132 138404 11188
rect 138460 11132 151060 11188
rect 151116 11132 151132 11188
rect 138388 11116 151132 11132
rect 151268 11188 185068 11204
rect 151268 11132 184996 11188
rect 185052 11132 185068 11188
rect 151268 11116 185068 11132
rect 189796 11188 208363 11204
rect 189796 11132 189812 11188
rect 189868 11132 190820 11188
rect 190876 11132 208363 11188
rect 189796 11116 208363 11132
rect 114980 11024 115068 11116
rect 22692 11008 63436 11024
rect 22692 10952 22708 11008
rect 22764 10952 63364 11008
rect 63420 10952 63436 11008
rect 22692 10936 63436 10952
rect 68612 11008 83932 11024
rect 68612 10952 68628 11008
rect 68684 10952 83860 11008
rect 83916 10952 83932 11008
rect 68612 10936 83932 10952
rect 84068 11008 85052 11024
rect 84068 10952 84084 11008
rect 84140 10952 84980 11008
rect 85036 10952 85052 11008
rect 84068 10936 85052 10952
rect 85188 11008 113164 11024
rect 85188 10952 85204 11008
rect 85260 10952 113092 11008
rect 113148 10952 113164 11008
rect 85188 10936 113164 10952
rect 113300 11008 114508 11024
rect 113300 10952 113316 11008
rect 113372 10952 114436 11008
rect 114492 10952 114508 11008
rect 113300 10936 114508 10952
rect 114980 11008 120668 11024
rect 114980 10952 120596 11008
rect 120652 10952 120668 11008
rect 114980 10936 120668 10952
rect 120804 11008 122572 11024
rect 120804 10952 120820 11008
rect 120876 10952 122500 11008
rect 122556 10952 122572 11008
rect 120804 10936 122572 10952
rect 122708 11008 150124 11024
rect 122708 10952 122724 11008
rect 122780 10952 150052 11008
rect 150108 10952 150124 11008
rect 122708 10936 150124 10952
rect 151156 11008 204556 11024
rect 151156 10952 151172 11008
rect 151228 10952 204484 11008
rect 204540 10952 204556 11008
rect 151156 10936 204556 10952
rect 10260 10828 86284 10844
rect 10260 10772 10276 10828
rect 10332 10772 86212 10828
rect 86268 10772 86284 10828
rect 10260 10756 86284 10772
rect 86420 10828 92332 10844
rect 86420 10772 86436 10828
rect 86492 10772 92260 10828
rect 92316 10772 92332 10828
rect 86420 10756 92332 10772
rect 92580 10828 100732 10844
rect 92580 10772 92596 10828
rect 92652 10772 100660 10828
rect 100716 10772 100732 10828
rect 92580 10756 100732 10772
rect 101092 10828 106108 10844
rect 101092 10772 101108 10828
rect 101164 10772 106036 10828
rect 106092 10772 106108 10828
rect 101092 10756 106108 10772
rect 106244 10828 113836 10844
rect 106244 10772 106260 10828
rect 106316 10772 113764 10828
rect 113820 10772 113836 10828
rect 106244 10756 113836 10772
rect 114308 10828 134892 10844
rect 114308 10772 114324 10828
rect 114380 10772 134820 10828
rect 134876 10772 134892 10828
rect 114308 10756 134892 10772
rect 136036 10828 193916 10844
rect 136036 10772 136052 10828
rect 136108 10772 193844 10828
rect 193900 10772 193916 10828
rect 136036 10756 193916 10772
rect 29972 10648 55820 10664
rect 29972 10592 29988 10648
rect 30044 10592 55748 10648
rect 55804 10592 55820 10648
rect 29972 10576 55820 10592
rect 55956 10648 56828 10664
rect 55956 10592 56756 10648
rect 56812 10592 56828 10648
rect 55956 10576 56828 10592
rect 56964 10648 115964 10664
rect 56964 10592 56980 10648
rect 57036 10592 115892 10648
rect 115948 10592 115964 10648
rect 56964 10576 115964 10592
rect 116324 10648 121340 10664
rect 116324 10592 116340 10648
rect 116396 10592 121268 10648
rect 121324 10592 121340 10648
rect 116324 10576 121340 10592
rect 122036 10648 122572 10664
rect 122036 10592 122052 10648
rect 122108 10592 122572 10648
rect 122036 10576 122572 10592
rect 131332 10648 138028 10664
rect 131332 10592 131348 10648
rect 131404 10592 137956 10648
rect 138012 10592 138028 10648
rect 131332 10576 138028 10592
rect 138164 10648 147884 10664
rect 138164 10592 138180 10648
rect 138236 10592 147812 10648
rect 147868 10592 147884 10648
rect 138164 10576 147884 10592
rect 150036 10648 162892 10664
rect 150036 10592 150052 10648
rect 150108 10592 162820 10648
rect 162876 10592 162892 10648
rect 150036 10576 162892 10592
rect 164596 10648 173420 10664
rect 164596 10592 164612 10648
rect 164668 10592 173348 10648
rect 173404 10592 173420 10648
rect 164596 10576 173420 10592
rect 182740 10648 196716 10664
rect 182740 10592 182756 10648
rect 182812 10592 196644 10648
rect 196700 10592 196716 10648
rect 182740 10576 196716 10592
rect 55956 10484 56044 10576
rect 122484 10484 122572 10576
rect 36804 10468 56044 10484
rect 36804 10412 36820 10468
rect 36876 10412 56044 10468
rect 36804 10396 56044 10412
rect 56180 10468 68252 10484
rect 56180 10412 68180 10468
rect 68236 10412 68252 10468
rect 56180 10396 68252 10412
rect 68388 10468 78220 10484
rect 68388 10412 68404 10468
rect 68460 10412 78148 10468
rect 78204 10412 78220 10468
rect 68388 10396 78220 10412
rect 78356 10468 87516 10484
rect 78356 10412 78372 10468
rect 78428 10412 87444 10468
rect 87500 10412 87516 10468
rect 78356 10396 87516 10412
rect 87652 10468 90428 10484
rect 87652 10412 87668 10468
rect 87724 10412 90356 10468
rect 90412 10412 90428 10468
rect 87652 10396 90428 10412
rect 90564 10468 94796 10484
rect 90564 10412 90580 10468
rect 90636 10412 94724 10468
rect 94780 10412 94796 10468
rect 90564 10396 94796 10412
rect 94932 10468 101964 10484
rect 94932 10412 94948 10468
rect 95004 10412 101892 10468
rect 101948 10412 101964 10468
rect 94932 10396 101964 10412
rect 102324 10468 113612 10484
rect 102324 10412 102340 10468
rect 102396 10412 113540 10468
rect 113596 10412 113612 10468
rect 102324 10396 113612 10412
rect 113748 10468 117868 10484
rect 113748 10412 113764 10468
rect 113820 10412 117796 10468
rect 117852 10412 117868 10468
rect 113748 10396 117868 10412
rect 118004 10468 120108 10484
rect 118004 10412 118020 10468
rect 118076 10412 120108 10468
rect 118004 10396 120108 10412
rect 120244 10468 122124 10484
rect 120244 10412 120260 10468
rect 120316 10412 122124 10468
rect 120244 10396 122124 10412
rect 122484 10396 135452 10484
rect 135924 10468 142844 10484
rect 135924 10412 135940 10468
rect 135996 10412 142772 10468
rect 142828 10412 142844 10468
rect 135924 10396 142844 10412
rect 144435 10468 147772 10484
rect 144435 10412 147700 10468
rect 147756 10412 147772 10468
rect 144435 10396 147772 10412
rect 150260 10468 166028 10484
rect 150260 10412 150276 10468
rect 150332 10412 165956 10468
rect 166012 10412 166028 10468
rect 150260 10396 166028 10412
rect 178148 10468 198284 10484
rect 178148 10412 178164 10468
rect 178220 10412 198212 10468
rect 198268 10412 198284 10468
rect 178148 10396 198284 10412
rect 56180 10304 56268 10396
rect 120020 10304 120108 10396
rect 122036 10304 122124 10396
rect 135364 10304 135452 10396
rect 144435 10304 144523 10396
rect 208275 10304 208363 11116
rect 16196 10288 56268 10304
rect 16196 10232 16212 10288
rect 16268 10232 56268 10288
rect 16196 10216 56268 10232
rect 56740 10288 67132 10304
rect 56740 10232 56756 10288
rect 56812 10232 67060 10288
rect 67116 10232 67132 10288
rect 56740 10216 67132 10232
rect 67268 10288 76316 10304
rect 67268 10232 76244 10288
rect 76300 10232 76316 10288
rect 67268 10216 76316 10232
rect 77572 10288 79116 10304
rect 77572 10232 77588 10288
rect 77644 10232 79044 10288
rect 79100 10232 79116 10288
rect 77572 10216 79116 10232
rect 79252 10288 88524 10304
rect 79252 10232 79268 10288
rect 79324 10232 88524 10288
rect 79252 10216 88524 10232
rect 88660 10288 115068 10304
rect 88660 10232 88676 10288
rect 88732 10232 114996 10288
rect 115052 10232 115068 10288
rect 88660 10216 115068 10232
rect 115204 10288 118316 10304
rect 115204 10232 115220 10288
rect 115276 10232 118244 10288
rect 118300 10232 118316 10288
rect 115204 10216 118316 10232
rect 118452 10288 119884 10304
rect 118452 10232 118468 10288
rect 118524 10232 119884 10288
rect 118452 10216 119884 10232
rect 120020 10288 121900 10304
rect 120020 10232 121828 10288
rect 121884 10232 121900 10288
rect 120020 10216 121900 10232
rect 122036 10288 134332 10304
rect 122036 10232 134260 10288
rect 134316 10232 134332 10288
rect 122036 10216 134332 10232
rect 135364 10288 138140 10304
rect 135364 10232 138068 10288
rect 138124 10232 138140 10288
rect 135364 10216 138140 10232
rect 138500 10216 144523 10304
rect 144884 10288 153036 10304
rect 144884 10232 144900 10288
rect 144956 10232 152964 10288
rect 153020 10232 153036 10288
rect 144884 10216 153036 10232
rect 153172 10288 161436 10304
rect 153172 10232 153188 10288
rect 153244 10232 161436 10288
rect 153172 10216 161436 10232
rect 162916 10288 184060 10304
rect 162916 10232 162932 10288
rect 162988 10232 183988 10288
rect 184044 10232 184060 10288
rect 162916 10216 184060 10232
rect 184980 10288 200412 10304
rect 184980 10232 184996 10288
rect 185052 10232 192164 10288
rect 192220 10232 200340 10288
rect 200396 10232 200412 10288
rect 184980 10216 200412 10232
rect 208275 10288 211276 10304
rect 208275 10232 211204 10288
rect 211260 10232 211276 10288
rect 208275 10216 211276 10232
rect 67268 10124 67356 10216
rect 88436 10124 88524 10216
rect 119796 10124 119884 10216
rect 138500 10124 138588 10216
rect 161348 10124 161436 10216
rect 46100 10108 56380 10124
rect 46100 10052 46116 10108
rect 46172 10052 56308 10108
rect 56364 10052 56380 10108
rect 46100 10036 56380 10052
rect 59540 10108 67356 10124
rect 59540 10052 59556 10108
rect 59612 10052 67356 10108
rect 59540 10036 67356 10052
rect 68612 10108 79228 10124
rect 68612 10052 68628 10108
rect 68684 10052 79156 10108
rect 79212 10052 79228 10108
rect 68612 10036 79228 10052
rect 80036 10108 88188 10124
rect 80036 10052 80052 10108
rect 80108 10052 88116 10108
rect 88172 10052 88188 10108
rect 80036 10036 88188 10052
rect 88436 10108 102524 10124
rect 88436 10052 102452 10108
rect 102508 10052 102524 10108
rect 88436 10036 102524 10052
rect 102660 10108 104652 10124
rect 102660 10052 102676 10108
rect 102732 10052 104580 10108
rect 104636 10052 104652 10108
rect 102660 10036 104652 10052
rect 105796 10108 119660 10124
rect 105796 10052 105812 10108
rect 105868 10052 119588 10108
rect 119644 10052 119660 10108
rect 105796 10036 119660 10052
rect 119796 10108 121004 10124
rect 119796 10052 120932 10108
rect 120988 10052 121004 10108
rect 119796 10036 121004 10052
rect 121364 10108 126156 10124
rect 121364 10052 121380 10108
rect 121436 10052 126084 10108
rect 126140 10052 126156 10108
rect 121364 10036 126156 10052
rect 126292 10108 138588 10124
rect 126292 10052 126308 10108
rect 126364 10052 138588 10108
rect 126292 10036 138588 10052
rect 138724 10108 141052 10124
rect 138724 10052 138740 10108
rect 138796 10052 140980 10108
rect 141036 10052 141052 10108
rect 138724 10036 141052 10052
rect 141636 10108 142956 10124
rect 141636 10052 141652 10108
rect 141708 10052 142884 10108
rect 142940 10052 142956 10108
rect 141636 10036 142956 10052
rect 144324 10108 150348 10124
rect 144324 10052 144340 10108
rect 144396 10052 150276 10108
rect 150332 10052 150348 10108
rect 144324 10036 150348 10052
rect 156084 10108 156283 10124
rect 156084 10052 156100 10108
rect 156156 10052 156283 10108
rect 156084 10036 156283 10052
rect 157988 10108 161212 10124
rect 157988 10052 158004 10108
rect 158060 10052 161140 10108
rect 161196 10052 161212 10108
rect 157988 10036 161212 10052
rect 161348 10108 164796 10124
rect 161348 10052 164724 10108
rect 164780 10052 164796 10108
rect 161348 10036 164796 10052
rect 173332 10108 186524 10124
rect 173332 10052 173348 10108
rect 173404 10052 186452 10108
rect 186508 10052 186524 10108
rect 173332 10036 186524 10052
rect 190916 10108 198060 10124
rect 190916 10052 190932 10108
rect 190988 10052 197988 10108
rect 198044 10052 198060 10108
rect 190916 10036 198060 10052
rect 156195 9944 156283 10036
rect 21684 9928 62988 9944
rect 21684 9872 21700 9928
rect 21756 9872 62916 9928
rect 62972 9872 62988 9928
rect 21684 9856 62988 9872
rect 63572 9928 73740 9944
rect 63572 9872 63588 9928
rect 63644 9872 73668 9928
rect 73724 9872 73740 9928
rect 63572 9856 73740 9872
rect 73876 9928 77660 9944
rect 73876 9872 73892 9928
rect 73948 9872 77588 9928
rect 77644 9872 77660 9928
rect 73876 9856 77660 9872
rect 77796 9928 82364 9944
rect 77796 9872 77812 9928
rect 77868 9872 82292 9928
rect 82348 9872 82364 9928
rect 77796 9856 82364 9872
rect 82500 9928 94572 9944
rect 82500 9872 82516 9928
rect 82572 9872 94500 9928
rect 94556 9872 94572 9928
rect 82500 9856 94572 9872
rect 94708 9928 120108 9944
rect 94708 9872 94724 9928
rect 94780 9872 120036 9928
rect 120092 9872 120108 9928
rect 94708 9856 120108 9872
rect 121140 9928 135004 9944
rect 121140 9872 121156 9928
rect 121212 9872 134932 9928
rect 134988 9872 135004 9928
rect 121140 9856 135004 9872
rect 147684 9928 156060 9944
rect 147684 9872 147700 9928
rect 147756 9872 155988 9928
rect 156044 9872 156060 9928
rect 147684 9856 156060 9872
rect 156195 9928 156384 9944
rect 156195 9872 156212 9928
rect 156268 9872 156384 9928
rect 156195 9856 156384 9872
rect 156532 9928 178908 9944
rect 156532 9872 156548 9928
rect 156604 9872 178836 9928
rect 178892 9872 178908 9928
rect 156532 9856 178908 9872
rect 179044 9928 193132 9944
rect 179044 9872 179060 9928
rect 179116 9872 193060 9928
rect 193116 9872 193132 9928
rect 179044 9856 193132 9872
rect 1284 9729 218684 9757
rect 1284 9673 28376 9729
rect 28432 9673 28480 9729
rect 28536 9673 28584 9729
rect 28640 9673 82704 9729
rect 82760 9673 82808 9729
rect 82864 9673 82912 9729
rect 82968 9673 137032 9729
rect 137088 9673 137136 9729
rect 137192 9673 137240 9729
rect 137296 9673 191360 9729
rect 191416 9673 191464 9729
rect 191520 9673 191568 9729
rect 191624 9673 218684 9729
rect 1284 9625 218684 9673
rect 1284 9569 28376 9625
rect 28432 9569 28480 9625
rect 28536 9569 28584 9625
rect 28640 9569 82704 9625
rect 82760 9569 82808 9625
rect 82864 9569 82912 9625
rect 82968 9569 137032 9625
rect 137088 9569 137136 9625
rect 137192 9569 137240 9625
rect 137296 9569 191360 9625
rect 191416 9569 191464 9625
rect 191520 9569 191568 9625
rect 191624 9569 218684 9625
rect 1284 9521 218684 9569
rect 1284 9465 28376 9521
rect 28432 9465 28480 9521
rect 28536 9465 28584 9521
rect 28640 9465 82704 9521
rect 82760 9465 82808 9521
rect 82864 9465 82912 9521
rect 82968 9465 137032 9521
rect 137088 9465 137136 9521
rect 137192 9465 137240 9521
rect 137296 9465 191360 9521
rect 191416 9465 191464 9521
rect 191520 9465 191568 9521
rect 191624 9465 218684 9521
rect 1284 9437 218684 9465
rect 78692 9324 81468 9340
rect 78692 9268 78708 9324
rect 78764 9268 81396 9324
rect 81452 9268 81468 9324
rect 78692 9252 81468 9268
rect 81828 9324 86956 9340
rect 81828 9268 81844 9324
rect 81900 9268 86884 9324
rect 86940 9268 86956 9324
rect 81828 9252 86956 9268
rect 88100 9324 89420 9340
rect 88100 9268 88116 9324
rect 88172 9268 89348 9324
rect 89404 9268 89420 9324
rect 88100 9252 89420 9268
rect 1284 9030 218684 9058
rect 1284 8974 55540 9030
rect 55596 8974 55644 9030
rect 55700 8974 55748 9030
rect 55804 8974 109868 9030
rect 109924 8974 109972 9030
rect 110028 8974 110076 9030
rect 110132 8974 164196 9030
rect 164252 8974 164300 9030
rect 164356 8974 164404 9030
rect 164460 8974 218684 9030
rect 1284 8926 218684 8974
rect 1284 8870 55540 8926
rect 55596 8870 55644 8926
rect 55700 8870 55748 8926
rect 55804 8870 109868 8926
rect 109924 8870 109972 8926
rect 110028 8870 110076 8926
rect 110132 8870 164196 8926
rect 164252 8870 164300 8926
rect 164356 8870 164404 8926
rect 164460 8870 218684 8926
rect 1284 8822 218684 8870
rect 1284 8766 55540 8822
rect 55596 8766 55644 8822
rect 55700 8766 55748 8822
rect 55804 8766 109868 8822
rect 109924 8766 109972 8822
rect 110028 8766 110076 8822
rect 110132 8766 164196 8822
rect 164252 8766 164300 8822
rect 164356 8766 164404 8822
rect 164460 8766 218684 8822
rect 1284 8738 218684 8766
rect 77012 8540 77323 8556
rect 77012 8484 77028 8540
rect 77084 8484 77251 8540
rect 77307 8484 77323 8540
rect 77012 8468 77323 8484
rect 77684 8540 79452 8556
rect 77684 8484 77700 8540
rect 77756 8484 79380 8540
rect 79436 8484 79452 8540
rect 77684 8468 79452 8484
rect 79812 8540 81580 8556
rect 79812 8484 79828 8540
rect 79884 8484 81508 8540
rect 81564 8484 81580 8540
rect 79812 8468 81580 8484
rect 82052 8540 87068 8556
rect 82052 8484 82068 8540
rect 82124 8484 86996 8540
rect 87052 8484 87068 8540
rect 82052 8468 87068 8484
rect 100420 8540 104652 8556
rect 100420 8484 100436 8540
rect 100492 8484 104580 8540
rect 104636 8484 104652 8540
rect 100420 8468 104652 8484
rect 113188 8540 118764 8556
rect 113188 8484 113204 8540
rect 113260 8484 118692 8540
rect 118748 8484 118764 8540
rect 113188 8468 118764 8484
rect 1284 8331 218684 8359
rect 1284 8275 28376 8331
rect 28432 8275 28480 8331
rect 28536 8275 28584 8331
rect 28640 8275 82704 8331
rect 82760 8275 82808 8331
rect 82864 8275 82912 8331
rect 82968 8275 137032 8331
rect 137088 8275 137136 8331
rect 137192 8275 137240 8331
rect 137296 8275 191360 8331
rect 191416 8275 191464 8331
rect 191520 8275 191568 8331
rect 191624 8275 218684 8331
rect 1284 8227 218684 8275
rect 1284 8171 28376 8227
rect 28432 8171 28480 8227
rect 28536 8171 28584 8227
rect 28640 8171 82704 8227
rect 82760 8171 82808 8227
rect 82864 8171 82912 8227
rect 82968 8171 137032 8227
rect 137088 8171 137136 8227
rect 137192 8171 137240 8227
rect 137296 8171 191360 8227
rect 191416 8171 191464 8227
rect 191520 8171 191568 8227
rect 191624 8171 218684 8227
rect 1284 8123 218684 8171
rect 1284 8067 28376 8123
rect 28432 8067 28480 8123
rect 28536 8067 28584 8123
rect 28640 8067 82704 8123
rect 82760 8067 82808 8123
rect 82864 8067 82912 8123
rect 82968 8067 137032 8123
rect 137088 8067 137136 8123
rect 137192 8067 137240 8123
rect 137296 8067 191360 8123
rect 191416 8067 191464 8123
rect 191520 8067 191568 8123
rect 191624 8067 218684 8123
rect 1284 8039 218684 8067
rect 74772 7868 79004 7884
rect 74772 7812 74788 7868
rect 74844 7812 78932 7868
rect 78988 7812 79004 7868
rect 74772 7796 79004 7812
rect 80148 7868 82588 7884
rect 80148 7812 80164 7868
rect 80220 7812 82516 7868
rect 82572 7812 82588 7868
rect 80148 7796 82588 7812
rect 114868 7868 117756 7884
rect 114868 7812 114884 7868
rect 114940 7812 117684 7868
rect 117740 7812 117756 7868
rect 114868 7796 117756 7812
rect 1284 7632 218684 7660
rect 1284 7576 55540 7632
rect 55596 7576 55644 7632
rect 55700 7576 55748 7632
rect 55804 7576 109868 7632
rect 109924 7576 109972 7632
rect 110028 7576 110076 7632
rect 110132 7576 164196 7632
rect 164252 7576 164300 7632
rect 164356 7576 164404 7632
rect 164460 7576 218684 7632
rect 1284 7528 218684 7576
rect 1284 7472 55540 7528
rect 55596 7472 55644 7528
rect 55700 7472 55748 7528
rect 55804 7472 109868 7528
rect 109924 7472 109972 7528
rect 110028 7472 110076 7528
rect 110132 7472 164196 7528
rect 164252 7472 164300 7528
rect 164356 7472 164404 7528
rect 164460 7472 218684 7528
rect 1284 7424 218684 7472
rect 1284 7368 55540 7424
rect 55596 7368 55644 7424
rect 55700 7368 55748 7424
rect 55804 7368 109868 7424
rect 109924 7368 109972 7424
rect 110028 7368 110076 7424
rect 110132 7368 164196 7424
rect 164252 7368 164300 7424
rect 164356 7368 164404 7424
rect 164460 7368 218684 7424
rect 1284 7340 218684 7368
rect 63348 7228 67356 7244
rect 63348 7172 63364 7228
rect 63420 7172 67284 7228
rect 67340 7172 67356 7228
rect 63348 7156 67356 7172
rect 68164 7228 86732 7244
rect 68164 7172 68180 7228
rect 68236 7172 86660 7228
rect 86716 7172 86732 7228
rect 68164 7156 86732 7172
rect 88324 7228 100732 7244
rect 88324 7172 88340 7228
rect 88396 7172 100660 7228
rect 100716 7172 100732 7228
rect 88324 7156 100732 7172
rect 101652 7228 103084 7244
rect 101652 7172 101668 7228
rect 101724 7172 103012 7228
rect 103068 7172 103084 7228
rect 101652 7156 103084 7172
rect 103220 7228 117532 7244
rect 103220 7172 103236 7228
rect 103292 7172 117460 7228
rect 117516 7172 117532 7228
rect 103220 7156 117532 7172
rect 118004 7228 120780 7244
rect 118004 7172 118020 7228
rect 118076 7172 120708 7228
rect 120764 7172 120780 7228
rect 118004 7156 120780 7172
rect 120916 7228 127836 7244
rect 120916 7172 120932 7228
rect 120988 7172 127764 7228
rect 127820 7172 127836 7228
rect 120916 7156 127836 7172
rect 134244 7228 139484 7244
rect 134244 7172 134260 7228
rect 134316 7172 139412 7228
rect 139468 7172 139484 7228
rect 134244 7156 139484 7172
rect 143988 7228 148108 7244
rect 143988 7172 144004 7228
rect 144060 7172 148036 7228
rect 148092 7172 148108 7228
rect 143988 7156 148108 7172
rect 1284 6933 218684 6961
rect 1284 6877 28376 6933
rect 28432 6877 28480 6933
rect 28536 6877 28584 6933
rect 28640 6877 82704 6933
rect 82760 6877 82808 6933
rect 82864 6877 82912 6933
rect 82968 6877 137032 6933
rect 137088 6877 137136 6933
rect 137192 6877 137240 6933
rect 137296 6877 191360 6933
rect 191416 6877 191464 6933
rect 191520 6877 191568 6933
rect 191624 6877 218684 6933
rect 1284 6829 218684 6877
rect 1284 6773 28376 6829
rect 28432 6773 28480 6829
rect 28536 6773 28584 6829
rect 28640 6773 82704 6829
rect 82760 6773 82808 6829
rect 82864 6773 82912 6829
rect 82968 6773 137032 6829
rect 137088 6773 137136 6829
rect 137192 6773 137240 6829
rect 137296 6773 191360 6829
rect 191416 6773 191464 6829
rect 191520 6773 191568 6829
rect 191624 6773 218684 6829
rect 1284 6725 218684 6773
rect 1284 6669 28376 6725
rect 28432 6669 28480 6725
rect 28536 6669 28584 6725
rect 28640 6669 82704 6725
rect 82760 6669 82808 6725
rect 82864 6669 82912 6725
rect 82968 6669 137032 6725
rect 137088 6669 137136 6725
rect 137192 6669 137240 6725
rect 137296 6669 191360 6725
rect 191416 6669 191464 6725
rect 191520 6669 191568 6725
rect 191624 6669 218684 6725
rect 1284 6641 218684 6669
rect 58420 6508 63660 6524
rect 58420 6452 58436 6508
rect 58492 6452 63588 6508
rect 63644 6452 63660 6508
rect 58420 6436 63660 6452
rect 66708 6508 85724 6524
rect 66708 6452 66724 6508
rect 66780 6452 85652 6508
rect 85708 6452 85724 6508
rect 66708 6436 85724 6452
rect 85860 6508 100732 6524
rect 85860 6452 85876 6508
rect 85932 6452 100660 6508
rect 100716 6452 100732 6508
rect 85860 6436 100732 6452
rect 101092 6508 113164 6524
rect 101092 6452 101108 6508
rect 101164 6452 113092 6508
rect 113148 6452 113164 6508
rect 101092 6436 113164 6452
rect 113524 6508 114172 6524
rect 113524 6452 113540 6508
rect 113596 6452 114100 6508
rect 114156 6452 114172 6508
rect 113524 6436 114172 6452
rect 114308 6508 114732 6524
rect 114308 6452 114324 6508
rect 114380 6452 114660 6508
rect 114716 6452 114732 6508
rect 114308 6436 114732 6452
rect 115316 6508 136012 6524
rect 115316 6452 115332 6508
rect 115388 6452 135940 6508
rect 135996 6452 136012 6508
rect 115316 6436 136012 6452
rect 142756 6508 162892 6524
rect 142756 6452 142772 6508
rect 142828 6452 162820 6508
rect 162876 6452 162892 6508
rect 142756 6436 162892 6452
rect 1284 6234 218684 6262
rect 1284 6178 55540 6234
rect 55596 6178 55644 6234
rect 55700 6178 55748 6234
rect 55804 6178 109868 6234
rect 109924 6178 109972 6234
rect 110028 6178 110076 6234
rect 110132 6178 164196 6234
rect 164252 6178 164300 6234
rect 164356 6178 164404 6234
rect 164460 6178 218684 6234
rect 1284 6130 218684 6178
rect 1284 6074 55540 6130
rect 55596 6074 55644 6130
rect 55700 6074 55748 6130
rect 55804 6074 109868 6130
rect 109924 6074 109972 6130
rect 110028 6074 110076 6130
rect 110132 6074 164196 6130
rect 164252 6074 164300 6130
rect 164356 6074 164404 6130
rect 164460 6074 218684 6130
rect 1284 6026 218684 6074
rect 1284 5970 55540 6026
rect 55596 5970 55644 6026
rect 55700 5970 55748 6026
rect 55804 5970 109868 6026
rect 109924 5970 109972 6026
rect 110028 5970 110076 6026
rect 110132 5970 164196 6026
rect 164252 5970 164300 6026
rect 164356 5970 164404 6026
rect 164460 5970 218684 6026
rect 1284 5942 218684 5970
rect 63684 5788 83260 5804
rect 63684 5732 63700 5788
rect 63756 5732 83188 5788
rect 83244 5732 83260 5788
rect 63684 5716 83260 5732
rect 83396 5788 85164 5804
rect 83396 5732 83412 5788
rect 83468 5732 85092 5788
rect 85148 5732 85164 5788
rect 83396 5716 85164 5732
rect 85748 5788 99276 5804
rect 85748 5732 85764 5788
rect 85820 5732 99204 5788
rect 99260 5732 99276 5788
rect 85748 5716 99276 5732
rect 99412 5788 101740 5804
rect 99412 5732 99428 5788
rect 99484 5732 101668 5788
rect 101724 5732 101740 5788
rect 99412 5716 101740 5732
rect 101988 5788 109468 5804
rect 101988 5732 102004 5788
rect 102060 5732 109396 5788
rect 109452 5732 109468 5788
rect 101988 5716 109468 5732
rect 109604 5788 112940 5804
rect 109604 5732 109620 5788
rect 109676 5732 112868 5788
rect 112924 5732 112940 5788
rect 109604 5716 112940 5732
rect 113076 5788 117084 5804
rect 113076 5732 113092 5788
rect 113148 5732 117012 5788
rect 117068 5732 117084 5788
rect 113076 5716 117084 5732
rect 117220 5788 134332 5804
rect 117220 5732 117236 5788
rect 117292 5732 134260 5788
rect 134316 5732 134332 5788
rect 117220 5716 134332 5732
rect 140292 5788 145196 5804
rect 140292 5732 140308 5788
rect 140364 5732 145124 5788
rect 145180 5732 145196 5788
rect 140292 5716 145196 5732
rect 1284 5535 218684 5563
rect 1284 5479 28376 5535
rect 28432 5479 28480 5535
rect 28536 5479 28584 5535
rect 28640 5479 82704 5535
rect 82760 5479 82808 5535
rect 82864 5479 82912 5535
rect 82968 5479 137032 5535
rect 137088 5479 137136 5535
rect 137192 5479 137240 5535
rect 137296 5479 191360 5535
rect 191416 5479 191464 5535
rect 191520 5479 191568 5535
rect 191624 5479 218684 5535
rect 1284 5431 218684 5479
rect 1284 5375 28376 5431
rect 28432 5375 28480 5431
rect 28536 5375 28584 5431
rect 28640 5375 82704 5431
rect 82760 5375 82808 5431
rect 82864 5375 82912 5431
rect 82968 5375 137032 5431
rect 137088 5375 137136 5431
rect 137192 5375 137240 5431
rect 137296 5375 191360 5431
rect 191416 5375 191464 5431
rect 191520 5375 191568 5431
rect 191624 5375 218684 5431
rect 1284 5327 218684 5375
rect 1284 5271 28376 5327
rect 28432 5271 28480 5327
rect 28536 5271 28584 5327
rect 28640 5271 82704 5327
rect 82760 5271 82808 5327
rect 82864 5271 82912 5327
rect 82968 5271 137032 5327
rect 137088 5271 137136 5327
rect 137192 5271 137240 5327
rect 137296 5271 191360 5327
rect 191416 5271 191464 5327
rect 191520 5271 191568 5327
rect 191624 5271 218684 5327
rect 1284 5243 218684 5271
rect 62788 5068 70156 5084
rect 62788 5012 62804 5068
rect 62860 5012 70084 5068
rect 70140 5012 70156 5068
rect 62788 4996 70156 5012
rect 70292 5068 80124 5084
rect 70292 5012 70308 5068
rect 70364 5012 80052 5068
rect 80108 5012 80124 5068
rect 70292 4996 80124 5012
rect 80708 5068 81580 5084
rect 80708 5012 81508 5068
rect 81564 5012 81580 5068
rect 80708 4996 81580 5012
rect 81716 5068 84716 5084
rect 81716 5012 81732 5068
rect 81788 5012 84644 5068
rect 84700 5012 84716 5068
rect 81716 4996 84716 5012
rect 84852 5068 95804 5084
rect 84852 5012 84868 5068
rect 84924 5012 95732 5068
rect 95788 5012 95804 5068
rect 84852 4996 95804 5012
rect 95940 5068 100620 5084
rect 95940 5012 95956 5068
rect 96012 5012 100548 5068
rect 100604 5012 100620 5068
rect 95940 4996 100620 5012
rect 100756 5068 115628 5084
rect 100756 5012 100772 5068
rect 100828 5012 115556 5068
rect 115612 5012 115628 5068
rect 100756 4996 115628 5012
rect 116436 5068 118316 5084
rect 116436 5012 116452 5068
rect 116508 5012 118244 5068
rect 118300 5012 118316 5068
rect 116436 4996 118316 5012
rect 118788 5068 131084 5084
rect 118788 5012 118804 5068
rect 118860 5012 131012 5068
rect 131068 5012 131084 5068
rect 118788 4996 131084 5012
rect 133460 5068 138476 5084
rect 133460 5012 133476 5068
rect 133532 5012 138404 5068
rect 138460 5012 138476 5068
rect 133460 4996 138476 5012
rect 142420 5068 144972 5084
rect 142420 5012 142436 5068
rect 142492 5012 144900 5068
rect 144956 5012 144972 5068
rect 142420 4996 144972 5012
rect 145108 5068 150908 5084
rect 145108 5012 148596 5068
rect 148652 5012 150836 5068
rect 150892 5012 150908 5068
rect 145108 4996 150908 5012
rect 159444 5068 166812 5084
rect 159444 5012 159460 5068
rect 159516 5012 166740 5068
rect 166796 5012 166812 5068
rect 159444 4996 166812 5012
rect 188900 5068 192236 5084
rect 188900 5012 188916 5068
rect 188972 5012 192236 5068
rect 188900 4996 192236 5012
rect 80708 4904 80796 4996
rect 145108 4904 145196 4996
rect 192148 4904 192236 4996
rect 51588 4888 63772 4904
rect 51588 4832 51604 4888
rect 51660 4832 63700 4888
rect 63756 4832 63772 4888
rect 51588 4816 63772 4832
rect 67492 4888 80796 4904
rect 67492 4832 67508 4888
rect 67564 4832 80796 4888
rect 67492 4816 80796 4832
rect 80932 4888 98156 4904
rect 80932 4832 80948 4888
rect 81004 4832 98084 4888
rect 98140 4832 98156 4888
rect 80932 4816 98156 4832
rect 98852 4888 102300 4904
rect 98852 4832 98868 4888
rect 98924 4832 102228 4888
rect 102284 4832 102300 4888
rect 98852 4816 102300 4832
rect 103220 4888 115852 4904
rect 103220 4832 115780 4888
rect 115836 4832 115852 4888
rect 103220 4816 115852 4832
rect 116212 4888 117756 4904
rect 116212 4832 116228 4888
rect 116284 4832 117684 4888
rect 117740 4832 117756 4888
rect 116212 4816 117756 4832
rect 118116 4888 119100 4904
rect 118116 4832 118132 4888
rect 118188 4832 119028 4888
rect 119084 4832 119100 4888
rect 118116 4816 119100 4832
rect 119348 4888 120332 4904
rect 119348 4832 119364 4888
rect 119420 4832 120332 4888
rect 119348 4816 120332 4832
rect 120468 4888 121340 4904
rect 120468 4832 120484 4888
rect 120540 4832 121268 4888
rect 121324 4832 121340 4888
rect 120468 4816 121340 4832
rect 121476 4888 131196 4904
rect 121476 4832 121492 4888
rect 121548 4832 131124 4888
rect 131180 4832 131196 4888
rect 121476 4816 131196 4832
rect 131444 4888 136012 4904
rect 131444 4832 131460 4888
rect 131516 4832 135940 4888
rect 135996 4832 136012 4888
rect 131444 4816 136012 4832
rect 136260 4888 138812 4904
rect 136260 4832 136276 4888
rect 136332 4832 138740 4888
rect 138796 4832 138812 4888
rect 136260 4816 138812 4832
rect 139508 4888 144412 4904
rect 139508 4832 139524 4888
rect 139580 4832 144340 4888
rect 144396 4832 144412 4888
rect 139508 4816 144412 4832
rect 144660 4888 145196 4904
rect 144660 4832 144676 4888
rect 144732 4832 145196 4888
rect 144660 4816 145196 4832
rect 148020 4888 149900 4904
rect 148020 4832 148036 4888
rect 148092 4832 149828 4888
rect 149884 4832 149900 4888
rect 148020 4816 149900 4832
rect 150932 4888 154828 4904
rect 150932 4832 150948 4888
rect 151004 4832 154756 4888
rect 154812 4832 154828 4888
rect 150932 4816 154828 4832
rect 161124 4888 164684 4904
rect 161124 4832 161140 4888
rect 161196 4832 164612 4888
rect 164668 4832 164684 4888
rect 161124 4816 164684 4832
rect 177700 4888 192012 4904
rect 177700 4832 177716 4888
rect 177772 4832 180628 4888
rect 180684 4832 191940 4888
rect 191996 4832 192012 4888
rect 177700 4816 192012 4832
rect 192148 4888 211836 4904
rect 192148 4832 203700 4888
rect 203756 4832 211764 4888
rect 211820 4832 211836 4888
rect 192148 4816 211836 4832
rect 103220 4724 103308 4816
rect 120244 4724 120332 4816
rect 35684 4708 68028 4724
rect 35684 4652 35700 4708
rect 35756 4652 68028 4708
rect 35684 4636 68028 4652
rect 68164 4708 70380 4724
rect 68164 4652 68180 4708
rect 68236 4652 70308 4708
rect 70364 4652 70380 4708
rect 68164 4636 70380 4652
rect 70516 4708 73180 4724
rect 70516 4652 70532 4708
rect 70588 4652 73108 4708
rect 73164 4652 73180 4708
rect 70516 4636 73180 4652
rect 73316 4708 79900 4724
rect 73316 4652 73332 4708
rect 73388 4652 79828 4708
rect 79884 4652 79900 4708
rect 73316 4636 79900 4652
rect 80036 4708 88188 4724
rect 80036 4652 80052 4708
rect 80108 4652 88116 4708
rect 88172 4652 88188 4708
rect 80036 4636 88188 4652
rect 88324 4708 103308 4724
rect 88324 4652 88340 4708
rect 88396 4652 103308 4708
rect 88324 4636 103308 4652
rect 103892 4708 109692 4724
rect 103892 4652 103908 4708
rect 103964 4652 109620 4708
rect 109676 4652 109692 4708
rect 103892 4636 109692 4652
rect 109828 4708 120108 4724
rect 109828 4652 120036 4708
rect 120092 4652 120108 4708
rect 109828 4636 120108 4652
rect 120244 4708 136236 4724
rect 120244 4652 136164 4708
rect 136220 4652 136236 4708
rect 120244 4636 136236 4652
rect 136372 4708 143292 4724
rect 136372 4652 136388 4708
rect 136444 4652 143220 4708
rect 143276 4652 143292 4708
rect 136372 4636 143292 4652
rect 143428 4708 149452 4724
rect 143428 4652 143444 4708
rect 143500 4652 149380 4708
rect 149436 4652 149452 4708
rect 143428 4636 149452 4652
rect 149700 4708 152812 4724
rect 149700 4652 149716 4708
rect 149772 4652 152740 4708
rect 152796 4652 152812 4708
rect 149700 4636 152812 4652
rect 152948 4708 170956 4724
rect 152948 4652 152964 4708
rect 153020 4652 170884 4708
rect 170940 4652 170956 4708
rect 152948 4636 170956 4652
rect 171428 4708 197948 4724
rect 171428 4652 171444 4708
rect 171500 4652 197876 4708
rect 197932 4652 197948 4708
rect 171428 4636 197948 4652
rect 67940 4544 68028 4636
rect 109828 4544 109916 4636
rect 54164 4528 67804 4544
rect 54164 4472 54180 4528
rect 54236 4472 67804 4528
rect 54164 4456 67804 4472
rect 67940 4528 80572 4544
rect 67940 4472 80500 4528
rect 80556 4472 80572 4528
rect 67940 4456 80572 4472
rect 81492 4528 85948 4544
rect 81492 4472 81508 4528
rect 81564 4472 85876 4528
rect 85932 4472 85948 4528
rect 81492 4456 85948 4472
rect 86084 4528 88748 4544
rect 86084 4472 86100 4528
rect 86156 4472 88676 4528
rect 88732 4472 88748 4528
rect 86084 4456 88748 4472
rect 88884 4528 105772 4544
rect 88884 4472 88900 4528
rect 88956 4472 105700 4528
rect 105756 4472 105772 4528
rect 88884 4456 105772 4472
rect 105908 4528 109580 4544
rect 105908 4472 105924 4528
rect 105980 4472 109580 4528
rect 105908 4456 109580 4472
rect 109716 4528 109916 4544
rect 109716 4472 109732 4528
rect 109788 4472 109916 4528
rect 109716 4456 109916 4472
rect 112516 4528 115740 4544
rect 112516 4472 112532 4528
rect 112588 4472 115668 4528
rect 115724 4472 115740 4528
rect 112516 4456 115740 4472
rect 115988 4528 121452 4544
rect 115988 4472 116004 4528
rect 116060 4472 121380 4528
rect 121436 4472 121452 4528
rect 115988 4456 121452 4472
rect 124276 4528 132763 4544
rect 124276 4472 124292 4528
rect 124348 4472 132763 4528
rect 124276 4456 132763 4472
rect 134356 4528 149676 4544
rect 134356 4472 134372 4528
rect 134428 4472 149604 4528
rect 149660 4472 149676 4528
rect 134356 4456 149676 4472
rect 151044 4528 161548 4544
rect 151044 4472 151060 4528
rect 151116 4472 161476 4528
rect 161532 4472 161548 4528
rect 151044 4456 161548 4472
rect 164820 4528 182268 4544
rect 164820 4472 164836 4528
rect 164892 4472 182196 4528
rect 182252 4472 182268 4528
rect 164820 4456 182268 4472
rect 183076 4528 188988 4544
rect 183076 4472 183092 4528
rect 183148 4472 188916 4528
rect 188972 4472 188988 4528
rect 183076 4456 188988 4472
rect 189236 4528 210044 4544
rect 189236 4472 189252 4528
rect 189308 4472 209972 4528
rect 210028 4472 210044 4528
rect 189236 4456 210044 4472
rect 67716 4364 67804 4456
rect 109492 4364 109580 4456
rect 132675 4364 132763 4456
rect 11604 4348 67580 4364
rect 11604 4292 11620 4348
rect 11676 4292 67508 4348
rect 67564 4292 67580 4348
rect 11604 4276 67580 4292
rect 67716 4348 74076 4364
rect 67716 4292 74004 4348
rect 74060 4292 74076 4348
rect 67716 4276 74076 4292
rect 74212 4348 79004 4364
rect 74212 4292 74228 4348
rect 74284 4292 78932 4348
rect 78988 4292 79004 4348
rect 74212 4276 79004 4292
rect 79140 4348 87516 4364
rect 79140 4292 79156 4348
rect 79212 4292 87444 4348
rect 87500 4292 87516 4348
rect 79140 4276 87516 4292
rect 88100 4348 92220 4364
rect 88100 4292 88116 4348
rect 88172 4292 92148 4348
rect 92204 4292 92220 4348
rect 88100 4276 92220 4292
rect 92356 4348 109356 4364
rect 92356 4292 92372 4348
rect 92428 4292 109284 4348
rect 109340 4292 109356 4348
rect 92356 4276 109356 4292
rect 109492 4348 117420 4364
rect 109492 4292 117348 4348
rect 117404 4292 117420 4348
rect 109492 4276 117420 4292
rect 119236 4348 126380 4364
rect 119236 4292 119252 4348
rect 119308 4292 126308 4348
rect 126364 4292 126380 4348
rect 119236 4276 126380 4292
rect 126516 4348 131756 4364
rect 126516 4292 131684 4348
rect 131740 4292 131756 4348
rect 126516 4276 131756 4292
rect 132675 4348 136124 4364
rect 132675 4292 136052 4348
rect 136108 4292 136124 4348
rect 132675 4276 136124 4292
rect 141076 4348 144412 4364
rect 141076 4292 141092 4348
rect 141148 4292 144340 4348
rect 144396 4292 144412 4348
rect 141076 4276 144412 4292
rect 152836 4348 174988 4364
rect 152836 4292 152852 4348
rect 152908 4292 174916 4348
rect 174972 4292 174988 4348
rect 152836 4276 174988 4292
rect 179380 4348 193244 4364
rect 179380 4292 179396 4348
rect 179452 4292 193172 4348
rect 193228 4292 193244 4348
rect 179380 4276 193244 4292
rect 126516 4184 126604 4276
rect 16420 4168 55372 4184
rect 16420 4112 16436 4168
rect 16492 4112 55300 4168
rect 55356 4112 55372 4168
rect 16420 4096 55372 4112
rect 55508 4168 67132 4184
rect 55508 4112 55524 4168
rect 55580 4112 67060 4168
rect 67116 4112 67132 4168
rect 55508 4096 67132 4112
rect 67940 4168 88412 4184
rect 67940 4112 67956 4168
rect 68012 4112 88340 4168
rect 88396 4112 88412 4168
rect 67940 4096 88412 4112
rect 88548 4168 99500 4184
rect 88548 4112 88564 4168
rect 88620 4112 99428 4168
rect 99484 4112 99500 4168
rect 88548 4096 99500 4112
rect 99636 4168 103980 4184
rect 99636 4112 99652 4168
rect 99708 4112 103980 4168
rect 99636 4096 103980 4112
rect 104116 4168 105996 4184
rect 104116 4112 104132 4168
rect 104188 4112 105924 4168
rect 105980 4112 105996 4168
rect 104116 4096 105996 4112
rect 106132 4168 116076 4184
rect 106132 4112 106148 4168
rect 106204 4112 116004 4168
rect 116060 4112 116076 4168
rect 106132 4096 116076 4112
rect 116212 4168 124252 4184
rect 116212 4112 124180 4168
rect 124236 4112 124252 4168
rect 116212 4096 124252 4112
rect 124388 4096 126604 4184
rect 126852 4168 140156 4184
rect 126852 4112 126868 4168
rect 126924 4112 140084 4168
rect 140140 4112 140156 4168
rect 126852 4096 140156 4112
rect 140292 4168 141612 4184
rect 140292 4112 140308 4168
rect 140364 4112 141540 4168
rect 141596 4112 141612 4168
rect 140292 4096 141612 4112
rect 147908 4168 160988 4184
rect 147908 4112 147924 4168
rect 147980 4112 160916 4168
rect 160972 4112 160988 4168
rect 147908 4096 160988 4112
rect 163140 4168 178348 4184
rect 163140 4112 163156 4168
rect 163212 4112 178276 4168
rect 178332 4112 178348 4168
rect 163140 4096 178348 4112
rect 180388 4168 186412 4184
rect 180388 4112 180404 4168
rect 180460 4112 186340 4168
rect 186396 4112 186412 4168
rect 180388 4096 186412 4112
rect 103892 4004 103980 4096
rect 116212 4004 116300 4096
rect 124388 4004 124476 4096
rect 9588 3988 75196 4004
rect 9588 3932 9604 3988
rect 9660 3932 75124 3988
rect 75180 3932 75196 3988
rect 9588 3916 75196 3932
rect 75332 3988 78332 4004
rect 75332 3932 75348 3988
rect 75404 3932 78260 3988
rect 78316 3932 78332 3988
rect 75332 3916 78332 3932
rect 78468 3988 79452 4004
rect 78468 3932 79380 3988
rect 79436 3932 79452 3988
rect 78468 3916 79452 3932
rect 80596 3988 92332 4004
rect 80596 3932 80612 3988
rect 80668 3932 92260 3988
rect 92316 3932 92332 3988
rect 80596 3916 92332 3932
rect 97396 3988 103756 4004
rect 97396 3932 97412 3988
rect 97468 3932 103684 3988
rect 103740 3932 103756 3988
rect 97396 3916 103756 3932
rect 103892 3988 107676 4004
rect 103892 3932 107604 3988
rect 107660 3932 107676 3988
rect 103892 3916 107676 3932
rect 109380 3988 113836 4004
rect 109380 3932 109396 3988
rect 109452 3932 113764 3988
rect 113820 3932 113836 3988
rect 109380 3916 113836 3932
rect 113972 3988 116300 4004
rect 113972 3932 113988 3988
rect 114044 3932 116300 3988
rect 113972 3916 116300 3932
rect 116436 3988 120668 4004
rect 116436 3932 116452 3988
rect 116508 3932 120596 3988
rect 120652 3932 120668 3988
rect 116436 3916 120668 3932
rect 120804 3988 124476 4004
rect 120804 3932 120820 3988
rect 120876 3932 124476 3988
rect 120804 3916 124476 3932
rect 126068 3988 131532 4004
rect 126068 3932 126084 3988
rect 126140 3932 131460 3988
rect 131516 3932 131532 3988
rect 126068 3916 131532 3932
rect 131668 3988 140604 4004
rect 131668 3932 131684 3988
rect 131740 3932 140532 3988
rect 140588 3932 140604 3988
rect 131668 3916 140604 3932
rect 141300 3988 142732 4004
rect 141300 3932 141316 3988
rect 141372 3932 142660 3988
rect 142716 3932 142732 3988
rect 141300 3916 142732 3932
rect 143988 3988 147660 4004
rect 143988 3932 144004 3988
rect 144060 3932 147660 3988
rect 143988 3916 147660 3932
rect 147796 3988 151132 4004
rect 147796 3932 147812 3988
rect 147868 3932 151060 3988
rect 151116 3932 151132 3988
rect 147796 3916 151132 3932
rect 153844 3988 162332 4004
rect 153844 3932 153860 3988
rect 153916 3932 162260 3988
rect 162316 3932 162332 3988
rect 153844 3916 162332 3932
rect 168068 3988 178124 4004
rect 168068 3932 168084 3988
rect 168140 3932 178052 3988
rect 178108 3932 178124 3988
rect 168068 3916 178124 3932
rect 181508 3988 194924 4004
rect 181508 3932 181524 3988
rect 181580 3932 182980 3988
rect 183036 3932 194852 3988
rect 194908 3932 194924 3988
rect 181508 3916 194924 3932
rect 78468 3824 78556 3916
rect 147572 3824 147660 3916
rect 49236 3808 55596 3824
rect 49236 3752 49252 3808
rect 49308 3752 55524 3808
rect 55580 3752 55596 3808
rect 49236 3736 55596 3752
rect 62116 3808 67020 3824
rect 62116 3752 62132 3808
rect 62188 3752 67020 3808
rect 62116 3736 67020 3752
rect 67156 3808 78556 3824
rect 67156 3752 67172 3808
rect 67228 3752 78556 3808
rect 67156 3736 78556 3752
rect 78692 3808 85723 3824
rect 78692 3752 78708 3808
rect 78764 3752 85723 3808
rect 78692 3736 85723 3752
rect 86196 3808 110364 3824
rect 86196 3752 86212 3808
rect 86268 3752 110292 3808
rect 110348 3752 110364 3808
rect 86196 3736 110364 3752
rect 110612 3808 117532 3824
rect 110612 3752 110628 3808
rect 110684 3752 117460 3808
rect 117516 3752 117532 3808
rect 110612 3736 117532 3752
rect 118900 3808 131084 3824
rect 118900 3752 118916 3808
rect 118972 3752 131012 3808
rect 131068 3752 131084 3808
rect 118900 3736 131084 3752
rect 132788 3808 137916 3824
rect 132788 3752 132804 3808
rect 132860 3752 137916 3808
rect 132788 3736 137916 3752
rect 142532 3808 147436 3824
rect 142532 3752 142548 3808
rect 142604 3752 147364 3808
rect 147420 3752 147436 3808
rect 142532 3736 147436 3752
rect 147572 3808 149452 3824
rect 147572 3752 149380 3808
rect 149436 3752 149452 3808
rect 147572 3736 149452 3752
rect 150932 3808 165692 3824
rect 150932 3752 150948 3808
rect 151004 3752 165620 3808
rect 165676 3752 165692 3808
rect 150932 3736 165692 3752
rect 175124 3808 209708 3824
rect 175124 3752 175140 3808
rect 175196 3752 209636 3808
rect 209692 3752 209708 3808
rect 175124 3736 209708 3752
rect 66932 3644 67020 3736
rect 85635 3644 85723 3736
rect 137828 3644 137916 3736
rect 35460 3628 65452 3644
rect 35460 3572 35476 3628
rect 35532 3572 65380 3628
rect 65436 3572 65452 3628
rect 35460 3556 65452 3572
rect 66932 3628 79900 3644
rect 66932 3572 79828 3628
rect 79884 3572 79900 3628
rect 66932 3556 79900 3572
rect 80820 3628 83484 3644
rect 80820 3572 80836 3628
rect 80892 3572 83412 3628
rect 83468 3572 83484 3628
rect 80820 3556 83484 3572
rect 83620 3628 85164 3644
rect 83620 3572 83636 3628
rect 83692 3572 85092 3628
rect 85148 3572 85164 3628
rect 83620 3556 85164 3572
rect 85635 3556 91324 3644
rect 91460 3628 94124 3644
rect 91460 3572 91476 3628
rect 91532 3572 94052 3628
rect 94108 3572 94124 3628
rect 91460 3556 94124 3572
rect 94260 3628 99724 3644
rect 94260 3572 94276 3628
rect 94332 3572 99652 3628
rect 99708 3572 99724 3628
rect 94260 3556 99724 3572
rect 100980 3628 112604 3644
rect 100980 3572 100996 3628
rect 101052 3572 112532 3628
rect 112588 3572 112604 3628
rect 100980 3556 112604 3572
rect 112740 3628 116412 3644
rect 112740 3572 112756 3628
rect 112812 3572 116340 3628
rect 116396 3572 116412 3628
rect 112740 3556 116412 3572
rect 117220 3628 122684 3644
rect 117220 3572 117236 3628
rect 117292 3572 122612 3628
rect 122668 3572 122684 3628
rect 117220 3556 122684 3572
rect 124276 3628 132092 3644
rect 124276 3572 124292 3628
rect 124348 3572 132020 3628
rect 132076 3572 132092 3628
rect 124276 3556 132092 3572
rect 132228 3628 137692 3644
rect 132228 3572 137620 3628
rect 137676 3572 137692 3628
rect 132228 3556 137692 3572
rect 137828 3628 143964 3644
rect 137828 3572 143892 3628
rect 143948 3572 143964 3628
rect 137828 3556 143964 3572
rect 150596 3628 154716 3644
rect 150596 3572 150612 3628
rect 150668 3572 154644 3628
rect 154700 3572 154716 3628
rect 150596 3556 154716 3572
rect 159556 3628 181484 3644
rect 159556 3572 159572 3628
rect 159628 3572 181412 3628
rect 181468 3572 181484 3628
rect 159556 3556 181484 3572
rect 183524 3628 195036 3644
rect 183524 3572 194964 3628
rect 195020 3572 195036 3628
rect 183524 3556 195036 3572
rect 91236 3464 91324 3556
rect 132228 3464 132316 3556
rect 183524 3464 183612 3556
rect 34228 3448 72284 3464
rect 34228 3392 34244 3448
rect 34300 3392 72212 3448
rect 72268 3392 72284 3448
rect 34228 3376 72284 3392
rect 72980 3448 82252 3464
rect 72980 3392 72996 3448
rect 73052 3392 82180 3448
rect 82236 3392 82252 3448
rect 72980 3376 82252 3392
rect 82388 3448 83484 3464
rect 82388 3392 82404 3448
rect 82460 3392 83412 3448
rect 83468 3392 83484 3448
rect 82388 3376 83484 3392
rect 83844 3448 85724 3464
rect 83844 3392 83860 3448
rect 83916 3392 85724 3448
rect 83844 3376 85724 3392
rect 86308 3448 90876 3464
rect 86308 3392 86324 3448
rect 86380 3392 90876 3448
rect 86308 3376 90876 3392
rect 91236 3448 98940 3464
rect 91236 3392 98868 3448
rect 98924 3392 98940 3448
rect 91236 3376 98940 3392
rect 99076 3448 107788 3464
rect 99076 3392 99092 3448
rect 99148 3392 107716 3448
rect 107772 3392 107788 3448
rect 99076 3376 107788 3392
rect 107924 3448 114508 3464
rect 107924 3392 107940 3448
rect 107996 3392 114508 3448
rect 107924 3376 114508 3392
rect 114756 3448 119436 3464
rect 114756 3392 114772 3448
rect 114828 3392 119364 3448
rect 119420 3392 119436 3448
rect 114756 3376 119436 3392
rect 120020 3448 120780 3464
rect 120020 3392 120036 3448
rect 120092 3392 120708 3448
rect 120764 3392 120780 3448
rect 120020 3376 120780 3392
rect 120916 3448 127164 3464
rect 120916 3392 120932 3448
rect 120988 3392 127092 3448
rect 127148 3392 127164 3448
rect 120916 3376 127164 3392
rect 127300 3376 132316 3464
rect 134356 3448 141052 3464
rect 134356 3392 140980 3448
rect 141036 3392 141052 3448
rect 134356 3376 141052 3392
rect 141188 3448 152700 3464
rect 141188 3392 141204 3448
rect 141260 3392 152628 3448
rect 152684 3392 152700 3448
rect 141188 3376 152700 3392
rect 152835 3448 154828 3464
rect 152835 3392 154756 3448
rect 154812 3392 154828 3448
rect 152835 3376 154828 3392
rect 162804 3448 166364 3464
rect 162804 3392 162820 3448
rect 162876 3392 166292 3448
rect 166348 3392 166364 3448
rect 162804 3376 166364 3392
rect 181284 3448 183612 3464
rect 181284 3392 181300 3448
rect 181356 3392 183612 3448
rect 181284 3376 183612 3392
rect 189572 3448 212844 3464
rect 189572 3392 189588 3448
rect 189644 3392 212772 3448
rect 212828 3392 212844 3448
rect 189572 3376 212844 3392
rect 85636 3284 85724 3376
rect 90788 3284 90876 3376
rect 114420 3284 114508 3376
rect 127300 3284 127388 3376
rect 33892 3268 49548 3284
rect 33892 3212 33908 3268
rect 33964 3212 49548 3268
rect 33892 3196 49548 3212
rect 49684 3268 55148 3284
rect 49684 3212 49700 3268
rect 49756 3212 55076 3268
rect 55132 3212 55148 3268
rect 49684 3196 55148 3212
rect 55284 3268 65564 3284
rect 55284 3212 55300 3268
rect 55356 3212 65492 3268
rect 65548 3212 65564 3268
rect 55284 3196 65564 3212
rect 67716 3268 74636 3284
rect 67716 3212 67732 3268
rect 67788 3212 74564 3268
rect 74620 3212 74636 3268
rect 67716 3196 74636 3212
rect 74884 3268 76988 3284
rect 74884 3212 74900 3268
rect 74956 3212 76916 3268
rect 76972 3212 76988 3268
rect 74884 3196 76988 3212
rect 77348 3268 77996 3284
rect 77348 3212 77364 3268
rect 77420 3212 77924 3268
rect 77980 3212 77996 3268
rect 77348 3196 77996 3212
rect 79028 3268 81580 3284
rect 79028 3212 79044 3268
rect 79100 3212 81508 3268
rect 81564 3212 81580 3268
rect 79028 3196 81580 3212
rect 81940 3268 85388 3284
rect 81940 3212 81956 3268
rect 82012 3212 85316 3268
rect 85372 3212 85388 3268
rect 81940 3196 85388 3212
rect 85636 3268 90652 3284
rect 85636 3212 90580 3268
rect 90636 3212 90652 3268
rect 85636 3196 90652 3212
rect 90788 3196 91772 3284
rect 95604 3268 102412 3284
rect 95604 3212 95620 3268
rect 95676 3212 102340 3268
rect 102396 3212 102412 3268
rect 95604 3196 102412 3212
rect 102548 3268 114284 3284
rect 102548 3212 102564 3268
rect 102620 3212 114212 3268
rect 114268 3212 114284 3268
rect 102548 3196 114284 3212
rect 114420 3268 124476 3284
rect 114420 3212 124404 3268
rect 124460 3212 124476 3268
rect 114420 3196 124476 3212
rect 124612 3268 127388 3284
rect 124612 3212 124628 3268
rect 124684 3212 127388 3268
rect 124612 3196 127388 3212
rect 129652 3268 132764 3284
rect 129652 3212 129668 3268
rect 129724 3212 132692 3268
rect 132748 3212 132764 3268
rect 129652 3196 132764 3212
rect 28740 3088 49324 3104
rect 28740 3032 28756 3088
rect 28812 3032 49252 3088
rect 49308 3032 49324 3088
rect 28740 3016 49324 3032
rect 49460 2924 49548 3196
rect 64132 3088 75196 3104
rect 64132 3032 64148 3088
rect 64204 3032 75124 3088
rect 75180 3032 75196 3088
rect 64132 3016 75196 3032
rect 75444 3088 91548 3104
rect 75444 3032 75460 3088
rect 75516 3032 91548 3088
rect 75444 3016 91548 3032
rect 17764 2908 49100 2924
rect 17764 2852 17780 2908
rect 17836 2852 49028 2908
rect 49084 2852 49100 2908
rect 17764 2836 49100 2852
rect 49460 2836 50220 2924
rect 59204 2908 82028 2924
rect 59204 2852 59220 2908
rect 59276 2852 81956 2908
rect 82012 2852 82028 2908
rect 59204 2836 82028 2852
rect 82164 2908 86620 2924
rect 82164 2852 82180 2908
rect 82236 2852 86548 2908
rect 86604 2852 86620 2908
rect 82164 2836 86620 2852
rect 86756 2908 91324 2924
rect 86756 2852 86772 2908
rect 86828 2852 91252 2908
rect 91308 2852 91324 2908
rect 86756 2836 91324 2852
rect 50132 2744 50220 2836
rect 91460 2744 91548 3016
rect 91684 2924 91772 3196
rect 134356 3104 134444 3376
rect 152835 3284 152923 3376
rect 138724 3268 145644 3284
rect 138724 3212 138740 3268
rect 138796 3212 145572 3268
rect 145628 3212 145644 3268
rect 138724 3196 145644 3212
rect 145780 3268 151132 3284
rect 145780 3212 151060 3268
rect 151116 3212 151132 3268
rect 145780 3196 151132 3212
rect 151268 3268 152923 3284
rect 151268 3212 151284 3268
rect 151340 3212 152923 3268
rect 151268 3196 152923 3212
rect 154516 3268 170508 3284
rect 154516 3212 154532 3268
rect 154588 3212 170436 3268
rect 170492 3212 170508 3268
rect 154516 3196 170508 3212
rect 172995 3268 186188 3284
rect 172995 3212 186116 3268
rect 186172 3212 186188 3268
rect 172995 3196 186188 3212
rect 187332 3268 201644 3284
rect 187332 3212 187348 3268
rect 187404 3212 201572 3268
rect 201628 3212 201644 3268
rect 187332 3196 201644 3212
rect 145780 3104 145868 3196
rect 172995 3104 173083 3196
rect 91908 3088 97932 3104
rect 91908 3032 91924 3088
rect 91980 3032 97860 3088
rect 97916 3032 97932 3088
rect 91908 3016 97932 3032
rect 98068 3088 106220 3104
rect 98068 3032 98084 3088
rect 98140 3032 106148 3088
rect 106204 3032 106220 3088
rect 98068 3016 106220 3032
rect 107364 3088 115740 3104
rect 107364 3032 107380 3088
rect 107436 3032 115668 3088
rect 115724 3032 115740 3088
rect 107364 3016 115740 3032
rect 115876 3088 118652 3104
rect 115876 3032 115892 3088
rect 115948 3032 118580 3088
rect 118636 3032 118652 3088
rect 115876 3016 118652 3032
rect 119236 3088 121788 3104
rect 119236 3032 119252 3088
rect 119308 3032 121716 3088
rect 121772 3032 121788 3088
rect 119236 3016 121788 3032
rect 121924 3088 134444 3104
rect 121924 3032 121940 3088
rect 121996 3032 134444 3088
rect 121924 3016 134444 3032
rect 136036 3088 145868 3104
rect 136036 3032 136052 3088
rect 136108 3032 145868 3088
rect 136036 3016 145868 3032
rect 146004 3088 148108 3104
rect 146004 3032 146020 3088
rect 146076 3032 148036 3088
rect 148092 3032 148108 3088
rect 146004 3016 148108 3032
rect 150260 3088 156283 3104
rect 150260 3032 150276 3088
rect 150332 3032 156283 3088
rect 150260 3016 156283 3032
rect 167844 3088 173083 3104
rect 167844 3032 167860 3088
rect 167916 3032 173083 3088
rect 167844 3016 173083 3032
rect 181396 3088 211388 3104
rect 181396 3032 181412 3088
rect 181468 3032 211316 3088
rect 211372 3032 211388 3088
rect 181396 3016 211388 3032
rect 156195 2924 156283 3016
rect 91684 2908 100060 2924
rect 91684 2852 99988 2908
rect 100044 2852 100060 2908
rect 91684 2836 100060 2852
rect 100196 2908 102636 2924
rect 100196 2852 100212 2908
rect 100268 2852 102564 2908
rect 102620 2852 102636 2908
rect 100196 2836 102636 2852
rect 102772 2908 117756 2924
rect 102772 2852 102788 2908
rect 102844 2852 117684 2908
rect 117740 2852 117756 2908
rect 102772 2836 117756 2852
rect 118116 2908 132763 2924
rect 118116 2852 118132 2908
rect 118188 2852 132763 2908
rect 118116 2836 132763 2852
rect 134580 2908 136012 2924
rect 134580 2852 134596 2908
rect 134652 2852 135940 2908
rect 135996 2852 136012 2908
rect 134580 2836 136012 2852
rect 136148 2908 154492 2924
rect 136148 2852 136164 2908
rect 136220 2852 154420 2908
rect 154476 2852 154492 2908
rect 136148 2836 154492 2852
rect 156195 2908 166700 2924
rect 156195 2852 166628 2908
rect 166684 2852 166700 2908
rect 156195 2836 166700 2852
rect 167060 2908 187980 2924
rect 167060 2852 167076 2908
rect 167132 2852 187908 2908
rect 187964 2852 187980 2908
rect 167060 2836 187980 2852
rect 188340 2908 189436 2924
rect 188340 2852 188356 2908
rect 188412 2852 189436 2908
rect 188340 2836 189436 2852
rect 190692 2908 198284 2924
rect 190692 2852 190708 2908
rect 190764 2852 198212 2908
rect 198268 2852 198284 2908
rect 190692 2836 198284 2852
rect 132675 2744 132763 2836
rect 189348 2744 189436 2836
rect 25156 2728 49996 2744
rect 25156 2672 25172 2728
rect 25228 2672 49924 2728
rect 49980 2672 49996 2728
rect 25156 2656 49996 2672
rect 50132 2728 67468 2744
rect 50132 2672 67396 2728
rect 67452 2672 67468 2728
rect 50132 2656 67468 2672
rect 68052 2728 73852 2744
rect 68052 2672 68068 2728
rect 68124 2672 73780 2728
rect 73836 2672 73852 2728
rect 68052 2656 73852 2672
rect 73988 2728 84940 2744
rect 73988 2672 74004 2728
rect 74060 2672 84868 2728
rect 84924 2672 84940 2728
rect 73988 2656 84940 2672
rect 85076 2656 91324 2744
rect 91460 2728 103532 2744
rect 91460 2672 103460 2728
rect 103516 2672 103532 2728
rect 91460 2656 103532 2672
rect 103668 2728 122012 2744
rect 103668 2672 103684 2728
rect 103740 2672 121940 2728
rect 121996 2672 122012 2728
rect 103668 2656 122012 2672
rect 122372 2728 129740 2744
rect 122372 2672 122388 2728
rect 122444 2672 129668 2728
rect 129724 2672 129740 2728
rect 122372 2656 129740 2672
rect 132675 2728 136908 2744
rect 132675 2672 136836 2728
rect 136892 2672 136908 2728
rect 132675 2656 136908 2672
rect 139060 2728 142956 2744
rect 139060 2672 142884 2728
rect 142940 2672 142956 2728
rect 139060 2656 142956 2672
rect 145556 2728 151356 2744
rect 145556 2672 145572 2728
rect 145628 2672 151284 2728
rect 151340 2672 151356 2728
rect 145556 2656 151356 2672
rect 151492 2728 163788 2744
rect 151492 2672 151508 2728
rect 151564 2672 163716 2728
rect 163772 2672 163788 2728
rect 151492 2656 163788 2672
rect 165604 2728 189212 2744
rect 165604 2672 165620 2728
rect 165676 2672 189140 2728
rect 189196 2672 189212 2728
rect 165604 2656 189212 2672
rect 189348 2728 197724 2744
rect 189348 2672 197652 2728
rect 197708 2672 197724 2728
rect 189348 2656 197724 2672
rect 85076 2564 85164 2656
rect 91236 2564 91324 2656
rect 139060 2564 139148 2656
rect 18436 2548 53468 2564
rect 18436 2492 18452 2548
rect 18508 2492 53468 2548
rect 18436 2476 53468 2492
rect 58756 2548 65116 2564
rect 58756 2492 58772 2548
rect 58828 2492 65044 2548
rect 65100 2492 65116 2548
rect 58756 2476 65116 2492
rect 65476 2548 80572 2564
rect 65476 2492 65492 2548
rect 65548 2492 80500 2548
rect 80556 2492 80572 2548
rect 65476 2476 80572 2492
rect 80708 2476 85164 2564
rect 85300 2548 88972 2564
rect 85300 2492 85316 2548
rect 85372 2492 88900 2548
rect 88956 2492 88972 2548
rect 85300 2476 88972 2492
rect 89108 2548 91100 2564
rect 89108 2492 89124 2548
rect 89180 2492 91028 2548
rect 91084 2492 91100 2548
rect 89108 2476 91100 2492
rect 91236 2548 95692 2564
rect 91236 2492 95620 2548
rect 95676 2492 95692 2548
rect 91236 2476 95692 2492
rect 95828 2548 104092 2564
rect 95828 2492 104020 2548
rect 104076 2492 104092 2548
rect 95828 2476 104092 2492
rect 106132 2548 108572 2564
rect 106132 2492 106148 2548
rect 106204 2492 108500 2548
rect 108556 2492 108572 2548
rect 106132 2476 108572 2492
rect 110388 2548 114844 2564
rect 110388 2492 110404 2548
rect 110460 2492 114772 2548
rect 114828 2492 114844 2548
rect 110388 2476 114844 2492
rect 114980 2548 121004 2564
rect 114980 2492 114996 2548
rect 115052 2492 120932 2548
rect 120988 2492 121004 2548
rect 114980 2476 121004 2492
rect 121140 2548 135788 2564
rect 121140 2492 121156 2548
rect 121212 2492 135716 2548
rect 135772 2492 135788 2548
rect 121140 2476 135788 2492
rect 135924 2548 139148 2564
rect 135924 2492 135940 2548
rect 135996 2492 139148 2548
rect 135924 2476 139148 2492
rect 142756 2548 146092 2564
rect 142756 2492 142772 2548
rect 142828 2492 146020 2548
rect 146076 2492 146092 2548
rect 142756 2476 146092 2492
rect 146228 2548 156060 2564
rect 146228 2492 146244 2548
rect 146300 2492 155988 2548
rect 156044 2492 156060 2548
rect 146228 2476 156060 2492
rect 156195 2548 181596 2564
rect 156195 2492 156211 2548
rect 156267 2492 181524 2548
rect 181580 2492 181596 2548
rect 156195 2476 181596 2492
rect 183076 2548 190780 2564
rect 183076 2492 183092 2548
rect 183148 2492 184436 2548
rect 184492 2492 190708 2548
rect 190764 2492 190780 2548
rect 183076 2476 190780 2492
rect 53380 2384 53468 2476
rect 80708 2384 80796 2476
rect 95828 2384 95916 2476
rect 49012 2368 53244 2384
rect 49012 2312 49028 2368
rect 49084 2312 53172 2368
rect 53228 2312 53244 2368
rect 49012 2296 53244 2312
rect 53380 2368 60412 2384
rect 53380 2312 60340 2368
rect 60396 2312 60412 2368
rect 53380 2296 60412 2312
rect 60548 2368 67804 2384
rect 60548 2312 67732 2368
rect 67788 2312 67804 2368
rect 60548 2296 67804 2312
rect 67940 2368 76540 2384
rect 67940 2312 76468 2368
rect 76524 2312 76540 2368
rect 67940 2296 76540 2312
rect 76900 2368 80796 2384
rect 76900 2312 76916 2368
rect 76972 2312 80796 2368
rect 76900 2296 80796 2312
rect 81044 2368 82812 2384
rect 81044 2312 81060 2368
rect 81116 2312 82740 2368
rect 82796 2312 82812 2368
rect 81044 2296 82812 2312
rect 83284 2368 91884 2384
rect 83284 2312 83300 2368
rect 83356 2312 91812 2368
rect 91868 2312 91884 2368
rect 83284 2296 91884 2312
rect 92020 2368 95916 2384
rect 92020 2312 92036 2368
rect 92092 2312 95916 2368
rect 92020 2296 95916 2312
rect 96500 2368 99163 2384
rect 96500 2312 96516 2368
rect 96572 2312 99163 2368
rect 96500 2296 99163 2312
rect 99300 2368 103980 2384
rect 99300 2312 99316 2368
rect 99372 2312 103908 2368
rect 103964 2312 103980 2368
rect 99300 2296 103980 2312
rect 104116 2368 117644 2384
rect 104116 2312 104132 2368
rect 104188 2312 117572 2368
rect 117628 2312 117644 2368
rect 104116 2296 117644 2312
rect 119124 2368 132763 2384
rect 119124 2312 119140 2368
rect 119196 2312 132763 2368
rect 119124 2296 132763 2312
rect 134244 2368 149564 2384
rect 134244 2312 134260 2368
rect 134316 2312 149492 2368
rect 149548 2312 149564 2368
rect 134244 2296 149564 2312
rect 150820 2368 178236 2384
rect 150820 2312 150836 2368
rect 150892 2312 178164 2368
rect 178220 2312 178236 2368
rect 150820 2296 178236 2312
rect 179604 2368 191676 2384
rect 179604 2312 179620 2368
rect 179676 2312 191604 2368
rect 191660 2312 191676 2368
rect 179604 2296 191676 2312
rect 60548 2204 60636 2296
rect 67940 2204 68028 2296
rect 99075 2204 99163 2296
rect 33668 2188 55372 2204
rect 33668 2132 33684 2188
rect 33740 2132 55300 2188
rect 55356 2132 55372 2188
rect 33668 2116 55372 2132
rect 55508 2188 60636 2204
rect 55508 2132 55524 2188
rect 55580 2132 60636 2188
rect 55508 2116 60636 2132
rect 60772 2188 68028 2204
rect 60772 2132 60788 2188
rect 60844 2132 68028 2188
rect 60772 2116 68028 2132
rect 70516 2188 81020 2204
rect 70516 2132 70532 2188
rect 70588 2132 80948 2188
rect 81004 2132 81020 2188
rect 70516 2116 81020 2132
rect 81156 2188 85388 2204
rect 81156 2132 81172 2188
rect 81228 2132 85316 2188
rect 85372 2132 85388 2188
rect 81156 2116 85388 2132
rect 85524 2188 86396 2204
rect 85524 2132 85540 2188
rect 85596 2132 86324 2188
rect 86380 2132 86396 2188
rect 85524 2116 86396 2132
rect 86532 2188 91212 2204
rect 86532 2132 86548 2188
rect 86604 2132 91140 2188
rect 91196 2132 91212 2188
rect 86532 2116 91212 2132
rect 91460 2188 98940 2204
rect 91460 2132 91476 2188
rect 91532 2132 98868 2188
rect 98924 2132 98940 2188
rect 91460 2116 98940 2132
rect 99075 2188 106780 2204
rect 99075 2132 106708 2188
rect 106764 2132 106780 2188
rect 99075 2116 106780 2132
rect 108820 2188 111036 2204
rect 108820 2132 108836 2188
rect 108892 2132 110964 2188
rect 111020 2132 111036 2188
rect 108820 2116 111036 2132
rect 111284 2188 113948 2204
rect 111284 2132 111300 2188
rect 111356 2132 113876 2188
rect 113932 2132 113948 2188
rect 111284 2116 113948 2132
rect 114196 2188 115516 2204
rect 114196 2132 114212 2188
rect 114268 2132 115516 2188
rect 114196 2116 115516 2132
rect 115764 2188 116860 2204
rect 115764 2132 115780 2188
rect 115836 2132 116788 2188
rect 116844 2132 116860 2188
rect 115764 2116 116860 2132
rect 116996 2188 122460 2204
rect 116996 2132 117012 2188
rect 117068 2132 122388 2188
rect 122444 2132 122460 2188
rect 116996 2116 122460 2132
rect 122596 2188 126044 2204
rect 122596 2132 122612 2188
rect 122668 2132 125972 2188
rect 126028 2132 126044 2188
rect 122596 2116 126044 2132
rect 115428 2024 115516 2116
rect 132675 2024 132763 2296
rect 137828 2188 157852 2204
rect 137828 2132 137844 2188
rect 137900 2132 157780 2188
rect 157836 2132 157852 2188
rect 137828 2116 157852 2132
rect 157988 2188 191564 2204
rect 157988 2132 158004 2188
rect 158060 2132 191492 2188
rect 191548 2132 191564 2188
rect 157988 2116 191564 2132
rect 191700 2188 197388 2204
rect 191700 2132 191716 2188
rect 191772 2132 197316 2188
rect 197372 2132 197388 2188
rect 191700 2116 197388 2132
rect 203235 2188 203660 2204
rect 203235 2132 203588 2188
rect 203644 2132 203660 2188
rect 203235 2116 203660 2132
rect 203235 2024 203323 2116
rect 53604 2008 62540 2024
rect 53604 1952 53620 2008
rect 53676 1952 62468 2008
rect 62524 1952 62540 2008
rect 53604 1936 62540 1952
rect 62788 2008 73516 2024
rect 62788 1952 62804 2008
rect 62860 1952 73444 2008
rect 73500 1952 73516 2008
rect 62788 1936 73516 1952
rect 73764 2008 82364 2024
rect 73764 1952 73780 2008
rect 73836 1952 82292 2008
rect 82348 1952 82364 2008
rect 73764 1936 82364 1952
rect 82724 2008 115292 2024
rect 82724 1952 82740 2008
rect 82796 1952 115220 2008
rect 115276 1952 115292 2008
rect 82724 1936 115292 1952
rect 115428 2008 117420 2024
rect 115428 1952 117348 2008
rect 117404 1952 117420 2008
rect 115428 1936 117420 1952
rect 117668 2008 126828 2024
rect 117668 1952 117684 2008
rect 117740 1952 126828 2008
rect 117668 1936 126828 1952
rect 132675 2008 138812 2024
rect 132675 1952 138740 2008
rect 138796 1952 138812 2008
rect 132675 1936 138812 1952
rect 145220 2008 147660 2024
rect 145220 1952 145236 2008
rect 145292 1952 147588 2008
rect 147644 1952 147660 2008
rect 145220 1936 147660 1952
rect 147796 2008 151132 2024
rect 147796 1952 147812 2008
rect 147868 1952 151060 2008
rect 151116 1952 151132 2008
rect 147796 1936 151132 1952
rect 151940 2008 185964 2024
rect 151940 1952 151956 2008
rect 152012 1952 185892 2008
rect 185948 1952 185964 2008
rect 151940 1936 185964 1952
rect 186436 2008 188540 2024
rect 186436 1952 186452 2008
rect 186508 1952 188468 2008
rect 188524 1952 188540 2008
rect 186436 1936 188540 1952
rect 188676 2008 203323 2024
rect 188676 1952 188692 2008
rect 188748 1952 203323 2008
rect 188676 1936 203323 1952
rect 126740 1844 126828 1936
rect 50132 1828 74412 1844
rect 50132 1772 50148 1828
rect 50204 1772 74340 1828
rect 74396 1772 74412 1828
rect 50132 1756 74412 1772
rect 74548 1828 83260 1844
rect 74548 1772 74564 1828
rect 74620 1772 83188 1828
rect 83244 1772 83260 1828
rect 74548 1756 83260 1772
rect 83956 1828 91548 1844
rect 83956 1772 91476 1828
rect 91532 1772 91548 1828
rect 83956 1756 91548 1772
rect 91684 1828 102300 1844
rect 91684 1772 91700 1828
rect 91756 1772 102228 1828
rect 102284 1772 102300 1828
rect 91684 1756 102300 1772
rect 102436 1828 122572 1844
rect 102436 1772 102452 1828
rect 102508 1772 122500 1828
rect 122556 1772 122572 1828
rect 102436 1756 122572 1772
rect 122708 1828 126268 1844
rect 122708 1772 122724 1828
rect 122780 1772 126196 1828
rect 126252 1772 126268 1828
rect 122708 1756 126268 1772
rect 126740 1828 147772 1844
rect 126740 1772 147700 1828
rect 147756 1772 147772 1828
rect 126740 1756 147772 1772
rect 147908 1828 151804 1844
rect 147908 1772 147924 1828
rect 147980 1772 151732 1828
rect 151788 1772 151804 1828
rect 147908 1756 151804 1772
rect 153732 1828 187420 1844
rect 153732 1772 153748 1828
rect 153804 1772 187348 1828
rect 187404 1772 187420 1828
rect 153732 1756 187420 1772
rect 187668 1828 198284 1844
rect 187668 1772 187684 1828
rect 187740 1772 198212 1828
rect 198268 1772 198284 1828
rect 187668 1756 198284 1772
rect 83956 1664 84044 1756
rect 59876 1648 71948 1664
rect 59876 1592 59892 1648
rect 59948 1592 71876 1648
rect 71932 1592 71948 1648
rect 59876 1576 71948 1592
rect 72084 1648 84044 1664
rect 72084 1592 72100 1648
rect 72156 1592 84044 1648
rect 72084 1576 84044 1592
rect 84180 1648 97820 1664
rect 84180 1592 97748 1648
rect 97804 1592 97820 1648
rect 84180 1576 97820 1592
rect 98964 1648 117196 1664
rect 98964 1592 98980 1648
rect 99036 1592 117124 1648
rect 117180 1592 117196 1648
rect 98964 1576 117196 1592
rect 117444 1648 124364 1664
rect 117444 1592 117460 1648
rect 117516 1592 124292 1648
rect 124348 1592 124364 1648
rect 117444 1576 124364 1592
rect 134132 1648 136012 1664
rect 134132 1592 134148 1648
rect 134204 1592 136012 1648
rect 134132 1576 136012 1592
rect 140404 1648 204444 1664
rect 140404 1592 140420 1648
rect 140476 1592 204372 1648
rect 204428 1592 204444 1648
rect 140404 1576 204444 1592
rect 84180 1484 84268 1576
rect 34564 1468 79788 1484
rect 34564 1412 34580 1468
rect 34636 1412 79716 1468
rect 79772 1412 79788 1468
rect 34564 1396 79788 1412
rect 79924 1468 81244 1484
rect 79924 1412 79940 1468
rect 79996 1412 81172 1468
rect 81228 1412 81244 1468
rect 79924 1396 81244 1412
rect 81380 1468 82364 1484
rect 81380 1412 81396 1468
rect 81452 1412 82292 1468
rect 82348 1412 82364 1468
rect 81380 1396 82364 1412
rect 82500 1468 82588 1484
rect 82500 1412 82516 1468
rect 82572 1412 82588 1468
rect 82500 1304 82588 1412
rect 82948 1468 84268 1484
rect 82948 1412 82964 1468
rect 83020 1412 84268 1468
rect 82948 1396 84268 1412
rect 84516 1468 86508 1484
rect 84516 1412 84532 1468
rect 84588 1412 86436 1468
rect 86492 1412 86508 1468
rect 84516 1396 86508 1412
rect 86980 1468 127612 1484
rect 86980 1412 86996 1468
rect 87052 1412 127540 1468
rect 127596 1412 127612 1468
rect 86980 1396 127612 1412
rect 128420 1468 135676 1484
rect 128420 1412 128436 1468
rect 128492 1412 135604 1468
rect 135660 1412 135676 1468
rect 128420 1396 135676 1412
rect 135924 1304 136012 1576
rect 136148 1468 168044 1484
rect 136148 1412 136164 1468
rect 136220 1412 167972 1468
rect 168028 1412 168044 1468
rect 136148 1396 168044 1412
rect 201556 1468 211164 1484
rect 201556 1412 201572 1468
rect 201628 1412 211092 1468
rect 211148 1412 211164 1468
rect 201556 1396 211164 1412
rect 2532 1288 23116 1304
rect 2532 1232 2548 1288
rect 2604 1232 23044 1288
rect 23100 1232 23116 1288
rect 2532 1216 23116 1232
rect 42404 1288 75868 1304
rect 42404 1232 42420 1288
rect 42476 1232 75796 1288
rect 75852 1232 75868 1288
rect 42404 1216 75868 1232
rect 76228 1288 79452 1304
rect 76228 1232 76244 1288
rect 76300 1232 79380 1288
rect 79436 1232 79452 1288
rect 76228 1216 79452 1232
rect 79588 1288 82364 1304
rect 79588 1232 82292 1288
rect 82348 1232 82364 1288
rect 79588 1216 82364 1232
rect 82500 1288 107676 1304
rect 82500 1232 107604 1288
rect 107660 1232 107676 1288
rect 82500 1216 107676 1232
rect 109044 1288 109468 1304
rect 109044 1232 109060 1288
rect 109116 1232 109396 1288
rect 109452 1232 109468 1288
rect 109044 1216 109468 1232
rect 109604 1288 115516 1304
rect 109604 1232 109620 1288
rect 109676 1232 115444 1288
rect 115500 1232 115516 1288
rect 109604 1216 115516 1232
rect 115652 1288 120668 1304
rect 115652 1232 115668 1288
rect 115724 1232 120668 1288
rect 115652 1216 120668 1232
rect 120804 1288 123580 1304
rect 120804 1232 120820 1288
rect 120876 1232 123508 1288
rect 123564 1232 123580 1288
rect 120804 1216 123580 1232
rect 123940 1288 134556 1304
rect 123940 1232 123956 1288
rect 124012 1232 134484 1288
rect 134540 1232 134556 1288
rect 123940 1216 134556 1232
rect 135924 1288 142284 1304
rect 135924 1232 142212 1288
rect 142268 1232 142284 1288
rect 135924 1216 142284 1232
rect 143988 1288 145084 1304
rect 143988 1232 144004 1288
rect 144060 1232 145012 1288
rect 145068 1232 145084 1288
rect 143988 1216 145084 1232
rect 194052 1288 203100 1304
rect 194052 1232 194068 1288
rect 194124 1232 203028 1288
rect 203084 1232 203100 1288
rect 194052 1216 203100 1232
rect 79588 1124 79676 1216
rect 120580 1124 120668 1216
rect 1300 1108 21212 1124
rect 1300 1052 1316 1108
rect 1372 1052 21140 1108
rect 21196 1052 21212 1108
rect 1300 1036 21212 1052
rect 26388 1108 60412 1124
rect 26388 1052 26404 1108
rect 26460 1052 60340 1108
rect 60396 1052 60412 1108
rect 26388 1036 60412 1052
rect 60548 1108 79676 1124
rect 60548 1052 60564 1108
rect 60620 1052 79676 1108
rect 60548 1036 79676 1052
rect 79812 1108 87068 1124
rect 79812 1052 79828 1108
rect 79884 1052 86996 1108
rect 87052 1052 87068 1108
rect 79812 1036 87068 1052
rect 87204 1108 97372 1124
rect 87204 1052 87220 1108
rect 87276 1052 97300 1108
rect 97356 1052 97372 1108
rect 87204 1036 97372 1052
rect 97508 1108 101628 1124
rect 97508 1052 97524 1108
rect 97580 1052 101556 1108
rect 101612 1052 101628 1108
rect 97508 1036 101628 1052
rect 101764 1108 120444 1124
rect 101764 1052 101780 1108
rect 101836 1052 120372 1108
rect 120428 1052 120444 1108
rect 101764 1036 120444 1052
rect 120580 1108 122348 1124
rect 120580 1052 122276 1108
rect 122332 1052 122348 1108
rect 120580 1036 122348 1052
rect 122820 1108 136012 1124
rect 122820 1052 122836 1108
rect 122892 1052 135940 1108
rect 135996 1052 136012 1108
rect 122820 1036 136012 1052
rect 145668 1108 195260 1124
rect 145668 1052 145684 1108
rect 145740 1052 195188 1108
rect 195244 1052 195260 1108
rect 145668 1036 195260 1052
rect 18212 928 40476 944
rect 18212 872 18228 928
rect 18284 872 40404 928
rect 40460 872 40476 928
rect 18212 856 40476 872
rect 50355 928 76428 944
rect 50355 872 76356 928
rect 76412 872 76428 928
rect 50355 856 76428 872
rect 76564 928 94124 944
rect 76564 872 94052 928
rect 94108 872 94124 928
rect 76564 856 94124 872
rect 97396 928 100396 944
rect 97396 872 97412 928
rect 97468 872 100324 928
rect 100380 872 100396 928
rect 97396 856 100396 872
rect 100532 928 106444 944
rect 100532 872 100548 928
rect 100604 872 106372 928
rect 106428 872 106444 928
rect 100532 856 106444 872
rect 107476 928 125932 944
rect 107476 872 107492 928
rect 107548 872 125860 928
rect 125916 872 125932 928
rect 107476 856 125932 872
rect 137716 928 192908 944
rect 137716 872 137732 928
rect 137788 872 192836 928
rect 192892 872 192908 928
rect 137716 856 192908 872
rect 198196 928 212956 944
rect 198196 872 198212 928
rect 198268 872 212884 928
rect 212940 872 212956 928
rect 198196 856 212956 872
rect 50355 764 50443 856
rect 76564 764 76652 856
rect 18100 748 41036 764
rect 18100 692 18116 748
rect 18172 692 40964 748
rect 41020 692 41036 748
rect 18100 676 41036 692
rect 48676 748 50443 764
rect 48676 692 48692 748
rect 48748 692 50443 748
rect 48676 676 50443 692
rect 68500 748 72060 764
rect 68500 692 68516 748
rect 68572 692 71988 748
rect 72044 692 72060 748
rect 68500 676 72060 692
rect 72196 748 76652 764
rect 72196 692 72212 748
rect 72268 692 76652 748
rect 72196 676 76652 692
rect 76788 748 101852 764
rect 76788 692 76804 748
rect 76860 692 101780 748
rect 101836 692 101852 748
rect 76788 676 101852 692
rect 101988 748 106108 764
rect 101988 692 102004 748
rect 102060 692 106036 748
rect 106092 692 106108 748
rect 101988 676 106108 692
rect 107588 748 151132 764
rect 107588 692 107604 748
rect 107660 692 151060 748
rect 151116 692 151132 748
rect 107588 676 151132 692
rect 1972 568 23452 584
rect 1972 512 1988 568
rect 2044 512 23380 568
rect 23436 512 23452 568
rect 1972 496 23452 512
rect 25940 568 52236 584
rect 25940 512 25956 568
rect 26012 512 52164 568
rect 52220 512 52236 568
rect 25940 496 52236 512
rect 57300 568 68140 584
rect 57300 512 57316 568
rect 57372 512 68140 568
rect 57300 496 68140 512
rect 72084 568 109468 584
rect 72084 512 72100 568
rect 72156 512 109396 568
rect 109452 512 109468 568
rect 72084 496 109468 512
rect 109604 568 111148 584
rect 109604 512 109620 568
rect 109676 512 111076 568
rect 111132 512 111148 568
rect 109604 496 111148 512
rect 111396 568 117868 584
rect 111396 512 111412 568
rect 111468 512 117796 568
rect 117852 512 117868 568
rect 111396 496 117868 512
rect 118788 568 124028 584
rect 118788 512 118804 568
rect 118860 512 123956 568
rect 124012 512 124028 568
rect 118788 496 124028 512
rect 124164 568 205676 584
rect 124164 512 124180 568
rect 124236 512 205604 568
rect 205660 512 205676 568
rect 124164 496 205676 512
rect 19668 388 67916 404
rect 19668 332 19684 388
rect 19740 332 67844 388
rect 67900 332 67916 388
rect 19668 316 67916 332
rect 68052 224 68140 496
rect 75220 388 78220 404
rect 75220 332 75236 388
rect 75292 332 78148 388
rect 78204 332 78220 388
rect 75220 316 78220 332
rect 78356 388 82252 404
rect 78356 332 78372 388
rect 78428 332 82180 388
rect 82236 332 82252 388
rect 78356 316 82252 332
rect 83284 388 197164 404
rect 83284 332 83300 388
rect 83356 332 197092 388
rect 197148 332 197164 388
rect 83284 316 197164 332
rect 197300 388 217212 404
rect 197300 332 197316 388
rect 197372 332 217140 388
rect 217196 332 217212 388
rect 197300 316 217212 332
rect 15972 208 49884 224
rect 15972 152 15988 208
rect 16044 152 49812 208
rect 49868 152 49884 208
rect 15972 136 49884 152
rect 63236 208 67804 224
rect 63236 152 63252 208
rect 63308 152 67732 208
rect 67788 152 67804 208
rect 63236 136 67804 152
rect 68052 208 77436 224
rect 68052 152 77364 208
rect 77420 152 77436 208
rect 68052 136 77436 152
rect 77572 208 206908 224
rect 77572 152 77588 208
rect 77644 152 206836 208
rect 206892 152 206908 208
rect 77572 136 206908 152
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__000__I pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 87920 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__001__I
timestamp 1654395037
transform -1 0 88592 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__002__I
timestamp 1654395037
transform 1 0 89040 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__003__I
timestamp 1654395037
transform 1 0 91728 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__004__I
timestamp 1654395037
transform 1 0 91056 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__005__I
timestamp 1654395037
transform -1 0 78064 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__006__I
timestamp 1654395037
transform 1 0 91616 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__007__I
timestamp 1654395037
transform 1 0 101248 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__008__I
timestamp 1654395037
transform 1 0 110880 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__009__I
timestamp 1654395037
transform 1 0 118944 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__010__I
timestamp 1654395037
transform 1 0 123760 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__011__I
timestamp 1654395037
transform 1 0 127232 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__012__I
timestamp 1654395037
transform 1 0 130928 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__013__I
timestamp 1654395037
transform 1 0 137088 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__014__I
timestamp 1654395037
transform 1 0 147616 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__015__I
timestamp 1654395037
transform -1 0 152768 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__016__I
timestamp 1654395037
transform 1 0 167776 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__017__I
timestamp 1654395037
transform 1 0 179648 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__018__I
timestamp 1654395037
transform 1 0 183680 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__019__I
timestamp 1654395037
transform 1 0 191744 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__020__I
timestamp 1654395037
transform 1 0 197344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__021__I
timestamp 1654395037
transform 1 0 198016 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__022__I
timestamp 1654395037
transform -1 0 200480 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__023__I
timestamp 1654395037
transform 1 0 212240 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__024__I
timestamp 1654395037
transform 1 0 212016 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__025__I
timestamp 1654395037
transform 1 0 213136 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__026__I
timestamp 1654395037
transform 1 0 212352 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__027__I
timestamp 1654395037
transform 1 0 197680 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__028__I
timestamp 1654395037
transform 1 0 201264 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__029__I
timestamp 1654395037
transform 1 0 212128 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__030__I
timestamp 1654395037
transform 1 0 213584 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__031__I
timestamp 1654395037
transform 1 0 212576 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__032__I
timestamp 1654395037
transform 1 0 213024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__033__I
timestamp 1654395037
transform 1 0 213696 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__034__I
timestamp 1654395037
transform 1 0 213696 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__035__I
timestamp 1654395037
transform 1 0 215040 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__036__I
timestamp 1654395037
transform 1 0 215040 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__037__I
timestamp 1654395037
transform 1 0 214592 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__038__I
timestamp 1654395037
transform 1 0 215376 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__039__I
timestamp 1654395037
transform 1 0 60144 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__040__I
timestamp 1654395037
transform 1 0 57680 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__041__I
timestamp 1654395037
transform 1 0 58352 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__042__I
timestamp 1654395037
transform 1 0 50960 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__043__I
timestamp 1654395037
transform 1 0 58800 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__044__I
timestamp 1654395037
transform -1 0 67088 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__045__I
timestamp 1654395037
transform 1 0 68656 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__046__I
timestamp 1654395037
transform -1 0 67536 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__047__I
timestamp 1654395037
transform -1 0 67536 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__048__I
timestamp 1654395037
transform -1 0 67984 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__049__I
timestamp 1654395037
transform -1 0 68432 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__050__I
timestamp 1654395037
transform -1 0 67984 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__051__I
timestamp 1654395037
transform -1 0 68880 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__052__I
timestamp 1654395037
transform -1 0 71680 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__053__I
timestamp 1654395037
transform -1 0 72688 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__054__I
timestamp 1654395037
transform 1 0 76272 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__055__I
timestamp 1654395037
transform 1 0 74592 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__056__I
timestamp 1654395037
transform 1 0 76048 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__057__I
timestamp 1654395037
transform 1 0 77504 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__058__I
timestamp 1654395037
transform 1 0 83888 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__059__I
timestamp 1654395037
transform -1 0 84560 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__060__I
timestamp 1654395037
transform 1 0 91728 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__061__I
timestamp 1654395037
transform 1 0 79744 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__062__I
timestamp 1654395037
transform -1 0 85344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__063__I
timestamp 1654395037
transform 1 0 86464 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__064__I
timestamp 1654395037
transform 1 0 76720 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__065__I
timestamp 1654395037
transform 1 0 77728 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__066__I
timestamp 1654395037
transform -1 0 78512 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__067__I
timestamp 1654395037
transform 1 0 78624 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__068__I
timestamp 1654395037
transform 1 0 83104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__069__I
timestamp 1654395037
transform -1 0 80192 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__070__I
timestamp 1654395037
transform 1 0 84672 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__071__I
timestamp 1654395037
transform -1 0 86016 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__072__I
timestamp 1654395037
transform 1 0 83888 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__073__I
timestamp 1654395037
transform 1 0 78848 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__074__I
timestamp 1654395037
transform 1 0 78176 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__075__I
timestamp 1654395037
transform -1 0 78960 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__076__I
timestamp 1654395037
transform 1 0 83776 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__077__I
timestamp 1654395037
transform 1 0 84224 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__078__I
timestamp 1654395037
transform 1 0 87024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__079__I
timestamp 1654395037
transform -1 0 89152 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__080__I
timestamp 1654395037
transform 1 0 89712 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__081__I
timestamp 1654395037
transform 1 0 92176 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__082__I
timestamp 1654395037
transform 1 0 95312 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__083__I
timestamp 1654395037
transform 1 0 100016 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__084__I
timestamp 1654395037
transform -1 0 103040 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__085__I
timestamp 1654395037
transform 1 0 104272 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__086__I
timestamp 1654395037
transform 1 0 109200 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__087__I
timestamp 1654395037
transform -1 0 106960 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__088__I
timestamp 1654395037
transform 1 0 108304 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__089__I
timestamp 1654395037
transform -1 0 110880 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__090__I
timestamp 1654395037
transform -1 0 114800 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__091__I
timestamp 1654395037
transform -1 0 120624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__092__I
timestamp 1654395037
transform -1 0 128464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__093__I
timestamp 1654395037
transform 1 0 144928 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__094__I
timestamp 1654395037
transform 1 0 129584 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__095__I
timestamp 1654395037
transform 1 0 130816 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__096__I
timestamp 1654395037
transform 1 0 132048 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__097__I
timestamp 1654395037
transform 1 0 141680 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__098__I
timestamp 1654395037
transform 1 0 139216 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__099__I
timestamp 1654395037
transform 1 0 147504 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__100__I
timestamp 1654395037
transform 1 0 147952 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__101__I
timestamp 1654395037
transform 1 0 148400 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__102__I
timestamp 1654395037
transform 1 0 151424 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__103__I
timestamp 1654395037
transform 1 0 155344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__104__I
timestamp 1654395037
transform 1 0 161728 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__105__I
timestamp 1654395037
transform 1 0 175728 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__106__I
timestamp 1654395037
transform 1 0 192192 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__107__I
timestamp 1654395037
transform 1 0 195552 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__108__I
timestamp 1654395037
transform 1 0 196000 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__109__I
timestamp 1654395037
transform 1 0 198912 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__110__I
timestamp 1654395037
transform 1 0 202832 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__111__I
timestamp 1654395037
transform 1 0 203280 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__112__I
timestamp 1654395037
transform 1 0 199584 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__113__I
timestamp 1654395037
transform -1 0 203728 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__114__I
timestamp 1654395037
transform 1 0 203728 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__115__I
timestamp 1654395037
transform 1 0 211232 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__116__I
timestamp 1654395037
transform 1 0 212240 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__117__I
timestamp 1654395037
transform 1 0 214144 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__118__I
timestamp 1654395037
transform 1 0 213472 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__119__I
timestamp 1654395037
transform 1 0 215040 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__120__I
timestamp 1654395037
transform 1 0 215488 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__121__I
timestamp 1654395037
transform 1 0 214816 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__122__I
timestamp 1654395037
transform 1 0 213472 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__123__I
timestamp 1654395037
transform 1 0 215264 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__124__I
timestamp 1654395037
transform 1 0 215936 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__125__I
timestamp 1654395037
transform 1 0 216384 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__126__I
timestamp 1654395037
transform 1 0 214816 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__127__I
timestamp 1654395037
transform 1 0 215824 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__128__I
timestamp 1654395037
transform 1 0 194320 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__129__I
timestamp 1654395037
transform 1 0 192864 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__130__I
timestamp 1654395037
transform 1 0 193648 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__131__I
timestamp 1654395037
transform 1 0 194656 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__132__I
timestamp 1654395037
transform 1 0 192416 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__133__I
timestamp 1654395037
transform 1 0 193760 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__134__I
timestamp 1654395037
transform 1 0 194544 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__135__I
timestamp 1654395037
transform 1 0 196336 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__136__I
timestamp 1654395037
transform 1 0 196336 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__137__I
timestamp 1654395037
transform 1 0 198464 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__138__I
timestamp 1654395037
transform 1 0 200816 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__139__I
timestamp 1654395037
transform 1 0 200816 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__140__I
timestamp 1654395037
transform 1 0 199808 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__141__I
timestamp 1654395037
transform -1 0 35840 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__142__I
timestamp 1654395037
transform -1 0 38192 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__143__I
timestamp 1654395037
transform 1 0 40096 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__144__I
timestamp 1654395037
transform -1 0 41552 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__145__I
timestamp 1654395037
transform 1 0 43904 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__146__I
timestamp 1654395037
transform -1 0 45472 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__147__I
timestamp 1654395037
transform -1 0 46928 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__148__I
timestamp 1654395037
transform -1 0 48944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__149__I
timestamp 1654395037
transform 1 0 43232 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__150__I
timestamp 1654395037
transform 1 0 42336 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__151__I
timestamp 1654395037
transform 1 0 44352 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__152__I
timestamp 1654395037
transform -1 0 46592 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__153__I
timestamp 1654395037
transform 1 0 49280 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__154__I
timestamp 1654395037
transform 1 0 51520 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__155__I
timestamp 1654395037
transform -1 0 53648 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__156__I
timestamp 1654395037
transform 1 0 59472 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__157__I
timestamp 1654395037
transform 1 0 63504 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__158__I
timestamp 1654395037
transform -1 0 67984 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__159__I
timestamp 1654395037
transform -1 0 72128 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__160__I
timestamp 1654395037
transform -1 0 9072 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__161__I
timestamp 1654395037
transform 1 0 213920 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__162__I
timestamp 1654395037
transform 1 0 213136 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__163__I
timestamp 1654395037
transform 1 0 213584 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__164__I
timestamp 1654395037
transform 1 0 214592 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__165__I
timestamp 1654395037
transform 1 0 214368 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__166__I
timestamp 1654395037
transform 1 0 18480 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__167__I
timestamp 1654395037
transform 1 0 20608 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__168__I
timestamp 1654395037
transform -1 0 22624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__169__I
timestamp 1654395037
transform 1 0 26320 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__170__I
timestamp 1654395037
transform -1 0 27552 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__171__I
timestamp 1654395037
transform -1 0 30464 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__172__I
timestamp 1654395037
transform -1 0 32480 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__173__I
timestamp 1654395037
transform 1 0 34496 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__174__I
timestamp 1654395037
transform -1 0 37072 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__175__I
timestamp 1654395037
transform 1 0 39200 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__176__I
timestamp 1654395037
transform -1 0 40880 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__177__I
timestamp 1654395037
transform -1 0 44016 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__178__I
timestamp 1654395037
transform 1 0 44576 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__179__I
timestamp 1654395037
transform -1 0 47152 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__180__I
timestamp 1654395037
transform 1 0 49840 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__181__I
timestamp 1654395037
transform -1 0 44128 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__182__I
timestamp 1654395037
transform -1 0 42672 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__183__I
timestamp 1654395037
transform -1 0 43568 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__184__I
timestamp 1654395037
transform -1 0 46144 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__185__I
timestamp 1654395037
transform -1 0 48048 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__186__I
timestamp 1654395037
transform -1 0 50624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__187__I
timestamp 1654395037
transform -1 0 52864 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__188__I
timestamp 1654395037
transform -1 0 58128 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__189__I
timestamp 1654395037
transform 1 0 61936 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__190__I
timestamp 1654395037
transform -1 0 66640 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__191__I
timestamp 1654395037
transform 1 0 70560 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__192__I
timestamp 1654395037
transform 1 0 74816 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__193__I
timestamp 1654395037
transform 1 0 189728 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__194__I
timestamp 1654395037
transform 1 0 191408 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__195__I
timestamp 1654395037
transform 1 0 191072 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__196__I
timestamp 1654395037
transform 1 0 192640 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__197__I
timestamp 1654395037
transform -1 0 8960 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__198__I
timestamp 1654395037
transform -1 0 12656 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__199__I
timestamp 1654395037
transform 1 0 10304 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__200__I
timestamp 1654395037
transform 1 0 216720 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__201__I
timestamp 1654395037
transform 1 0 8288 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[0\]_EN
timestamp 1654395037
transform 1 0 18592 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[0\]_I
timestamp 1654395037
transform -1 0 19264 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[1\]_EN
timestamp 1654395037
transform 1 0 18704 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[1\]_I
timestamp 1654395037
transform 1 0 19152 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[2\]_EN
timestamp 1654395037
transform -1 0 17696 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[2\]_I
timestamp 1654395037
transform -1 0 18144 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[3\]_EN
timestamp 1654395037
transform 1 0 17472 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[3\]_I
timestamp 1654395037
transform -1 0 18144 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[4\]_EN
timestamp 1654395037
transform -1 0 13664 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[4\]_I
timestamp 1654395037
transform 1 0 13888 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[5\]_EN
timestamp 1654395037
transform -1 0 14112 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[5\]_I
timestamp 1654395037
transform 1 0 13328 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[6\]_EN
timestamp 1654395037
transform 1 0 9520 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[6\]_I
timestamp 1654395037
transform 1 0 8736 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[7\]_EN
timestamp 1654395037
transform -1 0 15680 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[7\]_I
timestamp 1654395037
transform -1 0 16128 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[8\]_EN
timestamp 1654395037
transform -1 0 24640 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[8\]_I
timestamp 1654395037
transform -1 0 25648 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[9\]_EN
timestamp 1654395037
transform -1 0 30240 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[9\]_I
timestamp 1654395037
transform -1 0 30688 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[10\]_EN
timestamp 1654395037
transform 1 0 35056 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[10\]_I
timestamp 1654395037
transform 1 0 35504 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[11\]_EN
timestamp 1654395037
transform -1 0 39872 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[11\]_I
timestamp 1654395037
transform 1 0 38976 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[12\]_EN
timestamp 1654395037
transform 1 0 43792 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[12\]_I
timestamp 1654395037
transform 1 0 44240 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[13\]_EN
timestamp 1654395037
transform 1 0 48608 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[13\]_I
timestamp 1654395037
transform 1 0 48160 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[14\]_I
timestamp 1654395037
transform -1 0 52304 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[15\]_I
timestamp 1654395037
transform 1 0 61712 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[16\]_I
timestamp 1654395037
transform -1 0 68656 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[17\]_I
timestamp 1654395037
transform 1 0 78512 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[18\]_I
timestamp 1654395037
transform 1 0 86128 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[19\]_I
timestamp 1654395037
transform -1 0 92512 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[20\]_I
timestamp 1654395037
transform -1 0 97776 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[21\]_I
timestamp 1654395037
transform 1 0 101584 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[22\]_EN
timestamp 1654395037
transform 1 0 25424 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[22\]_I
timestamp 1654395037
transform 1 0 25872 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[23\]_EN
timestamp 1654395037
transform -1 0 57456 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[23\]_I
timestamp 1654395037
transform 1 0 58800 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[24\]_EN
timestamp 1654395037
transform -1 0 57456 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[24\]_I
timestamp 1654395037
transform 1 0 56560 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[25\]_EN
timestamp 1654395037
transform -1 0 57120 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[25\]_I
timestamp 1654395037
transform 1 0 57344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[26\]_EN
timestamp 1654395037
transform -1 0 59472 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[26\]_I
timestamp 1654395037
transform 1 0 58576 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[27\]_EN
timestamp 1654395037
transform -1 0 65408 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[27\]_I
timestamp 1654395037
transform 1 0 60480 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[28\]_I
timestamp 1654395037
transform 1 0 72352 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[29\]_EN
timestamp 1654395037
transform -1 0 73360 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[29\]_I
timestamp 1654395037
transform -1 0 68208 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[30\]_EN
timestamp 1654395037
transform -1 0 52752 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[30\]_I
timestamp 1654395037
transform 1 0 52528 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[31\]_I
timestamp 1654395037
transform 1 0 78288 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[32\]_I
timestamp 1654395037
transform 1 0 96208 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[33\]_I
timestamp 1654395037
transform -1 0 107632 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[34\]_I
timestamp 1654395037
transform 1 0 116144 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[35\]_I
timestamp 1654395037
transform -1 0 121744 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[36\]_I
timestamp 1654395037
transform -1 0 124880 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[37\]_I
timestamp 1654395037
transform -1 0 128352 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[38\]_I
timestamp 1654395037
transform 1 0 135072 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[39\]_I
timestamp 1654395037
transform 1 0 143696 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[40\]_I
timestamp 1654395037
transform 1 0 149968 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[41\]_I
timestamp 1654395037
transform -1 0 153664 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[42\]_I
timestamp 1654395037
transform 1 0 161056 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[43\]_I
timestamp 1654395037
transform 1 0 169120 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[44\]_I
timestamp 1654395037
transform 1 0 173264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[45\]_I
timestamp 1654395037
transform 1 0 177184 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[46\]_I
timestamp 1654395037
transform 1 0 181104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[47\]_I
timestamp 1654395037
transform 1 0 192416 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[48\]_I
timestamp 1654395037
transform 1 0 192416 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[49\]_I
timestamp 1654395037
transform 1 0 193312 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[50\]_I
timestamp 1654395037
transform 1 0 195104 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[51\]_I
timestamp 1654395037
transform 1 0 194768 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[52\]_I
timestamp 1654395037
transform 1 0 192864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[53\]_I
timestamp 1654395037
transform 1 0 191968 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[54\]_I
timestamp 1654395037
transform 1 0 195216 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[55\]_I
timestamp 1654395037
transform 1 0 197232 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[56\]_I
timestamp 1654395037
transform 1 0 212240 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[57\]_I
timestamp 1654395037
transform 1 0 214032 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[58\]_I
timestamp 1654395037
transform 1 0 214032 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[59\]_I
timestamp 1654395037
transform 1 0 213248 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[60\]_I
timestamp 1654395037
transform 1 0 214480 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[61\]_I
timestamp 1654395037
transform 1 0 214592 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[62\]_I
timestamp 1654395037
transform 1 0 214480 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_la_buf\[63\]_I
timestamp 1654395037
transform 1 0 213920 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_irq_gates\[0\]_A1
timestamp 1654395037
transform -1 0 215152 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_irq_gates\[0\]_A2
timestamp 1654395037
transform 1 0 214368 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_irq_gates\[1\]_A1
timestamp 1654395037
transform 1 0 215264 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_irq_gates\[1\]_A2
timestamp 1654395037
transform 1 0 214928 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_irq_gates\[2\]_A1
timestamp 1654395037
transform -1 0 215600 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_irq_gates\[2\]_A2
timestamp 1654395037
transform -1 0 217392 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_buffers\[0\]_I
timestamp 1654395037
transform -1 0 21840 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_buffers\[1\]_I
timestamp 1654395037
transform -1 0 25312 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_buffers\[2\]_I
timestamp 1654395037
transform -1 0 22400 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_buffers\[3\]_I
timestamp 1654395037
transform 1 0 25424 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_buffers\[4\]_I
timestamp 1654395037
transform -1 0 25088 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_buffers\[5\]_I
timestamp 1654395037
transform -1 0 21392 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_buffers\[6\]_I
timestamp 1654395037
transform -1 0 25312 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_buffers\[7\]_I
timestamp 1654395037
transform -1 0 28448 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_buffers\[8\]_I
timestamp 1654395037
transform -1 0 29232 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_buffers\[9\]_I
timestamp 1654395037
transform 1 0 30576 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_buffers\[10\]_I
timestamp 1654395037
transform 1 0 33376 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_buffers\[11\]_I
timestamp 1654395037
transform -1 0 35728 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_buffers\[12\]_I
timestamp 1654395037
transform 1 0 37520 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_buffers\[13\]_I
timestamp 1654395037
transform -1 0 10752 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_buffers\[14\]_I
timestamp 1654395037
transform -1 0 10640 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_buffers\[15\]_I
timestamp 1654395037
transform -1 0 13664 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_buffers\[16\]_I
timestamp 1654395037
transform -1 0 9632 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_buffers\[17\]_I
timestamp 1654395037
transform 1 0 9520 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_buffers\[18\]_I
timestamp 1654395037
transform -1 0 16464 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_buffers\[19\]_I
timestamp 1654395037
transform -1 0 21616 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_buffers\[20\]_I
timestamp 1654395037
transform 1 0 28672 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_buffers\[21\]_I
timestamp 1654395037
transform 1 0 33824 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_buffers\[22\]_I
timestamp 1654395037
transform -1 0 39312 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_buffers\[23\]_I
timestamp 1654395037
transform -1 0 43792 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_buffers\[24\]_I
timestamp 1654395037
transform 1 0 47040 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_buffers\[25\]_I
timestamp 1654395037
transform -1 0 48832 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_buffers\[26\]_I
timestamp 1654395037
transform 1 0 51520 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_buffers\[27\]_I
timestamp 1654395037
transform -1 0 52752 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_buffers\[28\]_I
timestamp 1654395037
transform -1 0 56672 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_buffers\[29\]_I
timestamp 1654395037
transform -1 0 60592 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_buffers\[30\]_I
timestamp 1654395037
transform -1 0 64512 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_buffers\[31\]_I
timestamp 1654395037
transform 1 0 66864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_buffers\[32\]_I
timestamp 1654395037
transform -1 0 68656 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_buffers\[33\]_I
timestamp 1654395037
transform -1 0 75264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_buffers\[34\]_I
timestamp 1654395037
transform -1 0 78176 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_buffers\[35\]_I
timestamp 1654395037
transform -1 0 80192 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_buffers\[36\]_I
timestamp 1654395037
transform -1 0 84560 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_buffers\[37\]_I
timestamp 1654395037
transform -1 0 85008 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_buffers\[38\]_I
timestamp 1654395037
transform 1 0 85792 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_buffers\[39\]_I
timestamp 1654395037
transform -1 0 88032 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_buffers\[40\]_I
timestamp 1654395037
transform -1 0 91280 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_buffers\[41\]_I
timestamp 1654395037
transform -1 0 94864 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_buffers\[42\]_I
timestamp 1654395037
transform -1 0 98112 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_buffers\[43\]_I
timestamp 1654395037
transform -1 0 101808 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_buffers\[44\]_I
timestamp 1654395037
transform -1 0 103712 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_buffers\[45\]_I
timestamp 1654395037
transform -1 0 107632 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_buffers\[46\]_I
timestamp 1654395037
transform -1 0 111552 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_buffers\[47\]_I
timestamp 1654395037
transform -1 0 114240 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_buffers\[48\]_I
timestamp 1654395037
transform -1 0 117712 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_buffers\[49\]_I
timestamp 1654395037
transform 1 0 119728 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_buffers\[50\]_I
timestamp 1654395037
transform 1 0 122416 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_buffers\[51\]_I
timestamp 1654395037
transform -1 0 125552 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_buffers\[52\]_I
timestamp 1654395037
transform -1 0 129472 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_buffers\[53\]_I
timestamp 1654395037
transform 1 0 131040 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_buffers\[54\]_I
timestamp 1654395037
transform -1 0 133504 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_buffers\[55\]_I
timestamp 1654395037
transform -1 0 132608 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_buffers\[56\]_I
timestamp 1654395037
transform -1 0 142240 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_buffers\[57\]_I
timestamp 1654395037
transform -1 0 142912 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_buffers\[58\]_I
timestamp 1654395037
transform -1 0 147728 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_buffers\[59\]_I
timestamp 1654395037
transform -1 0 151872 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_buffers\[60\]_I
timestamp 1654395037
transform -1 0 160832 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_buffers\[61\]_I
timestamp 1654395037
transform -1 0 185248 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_buffers\[62\]_I
timestamp 1654395037
transform 1 0 192864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[0\]_A1
timestamp 1654395037
transform -1 0 47488 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[0\]_A2
timestamp 1654395037
transform 1 0 49616 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[1\]_A1
timestamp 1654395037
transform -1 0 51856 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[1\]_A2
timestamp 1654395037
transform 1 0 52080 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[2\]_A1
timestamp 1654395037
transform -1 0 53648 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[2\]_A2
timestamp 1654395037
transform -1 0 56672 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[3\]_A1
timestamp 1654395037
transform -1 0 60032 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[3\]_A2
timestamp 1654395037
transform 1 0 59360 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[4\]_A1
timestamp 1654395037
transform 1 0 63840 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[4\]_A2
timestamp 1654395037
transform 1 0 63392 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[5\]_A1
timestamp 1654395037
transform -1 0 66640 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[5\]_A2
timestamp 1654395037
transform 1 0 67200 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[6\]_A1
timestamp 1654395037
transform 1 0 70896 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[6\]_A2
timestamp 1654395037
transform -1 0 71344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[7\]_A1
timestamp 1654395037
transform 1 0 75600 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[7\]_A2
timestamp 1654395037
transform 1 0 75152 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[8\]_A1
timestamp 1654395037
transform -1 0 78064 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[8\]_A2
timestamp 1654395037
transform 1 0 78288 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[9\]_A1
timestamp 1654395037
transform -1 0 84112 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[9\]_A2
timestamp 1654395037
transform 1 0 83440 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[10\]_A1
timestamp 1654395037
transform -1 0 85904 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[10\]_A2
timestamp 1654395037
transform 1 0 85344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[11\]_A1
timestamp 1654395037
transform 1 0 87696 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[11\]_A2
timestamp 1654395037
transform 1 0 87920 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[12\]_A1
timestamp 1654395037
transform -1 0 91504 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[12\]_A2
timestamp 1654395037
transform 1 0 91504 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[13\]_A1
timestamp 1654395037
transform 1 0 94864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[13\]_A2
timestamp 1654395037
transform -1 0 96096 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[14\]_A1
timestamp 1654395037
transform -1 0 98448 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[14\]_A2
timestamp 1654395037
transform -1 0 98000 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[15\]_A1
timestamp 1654395037
transform 1 0 98896 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[15\]_A2
timestamp 1654395037
transform -1 0 99792 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[16\]_A1
timestamp 1654395037
transform -1 0 101360 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[16\]_A2
timestamp 1654395037
transform -1 0 101136 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[17\]_A1
timestamp 1654395037
transform -1 0 104160 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[17\]_A2
timestamp 1654395037
transform -1 0 103712 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[18\]_A1
timestamp 1654395037
transform 1 0 104496 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[18\]_A2
timestamp 1654395037
transform 1 0 104944 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[19\]_A1
timestamp 1654395037
transform 1 0 107856 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[19\]_A2
timestamp 1654395037
transform 1 0 107632 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[20\]_A1
timestamp 1654395037
transform -1 0 111552 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[20\]_A2
timestamp 1654395037
transform 1 0 110880 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[21\]_A1
timestamp 1654395037
transform -1 0 113344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[21\]_A2
timestamp 1654395037
transform -1 0 113792 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[22\]_A1
timestamp 1654395037
transform 1 0 115920 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[22\]_A2
timestamp 1654395037
transform 1 0 115920 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[23\]_A1
timestamp 1654395037
transform -1 0 118496 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[23\]_A2
timestamp 1654395037
transform 1 0 118720 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[24\]_A1
timestamp 1654395037
transform 1 0 120848 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[24\]_A2
timestamp 1654395037
transform 1 0 121296 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[25\]_A1
timestamp 1654395037
transform -1 0 123200 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[25\]_A2
timestamp 1654395037
transform -1 0 123648 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[26\]_A1
timestamp 1654395037
transform -1 0 126784 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[26\]_A2
timestamp 1654395037
transform 1 0 127008 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[27\]_A1
timestamp 1654395037
transform -1 0 128352 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[27\]_A2
timestamp 1654395037
transform -1 0 129136 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[28\]_A1
timestamp 1654395037
transform -1 0 131488 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[28\]_A2
timestamp 1654395037
transform -1 0 131936 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[29\]_A1
timestamp 1654395037
transform -1 0 134400 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[29\]_A2
timestamp 1654395037
transform -1 0 133952 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[30\]_A1
timestamp 1654395037
transform -1 0 138208 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[30\]_A2
timestamp 1654395037
transform -1 0 131712 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[31\]_A1
timestamp 1654395037
transform -1 0 143472 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[31\]_A2
timestamp 1654395037
transform -1 0 132160 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[32\]_A1
timestamp 1654395037
transform -1 0 143360 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[32\]_A2
timestamp 1654395037
transform 1 0 141568 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[33\]_A1
timestamp 1654395037
transform -1 0 145376 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[33\]_A2
timestamp 1654395037
transform 1 0 141120 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[34\]_A1
timestamp 1654395037
transform -1 0 146832 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[34\]_A2
timestamp 1654395037
transform 1 0 143584 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[35\]_A1
timestamp 1654395037
transform -1 0 148176 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[35\]_A2
timestamp 1654395037
transform 1 0 147168 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[36\]_A1
timestamp 1654395037
transform 1 0 147056 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[36\]_A2
timestamp 1654395037
transform 1 0 146720 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[37\]_A1
timestamp 1654395037
transform 1 0 148736 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[37\]_A2
timestamp 1654395037
transform 1 0 147056 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[38\]_A1
timestamp 1654395037
transform -1 0 148624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[38\]_A2
timestamp 1654395037
transform 1 0 147952 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[39\]_A1
timestamp 1654395037
transform -1 0 150864 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[39\]_A2
timestamp 1654395037
transform 1 0 149184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[40\]_A1
timestamp 1654395037
transform -1 0 149520 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[40\]_A2
timestamp 1654395037
transform 1 0 148848 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[41\]_A1
timestamp 1654395037
transform 1 0 151760 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[41\]_A2
timestamp 1654395037
transform 1 0 149744 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[42\]_A1
timestamp 1654395037
transform -1 0 153776 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[42\]_A2
timestamp 1654395037
transform 1 0 151088 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[43\]_A1
timestamp 1654395037
transform 1 0 154672 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[43\]_A2
timestamp 1654395037
transform 1 0 153104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[44\]_A1
timestamp 1654395037
transform 1 0 160608 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[44\]_A2
timestamp 1654395037
transform 1 0 154448 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[45\]_A1
timestamp 1654395037
transform -1 0 163408 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[45\]_A2
timestamp 1654395037
transform 1 0 155344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[46\]_A1
timestamp 1654395037
transform -1 0 165200 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[46\]_A2
timestamp 1654395037
transform 1 0 163632 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[47\]_A1
timestamp 1654395037
transform -1 0 161504 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[47\]_A2
timestamp 1654395037
transform 1 0 159152 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[48\]_A1
timestamp 1654395037
transform 1 0 157136 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[48\]_A2
timestamp 1654395037
transform 1 0 156688 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[49\]_A1
timestamp 1654395037
transform 1 0 190624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[49\]_A2
timestamp 1654395037
transform 1 0 191408 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[50\]_A1
timestamp 1654395037
transform 1 0 195664 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[50\]_A2
timestamp 1654395037
transform 1 0 194208 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[51\]_A1
timestamp 1654395037
transform 1 0 196448 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[51\]_A2
timestamp 1654395037
transform 1 0 198464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[52\]_A1
timestamp 1654395037
transform 1 0 196784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[52\]_A2
timestamp 1654395037
transform 1 0 195552 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[53\]_A1
timestamp 1654395037
transform 1 0 199360 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[53\]_A2
timestamp 1654395037
transform 1 0 198464 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[54\]_A1
timestamp 1654395037
transform 1 0 198688 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[54\]_A2
timestamp 1654395037
transform 1 0 195440 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[55\]_A1
timestamp 1654395037
transform 1 0 200256 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[55\]_A2
timestamp 1654395037
transform 1 0 198912 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[56\]_A1
timestamp 1654395037
transform -1 0 200592 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[56\]_A2
timestamp 1654395037
transform 1 0 199136 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[57\]_A1
timestamp 1654395037
transform -1 0 201488 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[57\]_A2
timestamp 1654395037
transform 1 0 198128 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[58\]_A1
timestamp 1654395037
transform 1 0 203056 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[58\]_A2
timestamp 1654395037
transform 1 0 201712 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[59\]_A1
timestamp 1654395037
transform 1 0 204288 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[59\]_A2
timestamp 1654395037
transform 1 0 200704 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[60\]_A1
timestamp 1654395037
transform 1 0 207536 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[60\]_A2
timestamp 1654395037
transform 1 0 202608 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[61\]_A1
timestamp 1654395037
transform 1 0 212688 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[61\]_A2
timestamp 1654395037
transform 1 0 203616 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[62\]_A1
timestamp 1654395037
transform 1 0 211680 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[62\]_A2
timestamp 1654395037
transform 1 0 202608 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[63\]_A1
timestamp 1654395037
transform 1 0 212800 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_to_mprj_in_gates\[63\]_A2
timestamp 1654395037
transform 1 0 211568 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_ack_gate_A1
timestamp 1654395037
transform 1 0 216272 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_ack_gate_A2
timestamp 1654395037
transform 1 0 216272 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_buffers\[0\]_I
timestamp 1654395037
transform 1 0 164528 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_buffers\[1\]_I
timestamp 1654395037
transform 1 0 173376 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_buffers\[2\]_I
timestamp 1654395037
transform 1 0 165424 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_buffers\[3\]_I
timestamp 1654395037
transform 1 0 164976 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_buffers\[4\]_I
timestamp 1654395037
transform 1 0 183680 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_buffers\[5\]_I
timestamp 1654395037
transform 1 0 190176 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_buffers\[6\]_I
timestamp 1654395037
transform 1 0 191520 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_buffers\[7\]_I
timestamp 1654395037
transform 1 0 180432 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_buffers\[8\]_I
timestamp 1654395037
transform 1 0 191296 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_buffers\[9\]_I
timestamp 1654395037
transform 1 0 194096 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_buffers\[10\]_I
timestamp 1654395037
transform 1 0 193536 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_buffers\[11\]_I
timestamp 1654395037
transform 1 0 194992 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_buffers\[12\]_I
timestamp 1654395037
transform 1 0 193088 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_buffers\[13\]_I
timestamp 1654395037
transform 1 0 195888 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_buffers\[14\]_I
timestamp 1654395037
transform 1 0 196784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_buffers\[15\]_I
timestamp 1654395037
transform 1 0 197792 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_buffers\[16\]_I
timestamp 1654395037
transform 1 0 199360 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_buffers\[24\]_I
timestamp 1654395037
transform 1 0 212464 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_buffers\[26\]_I
timestamp 1654395037
transform 1 0 213248 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_buffers\[28\]_I
timestamp 1654395037
transform 1 0 214144 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_buffers\[29\]_I
timestamp 1654395037
transform 1 0 214144 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_buffers\[31\]_I
timestamp 1654395037
transform 1 0 215488 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_gates\[0\]_A1
timestamp 1654395037
transform -1 0 131712 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_gates\[0\]_A2
timestamp 1654395037
transform 1 0 133952 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_gates\[1\]_A1
timestamp 1654395037
transform -1 0 131488 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_gates\[1\]_A2
timestamp 1654395037
transform -1 0 134176 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_gates\[2\]_A1
timestamp 1654395037
transform 1 0 135744 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_gates\[2\]_A2
timestamp 1654395037
transform 1 0 135520 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_gates\[3\]_A1
timestamp 1654395037
transform 1 0 135184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_gates\[3\]_A2
timestamp 1654395037
transform 1 0 135968 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_gates\[4\]_A1
timestamp 1654395037
transform 1 0 137760 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_gates\[4\]_A2
timestamp 1654395037
transform 1 0 138768 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_gates\[5\]_A1
timestamp 1654395037
transform 1 0 141680 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_gates\[5\]_A2
timestamp 1654395037
transform 1 0 139664 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_gates\[6\]_A1
timestamp 1654395037
transform 1 0 137536 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_gates\[6\]_A2
timestamp 1654395037
transform 1 0 144704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_gates\[7\]_A1
timestamp 1654395037
transform 1 0 142800 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_gates\[7\]_A2
timestamp 1654395037
transform -1 0 145600 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_gates\[8\]_A1
timestamp 1654395037
transform 1 0 144480 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_gates\[8\]_A2
timestamp 1654395037
transform -1 0 146048 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_gates\[9\]_A1
timestamp 1654395037
transform 1 0 146944 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_gates\[9\]_A2
timestamp 1654395037
transform 1 0 147392 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_gates\[10\]_A1
timestamp 1654395037
transform 1 0 148848 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_gates\[10\]_A2
timestamp 1654395037
transform 1 0 150640 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_gates\[11\]_A1
timestamp 1654395037
transform 1 0 151088 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_gates\[11\]_A2
timestamp 1654395037
transform 1 0 151312 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_gates\[12\]_A1
timestamp 1654395037
transform 1 0 153552 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_gates\[12\]_A2
timestamp 1654395037
transform 1 0 154896 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_gates\[13\]_A1
timestamp 1654395037
transform 1 0 157584 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_gates\[13\]_A2
timestamp 1654395037
transform 1 0 161504 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_gates\[14\]_A1
timestamp 1654395037
transform 1 0 164528 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_gates\[14\]_A2
timestamp 1654395037
transform 1 0 169456 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_gates\[15\]_A1
timestamp 1654395037
transform 1 0 168672 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_gates\[15\]_A2
timestamp 1654395037
transform -1 0 174272 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_gates\[16\]_A1
timestamp 1654395037
transform 1 0 188720 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_gates\[16\]_A2
timestamp 1654395037
transform -1 0 192864 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_gates\[17\]_A1
timestamp 1654395037
transform 1 0 147504 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_gates\[17\]_A2
timestamp 1654395037
transform -1 0 149520 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_gates\[18\]_A1
timestamp 1654395037
transform 1 0 149744 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_gates\[18\]_A2
timestamp 1654395037
transform 1 0 150416 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_gates\[19\]_A1
timestamp 1654395037
transform -1 0 151088 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_gates\[19\]_A2
timestamp 1654395037
transform -1 0 152320 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_gates\[20\]_A1
timestamp 1654395037
transform 1 0 152992 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_gates\[20\]_A2
timestamp 1654395037
transform 1 0 156576 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_gates\[21\]_A1
timestamp 1654395037
transform -1 0 155344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_gates\[21\]_A2
timestamp 1654395037
transform 1 0 159600 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_gates\[22\]_A1
timestamp 1654395037
transform 1 0 161280 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_gates\[22\]_A2
timestamp 1654395037
transform 1 0 166432 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_gates\[23\]_A1
timestamp 1654395037
transform 1 0 164304 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_gates\[23\]_A2
timestamp 1654395037
transform 1 0 166880 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_gates\[24\]_A1
timestamp 1654395037
transform 1 0 196896 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_gates\[24\]_A2
timestamp 1654395037
transform -1 0 200032 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_gates\[25\]_A1
timestamp 1654395037
transform 1 0 198240 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_gates\[25\]_A2
timestamp 1654395037
transform 1 0 200368 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_gates\[26\]_A1
timestamp 1654395037
transform 1 0 200816 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_gates\[26\]_A2
timestamp 1654395037
transform 1 0 201712 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_gates\[27\]_A1
timestamp 1654395037
transform 1 0 200704 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_gates\[27\]_A2
timestamp 1654395037
transform 1 0 200368 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_gates\[28\]_A1
timestamp 1654395037
transform 1 0 202160 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_gates\[28\]_A2
timestamp 1654395037
transform 1 0 203056 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_gates\[29\]_A1
timestamp 1654395037
transform 1 0 202160 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_gates\[29\]_A2
timestamp 1654395037
transform 1 0 203504 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_gates\[30\]_A1
timestamp 1654395037
transform 1 0 202384 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_gates\[30\]_A2
timestamp 1654395037
transform -1 0 203952 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_gates\[31\]_A1
timestamp 1654395037
transform 1 0 211232 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_user_wb_dat_gates\[31\]_A2
timestamp 1654395037
transform 1 0 212688 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2 pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34 pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 5152 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37 pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 5488 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45 pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 6384 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49
timestamp 1654395037
transform 1 0 6832 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_68 pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 8960 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74
timestamp 1654395037
transform 1 0 9632 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_78
timestamp 1654395037
transform 1 0 10080 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80
timestamp 1654395037
transform 1 0 10304 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_83
timestamp 1654395037
transform 1 0 10640 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_103
timestamp 1654395037
transform 1 0 12880 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_109
timestamp 1654395037
transform 1 0 13552 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_131
timestamp 1654395037
transform 1 0 16016 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_135
timestamp 1654395037
transform 1 0 16464 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_139
timestamp 1654395037
transform 1 0 16912 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_142
timestamp 1654395037
transform 1 0 17248 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_150
timestamp 1654395037
transform 1 0 18144 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_154
timestamp 1654395037
transform 1 0 18592 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_173
timestamp 1654395037
transform 1 0 20720 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_179
timestamp 1654395037
transform 1 0 21392 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_183
timestamp 1654395037
transform 1 0 21840 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_185
timestamp 1654395037
transform 1 0 22064 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_188
timestamp 1654395037
transform 1 0 22400 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_208
timestamp 1654395037
transform 1 0 24640 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_214
timestamp 1654395037
transform 1 0 25312 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_222
timestamp 1654395037
transform 1 0 26208 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_224
timestamp 1654395037
transform 1 0 26432 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_243
timestamp 1654395037
transform 1 0 28560 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_249
timestamp 1654395037
transform 1 0 29232 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_257
timestamp 1654395037
transform 1 0 30128 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_259
timestamp 1654395037
transform 1 0 30352 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_278
timestamp 1654395037
transform 1 0 32480 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_282
timestamp 1654395037
transform 1 0 32928 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_284
timestamp 1654395037
transform 1 0 33152 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_303
timestamp 1654395037
transform 1 0 35280 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_307
timestamp 1654395037
transform 1 0 35728 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_335
timestamp 1654395037
transform 1 0 38864 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_339
timestamp 1654395037
transform 1 0 39312 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_347
timestamp 1654395037
transform 1 0 40208 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_349
timestamp 1654395037
transform 1 0 40432 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_352
timestamp 1654395037
transform 1 0 40768 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_356
timestamp 1654395037
transform 1 0 41216 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_375
timestamp 1654395037
transform 1 0 43344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_379
timestamp 1654395037
transform 1 0 43792 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_383
timestamp 1654395037
transform 1 0 44240 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_387
timestamp 1654395037
transform 1 0 44688 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_395
timestamp 1654395037
transform 1 0 45584 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_399
timestamp 1654395037
transform 1 0 46032 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_418
timestamp 1654395037
transform 1 0 48160 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_424
timestamp 1654395037
transform 1 0 48832 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_428
timestamp 1654395037
transform 1 0 49280 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_430
timestamp 1654395037
transform 1 0 49504 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_433
timestamp 1654395037
transform 1 0 49840 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_453
timestamp 1654395037
transform 1 0 52080 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_459
timestamp 1654395037
transform 1 0 52752 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_467
timestamp 1654395037
transform 1 0 53648 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_469
timestamp 1654395037
transform 1 0 53872 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_488
timestamp 1654395037
transform 1 0 56000 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_494
timestamp 1654395037
transform 1 0 56672 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_498
timestamp 1654395037
transform 1 0 57120 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_501
timestamp 1654395037
transform 1 0 57456 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_523
timestamp 1654395037
transform 1 0 59920 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_529
timestamp 1654395037
transform 1 0 60592 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_537
timestamp 1654395037
transform 1 0 61488 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_539
timestamp 1654395037
transform 1 0 61712 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_558
timestamp 1654395037
transform 1 0 63840 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_564
timestamp 1654395037
transform 1 0 64512 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_572
timestamp 1654395037
transform 1 0 65408 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_592
timestamp 1654395037
transform 1 0 67648 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_594
timestamp 1654395037
transform 1 0 67872 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_597
timestamp 1654395037
transform 1 0 68208 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_601
timestamp 1654395037
transform 1 0 68656 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_621
timestamp 1654395037
transform 1 0 70896 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_625
timestamp 1654395037
transform 1 0 71344 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_628
timestamp 1654395037
transform 1 0 71680 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_650
timestamp 1654395037
transform 1 0 74144 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_656
timestamp 1654395037
transform 1 0 74816 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_660
timestamp 1654395037
transform 1 0 75264 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_664
timestamp 1654395037
transform 1 0 75712 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_667
timestamp 1654395037
transform 1 0 76048 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_675
timestamp 1654395037
transform 1 0 76944 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_679
timestamp 1654395037
transform 1 0 77392 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_698
timestamp 1654395037
transform 1 0 79520 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_704
timestamp 1654395037
transform 1 0 80192 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_712
timestamp 1654395037
transform 1 0 81088 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_714
timestamp 1654395037
transform 1 0 81312 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_733
timestamp 1654395037
transform 1 0 83440 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_739
timestamp 1654395037
transform 1 0 84112 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_743
timestamp 1654395037
transform 1 0 84560 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_747
timestamp 1654395037
transform 1 0 85008 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_749
timestamp 1654395037
transform 1 0 85232 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_768
timestamp 1654395037
transform 1 0 87360 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_774
timestamp 1654395037
transform 1 0 88032 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_778
timestamp 1654395037
transform 1 0 88480 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_780
timestamp 1654395037
transform 1 0 88704 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_799
timestamp 1654395037
transform 1 0 90832 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_803
timestamp 1654395037
transform 1 0 91280 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_807
timestamp 1654395037
transform 1 0 91728 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_811
timestamp 1654395037
transform 1 0 92176 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_831
timestamp 1654395037
transform 1 0 94416 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_835
timestamp 1654395037
transform 1 0 94864 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_839
timestamp 1654395037
transform 1 0 95312 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_860
timestamp 1654395037
transform 1 0 97664 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_864
timestamp 1654395037
transform 1 0 98112 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_872
timestamp 1654395037
transform 1 0 99008 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_874
timestamp 1654395037
transform 1 0 99232 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_877
timestamp 1654395037
transform 1 0 99568 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_885
timestamp 1654395037
transform 1 0 100464 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_889
timestamp 1654395037
transform 1 0 100912 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_908
timestamp 1654395037
transform 1 0 103040 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_914
timestamp 1654395037
transform 1 0 103712 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_922
timestamp 1654395037
transform 1 0 104608 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_924
timestamp 1654395037
transform 1 0 104832 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_943
timestamp 1654395037
transform 1 0 106960 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_949
timestamp 1654395037
transform 1 0 107632 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_975
timestamp 1654395037
transform 1 0 110544 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_979
timestamp 1654395037
transform 1 0 110992 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_984
timestamp 1654395037
transform 1 0 111552 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1004
timestamp 1654395037
transform 1 0 113792 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1008
timestamp 1654395037
transform 1 0 114240 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1012
timestamp 1654395037
transform 1 0 114688 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1014
timestamp 1654395037
transform 1 0 114912 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1035
timestamp 1654395037
transform 1 0 117264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1039
timestamp 1654395037
transform 1 0 117712 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1047
timestamp 1654395037
transform 1 0 118608 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1049
timestamp 1654395037
transform 1 0 118832 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1052
timestamp 1654395037
transform 1 0 119168 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1060
timestamp 1654395037
transform 1 0 120064 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1062
timestamp 1654395037
transform 1 0 120288 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1081
timestamp 1654395037
transform 1 0 122416 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1105
timestamp 1654395037
transform 1 0 125104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1109
timestamp 1654395037
transform 1 0 125552 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1117
timestamp 1654395037
transform 1 0 126448 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1119
timestamp 1654395037
transform 1 0 126672 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1140
timestamp 1654395037
transform 1 0 129024 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1144
timestamp 1654395037
transform 1 0 129472 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1152
timestamp 1654395037
transform 1 0 130368 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1154
timestamp 1654395037
transform 1 0 130592 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1157
timestamp 1654395037
transform 1 0 130928 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1176
timestamp 1654395037
transform 1 0 133056 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1180
timestamp 1654395037
transform 1 0 133504 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1184
timestamp 1654395037
transform 1 0 133952 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1188
timestamp 1654395037
transform 1 0 134400 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1210
timestamp 1654395037
transform 1 0 136864 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1214
timestamp 1654395037
transform 1 0 137312 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1218
timestamp 1654395037
transform 1 0 137760 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1222
timestamp 1654395037
transform 1 0 138208 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1224
timestamp 1654395037
transform 1 0 138432 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1227
timestamp 1654395037
transform 1 0 138768 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1246
timestamp 1654395037
transform 1 0 140896 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1250
timestamp 1654395037
transform 1 0 141344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1254
timestamp 1654395037
transform 1 0 141792 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1258
timestamp 1654395037
transform 1 0 142240 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1264
timestamp 1654395037
transform 1 0 142912 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1268
timestamp 1654395037
transform 1 0 143360 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1272
timestamp 1654395037
transform 1 0 143808 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1274
timestamp 1654395037
transform 1 0 144032 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1293
timestamp 1654395037
transform 1 0 146160 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1299
timestamp 1654395037
transform 1 0 146832 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1303
timestamp 1654395037
transform 1 0 147280 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1307
timestamp 1654395037
transform 1 0 147728 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1311
timestamp 1654395037
transform 1 0 148176 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1315
timestamp 1654395037
transform 1 0 148624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1319
timestamp 1654395037
transform 1 0 149072 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1323
timestamp 1654395037
transform 1 0 149520 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1327
timestamp 1654395037
transform 1 0 149968 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1329
timestamp 1654395037
transform 1 0 150192 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1332
timestamp 1654395037
transform 1 0 150528 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1334
timestamp 1654395037
transform 1 0 150752 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1353
timestamp 1654395037
transform 1 0 152880 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1357
timestamp 1654395037
transform 1 0 153328 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1361
timestamp 1654395037
transform 1 0 153776 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1369
timestamp 1654395037
transform 1 0 154672 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1373
timestamp 1654395037
transform 1 0 155120 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1377
timestamp 1654395037
transform 1 0 155568 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1379
timestamp 1654395037
transform 1 0 155792 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1398
timestamp 1654395037
transform 1 0 157920 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1420
timestamp 1654395037
transform 1 0 160384 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1424
timestamp 1654395037
transform 1 0 160832 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1428
timestamp 1654395037
transform 1 0 161280 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1432
timestamp 1654395037
transform 1 0 161728 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1434
timestamp 1654395037
transform 1 0 161952 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1455
timestamp 1654395037
transform 1 0 164304 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1459
timestamp 1654395037
transform 1 0 164752 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1463
timestamp 1654395037
transform 1 0 165200 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1467
timestamp 1654395037
transform 1 0 165648 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1469
timestamp 1654395037
transform 1 0 165872 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1490
timestamp 1654395037
transform 1 0 168224 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1492
timestamp 1654395037
transform 1 0 168448 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1499
timestamp 1654395037
transform 1 0 169232 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1503
timestamp 1654395037
transform 1 0 169680 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1525
timestamp 1654395037
transform 1 0 172144 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1535
timestamp 1654395037
transform 1 0 173264 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1539
timestamp 1654395037
transform 1 0 173712 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1560
timestamp 1654395037
transform 1 0 176064 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1568
timestamp 1654395037
transform 1 0 176960 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1572
timestamp 1654395037
transform 1 0 177408 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1574
timestamp 1654395037
transform 1 0 177632 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1595
timestamp 1654395037
transform 1 0 179984 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1603
timestamp 1654395037
transform 1 0 180880 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1607
timestamp 1654395037
transform 1 0 181328 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1609
timestamp 1654395037
transform 1 0 181552 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1630
timestamp 1654395037
transform 1 0 183904 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1638
timestamp 1654395037
transform 1 0 184800 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1642
timestamp 1654395037
transform 1 0 185248 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1644
timestamp 1654395037
transform 1 0 185472 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1663
timestamp 1654395037
transform 1 0 187600 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1671
timestamp 1654395037
transform 1 0 188496 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1677
timestamp 1654395037
transform 1 0 189168 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1679
timestamp 1654395037
transform 1 0 189392 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1684
timestamp 1654395037
transform 1 0 189952 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1688
timestamp 1654395037
transform 1 0 190400 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1692
timestamp 1654395037
transform 1 0 190848 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1696
timestamp 1654395037
transform 1 0 191296 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1700
timestamp 1654395037
transform 1 0 191744 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1704
timestamp 1654395037
transform 1 0 192192 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1708
timestamp 1654395037
transform 1 0 192640 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1712
timestamp 1654395037
transform 1 0 193088 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1714
timestamp 1654395037
transform 1 0 193312 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1719
timestamp 1654395037
transform 1 0 193872 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1723
timestamp 1654395037
transform 1 0 194320 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1727
timestamp 1654395037
transform 1 0 194768 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1731
timestamp 1654395037
transform 1 0 195216 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1735
timestamp 1654395037
transform 1 0 195664 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1739
timestamp 1654395037
transform 1 0 196112 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1743
timestamp 1654395037
transform 1 0 196560 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1747
timestamp 1654395037
transform 1 0 197008 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1749
timestamp 1654395037
transform 1 0 197232 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1770
timestamp 1654395037
transform 1 0 199584 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1774
timestamp 1654395037
transform 1 0 200032 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1778
timestamp 1654395037
transform 1 0 200480 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1782
timestamp 1654395037
transform 1 0 200928 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1784
timestamp 1654395037
transform 1 0 201152 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1805
timestamp 1654395037
transform 1 0 203504 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1809
timestamp 1654395037
transform 1 0 203952 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1813
timestamp 1654395037
transform 1 0 204400 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1818
timestamp 1654395037
transform 1 0 204960 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1840
timestamp 1654395037
transform 1 0 207424 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1846
timestamp 1654395037
transform 1 0 208096 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1852
timestamp 1654395037
transform 1 0 208768 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1854
timestamp 1654395037
transform 1 0 208992 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1875
timestamp 1654395037
transform 1 0 211344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1879
timestamp 1654395037
transform 1 0 211792 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1883
timestamp 1654395037
transform 1 0 212240 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1887
timestamp 1654395037
transform 1 0 212688 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1889
timestamp 1654395037
transform 1 0 212912 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1894
timestamp 1654395037
transform 1 0 213472 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1898
timestamp 1654395037
transform 1 0 213920 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1902
timestamp 1654395037
transform 1 0 214368 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1906
timestamp 1654395037
transform 1 0 214816 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1910
timestamp 1654395037
transform 1 0 215264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1914
timestamp 1654395037
transform 1 0 215712 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1922
timestamp 1654395037
transform 1 0 216608 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1924
timestamp 1654395037
transform 1 0 216832 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1927
timestamp 1654395037
transform 1 0 217168 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_1935
timestamp 1654395037
transform 1 0 218064 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1937
timestamp 1654395037
transform 1 0 218288 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_2
timestamp 1654395037
transform 1 0 1568 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_34 pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 5152 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_50
timestamp 1654395037
transform 1 0 6944 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_69
timestamp 1654395037
transform 1 0 9072 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_75
timestamp 1654395037
transform 1 0 9744 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_79
timestamp 1654395037
transform 1 0 10192 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_81
timestamp 1654395037
transform 1 0 10416 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_84
timestamp 1654395037
transform 1 0 10752 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_104
timestamp 1654395037
transform 1 0 12992 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_140
timestamp 1654395037
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_146
timestamp 1654395037
transform 1 0 17696 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_150
timestamp 1654395037
transform 1 0 18144 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_152
timestamp 1654395037
transform 1 0 18368 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_171
timestamp 1654395037
transform 1 0 20496 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_191
timestamp 1654395037
transform 1 0 22736 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_211
timestamp 1654395037
transform 1 0 24976 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_217
timestamp 1654395037
transform 1 0 25648 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_221
timestamp 1654395037
transform 1 0 26096 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_223
timestamp 1654395037
transform 1 0 26320 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_242
timestamp 1654395037
transform 1 0 28448 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_262
timestamp 1654395037
transform 1 0 30688 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_282
timestamp 1654395037
transform 1 0 32928 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_288
timestamp 1654395037
transform 1 0 33600 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_292
timestamp 1654395037
transform 1 0 34048 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_300
timestamp 1654395037
transform 1 0 34944 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_302
timestamp 1654395037
transform 1 0 35168 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_321
timestamp 1654395037
transform 1 0 37296 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_325
timestamp 1654395037
transform 1 0 37744 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_341
timestamp 1654395037
transform 1 0 39536 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_349
timestamp 1654395037
transform 1 0 40432 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_353
timestamp 1654395037
transform 1 0 40880 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_357
timestamp 1654395037
transform 1 0 41328 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_365
timestamp 1654395037
transform 1 0 42224 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_368
timestamp 1654395037
transform 1 0 42560 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_372
timestamp 1654395037
transform 1 0 43008 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_376
timestamp 1654395037
transform 1 0 43456 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_378
timestamp 1654395037
transform 1 0 43680 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_381
timestamp 1654395037
transform 1 0 44016 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_385
timestamp 1654395037
transform 1 0 44464 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_387
timestamp 1654395037
transform 1 0 44688 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_406
timestamp 1654395037
transform 1 0 46816 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_410
timestamp 1654395037
transform 1 0 47264 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_420
timestamp 1654395037
transform 1 0 48384 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_424
timestamp 1654395037
transform 1 0 48832 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_446
timestamp 1654395037
transform 1 0 51296 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_450
timestamp 1654395037
transform 1 0 51744 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_452
timestamp 1654395037
transform 1 0 51968 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_455
timestamp 1654395037
transform 1 0 52304 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_491
timestamp 1654395037
transform 1 0 56336 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_495
timestamp 1654395037
transform 1 0 56784 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_501
timestamp 1654395037
transform 1 0 57456 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_505
timestamp 1654395037
transform 1 0 57904 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_511
timestamp 1654395037
transform 1 0 58576 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_515
timestamp 1654395037
transform 1 0 59024 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_547
timestamp 1654395037
transform 1 0 62608 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_563
timestamp 1654395037
transform 1 0 64400 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_567
timestamp 1654395037
transform 1 0 64848 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_570
timestamp 1654395037
transform 1 0 65184 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_578
timestamp 1654395037
transform 1 0 66080 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_582
timestamp 1654395037
transform 1 0 66528 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_584
timestamp 1654395037
transform 1 0 66752 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_587
timestamp 1654395037
transform 1 0 67088 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_591
timestamp 1654395037
transform 1 0 67536 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_595
timestamp 1654395037
transform 1 0 67984 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_599
timestamp 1654395037
transform 1 0 68432 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_603
timestamp 1654395037
transform 1 0 68880 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_609
timestamp 1654395037
transform 1 0 69552 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_615
timestamp 1654395037
transform 1 0 70224 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_621
timestamp 1654395037
transform 1 0 70896 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_627
timestamp 1654395037
transform 1 0 71568 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_633
timestamp 1654395037
transform 1 0 72240 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_637
timestamp 1654395037
transform 1 0 72688 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_645
timestamp 1654395037
transform 1 0 73584 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_649
timestamp 1654395037
transform 1 0 74032 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_654
timestamp 1654395037
transform 1 0 74592 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_658
timestamp 1654395037
transform 1 0 75040 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_677
timestamp 1654395037
transform 1 0 77168 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_679
timestamp 1654395037
transform 1 0 77392 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_682
timestamp 1654395037
transform 1 0 77728 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_686
timestamp 1654395037
transform 1 0 78176 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_688
timestamp 1654395037
transform 1 0 78400 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_691
timestamp 1654395037
transform 1 0 78736 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_699
timestamp 1654395037
transform 1 0 79632 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_702
timestamp 1654395037
transform 1 0 79968 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_730
timestamp 1654395037
transform 1 0 83104 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_752
timestamp 1654395037
transform 1 0 85568 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_756
timestamp 1654395037
transform 1 0 86016 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_772
timestamp 1654395037
transform 1 0 87808 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_775
timestamp 1654395037
transform 1 0 88144 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_779
timestamp 1654395037
transform 1 0 88592 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_783 pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 89040 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_847
timestamp 1654395037
transform 1 0 96208 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_851
timestamp 1654395037
transform 1 0 96656 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_854
timestamp 1654395037
transform 1 0 96992 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_870
timestamp 1654395037
transform 1 0 98784 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_889
timestamp 1654395037
transform 1 0 100912 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_893
timestamp 1654395037
transform 1 0 101360 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_897
timestamp 1654395037
transform 1 0 101808 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_913
timestamp 1654395037
transform 1 0 103600 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_921
timestamp 1654395037
transform 1 0 104496 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_925
timestamp 1654395037
transform 1 0 104944 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_957
timestamp 1654395037
transform 1 0 108528 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_973
timestamp 1654395037
transform 1 0 110320 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_977
timestamp 1654395037
transform 1 0 110768 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_980
timestamp 1654395037
transform 1 0 111104 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_984
timestamp 1654395037
transform 1 0 111552 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_992
timestamp 1654395037
transform 1 0 112448 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_996
timestamp 1654395037
transform 1 0 112896 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_1028
timestamp 1654395037
transform 1 0 116480 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1036
timestamp 1654395037
transform 1 0 117376 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1055
timestamp 1654395037
transform 1 0 119504 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_1059
timestamp 1654395037
transform 1 0 119952 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1063
timestamp 1654395037
transform 1 0 120400 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_1067
timestamp 1654395037
transform 1 0 120848 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_1075
timestamp 1654395037
transform 1 0 121744 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1079
timestamp 1654395037
transform 1 0 122192 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_1083
timestamp 1654395037
transform 1 0 122640 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1115
timestamp 1654395037
transform 1 0 126224 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1117
timestamp 1654395037
transform 1 0 126448 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1120
timestamp 1654395037
transform 1 0 126784 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_1124
timestamp 1654395037
transform 1 0 127232 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1134
timestamp 1654395037
transform 1 0 128352 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1156
timestamp 1654395037
transform 1 0 130816 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1160
timestamp 1654395037
transform 1 0 131264 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1164
timestamp 1654395037
transform 1 0 131712 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1168
timestamp 1654395037
transform 1 0 132160 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1172
timestamp 1654395037
transform 1 0 132608 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1192
timestamp 1654395037
transform 1 0 134848 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1196
timestamp 1654395037
transform 1 0 135296 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1200
timestamp 1654395037
transform 1 0 135744 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1204
timestamp 1654395037
transform 1 0 136192 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1206
timestamp 1654395037
transform 1 0 136416 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1209
timestamp 1654395037
transform 1 0 136752 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1229
timestamp 1654395037
transform 1 0 138992 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1247
timestamp 1654395037
transform 1 0 141008 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1265
timestamp 1654395037
transform 1 0 143024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1269
timestamp 1654395037
transform 1 0 143472 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_1273
timestamp 1654395037
transform 1 0 143920 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1277
timestamp 1654395037
transform 1 0 144368 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1296
timestamp 1654395037
transform 1 0 146496 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1314
timestamp 1654395037
transform 1 0 148512 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1318
timestamp 1654395037
transform 1 0 148960 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1322
timestamp 1654395037
transform 1 0 149408 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1340
timestamp 1654395037
transform 1 0 151424 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_1344
timestamp 1654395037
transform 1 0 151872 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1348
timestamp 1654395037
transform 1 0 152320 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1367
timestamp 1654395037
transform 1 0 154448 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1371
timestamp 1654395037
transform 1 0 154896 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_1375
timestamp 1654395037
transform 1 0 155344 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1379
timestamp 1654395037
transform 1 0 155792 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1396
timestamp 1654395037
transform 1 0 157696 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_1416
timestamp 1654395037
transform 1 0 159936 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1424
timestamp 1654395037
transform 1 0 160832 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1426
timestamp 1654395037
transform 1 0 161056 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1461
timestamp 1654395037
transform 1 0 164976 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1481
timestamp 1654395037
transform 1 0 167216 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1489
timestamp 1654395037
transform 1 0 168112 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_1511
timestamp 1654395037
transform 1 0 170576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1549
timestamp 1654395037
transform 1 0 174832 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_1557
timestamp 1654395037
transform 1 0 175728 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1561
timestamp 1654395037
transform 1 0 176176 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1598
timestamp 1654395037
transform 1 0 180320 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1618
timestamp 1654395037
transform 1 0 182560 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1626
timestamp 1654395037
transform 1 0 183456 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1630
timestamp 1654395037
transform 1 0 183904 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1632
timestamp 1654395037
transform 1 0 184128 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1653
timestamp 1654395037
transform 1 0 186480 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1671
timestamp 1654395037
transform 1 0 188496 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1689
timestamp 1654395037
transform 1 0 190512 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1695
timestamp 1654395037
transform 1 0 191184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_1699
timestamp 1654395037
transform 1 0 191632 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1703
timestamp 1654395037
transform 1 0 192080 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1708
timestamp 1654395037
transform 1 0 192640 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1712
timestamp 1654395037
transform 1 0 193088 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1716
timestamp 1654395037
transform 1 0 193536 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1720
timestamp 1654395037
transform 1 0 193984 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1724
timestamp 1654395037
transform 1 0 194432 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1728
timestamp 1654395037
transform 1 0 194880 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1732
timestamp 1654395037
transform 1 0 195328 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_1736
timestamp 1654395037
transform 1 0 195776 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1758
timestamp 1654395037
transform 1 0 198240 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1762
timestamp 1654395037
transform 1 0 198688 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1766
timestamp 1654395037
transform 1 0 199136 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_1770
timestamp 1654395037
transform 1 0 199584 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1774
timestamp 1654395037
transform 1 0 200032 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1779
timestamp 1654395037
transform 1 0 200592 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1783
timestamp 1654395037
transform 1 0 201040 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1819
timestamp 1654395037
transform 1 0 205072 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1839
timestamp 1654395037
transform 1 0 207312 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1843
timestamp 1654395037
transform 1 0 207760 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1845
timestamp 1654395037
transform 1 0 207984 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1882
timestamp 1654395037
transform 1 0 212128 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1886
timestamp 1654395037
transform 1 0 212576 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1890
timestamp 1654395037
transform 1 0 213024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1894
timestamp 1654395037
transform 1 0 213472 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1898
timestamp 1654395037
transform 1 0 213920 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1902
timestamp 1654395037
transform 1 0 214368 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1906
timestamp 1654395037
transform 1 0 214816 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_1910
timestamp 1654395037
transform 1 0 215264 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1914
timestamp 1654395037
transform 1 0 215712 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1916
timestamp 1654395037
transform 1 0 215936 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_1919
timestamp 1654395037
transform 1 0 216272 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_1935
timestamp 1654395037
transform 1 0 218064 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1937
timestamp 1654395037
transform 1 0 218288 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_2
timestamp 1654395037
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_34
timestamp 1654395037
transform 1 0 5152 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_37
timestamp 1654395037
transform 1 0 5488 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_53
timestamp 1654395037
transform 1 0 7280 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_61
timestamp 1654395037
transform 1 0 8176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_65
timestamp 1654395037
transform 1 0 8624 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_68
timestamp 1654395037
transform 1 0 8960 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_104
timestamp 1654395037
transform 1 0 12992 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_110
timestamp 1654395037
transform 1 0 13664 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_114
timestamp 1654395037
transform 1 0 14112 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_152
timestamp 1654395037
transform 1 0 18368 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_156
timestamp 1654395037
transform 1 0 18816 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_175
timestamp 1654395037
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_181
timestamp 1654395037
transform 1 0 21616 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_189
timestamp 1654395037
transform 1 0 22512 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_208
timestamp 1654395037
transform 1 0 24640 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_212
timestamp 1654395037
transform 1 0 25088 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_238
timestamp 1654395037
transform 1 0 28000 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_242
timestamp 1654395037
transform 1 0 28448 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_246
timestamp 1654395037
transform 1 0 28896 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_250
timestamp 1654395037
transform 1 0 29344 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_258
timestamp 1654395037
transform 1 0 30240 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_260
timestamp 1654395037
transform 1 0 30464 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_263
timestamp 1654395037
transform 1 0 30800 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_299
timestamp 1654395037
transform 1 0 34832 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_303
timestamp 1654395037
transform 1 0 35280 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_307
timestamp 1654395037
transform 1 0 35728 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_315
timestamp 1654395037
transform 1 0 36624 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_321
timestamp 1654395037
transform 1 0 37296 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_329
timestamp 1654395037
transform 1 0 38192 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_333
timestamp 1654395037
transform 1 0 38640 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_335
timestamp 1654395037
transform 1 0 38864 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_338
timestamp 1654395037
transform 1 0 39200 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_342
timestamp 1654395037
transform 1 0 39648 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_377
timestamp 1654395037
transform 1 0 43568 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_379
timestamp 1654395037
transform 1 0 43792 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_382
timestamp 1654395037
transform 1 0 44128 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_386
timestamp 1654395037
transform 1 0 44576 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_392
timestamp 1654395037
transform 1 0 45248 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_408
timestamp 1654395037
transform 1 0 47040 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_412
timestamp 1654395037
transform 1 0 47488 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_430
timestamp 1654395037
transform 1 0 49504 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_432
timestamp 1654395037
transform 1 0 49728 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_435
timestamp 1654395037
transform 1 0 50064 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_441
timestamp 1654395037
transform 1 0 50736 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_445
timestamp 1654395037
transform 1 0 51184 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_451
timestamp 1654395037
transform 1 0 51856 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_455
timestamp 1654395037
transform 1 0 52304 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_459
timestamp 1654395037
transform 1 0 52752 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_497
timestamp 1654395037
transform 1 0 57008 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_503
timestamp 1654395037
transform 1 0 57680 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_509
timestamp 1654395037
transform 1 0 58352 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_513
timestamp 1654395037
transform 1 0 58800 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_517
timestamp 1654395037
transform 1 0 59248 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_520
timestamp 1654395037
transform 1 0 59584 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_524
timestamp 1654395037
transform 1 0 60032 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_534
timestamp 1654395037
transform 1 0 61152 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_538
timestamp 1654395037
transform 1 0 61600 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_541
timestamp 1654395037
transform 1 0 61936 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_577
timestamp 1654395037
transform 1 0 65968 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_583
timestamp 1654395037
transform 1 0 66640 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_587
timestamp 1654395037
transform 1 0 67088 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_591
timestamp 1654395037
transform 1 0 67536 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_595
timestamp 1654395037
transform 1 0 67984 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_601
timestamp 1654395037
transform 1 0 68656 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_605
timestamp 1654395037
transform 1 0 69104 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_610
timestamp 1654395037
transform 1 0 69664 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_616
timestamp 1654395037
transform 1 0 70336 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_652
timestamp 1654395037
transform 1 0 74368 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_656
timestamp 1654395037
transform 1 0 74816 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_661
timestamp 1654395037
transform 1 0 75376 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_667
timestamp 1654395037
transform 1 0 76048 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_671
timestamp 1654395037
transform 1 0 76496 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_673
timestamp 1654395037
transform 1 0 76720 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_680
timestamp 1654395037
transform 1 0 77504 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_682
timestamp 1654395037
transform 1 0 77728 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_685
timestamp 1654395037
transform 1 0 78064 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_689
timestamp 1654395037
transform 1 0 78512 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_725
timestamp 1654395037
transform 1 0 82544 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_731
timestamp 1654395037
transform 1 0 83216 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_735
timestamp 1654395037
transform 1 0 83664 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_739
timestamp 1654395037
transform 1 0 84112 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_743
timestamp 1654395037
transform 1 0 84560 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_751
timestamp 1654395037
transform 1 0 85456 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_755
timestamp 1654395037
transform 1 0 85904 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_759
timestamp 1654395037
transform 1 0 86352 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_795
timestamp 1654395037
transform 1 0 90384 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_801
timestamp 1654395037
transform 1 0 91056 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_805
timestamp 1654395037
transform 1 0 91504 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_809
timestamp 1654395037
transform 1 0 91952 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_813
timestamp 1654395037
transform 1 0 92400 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_815
timestamp 1654395037
transform 1 0 92624 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_818
timestamp 1654395037
transform 1 0 92960 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_834
timestamp 1654395037
transform 1 0 94752 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_842
timestamp 1654395037
transform 1 0 95648 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_859
timestamp 1654395037
transform 1 0 97552 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_863
timestamp 1654395037
transform 1 0 98000 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_867
timestamp 1654395037
transform 1 0 98448 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_885
timestamp 1654395037
transform 1 0 100464 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_891
timestamp 1654395037
transform 1 0 101136 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_897
timestamp 1654395037
transform 1 0 101808 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_933
timestamp 1654395037
transform 1 0 105840 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_951
timestamp 1654395037
transform 1 0 107856 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_955
timestamp 1654395037
transform 1 0 108304 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_957
timestamp 1654395037
transform 1 0 108528 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_976
timestamp 1654395037
transform 1 0 110656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_996
timestamp 1654395037
transform 1 0 112896 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1000
timestamp 1654395037
transform 1 0 113344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_1004
timestamp 1654395037
transform 1 0 113792 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1020
timestamp 1654395037
transform 1 0 115584 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1022
timestamp 1654395037
transform 1 0 115808 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1025
timestamp 1654395037
transform 1 0 116144 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_1031
timestamp 1654395037
transform 1 0 116816 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1039
timestamp 1654395037
transform 1 0 117712 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1043
timestamp 1654395037
transform 1 0 118160 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1046
timestamp 1654395037
transform 1 0 118496 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_1050
timestamp 1654395037
transform 1 0 118944 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1066
timestamp 1654395037
transform 1 0 120736 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1084
timestamp 1654395037
transform 1 0 122752 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1088
timestamp 1654395037
transform 1 0 123200 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_1092
timestamp 1654395037
transform 1 0 123648 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1118
timestamp 1654395037
transform 1 0 126560 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1120
timestamp 1654395037
transform 1 0 126784 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1137
timestamp 1654395037
transform 1 0 128688 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1141
timestamp 1654395037
transform 1 0 129136 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1158
timestamp 1654395037
transform 1 0 131040 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1162
timestamp 1654395037
transform 1 0 131488 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1166
timestamp 1654395037
transform 1 0 131936 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1170
timestamp 1654395037
transform 1 0 132384 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1189
timestamp 1654395037
transform 1 0 134512 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1207
timestamp 1654395037
transform 1 0 136528 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1225
timestamp 1654395037
transform 1 0 138544 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1229
timestamp 1654395037
transform 1 0 138992 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1233
timestamp 1654395037
transform 1 0 139440 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1237
timestamp 1654395037
transform 1 0 139888 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1241
timestamp 1654395037
transform 1 0 140336 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1260
timestamp 1654395037
transform 1 0 142464 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1278
timestamp 1654395037
transform 1 0 144480 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1296
timestamp 1654395037
transform 1 0 146496 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1300
timestamp 1654395037
transform 1 0 146944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1304
timestamp 1654395037
transform 1 0 147392 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1308
timestamp 1654395037
transform 1 0 147840 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1312
timestamp 1654395037
transform 1 0 148288 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1331
timestamp 1654395037
transform 1 0 150416 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1335
timestamp 1654395037
transform 1 0 150864 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1339
timestamp 1654395037
transform 1 0 151312 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1357
timestamp 1654395037
transform 1 0 153328 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1361
timestamp 1654395037
transform 1 0 153776 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1365
timestamp 1654395037
transform 1 0 154224 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1382
timestamp 1654395037
transform 1 0 156128 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1386
timestamp 1654395037
transform 1 0 156576 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1403
timestamp 1654395037
transform 1 0 158480 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1423
timestamp 1654395037
transform 1 0 160720 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1443
timestamp 1654395037
transform 1 0 162960 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1447
timestamp 1654395037
transform 1 0 163408 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1451
timestamp 1654395037
transform 1 0 163856 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1459
timestamp 1654395037
transform 1 0 164752 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1463
timestamp 1654395037
transform 1 0 165200 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1501
timestamp 1654395037
transform 1 0 169456 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1521
timestamp 1654395037
transform 1 0 171696 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1525
timestamp 1654395037
transform 1 0 172144 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1562
timestamp 1654395037
transform 1 0 176288 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1582
timestamp 1654395037
transform 1 0 178528 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1590
timestamp 1654395037
transform 1 0 179424 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1594
timestamp 1654395037
transform 1 0 179872 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1596
timestamp 1654395037
transform 1 0 180096 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1601
timestamp 1654395037
transform 1 0 180656 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1603
timestamp 1654395037
transform 1 0 180880 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1638
timestamp 1654395037
transform 1 0 184800 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1656
timestamp 1654395037
transform 1 0 186816 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1664
timestamp 1654395037
transform 1 0 187712 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1686
timestamp 1654395037
transform 1 0 190176 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1692
timestamp 1654395037
transform 1 0 190848 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1698
timestamp 1654395037
transform 1 0 191520 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1702
timestamp 1654395037
transform 1 0 191968 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1706
timestamp 1654395037
transform 1 0 192416 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1710
timestamp 1654395037
transform 1 0 192864 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1714
timestamp 1654395037
transform 1 0 193312 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1718
timestamp 1654395037
transform 1 0 193760 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1720
timestamp 1654395037
transform 1 0 193984 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1725
timestamp 1654395037
transform 1 0 194544 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1729
timestamp 1654395037
transform 1 0 194992 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1733
timestamp 1654395037
transform 1 0 195440 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1737
timestamp 1654395037
transform 1 0 195888 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1743
timestamp 1654395037
transform 1 0 196560 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1747
timestamp 1654395037
transform 1 0 197008 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1751
timestamp 1654395037
transform 1 0 197456 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1755
timestamp 1654395037
transform 1 0 197904 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1759
timestamp 1654395037
transform 1 0 198352 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1763
timestamp 1654395037
transform 1 0 198800 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1798
timestamp 1654395037
transform 1 0 202720 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1804
timestamp 1654395037
transform 1 0 203392 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1808
timestamp 1654395037
transform 1 0 203840 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1846
timestamp 1654395037
transform 1 0 208096 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1866
timestamp 1654395037
transform 1 0 210336 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1872
timestamp 1654395037
transform 1 0 211008 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1878
timestamp 1654395037
transform 1 0 211680 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1880
timestamp 1654395037
transform 1 0 211904 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1885
timestamp 1654395037
transform 1 0 212464 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1889
timestamp 1654395037
transform 1 0 212912 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1893
timestamp 1654395037
transform 1 0 213360 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1897
timestamp 1654395037
transform 1 0 213808 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1901
timestamp 1654395037
transform 1 0 214256 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1905
timestamp 1654395037
transform 1 0 214704 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_1909
timestamp 1654395037
transform 1 0 215152 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_1913
timestamp 1654395037
transform 1 0 215600 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_1929
timestamp 1654395037
transform 1 0 217392 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1937
timestamp 1654395037
transform 1 0 218288 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_2
timestamp 1654395037
transform 1 0 1568 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_34
timestamp 1654395037
transform 1 0 5152 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_69
timestamp 1654395037
transform 1 0 9072 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_75
timestamp 1654395037
transform 1 0 9744 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_79
timestamp 1654395037
transform 1 0 10192 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_82
timestamp 1654395037
transform 1 0 10528 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_104
timestamp 1654395037
transform 1 0 12992 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_140
timestamp 1654395037
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_146
timestamp 1654395037
transform 1 0 17696 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_150
timestamp 1654395037
transform 1 0 18144 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_156
timestamp 1654395037
transform 1 0 18816 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_160
timestamp 1654395037
transform 1 0 19264 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_168
timestamp 1654395037
transform 1 0 20160 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_204
timestamp 1654395037
transform 1 0 24192 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_208
timestamp 1654395037
transform 1 0 24640 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_212
timestamp 1654395037
transform 1 0 25088 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_217
timestamp 1654395037
transform 1 0 25648 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_219
timestamp 1654395037
transform 1 0 25872 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_254
timestamp 1654395037
transform 1 0 29792 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_258
timestamp 1654395037
transform 1 0 30240 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_262
timestamp 1654395037
transform 1 0 30688 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_278
timestamp 1654395037
transform 1 0 32480 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_282
timestamp 1654395037
transform 1 0 32928 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_286
timestamp 1654395037
transform 1 0 33376 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_294
timestamp 1654395037
transform 1 0 34272 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_298
timestamp 1654395037
transform 1 0 34720 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_336
timestamp 1654395037
transform 1 0 38976 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_340
timestamp 1654395037
transform 1 0 39424 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_344
timestamp 1654395037
transform 1 0 39872 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_348
timestamp 1654395037
transform 1 0 40320 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_350
timestamp 1654395037
transform 1 0 40544 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_353
timestamp 1654395037
transform 1 0 40880 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_357
timestamp 1654395037
transform 1 0 41328 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_359
timestamp 1654395037
transform 1 0 41552 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_366
timestamp 1654395037
transform 1 0 42336 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_374
timestamp 1654395037
transform 1 0 43232 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_382
timestamp 1654395037
transform 1 0 44128 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_388
timestamp 1654395037
transform 1 0 44800 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_424
timestamp 1654395037
transform 1 0 48832 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_434
timestamp 1654395037
transform 1 0 49952 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_438
timestamp 1654395037
transform 1 0 50400 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_455
timestamp 1654395037
transform 1 0 52304 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_459
timestamp 1654395037
transform 1 0 52752 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_495
timestamp 1654395037
transform 1 0 56784 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_499
timestamp 1654395037
transform 1 0 57232 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_516
timestamp 1654395037
transform 1 0 59136 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_518
timestamp 1654395037
transform 1 0 59360 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_521
timestamp 1654395037
transform 1 0 59696 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_527
timestamp 1654395037
transform 1 0 60368 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_535
timestamp 1654395037
transform 1 0 61264 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_552
timestamp 1654395037
transform 1 0 63168 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_556
timestamp 1654395037
transform 1 0 63616 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_560
timestamp 1654395037
transform 1 0 64064 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_586
timestamp 1654395037
transform 1 0 66976 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_590
timestamp 1654395037
transform 1 0 67424 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_594
timestamp 1654395037
transform 1 0 67872 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_597
timestamp 1654395037
transform 1 0 68208 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_601
timestamp 1654395037
transform 1 0 68656 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_637
timestamp 1654395037
transform 1 0 72688 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_657
timestamp 1654395037
transform 1 0 74928 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_661
timestamp 1654395037
transform 1 0 75376 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_665
timestamp 1654395037
transform 1 0 75824 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_669
timestamp 1654395037
transform 1 0 76272 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_673
timestamp 1654395037
transform 1 0 76720 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_690
timestamp 1654395037
transform 1 0 78624 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_694
timestamp 1654395037
transform 1 0 79072 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_700
timestamp 1654395037
transform 1 0 79744 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_708
timestamp 1654395037
transform 1 0 80640 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_728
timestamp 1654395037
transform 1 0 82880 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_748
timestamp 1654395037
transform 1 0 85120 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_752
timestamp 1654395037
transform 1 0 85568 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_754
timestamp 1654395037
transform 1 0 85792 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_771
timestamp 1654395037
transform 1 0 87696 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_775
timestamp 1654395037
transform 1 0 88144 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_779
timestamp 1654395037
transform 1 0 88592 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_799
timestamp 1654395037
transform 1 0 90832 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_803
timestamp 1654395037
transform 1 0 91280 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_807
timestamp 1654395037
transform 1 0 91728 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_811
timestamp 1654395037
transform 1 0 92176 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_814
timestamp 1654395037
transform 1 0 92512 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_850
timestamp 1654395037
transform 1 0 96544 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_854
timestamp 1654395037
transform 1 0 96992 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_858
timestamp 1654395037
transform 1 0 97440 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_861
timestamp 1654395037
transform 1 0 97776 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_897
timestamp 1654395037
transform 1 0 101808 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_921
timestamp 1654395037
transform 1 0 104496 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_927
timestamp 1654395037
transform 1 0 105168 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_947
timestamp 1654395037
transform 1 0 107408 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_983
timestamp 1654395037
transform 1 0 111440 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_991
timestamp 1654395037
transform 1 0 112336 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_993
timestamp 1654395037
transform 1 0 112560 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_996
timestamp 1654395037
transform 1 0 112896 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1004
timestamp 1654395037
transform 1 0 113792 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1021
timestamp 1654395037
transform 1 0 115696 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1025
timestamp 1654395037
transform 1 0 116144 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1027
timestamp 1654395037
transform 1 0 116368 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1044
timestamp 1654395037
transform 1 0 118272 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1046
timestamp 1654395037
transform 1 0 118496 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1063
timestamp 1654395037
transform 1 0 120400 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1069
timestamp 1654395037
transform 1 0 121072 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1073
timestamp 1654395037
transform 1 0 121520 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_1109
timestamp 1654395037
transform 1 0 125552 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1117
timestamp 1654395037
transform 1 0 126448 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1122
timestamp 1654395037
transform 1 0 127008 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_1126
timestamp 1654395037
transform 1 0 127456 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1130
timestamp 1654395037
transform 1 0 127904 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1134
timestamp 1654395037
transform 1 0 128352 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1138
timestamp 1654395037
transform 1 0 128800 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1140
timestamp 1654395037
transform 1 0 129024 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1175
timestamp 1654395037
transform 1 0 132944 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1193
timestamp 1654395037
transform 1 0 134960 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_1197
timestamp 1654395037
transform 1 0 135408 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1205
timestamp 1654395037
transform 1 0 136304 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1225
timestamp 1654395037
transform 1 0 138544 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1243
timestamp 1654395037
transform 1 0 140560 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1261
timestamp 1654395037
transform 1 0 142576 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_1265
timestamp 1654395037
transform 1 0 143024 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_1273
timestamp 1654395037
transform 1 0 143920 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1277
timestamp 1654395037
transform 1 0 144368 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1282
timestamp 1654395037
transform 1 0 144928 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_1286
timestamp 1654395037
transform 1 0 145376 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1290
timestamp 1654395037
transform 1 0 145824 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1325
timestamp 1654395037
transform 1 0 149744 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1329
timestamp 1654395037
transform 1 0 150192 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1333
timestamp 1654395037
transform 1 0 150640 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1337
timestamp 1654395037
transform 1 0 151088 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1341
timestamp 1654395037
transform 1 0 151536 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_1345
timestamp 1654395037
transform 1 0 151984 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1367
timestamp 1654395037
transform 1 0 154448 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1385
timestamp 1654395037
transform 1 0 156464 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1389
timestamp 1654395037
transform 1 0 156912 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1393
timestamp 1654395037
transform 1 0 157360 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1397
timestamp 1654395037
transform 1 0 157808 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1399
timestamp 1654395037
transform 1 0 158032 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1418
timestamp 1654395037
transform 1 0 160160 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1456
timestamp 1654395037
transform 1 0 164416 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1476
timestamp 1654395037
transform 1 0 166656 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1484
timestamp 1654395037
transform 1 0 167552 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1488
timestamp 1654395037
transform 1 0 168000 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1490
timestamp 1654395037
transform 1 0 168224 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1527
timestamp 1654395037
transform 1 0 172368 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1547
timestamp 1654395037
transform 1 0 174608 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1555
timestamp 1654395037
transform 1 0 175504 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1559
timestamp 1654395037
transform 1 0 175952 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1561
timestamp 1654395037
transform 1 0 176176 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1598
timestamp 1654395037
transform 1 0 180320 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1604
timestamp 1654395037
transform 1 0 180992 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1606
timestamp 1654395037
transform 1 0 181216 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1625
timestamp 1654395037
transform 1 0 183344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1631
timestamp 1654395037
transform 1 0 184016 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1651
timestamp 1654395037
transform 1 0 186256 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1669
timestamp 1654395037
transform 1 0 188272 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1687
timestamp 1654395037
transform 1 0 190288 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1695
timestamp 1654395037
transform 1 0 191184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1697
timestamp 1654395037
transform 1 0 191408 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1702
timestamp 1654395037
transform 1 0 191968 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1708
timestamp 1654395037
transform 1 0 192640 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_1712
timestamp 1654395037
transform 1 0 193088 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1716
timestamp 1654395037
transform 1 0 193536 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1721
timestamp 1654395037
transform 1 0 194096 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1725
timestamp 1654395037
transform 1 0 194544 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1727
timestamp 1654395037
transform 1 0 194768 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1732
timestamp 1654395037
transform 1 0 195328 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1736
timestamp 1654395037
transform 1 0 195776 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1740
timestamp 1654395037
transform 1 0 196224 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1744
timestamp 1654395037
transform 1 0 196672 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1748
timestamp 1654395037
transform 1 0 197120 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1752
timestamp 1654395037
transform 1 0 197568 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1756
timestamp 1654395037
transform 1 0 198016 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1760
timestamp 1654395037
transform 1 0 198464 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1764
timestamp 1654395037
transform 1 0 198912 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1768
timestamp 1654395037
transform 1 0 199360 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1772
timestamp 1654395037
transform 1 0 199808 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1774
timestamp 1654395037
transform 1 0 200032 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1795
timestamp 1654395037
transform 1 0 202384 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1799
timestamp 1654395037
transform 1 0 202832 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1803
timestamp 1654395037
transform 1 0 203280 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1807
timestamp 1654395037
transform 1 0 203728 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1809
timestamp 1654395037
transform 1 0 203952 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1844
timestamp 1654395037
transform 1 0 207872 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1864
timestamp 1654395037
transform 1 0 210112 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1872
timestamp 1654395037
transform 1 0 211008 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1876
timestamp 1654395037
transform 1 0 211456 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1880
timestamp 1654395037
transform 1 0 211904 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1884
timestamp 1654395037
transform 1 0 212352 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1888
timestamp 1654395037
transform 1 0 212800 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1892
timestamp 1654395037
transform 1 0 213248 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1896
timestamp 1654395037
transform 1 0 213696 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1900
timestamp 1654395037
transform 1 0 214144 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1904
timestamp 1654395037
transform 1 0 214592 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1908
timestamp 1654395037
transform 1 0 215040 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_1912
timestamp 1654395037
transform 1 0 215488 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1916
timestamp 1654395037
transform 1 0 215936 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_1919
timestamp 1654395037
transform 1 0 216272 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_1935
timestamp 1654395037
transform 1 0 218064 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1937
timestamp 1654395037
transform 1 0 218288 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_2
timestamp 1654395037
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_34
timestamp 1654395037
transform 1 0 5152 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_37
timestamp 1654395037
transform 1 0 5488 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_69
timestamp 1654395037
transform 1 0 9072 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_104
timestamp 1654395037
transform 1 0 12992 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_110
timestamp 1654395037
transform 1 0 13664 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_114
timestamp 1654395037
transform 1 0 14112 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_118
timestamp 1654395037
transform 1 0 14560 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_153
timestamp 1654395037
transform 1 0 18480 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_157
timestamp 1654395037
transform 1 0 18928 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_161
timestamp 1654395037
transform 1 0 19376 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_213
timestamp 1654395037
transform 1 0 25200 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_217
timestamp 1654395037
transform 1 0 25648 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_221
timestamp 1654395037
transform 1 0 26096 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_223
timestamp 1654395037
transform 1 0 26320 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_230
timestamp 1654395037
transform 1 0 27104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_234
timestamp 1654395037
transform 1 0 27552 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_242
timestamp 1654395037
transform 1 0 28448 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_246
timestamp 1654395037
transform 1 0 28896 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_256
timestamp 1654395037
transform 1 0 30016 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_260
timestamp 1654395037
transform 1 0 30464 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_274
timestamp 1654395037
transform 1 0 32032 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_278
timestamp 1654395037
transform 1 0 32480 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_286
timestamp 1654395037
transform 1 0 33376 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_296
timestamp 1654395037
transform 1 0 34496 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_304
timestamp 1654395037
transform 1 0 35392 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_308
timestamp 1654395037
transform 1 0 35840 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_310
timestamp 1654395037
transform 1 0 36064 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_317
timestamp 1654395037
transform 1 0 36848 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_327
timestamp 1654395037
transform 1 0 37968 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_331
timestamp 1654395037
transform 1 0 38416 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_338
timestamp 1654395037
transform 1 0 39200 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_346
timestamp 1654395037
transform 1 0 40096 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_356
timestamp 1654395037
transform 1 0 41216 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_364
timestamp 1654395037
transform 1 0 42112 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_372
timestamp 1654395037
transform 1 0 43008 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_380
timestamp 1654395037
transform 1 0 43904 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_388
timestamp 1654395037
transform 1 0 44800 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_392
timestamp 1654395037
transform 1 0 45248 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_399
timestamp 1654395037
transform 1 0 46032 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_407
timestamp 1654395037
transform 1 0 46928 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_415
timestamp 1654395037
transform 1 0 47824 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_423
timestamp 1654395037
transform 1 0 48720 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_459
timestamp 1654395037
transform 1 0 52752 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_463
timestamp 1654395037
transform 1 0 53200 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_467
timestamp 1654395037
transform 1 0 53648 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_475
timestamp 1654395037
transform 1 0 54544 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_511
timestamp 1654395037
transform 1 0 58576 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_519
timestamp 1654395037
transform 1 0 59472 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_525
timestamp 1654395037
transform 1 0 60144 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_527
timestamp 1654395037
transform 1 0 60368 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_530
timestamp 1654395037
transform 1 0 60704 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_534
timestamp 1654395037
transform 1 0 61152 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_569
timestamp 1654395037
transform 1 0 65072 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_579
timestamp 1654395037
transform 1 0 66192 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_583
timestamp 1654395037
transform 1 0 66640 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_591
timestamp 1654395037
transform 1 0 67536 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_595
timestamp 1654395037
transform 1 0 67984 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_601
timestamp 1654395037
transform 1 0 68656 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_621
timestamp 1654395037
transform 1 0 70896 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_623
timestamp 1654395037
transform 1 0 71120 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_630
timestamp 1654395037
transform 1 0 71904 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_636
timestamp 1654395037
transform 1 0 72576 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_672
timestamp 1654395037
transform 1 0 76608 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_676
timestamp 1654395037
transform 1 0 77056 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_680
timestamp 1654395037
transform 1 0 77504 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_682
timestamp 1654395037
transform 1 0 77728 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_685
timestamp 1654395037
transform 1 0 78064 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_689
timestamp 1654395037
transform 1 0 78512 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_693
timestamp 1654395037
transform 1 0 78960 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_699
timestamp 1654395037
transform 1 0 79632 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_707
timestamp 1654395037
transform 1 0 80528 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_743
timestamp 1654395037
transform 1 0 84560 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_747
timestamp 1654395037
transform 1 0 85008 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_750
timestamp 1654395037
transform 1 0 85344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_756
timestamp 1654395037
transform 1 0 86016 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_758
timestamp 1654395037
transform 1 0 86240 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_765
timestamp 1654395037
transform 1 0 87024 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_769
timestamp 1654395037
transform 1 0 87472 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_774
timestamp 1654395037
transform 1 0 88032 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_780
timestamp 1654395037
transform 1 0 88704 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_784
timestamp 1654395037
transform 1 0 89152 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_792
timestamp 1654395037
transform 1 0 90048 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_798
timestamp 1654395037
transform 1 0 90720 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_804
timestamp 1654395037
transform 1 0 91392 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_808
timestamp 1654395037
transform 1 0 91840 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_818
timestamp 1654395037
transform 1 0 92960 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_842
timestamp 1654395037
transform 1 0 95648 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_846
timestamp 1654395037
transform 1 0 96096 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_849
timestamp 1654395037
transform 1 0 96432 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_885
timestamp 1654395037
transform 1 0 100464 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_889
timestamp 1654395037
transform 1 0 100912 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_893
timestamp 1654395037
transform 1 0 101360 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_910
timestamp 1654395037
transform 1 0 103264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_914
timestamp 1654395037
transform 1 0 103712 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_918
timestamp 1654395037
transform 1 0 104160 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_920
timestamp 1654395037
transform 1 0 104384 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_923
timestamp 1654395037
transform 1 0 104720 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_939
timestamp 1654395037
transform 1 0 106512 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_949
timestamp 1654395037
transform 1 0 107632 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_953
timestamp 1654395037
transform 1 0 108080 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_957
timestamp 1654395037
transform 1 0 108528 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_960
timestamp 1654395037
transform 1 0 108864 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_968
timestamp 1654395037
transform 1 0 109760 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_976
timestamp 1654395037
transform 1 0 110656 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_980
timestamp 1654395037
transform 1 0 111104 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_1012
timestamp 1654395037
transform 1 0 114688 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_1020
timestamp 1654395037
transform 1 0 115584 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1024
timestamp 1654395037
transform 1 0 116032 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_1027
timestamp 1654395037
transform 1 0 116368 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_1065
timestamp 1654395037
transform 1 0 120624 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_1075
timestamp 1654395037
transform 1 0 121744 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_1083
timestamp 1654395037
transform 1 0 122640 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_1091
timestamp 1654395037
transform 1 0 123536 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_1095
timestamp 1654395037
transform 1 0 123984 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1099
timestamp 1654395037
transform 1 0 124432 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1102
timestamp 1654395037
transform 1 0 124768 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_1137
timestamp 1654395037
transform 1 0 128688 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_1141
timestamp 1654395037
transform 1 0 129136 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_1149
timestamp 1654395037
transform 1 0 130032 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_1155
timestamp 1654395037
transform 1 0 130704 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_1159
timestamp 1654395037
transform 1 0 131152 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1161
timestamp 1654395037
transform 1 0 131376 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_1164
timestamp 1654395037
transform 1 0 131712 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1166
timestamp 1654395037
transform 1 0 131936 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_1169
timestamp 1654395037
transform 1 0 132272 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_1173
timestamp 1654395037
transform 1 0 132720 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1175
timestamp 1654395037
transform 1 0 132944 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_1182
timestamp 1654395037
transform 1 0 133728 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_1186
timestamp 1654395037
transform 1 0 134176 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_1222
timestamp 1654395037
transform 1 0 138208 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_1240
timestamp 1654395037
transform 1 0 140224 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_1278
timestamp 1654395037
transform 1 0 144480 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1282
timestamp 1654395037
transform 1 0 144928 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_1299
timestamp 1654395037
transform 1 0 146832 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_1303
timestamp 1654395037
transform 1 0 147280 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_1307
timestamp 1654395037
transform 1 0 147728 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_1311
timestamp 1654395037
transform 1 0 148176 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_1331
timestamp 1654395037
transform 1 0 150416 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_1335
timestamp 1654395037
transform 1 0 150864 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_1339
timestamp 1654395037
transform 1 0 151312 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1341
timestamp 1654395037
transform 1 0 151536 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_1346
timestamp 1654395037
transform 1 0 152096 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_1382
timestamp 1654395037
transform 1 0 156128 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_1388
timestamp 1654395037
transform 1 0 156800 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_1426
timestamp 1654395037
transform 1 0 161056 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_1446
timestamp 1654395037
transform 1 0 163296 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1448
timestamp 1654395037
transform 1 0 163520 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_1453
timestamp 1654395037
transform 1 0 164080 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_1475
timestamp 1654395037
transform 1 0 166544 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_1495
timestamp 1654395037
transform 1 0 168784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_1515
timestamp 1654395037
transform 1 0 171024 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_1523
timestamp 1654395037
transform 1 0 171920 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1525
timestamp 1654395037
transform 1 0 172144 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_1534
timestamp 1654395037
transform 1 0 173152 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_1538
timestamp 1654395037
transform 1 0 173600 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1540
timestamp 1654395037
transform 1 0 173824 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_1575
timestamp 1654395037
transform 1 0 177744 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_1593
timestamp 1654395037
transform 1 0 179760 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_1615
timestamp 1654395037
transform 1 0 182224 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_1633
timestamp 1654395037
transform 1 0 184240 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_1651
timestamp 1654395037
transform 1 0 186256 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_1659
timestamp 1654395037
transform 1 0 187152 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_1665
timestamp 1654395037
transform 1 0 187824 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1667
timestamp 1654395037
transform 1 0 188048 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_1686
timestamp 1654395037
transform 1 0 190176 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_1694
timestamp 1654395037
transform 1 0 191072 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_1698
timestamp 1654395037
transform 1 0 191520 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1702
timestamp 1654395037
transform 1 0 191968 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_1737
timestamp 1654395037
transform 1 0 195888 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_1775
timestamp 1654395037
transform 1 0 200144 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_1779
timestamp 1654395037
transform 1 0 200592 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_1783
timestamp 1654395037
transform 1 0 201040 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_1787
timestamp 1654395037
transform 1 0 201488 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_1791
timestamp 1654395037
transform 1 0 201936 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_1795
timestamp 1654395037
transform 1 0 202384 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_1799
timestamp 1654395037
transform 1 0 202832 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_1803
timestamp 1654395037
transform 1 0 203280 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_1807
timestamp 1654395037
transform 1 0 203728 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1809
timestamp 1654395037
transform 1 0 203952 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_1814
timestamp 1654395037
transform 1 0 204512 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_1852
timestamp 1654395037
transform 1 0 208768 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_1872
timestamp 1654395037
transform 1 0 211008 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_1876
timestamp 1654395037
transform 1 0 211456 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1880
timestamp 1654395037
transform 1 0 211904 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_1885
timestamp 1654395037
transform 1 0 212464 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_1889
timestamp 1654395037
transform 1 0 212912 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_1893
timestamp 1654395037
transform 1 0 213360 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_1897
timestamp 1654395037
transform 1 0 213808 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_1901
timestamp 1654395037
transform 1 0 214256 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_1905
timestamp 1654395037
transform 1 0 214704 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_1909
timestamp 1654395037
transform 1 0 215152 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_1913
timestamp 1654395037
transform 1 0 215600 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_1917
timestamp 1654395037
transform 1 0 216048 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_1921
timestamp 1654395037
transform 1 0 216496 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1937
timestamp 1654395037
transform 1 0 218288 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_2
timestamp 1654395037
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_66
timestamp 1654395037
transform 1 0 8736 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_69
timestamp 1654395037
transform 1 0 9072 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_73
timestamp 1654395037
transform 1 0 9520 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_80
timestamp 1654395037
transform 1 0 10304 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_88
timestamp 1654395037
transform 1 0 11200 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_124
timestamp 1654395037
transform 1 0 15232 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_128
timestamp 1654395037
transform 1 0 15680 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_132
timestamp 1654395037
transform 1 0 16128 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_140
timestamp 1654395037
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_144
timestamp 1654395037
transform 1 0 17472 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_151
timestamp 1654395037
transform 1 0 18256 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_155
timestamp 1654395037
transform 1 0 18704 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_163
timestamp 1654395037
transform 1 0 19600 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_170
timestamp 1654395037
transform 1 0 20384 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_174
timestamp 1654395037
transform 1 0 20832 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_188
timestamp 1654395037
transform 1 0 22400 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_208
timestamp 1654395037
transform 1 0 24640 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_212
timestamp 1654395037
transform 1 0 25088 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_221
timestamp 1654395037
transform 1 0 26096 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_225
timestamp 1654395037
transform 1 0 26544 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_257
timestamp 1654395037
transform 1 0 30128 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_273
timestamp 1654395037
transform 1 0 31920 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_281
timestamp 1654395037
transform 1 0 32816 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_283
timestamp 1654395037
transform 1 0 33040 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_286
timestamp 1654395037
transform 1 0 33376 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_302
timestamp 1654395037
transform 1 0 35168 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_310
timestamp 1654395037
transform 1 0 36064 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_314
timestamp 1654395037
transform 1 0 36512 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_316
timestamp 1654395037
transform 1 0 36736 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_319
timestamp 1654395037
transform 1 0 37072 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_329
timestamp 1654395037
transform 1 0 38192 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_345
timestamp 1654395037
transform 1 0 39984 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_353
timestamp 1654395037
transform 1 0 40880 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_359
timestamp 1654395037
transform 1 0 41552 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_367
timestamp 1654395037
transform 1 0 42448 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_375
timestamp 1654395037
transform 1 0 43344 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_379
timestamp 1654395037
transform 1 0 43792 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_382
timestamp 1654395037
transform 1 0 44128 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_390
timestamp 1654395037
transform 1 0 45024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_394
timestamp 1654395037
transform 1 0 45472 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_402
timestamp 1654395037
transform 1 0 46368 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_404
timestamp 1654395037
transform 1 0 46592 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_407
timestamp 1654395037
transform 1 0 46928 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_415
timestamp 1654395037
transform 1 0 47824 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_423
timestamp 1654395037
transform 1 0 48720 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_425
timestamp 1654395037
transform 1 0 48944 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_430
timestamp 1654395037
transform 1 0 49504 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_438
timestamp 1654395037
transform 1 0 50400 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_446
timestamp 1654395037
transform 1 0 51296 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_450
timestamp 1654395037
transform 1 0 51744 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_458
timestamp 1654395037
transform 1 0 52640 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_494
timestamp 1654395037
transform 1 0 56672 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_496
timestamp 1654395037
transform 1 0 56896 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_505
timestamp 1654395037
transform 1 0 57904 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_511
timestamp 1654395037
transform 1 0 58576 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_515
timestamp 1654395037
transform 1 0 59024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_519
timestamp 1654395037
transform 1 0 59472 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_527
timestamp 1654395037
transform 1 0 60368 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_531
timestamp 1654395037
transform 1 0 60816 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_539
timestamp 1654395037
transform 1 0 61712 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_543
timestamp 1654395037
transform 1 0 62160 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_553
timestamp 1654395037
transform 1 0 63280 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_557
timestamp 1654395037
transform 1 0 63728 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_565
timestamp 1654395037
transform 1 0 64624 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_567
timestamp 1654395037
transform 1 0 64848 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_572
timestamp 1654395037
transform 1 0 65408 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_588
timestamp 1654395037
transform 1 0 67200 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_596
timestamp 1654395037
transform 1 0 68096 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_600
timestamp 1654395037
transform 1 0 68544 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_603
timestamp 1654395037
transform 1 0 68880 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_607
timestamp 1654395037
transform 1 0 69328 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_609
timestamp 1654395037
transform 1 0 69552 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_616
timestamp 1654395037
transform 1 0 70336 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_620
timestamp 1654395037
transform 1 0 70784 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_622
timestamp 1654395037
transform 1 0 71008 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_625
timestamp 1654395037
transform 1 0 71344 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_629
timestamp 1654395037
transform 1 0 71792 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_632
timestamp 1654395037
transform 1 0 72128 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_636
timestamp 1654395037
transform 1 0 72576 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_638
timestamp 1654395037
transform 1 0 72800 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_643
timestamp 1654395037
transform 1 0 73360 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_647
timestamp 1654395037
transform 1 0 73808 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_654
timestamp 1654395037
transform 1 0 74592 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_658
timestamp 1654395037
transform 1 0 75040 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_666
timestamp 1654395037
transform 1 0 75936 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_670
timestamp 1654395037
transform 1 0 76384 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_672
timestamp 1654395037
transform 1 0 76608 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_675
timestamp 1654395037
transform 1 0 76944 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_679
timestamp 1654395037
transform 1 0 77392 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_681
timestamp 1654395037
transform 1 0 77616 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_684
timestamp 1654395037
transform 1 0 77952 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_688
timestamp 1654395037
transform 1 0 78400 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_692
timestamp 1654395037
transform 1 0 78848 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_700
timestamp 1654395037
transform 1 0 79744 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_708
timestamp 1654395037
transform 1 0 80640 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_718
timestamp 1654395037
transform 1 0 81760 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_726
timestamp 1654395037
transform 1 0 82656 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_734
timestamp 1654395037
transform 1 0 83552 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_738
timestamp 1654395037
transform 1 0 84000 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_742
timestamp 1654395037
transform 1 0 84448 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_746
timestamp 1654395037
transform 1 0 84896 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_758
timestamp 1654395037
transform 1 0 86240 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_762
timestamp 1654395037
transform 1 0 86688 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_764
timestamp 1654395037
transform 1 0 86912 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_767
timestamp 1654395037
transform 1 0 87248 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_773
timestamp 1654395037
transform 1 0 87920 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_779
timestamp 1654395037
transform 1 0 88592 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_785
timestamp 1654395037
transform 1 0 89264 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_791
timestamp 1654395037
transform 1 0 89936 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_799
timestamp 1654395037
transform 1 0 90832 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_805
timestamp 1654395037
transform 1 0 91504 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_809
timestamp 1654395037
transform 1 0 91952 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_813
timestamp 1654395037
transform 1 0 92400 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_821
timestamp 1654395037
transform 1 0 93296 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_829
timestamp 1654395037
transform 1 0 94192 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_833
timestamp 1654395037
transform 1 0 94640 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_837
timestamp 1654395037
transform 1 0 95088 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_841
timestamp 1654395037
transform 1 0 95536 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_849
timestamp 1654395037
transform 1 0 96432 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_851
timestamp 1654395037
transform 1 0 96656 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_854
timestamp 1654395037
transform 1 0 96992 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_858
timestamp 1654395037
transform 1 0 97440 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_875
timestamp 1654395037
transform 1 0 99344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_883
timestamp 1654395037
transform 1 0 100240 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_885
timestamp 1654395037
transform 1 0 100464 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_890
timestamp 1654395037
transform 1 0 101024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_894
timestamp 1654395037
transform 1 0 101472 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_910
timestamp 1654395037
transform 1 0 103264 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_918
timestamp 1654395037
transform 1 0 104160 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_921
timestamp 1654395037
transform 1 0 104496 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_931
timestamp 1654395037
transform 1 0 105616 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_947
timestamp 1654395037
transform 1 0 107408 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_957
timestamp 1654395037
transform 1 0 108528 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_961
timestamp 1654395037
transform 1 0 108976 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_965
timestamp 1654395037
transform 1 0 109424 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_981
timestamp 1654395037
transform 1 0 111216 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_989
timestamp 1654395037
transform 1 0 112112 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_993
timestamp 1654395037
transform 1 0 112560 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_996
timestamp 1654395037
transform 1 0 112896 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_1028
timestamp 1654395037
transform 1 0 116480 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_1048
timestamp 1654395037
transform 1 0 118720 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_1052
timestamp 1654395037
transform 1 0 119168 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_1060
timestamp 1654395037
transform 1 0 120064 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1064
timestamp 1654395037
transform 1 0 120512 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_1067
timestamp 1654395037
transform 1 0 120848 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_1099
timestamp 1654395037
transform 1 0 124432 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_1103
timestamp 1654395037
transform 1 0 124880 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1135
timestamp 1654395037
transform 1 0 128464 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_1138
timestamp 1654395037
transform 1 0 128800 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_1142
timestamp 1654395037
transform 1 0 129248 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1144
timestamp 1654395037
transform 1 0 129472 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_1147
timestamp 1654395037
transform 1 0 129808 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1155
timestamp 1654395037
transform 1 0 130704 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_1158
timestamp 1654395037
transform 1 0 131040 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_1162
timestamp 1654395037
transform 1 0 131488 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_1180
timestamp 1654395037
transform 1 0 133504 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_1198
timestamp 1654395037
transform 1 0 135520 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_1202
timestamp 1654395037
transform 1 0 135968 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1206
timestamp 1654395037
transform 1 0 136416 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_1225
timestamp 1654395037
transform 1 0 138544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_1243
timestamp 1654395037
transform 1 0 140560 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_1251
timestamp 1654395037
transform 1 0 141456 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_1255
timestamp 1654395037
transform 1 0 141904 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1257
timestamp 1654395037
transform 1 0 142128 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_1274
timestamp 1654395037
transform 1 0 144032 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_1280
timestamp 1654395037
transform 1 0 144704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_1298
timestamp 1654395037
transform 1 0 146720 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_1302
timestamp 1654395037
transform 1 0 147168 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_1306
timestamp 1654395037
transform 1 0 147616 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1308
timestamp 1654395037
transform 1 0 147840 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_1325
timestamp 1654395037
transform 1 0 149744 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1329
timestamp 1654395037
transform 1 0 150192 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_1346
timestamp 1654395037
transform 1 0 152096 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1348
timestamp 1654395037
transform 1 0 152320 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1351
timestamp 1654395037
transform 1 0 152656 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_1368
timestamp 1654395037
transform 1 0 154560 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_1386
timestamp 1654395037
transform 1 0 156576 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1390
timestamp 1654395037
transform 1 0 157024 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_1407
timestamp 1654395037
transform 1 0 158928 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_1411
timestamp 1654395037
transform 1 0 159376 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_1415
timestamp 1654395037
transform 1 0 159824 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1419
timestamp 1654395037
transform 1 0 160272 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_1426
timestamp 1654395037
transform 1 0 161056 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_1430
timestamp 1654395037
transform 1 0 161504 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_1434
timestamp 1654395037
transform 1 0 161952 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_1472
timestamp 1654395037
transform 1 0 166208 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_1476
timestamp 1654395037
transform 1 0 166656 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_1480
timestamp 1654395037
transform 1 0 167104 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1484
timestamp 1654395037
transform 1 0 167552 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_1489
timestamp 1654395037
transform 1 0 168112 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_1509
timestamp 1654395037
transform 1 0 170352 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1511
timestamp 1654395037
transform 1 0 170576 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_1516
timestamp 1654395037
transform 1 0 171136 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_1552
timestamp 1654395037
transform 1 0 175168 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_1560
timestamp 1654395037
transform 1 0 176064 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_1570
timestamp 1654395037
transform 1 0 177184 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_1608
timestamp 1654395037
transform 1 0 181440 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_1626
timestamp 1654395037
transform 1 0 183456 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_1630
timestamp 1654395037
transform 1 0 183904 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1632
timestamp 1654395037
transform 1 0 184128 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_1651
timestamp 1654395037
transform 1 0 186256 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_1669
timestamp 1654395037
transform 1 0 188272 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_1687
timestamp 1654395037
transform 1 0 190288 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_1695
timestamp 1654395037
transform 1 0 191184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_1699
timestamp 1654395037
transform 1 0 191632 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1703
timestamp 1654395037
transform 1 0 192080 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_1722
timestamp 1654395037
transform 1 0 194208 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_1730
timestamp 1654395037
transform 1 0 195104 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_1738
timestamp 1654395037
transform 1 0 196000 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_1746
timestamp 1654395037
transform 1 0 196896 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_1754
timestamp 1654395037
transform 1 0 197792 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_1758
timestamp 1654395037
transform 1 0 198240 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_1762
timestamp 1654395037
transform 1 0 198688 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_1766
timestamp 1654395037
transform 1 0 199136 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_1770
timestamp 1654395037
transform 1 0 199584 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1774
timestamp 1654395037
transform 1 0 200032 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_1779
timestamp 1654395037
transform 1 0 200592 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_1783
timestamp 1654395037
transform 1 0 201040 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_1787
timestamp 1654395037
transform 1 0 201488 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_1791
timestamp 1654395037
transform 1 0 201936 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_1795
timestamp 1654395037
transform 1 0 202384 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1797
timestamp 1654395037
transform 1 0 202608 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_1804
timestamp 1654395037
transform 1 0 203392 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_1824
timestamp 1654395037
transform 1 0 205632 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_1844
timestamp 1654395037
transform 1 0 207872 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_1866
timestamp 1654395037
transform 1 0 210336 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_1884
timestamp 1654395037
transform 1 0 212352 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_1892
timestamp 1654395037
transform 1 0 213248 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_1896
timestamp 1654395037
transform 1 0 213696 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_1900
timestamp 1654395037
transform 1 0 214144 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_1904
timestamp 1654395037
transform 1 0 214592 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_1908
timestamp 1654395037
transform 1 0 215040 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_1912
timestamp 1654395037
transform 1 0 215488 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1916
timestamp 1654395037
transform 1 0 215936 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_1921
timestamp 1654395037
transform 1 0 216496 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_1925
timestamp 1654395037
transform 1 0 216944 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_1933
timestamp 1654395037
transform 1 0 217840 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1937
timestamp 1654395037
transform 1 0 218288 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_2
timestamp 1654395037
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_34
timestamp 1654395037
transform 1 0 5152 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_37
timestamp 1654395037
transform 1 0 5488 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_53
timestamp 1654395037
transform 1 0 7280 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_61
timestamp 1654395037
transform 1 0 8176 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_64
timestamp 1654395037
transform 1 0 8512 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_68
timestamp 1654395037
transform 1 0 8960 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_72
timestamp 1654395037
transform 1 0 9408 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_74
timestamp 1654395037
transform 1 0 9632 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_81
timestamp 1654395037
transform 1 0 10416 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_89
timestamp 1654395037
transform 1 0 11312 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_97
timestamp 1654395037
transform 1 0 12208 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_101
timestamp 1654395037
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_107
timestamp 1654395037
transform 1 0 13328 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_139
timestamp 1654395037
transform 1 0 16912 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_142
timestamp 1654395037
transform 1 0 17248 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_174
timestamp 1654395037
transform 1 0 20832 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_177
timestamp 1654395037
transform 1 0 21168 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_185
timestamp 1654395037
transform 1 0 22064 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_187
timestamp 1654395037
transform 1 0 22288 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_190
timestamp 1654395037
transform 1 0 22624 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_206
timestamp 1654395037
transform 1 0 24416 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_214
timestamp 1654395037
transform 1 0 25312 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_230
timestamp 1654395037
transform 1 0 27104 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_238
timestamp 1654395037
transform 1 0 28000 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_242
timestamp 1654395037
transform 1 0 28448 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_244
timestamp 1654395037
transform 1 0 28672 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_247
timestamp 1654395037
transform 1 0 29008 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_279
timestamp 1654395037
transform 1 0 32592 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_282
timestamp 1654395037
transform 1 0 32928 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_314
timestamp 1654395037
transform 1 0 36512 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_317
timestamp 1654395037
transform 1 0 36848 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_349
timestamp 1654395037
transform 1 0 40432 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_352
timestamp 1654395037
transform 1 0 40768 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_360
timestamp 1654395037
transform 1 0 41664 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_364
timestamp 1654395037
transform 1 0 42112 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_366
timestamp 1654395037
transform 1 0 42336 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_369
timestamp 1654395037
transform 1 0 42672 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_373
timestamp 1654395037
transform 1 0 43120 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_377
timestamp 1654395037
transform 1 0 43568 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_381
timestamp 1654395037
transform 1 0 44016 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_387
timestamp 1654395037
transform 1 0 44688 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_389
timestamp 1654395037
transform 1 0 44912 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_396
timestamp 1654395037
transform 1 0 45696 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_400
timestamp 1654395037
transform 1 0 46144 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_404
timestamp 1654395037
transform 1 0 46592 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_406
timestamp 1654395037
transform 1 0 46816 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_409
timestamp 1654395037
transform 1 0 47152 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_413
timestamp 1654395037
transform 1 0 47600 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_417
timestamp 1654395037
transform 1 0 48048 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_419
timestamp 1654395037
transform 1 0 48272 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_422
timestamp 1654395037
transform 1 0 48608 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_425
timestamp 1654395037
transform 1 0 48944 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_433
timestamp 1654395037
transform 1 0 49840 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_437
timestamp 1654395037
transform 1 0 50288 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_440
timestamp 1654395037
transform 1 0 50624 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_448
timestamp 1654395037
transform 1 0 51520 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_452
timestamp 1654395037
transform 1 0 51968 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_454
timestamp 1654395037
transform 1 0 52192 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_457
timestamp 1654395037
transform 1 0 52528 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_460
timestamp 1654395037
transform 1 0 52864 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_464
timestamp 1654395037
transform 1 0 53312 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_467
timestamp 1654395037
transform 1 0 53648 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_485
timestamp 1654395037
transform 1 0 55664 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_489
timestamp 1654395037
transform 1 0 56112 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_494
timestamp 1654395037
transform 1 0 56672 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_498
timestamp 1654395037
transform 1 0 57120 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_502
timestamp 1654395037
transform 1 0 57568 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_504
timestamp 1654395037
transform 1 0 57792 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_507
timestamp 1654395037
transform 1 0 58128 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_523
timestamp 1654395037
transform 1 0 59920 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_527
timestamp 1654395037
transform 1 0 60368 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_559
timestamp 1654395037
transform 1 0 63952 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_562
timestamp 1654395037
transform 1 0 64288 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_594
timestamp 1654395037
transform 1 0 67872 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_597
timestamp 1654395037
transform 1 0 68208 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_613
timestamp 1654395037
transform 1 0 70000 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_623
timestamp 1654395037
transform 1 0 71120 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_627
timestamp 1654395037
transform 1 0 71568 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_629
timestamp 1654395037
transform 1 0 71792 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_632
timestamp 1654395037
transform 1 0 72128 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_664
timestamp 1654395037
transform 1 0 75712 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_673
timestamp 1654395037
transform 1 0 76720 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_675
timestamp 1654395037
transform 1 0 76944 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_682
timestamp 1654395037
transform 1 0 77728 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_686
timestamp 1654395037
transform 1 0 78176 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_689
timestamp 1654395037
transform 1 0 78512 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_697
timestamp 1654395037
transform 1 0 79408 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_699
timestamp 1654395037
transform 1 0 79632 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_704
timestamp 1654395037
transform 1 0 80192 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_712
timestamp 1654395037
transform 1 0 81088 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_720
timestamp 1654395037
transform 1 0 81984 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_728
timestamp 1654395037
transform 1 0 82880 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_732
timestamp 1654395037
transform 1 0 83328 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_734
timestamp 1654395037
transform 1 0 83552 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_739
timestamp 1654395037
transform 1 0 84112 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_747
timestamp 1654395037
transform 1 0 85008 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_751
timestamp 1654395037
transform 1 0 85456 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_753
timestamp 1654395037
transform 1 0 85680 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_756
timestamp 1654395037
transform 1 0 86016 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_764
timestamp 1654395037
transform 1 0 86912 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_768
timestamp 1654395037
transform 1 0 87360 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_772
timestamp 1654395037
transform 1 0 87808 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_804
timestamp 1654395037
transform 1 0 91392 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_807
timestamp 1654395037
transform 1 0 91728 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_839
timestamp 1654395037
transform 1 0 95312 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_842
timestamp 1654395037
transform 1 0 95648 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_846
timestamp 1654395037
transform 1 0 96096 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_862
timestamp 1654395037
transform 1 0 97888 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_870
timestamp 1654395037
transform 1 0 98784 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_873
timestamp 1654395037
transform 1 0 99120 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_879
timestamp 1654395037
transform 1 0 99792 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_883
timestamp 1654395037
transform 1 0 100240 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_899
timestamp 1654395037
transform 1 0 102032 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_903
timestamp 1654395037
transform 1 0 102480 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_905
timestamp 1654395037
transform 1 0 102704 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_908
timestamp 1654395037
transform 1 0 103040 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_918
timestamp 1654395037
transform 1 0 104160 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_934
timestamp 1654395037
transform 1 0 105952 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_938
timestamp 1654395037
transform 1 0 106400 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_940
timestamp 1654395037
transform 1 0 106624 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_943
timestamp 1654395037
transform 1 0 106960 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_947
timestamp 1654395037
transform 1 0 107408 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_955
timestamp 1654395037
transform 1 0 108304 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_963
timestamp 1654395037
transform 1 0 109200 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_971
timestamp 1654395037
transform 1 0 110096 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_975
timestamp 1654395037
transform 1 0 110544 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_978
timestamp 1654395037
transform 1 0 110880 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_988
timestamp 1654395037
transform 1 0 112000 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1004
timestamp 1654395037
transform 1 0 113792 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1008
timestamp 1654395037
transform 1 0 114240 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1010
timestamp 1654395037
transform 1 0 114464 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1013
timestamp 1654395037
transform 1 0 114800 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_1023
timestamp 1654395037
transform 1 0 115920 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_1039
timestamp 1654395037
transform 1 0 117712 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1047
timestamp 1654395037
transform 1 0 118608 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1049
timestamp 1654395037
transform 1 0 118832 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_1052
timestamp 1654395037
transform 1 0 119168 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1060
timestamp 1654395037
transform 1 0 120064 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1062
timestamp 1654395037
transform 1 0 120288 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1065
timestamp 1654395037
transform 1 0 120624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_1073
timestamp 1654395037
transform 1 0 121520 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1081
timestamp 1654395037
transform 1 0 122416 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_1087
timestamp 1654395037
transform 1 0 123088 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1119
timestamp 1654395037
transform 1 0 126672 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_1122
timestamp 1654395037
transform 1 0 127008 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1130
timestamp 1654395037
transform 1 0 127904 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1132
timestamp 1654395037
transform 1 0 128128 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1135
timestamp 1654395037
transform 1 0 128464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1143
timestamp 1654395037
transform 1 0 129360 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1153
timestamp 1654395037
transform 1 0 130480 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1157
timestamp 1654395037
transform 1 0 130928 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1164
timestamp 1654395037
transform 1 0 131712 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1182
timestamp 1654395037
transform 1 0 133728 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1186
timestamp 1654395037
transform 1 0 134176 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1208
timestamp 1654395037
transform 1 0 136640 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1216
timestamp 1654395037
transform 1 0 137536 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1220
timestamp 1654395037
transform 1 0 137984 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1224
timestamp 1654395037
transform 1 0 138432 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1233
timestamp 1654395037
transform 1 0 139440 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1251
timestamp 1654395037
transform 1 0 141456 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1255
timestamp 1654395037
transform 1 0 141904 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1259
timestamp 1654395037
transform 1 0 142352 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1268
timestamp 1654395037
transform 1 0 143360 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1276
timestamp 1654395037
transform 1 0 144256 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1280
timestamp 1654395037
transform 1 0 144704 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1284
timestamp 1654395037
transform 1 0 145152 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1288
timestamp 1654395037
transform 1 0 145600 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1292
timestamp 1654395037
transform 1 0 146048 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1294
timestamp 1654395037
transform 1 0 146272 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1303
timestamp 1654395037
transform 1 0 147280 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1307
timestamp 1654395037
transform 1 0 147728 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1311
timestamp 1654395037
transform 1 0 148176 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1315
timestamp 1654395037
transform 1 0 148624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1319
timestamp 1654395037
transform 1 0 149072 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1323
timestamp 1654395037
transform 1 0 149520 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1327
timestamp 1654395037
transform 1 0 149968 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1329
timestamp 1654395037
transform 1 0 150192 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1338
timestamp 1654395037
transform 1 0 151200 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1342
timestamp 1654395037
transform 1 0 151648 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1348
timestamp 1654395037
transform 1 0 152320 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1352
timestamp 1654395037
transform 1 0 152768 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1356
timestamp 1654395037
transform 1 0 153216 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1360
timestamp 1654395037
transform 1 0 153664 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1364
timestamp 1654395037
transform 1 0 154112 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1373
timestamp 1654395037
transform 1 0 155120 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1377
timestamp 1654395037
transform 1 0 155568 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1381
timestamp 1654395037
transform 1 0 156016 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1398
timestamp 1654395037
transform 1 0 157920 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1408
timestamp 1654395037
transform 1 0 159040 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1426
timestamp 1654395037
transform 1 0 161056 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1430
timestamp 1654395037
transform 1 0 161504 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1434
timestamp 1654395037
transform 1 0 161952 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1453
timestamp 1654395037
transform 1 0 164080 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1457
timestamp 1654395037
transform 1 0 164528 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1461
timestamp 1654395037
transform 1 0 164976 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1468
timestamp 1654395037
transform 1 0 165760 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1472
timestamp 1654395037
transform 1 0 166208 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1492
timestamp 1654395037
transform 1 0 168448 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1496
timestamp 1654395037
transform 1 0 168896 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1500
timestamp 1654395037
transform 1 0 169344 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1504
timestamp 1654395037
transform 1 0 169792 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1523
timestamp 1654395037
transform 1 0 171920 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1533
timestamp 1654395037
transform 1 0 173040 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1537
timestamp 1654395037
transform 1 0 173488 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1539
timestamp 1654395037
transform 1 0 173712 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1544
timestamp 1654395037
transform 1 0 174272 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1546
timestamp 1654395037
transform 1 0 174496 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1565
timestamp 1654395037
transform 1 0 176624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1573
timestamp 1654395037
transform 1 0 177520 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1593
timestamp 1654395037
transform 1 0 179760 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1601
timestamp 1654395037
transform 1 0 180656 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1607
timestamp 1654395037
transform 1 0 181328 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1609
timestamp 1654395037
transform 1 0 181552 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1628
timestamp 1654395037
transform 1 0 183680 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1636
timestamp 1654395037
transform 1 0 184576 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1642
timestamp 1654395037
transform 1 0 185248 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1644
timestamp 1654395037
transform 1 0 185472 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1663
timestamp 1654395037
transform 1 0 187600 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1671
timestamp 1654395037
transform 1 0 188496 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1675
timestamp 1654395037
transform 1 0 188944 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1679
timestamp 1654395037
transform 1 0 189392 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1698
timestamp 1654395037
transform 1 0 191520 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1706
timestamp 1654395037
transform 1 0 192416 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1710
timestamp 1654395037
transform 1 0 192864 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1714
timestamp 1654395037
transform 1 0 193312 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1723
timestamp 1654395037
transform 1 0 194320 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1731
timestamp 1654395037
transform 1 0 195216 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1739
timestamp 1654395037
transform 1 0 196112 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1747
timestamp 1654395037
transform 1 0 197008 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1749
timestamp 1654395037
transform 1 0 197232 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1758
timestamp 1654395037
transform 1 0 198240 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1762
timestamp 1654395037
transform 1 0 198688 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1770
timestamp 1654395037
transform 1 0 199584 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1774
timestamp 1654395037
transform 1 0 200032 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1778
timestamp 1654395037
transform 1 0 200480 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1782
timestamp 1654395037
transform 1 0 200928 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1784
timestamp 1654395037
transform 1 0 201152 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1793
timestamp 1654395037
transform 1 0 202160 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1797
timestamp 1654395037
transform 1 0 202608 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1801
timestamp 1654395037
transform 1 0 203056 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1805
timestamp 1654395037
transform 1 0 203504 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1809
timestamp 1654395037
transform 1 0 203952 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1811
timestamp 1654395037
transform 1 0 204176 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1818
timestamp 1654395037
transform 1 0 204960 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1822
timestamp 1654395037
transform 1 0 205408 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1830
timestamp 1654395037
transform 1 0 206304 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1834
timestamp 1654395037
transform 1 0 206752 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1853
timestamp 1654395037
transform 1 0 208880 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1873
timestamp 1654395037
transform 1 0 211120 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1881
timestamp 1654395037
transform 1 0 212016 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1885
timestamp 1654395037
transform 1 0 212464 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1889
timestamp 1654395037
transform 1 0 212912 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1898
timestamp 1654395037
transform 1 0 213920 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1902
timestamp 1654395037
transform 1 0 214368 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1906
timestamp 1654395037
transform 1 0 214816 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1910
timestamp 1654395037
transform 1 0 215264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1914
timestamp 1654395037
transform 1 0 215712 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1918
timestamp 1654395037
transform 1 0 216160 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_1922
timestamp 1654395037
transform 1 0 216608 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1924
timestamp 1654395037
transform 1 0 216832 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_1929
timestamp 1654395037
transform 1 0 217392 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1937
timestamp 1654395037
transform 1 0 218288 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_0 pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_1
timestamp 1654395037
transform -1 0 218624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_2
timestamp 1654395037
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_3
timestamp 1654395037
transform -1 0 218624 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_4
timestamp 1654395037
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_5
timestamp 1654395037
transform -1 0 218624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_6
timestamp 1654395037
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_7
timestamp 1654395037
transform -1 0 218624 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_8
timestamp 1654395037
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_9
timestamp 1654395037
transform -1 0 218624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_10
timestamp 1654395037
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_11
timestamp 1654395037
transform -1 0 218624 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_12
timestamp 1654395037
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_13
timestamp 1654395037
transform -1 0 218624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_14
timestamp 1654395037
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_15
timestamp 1654395037
transform 1 0 9184 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_16
timestamp 1654395037
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_17
timestamp 1654395037
transform 1 0 17024 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_18
timestamp 1654395037
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_19
timestamp 1654395037
transform 1 0 24864 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_20
timestamp 1654395037
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_21
timestamp 1654395037
transform 1 0 32704 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_22
timestamp 1654395037
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_23
timestamp 1654395037
transform 1 0 40544 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_24
timestamp 1654395037
transform 1 0 44464 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_25
timestamp 1654395037
transform 1 0 48384 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_26
timestamp 1654395037
transform 1 0 52304 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_27
timestamp 1654395037
transform 1 0 56224 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_28
timestamp 1654395037
transform 1 0 60144 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_29
timestamp 1654395037
transform 1 0 64064 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_30
timestamp 1654395037
transform 1 0 67984 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_31
timestamp 1654395037
transform 1 0 71904 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_32
timestamp 1654395037
transform 1 0 75824 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_33
timestamp 1654395037
transform 1 0 79744 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_34
timestamp 1654395037
transform 1 0 83664 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_35
timestamp 1654395037
transform 1 0 87584 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_36
timestamp 1654395037
transform 1 0 91504 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_37
timestamp 1654395037
transform 1 0 95424 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_38
timestamp 1654395037
transform 1 0 99344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_39
timestamp 1654395037
transform 1 0 103264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_40
timestamp 1654395037
transform 1 0 107184 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_41
timestamp 1654395037
transform 1 0 111104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_42
timestamp 1654395037
transform 1 0 115024 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_43
timestamp 1654395037
transform 1 0 118944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_44
timestamp 1654395037
transform 1 0 122864 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_45
timestamp 1654395037
transform 1 0 126784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_46
timestamp 1654395037
transform 1 0 130704 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_47
timestamp 1654395037
transform 1 0 134624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_48
timestamp 1654395037
transform 1 0 138544 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_49
timestamp 1654395037
transform 1 0 142464 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_50
timestamp 1654395037
transform 1 0 146384 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_51
timestamp 1654395037
transform 1 0 150304 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_52
timestamp 1654395037
transform 1 0 154224 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_53
timestamp 1654395037
transform 1 0 158144 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_54
timestamp 1654395037
transform 1 0 162064 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_55
timestamp 1654395037
transform 1 0 165984 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_56
timestamp 1654395037
transform 1 0 169904 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_57
timestamp 1654395037
transform 1 0 173824 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_58
timestamp 1654395037
transform 1 0 177744 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_59
timestamp 1654395037
transform 1 0 181664 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_60
timestamp 1654395037
transform 1 0 185584 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_61
timestamp 1654395037
transform 1 0 189504 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_62
timestamp 1654395037
transform 1 0 193424 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_63
timestamp 1654395037
transform 1 0 197344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_64
timestamp 1654395037
transform 1 0 201264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_65
timestamp 1654395037
transform 1 0 205184 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_66
timestamp 1654395037
transform 1 0 209104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_67
timestamp 1654395037
transform 1 0 213024 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_68
timestamp 1654395037
transform 1 0 216944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_69
timestamp 1654395037
transform 1 0 9296 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_70
timestamp 1654395037
transform 1 0 17248 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_71
timestamp 1654395037
transform 1 0 25200 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_72
timestamp 1654395037
transform 1 0 33152 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_73
timestamp 1654395037
transform 1 0 41104 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_74
timestamp 1654395037
transform 1 0 49056 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_75
timestamp 1654395037
transform 1 0 57008 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_76
timestamp 1654395037
transform 1 0 64960 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_77
timestamp 1654395037
transform 1 0 72912 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_78
timestamp 1654395037
transform 1 0 80864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_79
timestamp 1654395037
transform 1 0 88816 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_80
timestamp 1654395037
transform 1 0 96768 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_81
timestamp 1654395037
transform 1 0 104720 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_82
timestamp 1654395037
transform 1 0 112672 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_83
timestamp 1654395037
transform 1 0 120624 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_84
timestamp 1654395037
transform 1 0 128576 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_85
timestamp 1654395037
transform 1 0 136528 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_86
timestamp 1654395037
transform 1 0 144480 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_87
timestamp 1654395037
transform 1 0 152432 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_88
timestamp 1654395037
transform 1 0 160384 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_89
timestamp 1654395037
transform 1 0 168336 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_90
timestamp 1654395037
transform 1 0 176288 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_91
timestamp 1654395037
transform 1 0 184240 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_92
timestamp 1654395037
transform 1 0 192192 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_93
timestamp 1654395037
transform 1 0 200144 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_94
timestamp 1654395037
transform 1 0 208096 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_95
timestamp 1654395037
transform 1 0 216048 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_96
timestamp 1654395037
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_97
timestamp 1654395037
transform 1 0 13216 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_98
timestamp 1654395037
transform 1 0 21168 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_99
timestamp 1654395037
transform 1 0 29120 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_100
timestamp 1654395037
transform 1 0 37072 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_101
timestamp 1654395037
transform 1 0 45024 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_102
timestamp 1654395037
transform 1 0 52976 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_103
timestamp 1654395037
transform 1 0 60928 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_104
timestamp 1654395037
transform 1 0 68880 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_105
timestamp 1654395037
transform 1 0 76832 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_106
timestamp 1654395037
transform 1 0 84784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_107
timestamp 1654395037
transform 1 0 92736 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_108
timestamp 1654395037
transform 1 0 100688 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_109
timestamp 1654395037
transform 1 0 108640 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_110
timestamp 1654395037
transform 1 0 116592 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_111
timestamp 1654395037
transform 1 0 124544 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_112
timestamp 1654395037
transform 1 0 132496 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_113
timestamp 1654395037
transform 1 0 140448 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_114
timestamp 1654395037
transform 1 0 148400 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_115
timestamp 1654395037
transform 1 0 156352 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_116
timestamp 1654395037
transform 1 0 164304 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_117
timestamp 1654395037
transform 1 0 172256 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_118
timestamp 1654395037
transform 1 0 180208 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_119
timestamp 1654395037
transform 1 0 188160 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_120
timestamp 1654395037
transform 1 0 196112 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_121
timestamp 1654395037
transform 1 0 204064 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_122
timestamp 1654395037
transform 1 0 212016 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_123
timestamp 1654395037
transform 1 0 9296 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_124
timestamp 1654395037
transform 1 0 17248 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_125
timestamp 1654395037
transform 1 0 25200 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_126
timestamp 1654395037
transform 1 0 33152 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_127
timestamp 1654395037
transform 1 0 41104 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_128
timestamp 1654395037
transform 1 0 49056 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_129
timestamp 1654395037
transform 1 0 57008 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_130
timestamp 1654395037
transform 1 0 64960 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_131
timestamp 1654395037
transform 1 0 72912 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_132
timestamp 1654395037
transform 1 0 80864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_133
timestamp 1654395037
transform 1 0 88816 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_134
timestamp 1654395037
transform 1 0 96768 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_135
timestamp 1654395037
transform 1 0 104720 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_136
timestamp 1654395037
transform 1 0 112672 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_137
timestamp 1654395037
transform 1 0 120624 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_138
timestamp 1654395037
transform 1 0 128576 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_139
timestamp 1654395037
transform 1 0 136528 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_140
timestamp 1654395037
transform 1 0 144480 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_141
timestamp 1654395037
transform 1 0 152432 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_142
timestamp 1654395037
transform 1 0 160384 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_143
timestamp 1654395037
transform 1 0 168336 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_144
timestamp 1654395037
transform 1 0 176288 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_145
timestamp 1654395037
transform 1 0 184240 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_146
timestamp 1654395037
transform 1 0 192192 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_147
timestamp 1654395037
transform 1 0 200144 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_148
timestamp 1654395037
transform 1 0 208096 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_149
timestamp 1654395037
transform 1 0 216048 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_150
timestamp 1654395037
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_151
timestamp 1654395037
transform 1 0 13216 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_152
timestamp 1654395037
transform 1 0 21168 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_153
timestamp 1654395037
transform 1 0 29120 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_154
timestamp 1654395037
transform 1 0 37072 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_155
timestamp 1654395037
transform 1 0 45024 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_156
timestamp 1654395037
transform 1 0 52976 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_157
timestamp 1654395037
transform 1 0 60928 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_158
timestamp 1654395037
transform 1 0 68880 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_159
timestamp 1654395037
transform 1 0 76832 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_160
timestamp 1654395037
transform 1 0 84784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_161
timestamp 1654395037
transform 1 0 92736 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_162
timestamp 1654395037
transform 1 0 100688 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_163
timestamp 1654395037
transform 1 0 108640 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_164
timestamp 1654395037
transform 1 0 116592 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_165
timestamp 1654395037
transform 1 0 124544 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_166
timestamp 1654395037
transform 1 0 132496 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_167
timestamp 1654395037
transform 1 0 140448 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_168
timestamp 1654395037
transform 1 0 148400 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_169
timestamp 1654395037
transform 1 0 156352 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_170
timestamp 1654395037
transform 1 0 164304 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_171
timestamp 1654395037
transform 1 0 172256 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_172
timestamp 1654395037
transform 1 0 180208 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_173
timestamp 1654395037
transform 1 0 188160 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_174
timestamp 1654395037
transform 1 0 196112 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_175
timestamp 1654395037
transform 1 0 204064 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_176
timestamp 1654395037
transform 1 0 212016 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_177
timestamp 1654395037
transform 1 0 9296 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_178
timestamp 1654395037
transform 1 0 17248 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_179
timestamp 1654395037
transform 1 0 25200 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_180
timestamp 1654395037
transform 1 0 33152 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_181
timestamp 1654395037
transform 1 0 41104 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_182
timestamp 1654395037
transform 1 0 49056 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_183
timestamp 1654395037
transform 1 0 57008 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_184
timestamp 1654395037
transform 1 0 64960 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_185
timestamp 1654395037
transform 1 0 72912 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_186
timestamp 1654395037
transform 1 0 80864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_187
timestamp 1654395037
transform 1 0 88816 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_188
timestamp 1654395037
transform 1 0 96768 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_189
timestamp 1654395037
transform 1 0 104720 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_190
timestamp 1654395037
transform 1 0 112672 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_191
timestamp 1654395037
transform 1 0 120624 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_192
timestamp 1654395037
transform 1 0 128576 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_193
timestamp 1654395037
transform 1 0 136528 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_194
timestamp 1654395037
transform 1 0 144480 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_195
timestamp 1654395037
transform 1 0 152432 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_196
timestamp 1654395037
transform 1 0 160384 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_197
timestamp 1654395037
transform 1 0 168336 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_198
timestamp 1654395037
transform 1 0 176288 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_199
timestamp 1654395037
transform 1 0 184240 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_200
timestamp 1654395037
transform 1 0 192192 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_201
timestamp 1654395037
transform 1 0 200144 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_202
timestamp 1654395037
transform 1 0 208096 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_203
timestamp 1654395037
transform 1 0 216048 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_204
timestamp 1654395037
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_205
timestamp 1654395037
transform 1 0 9184 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_206
timestamp 1654395037
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_207
timestamp 1654395037
transform 1 0 17024 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_208
timestamp 1654395037
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_209
timestamp 1654395037
transform 1 0 24864 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_210
timestamp 1654395037
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_211
timestamp 1654395037
transform 1 0 32704 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_212
timestamp 1654395037
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_213
timestamp 1654395037
transform 1 0 40544 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_214
timestamp 1654395037
transform 1 0 44464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_215
timestamp 1654395037
transform 1 0 48384 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_216
timestamp 1654395037
transform 1 0 52304 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_217
timestamp 1654395037
transform 1 0 56224 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_218
timestamp 1654395037
transform 1 0 60144 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_219
timestamp 1654395037
transform 1 0 64064 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_220
timestamp 1654395037
transform 1 0 67984 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_221
timestamp 1654395037
transform 1 0 71904 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_222
timestamp 1654395037
transform 1 0 75824 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_223
timestamp 1654395037
transform 1 0 79744 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_224
timestamp 1654395037
transform 1 0 83664 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_225
timestamp 1654395037
transform 1 0 87584 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_226
timestamp 1654395037
transform 1 0 91504 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_227
timestamp 1654395037
transform 1 0 95424 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_228
timestamp 1654395037
transform 1 0 99344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_229
timestamp 1654395037
transform 1 0 103264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_230
timestamp 1654395037
transform 1 0 107184 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_231
timestamp 1654395037
transform 1 0 111104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_232
timestamp 1654395037
transform 1 0 115024 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_233
timestamp 1654395037
transform 1 0 118944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_234
timestamp 1654395037
transform 1 0 122864 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_235
timestamp 1654395037
transform 1 0 126784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_236
timestamp 1654395037
transform 1 0 130704 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_237
timestamp 1654395037
transform 1 0 134624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_238
timestamp 1654395037
transform 1 0 138544 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_239
timestamp 1654395037
transform 1 0 142464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_240
timestamp 1654395037
transform 1 0 146384 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_241
timestamp 1654395037
transform 1 0 150304 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_242
timestamp 1654395037
transform 1 0 154224 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_243
timestamp 1654395037
transform 1 0 158144 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_244
timestamp 1654395037
transform 1 0 162064 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_245
timestamp 1654395037
transform 1 0 165984 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_246
timestamp 1654395037
transform 1 0 169904 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_247
timestamp 1654395037
transform 1 0 173824 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_248
timestamp 1654395037
transform 1 0 177744 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_249
timestamp 1654395037
transform 1 0 181664 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_250
timestamp 1654395037
transform 1 0 185584 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_251
timestamp 1654395037
transform 1 0 189504 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_252
timestamp 1654395037
transform 1 0 193424 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_253
timestamp 1654395037
transform 1 0 197344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_254
timestamp 1654395037
transform 1 0 201264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_255
timestamp 1654395037
transform 1 0 205184 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_256
timestamp 1654395037
transform 1 0 209104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_257
timestamp 1654395037
transform 1 0 213024 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_258
timestamp 1654395037
transform 1 0 216944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _000_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform -1 0 88032 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _001_
timestamp 1654395037
transform -1 0 88704 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _002_
timestamp 1654395037
transform -1 0 88592 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _003_
timestamp 1654395037
transform -1 0 91504 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _004_
timestamp 1654395037
transform -1 0 90720 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _005_
timestamp 1654395037
transform -1 0 79632 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _006_
timestamp 1654395037
transform -1 0 91392 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _007_
timestamp 1654395037
transform -1 0 101024 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _008_
timestamp 1654395037
transform -1 0 110656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _009_
timestamp 1654395037
transform -1 0 118720 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _010_
timestamp 1654395037
transform -1 0 123536 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _011_
timestamp 1654395037
transform -1 0 127008 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _012_
timestamp 1654395037
transform -1 0 130704 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _013_
timestamp 1654395037
transform -1 0 136304 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _014_
timestamp 1654395037
transform 1 0 143472 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _015_
timestamp 1654395037
transform -1 0 152096 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _016_
timestamp 1654395037
transform -1 0 161056 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _017_
timestamp 1654395037
transform -1 0 164080 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _018_
timestamp 1654395037
transform -1 0 168112 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _019_
timestamp 1654395037
transform -1 0 171136 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _020_
timestamp 1654395037
transform -1 0 180992 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _021_
timestamp 1654395037
transform -1 0 181328 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _022_
timestamp 1654395037
transform -1 0 185248 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _023_
timestamp 1654395037
transform -1 0 190848 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _024_
timestamp 1654395037
transform -1 0 189168 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _025_
timestamp 1654395037
transform -1 0 191520 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _026_
timestamp 1654395037
transform -1 0 191184 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _027_
timestamp 1654395037
transform -1 0 184016 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _028_
timestamp 1654395037
transform -1 0 187824 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _029_
timestamp 1654395037
transform -1 0 191968 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _030_
timestamp 1654395037
transform -1 0 194544 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _031_
timestamp 1654395037
transform -1 0 194096 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _032_
timestamp 1654395037
transform 1 0 194880 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _033_
timestamp 1654395037
transform -1 0 203392 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _034_
timestamp 1654395037
transform 1 0 204512 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _035_
timestamp 1654395037
transform -1 0 208768 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _036_
timestamp 1654395037
transform 1 0 211232 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _037_
timestamp 1654395037
transform 1 0 207648 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _038_
timestamp 1654395037
transform -1 0 211008 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _039_
timestamp 1654395037
transform -1 0 60144 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _040_
timestamp 1654395037
transform -1 0 57680 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _041_
timestamp 1654395037
transform -1 0 58352 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _042_
timestamp 1654395037
transform -1 0 50736 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _043_
timestamp 1654395037
transform -1 0 58576 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _044_
timestamp 1654395037
transform -1 0 68656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _045_
timestamp 1654395037
transform -1 0 68656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _046_
timestamp 1654395037
transform -1 0 69664 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _047_
timestamp 1654395037
transform -1 0 69552 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _048_
timestamp 1654395037
transform -1 0 70224 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _049_
timestamp 1654395037
transform -1 0 70896 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _050_
timestamp 1654395037
transform -1 0 70336 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _051_
timestamp 1654395037
transform -1 0 71568 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _052_
timestamp 1654395037
transform -1 0 72240 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _053_
timestamp 1654395037
transform -1 0 73584 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _054_
timestamp 1654395037
transform -1 0 76048 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _055_
timestamp 1654395037
transform -1 0 74592 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _056_
timestamp 1654395037
transform 1 0 74928 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _057_
timestamp 1654395037
transform 1 0 77056 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _058_
timestamp 1654395037
transform 1 0 82768 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _059_
timestamp 1654395037
transform 1 0 85008 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _060_
timestamp 1654395037
transform 1 0 90608 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _061_
timestamp 1654395037
transform -1 0 79744 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _062_
timestamp 1654395037
transform -1 0 86016 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _063_
timestamp 1654395037
transform -1 0 86240 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _064_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 76048 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _065_
timestamp 1654395037
transform 1 0 77056 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _066_
timestamp 1654395037
transform 1 0 78736 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _067_
timestamp 1654395037
transform 1 0 79968 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _068_
timestamp 1654395037
transform 1 0 82208 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _069_
timestamp 1654395037
transform 1 0 80416 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _070_
timestamp 1654395037
transform 1 0 81088 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _071_
timestamp 1654395037
transform 1 0 86240 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _072_
timestamp 1654395037
transform 1 0 81312 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _073_
timestamp 1654395037
transform 1 0 79968 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _074_
timestamp 1654395037
transform 1 0 79072 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _075_
timestamp 1654395037
transform 1 0 79856 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _076_
timestamp 1654395037
transform 1 0 82880 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _077_
timestamp 1654395037
transform 1 0 81984 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _078_
timestamp 1654395037
transform 1 0 86352 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _079_
timestamp 1654395037
transform 1 0 89376 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _080_
timestamp 1654395037
transform 1 0 90160 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _081_
timestamp 1654395037
transform 1 0 92624 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _082_
timestamp 1654395037
transform 1 0 95760 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _083_
timestamp 1654395037
transform 1 0 99568 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _084_
timestamp 1654395037
transform 1 0 103488 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _085_
timestamp 1654395037
transform 1 0 104944 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _086_
timestamp 1654395037
transform 1 0 109424 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _087_
timestamp 1654395037
transform 1 0 107632 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _088_
timestamp 1654395037
transform 1 0 108528 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _089_
timestamp 1654395037
transform 1 0 111328 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _090_
timestamp 1654395037
transform 1 0 115248 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _091_
timestamp 1654395037
transform 1 0 120848 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _092_
timestamp 1654395037
transform 1 0 128688 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _093_
timestamp 1654395037
transform 1 0 140784 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _094_
timestamp 1654395037
transform 1 0 129808 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _095_
timestamp 1654395037
transform 1 0 131040 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _096_
timestamp 1654395037
transform 1 0 133056 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _097_
timestamp 1654395037
transform 1 0 136864 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _098_
timestamp 1654395037
transform 1 0 138768 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _099_
timestamp 1654395037
transform 1 0 142688 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _100_
timestamp 1654395037
transform 1 0 143584 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _101_
timestamp 1654395037
transform 1 0 146608 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _102_
timestamp 1654395037
transform 1 0 150528 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _103_
timestamp 1654395037
transform 1 0 154448 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _104_
timestamp 1654395037
transform 1 0 158368 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _105_
timestamp 1654395037
transform 1 0 165088 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _106_
timestamp 1654395037
transform -1 0 173040 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _107_
timestamp 1654395037
transform -1 0 177520 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _108_
timestamp 1654395037
transform -1 0 180656 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _109_
timestamp 1654395037
transform -1 0 184576 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _110_
timestamp 1654395037
transform -1 0 191184 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _111_
timestamp 1654395037
transform -1 0 192416 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _112_
timestamp 1654395037
transform -1 0 188496 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _113_
timestamp 1654395037
transform -1 0 191072 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _114_
timestamp 1654395037
transform 1 0 187824 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _115_
timestamp 1654395037
transform -1 0 191184 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _116_
timestamp 1654395037
transform -1 0 194320 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _117_
timestamp 1654395037
transform 1 0 194544 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _118_
timestamp 1654395037
transform 1 0 195440 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _119_
timestamp 1654395037
transform 1 0 197568 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _120_
timestamp 1654395037
transform 1 0 198912 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _121_
timestamp 1654395037
transform 1 0 201488 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _122_
timestamp 1654395037
transform 1 0 202720 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _123_
timestamp 1654395037
transform 1 0 205632 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _124_
timestamp 1654395037
transform 1 0 204288 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _125_
timestamp 1654395037
transform 1 0 211344 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _126_
timestamp 1654395037
transform 1 0 210336 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _127_
timestamp 1654395037
transform 1 0 213248 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _128_
timestamp 1654395037
transform -1 0 173152 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _129_
timestamp 1654395037
transform -1 0 175504 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _130_
timestamp 1654395037
transform -1 0 173264 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _131_
timestamp 1654395037
transform -1 0 175728 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _132_
timestamp 1654395037
transform -1 0 176064 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _133_
timestamp 1654395037
transform -1 0 177184 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _134_
timestamp 1654395037
transform -1 0 176960 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _135_
timestamp 1654395037
transform -1 0 179424 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _136_
timestamp 1654395037
transform -1 0 180880 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _137_
timestamp 1654395037
transform -1 0 183456 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _138_
timestamp 1654395037
transform -1 0 187152 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _139_
timestamp 1654395037
transform -1 0 187712 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _140_
timestamp 1654395037
transform -1 0 184800 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _141_
timestamp 1654395037
transform 1 0 34720 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _142_
timestamp 1654395037
transform 1 0 37296 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _143_
timestamp 1654395037
transform 1 0 39424 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _144_
timestamp 1654395037
transform 1 0 41440 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _145_
timestamp 1654395037
transform 1 0 43232 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _146_
timestamp 1654395037
transform 1 0 45360 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _147_
timestamp 1654395037
transform 1 0 47152 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _148_
timestamp 1654395037
transform 1 0 48048 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _149_
timestamp 1654395037
transform 1 0 42560 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _150_
timestamp 1654395037
transform 1 0 41664 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _151_
timestamp 1654395037
transform 1 0 43456 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _152_
timestamp 1654395037
transform 1 0 45696 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _153_
timestamp 1654395037
transform 1 0 48048 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _154_
timestamp 1654395037
transform 1 0 50624 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _155_
timestamp 1654395037
transform 1 0 53872 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _156_
timestamp 1654395037
transform 1 0 58800 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _157_
timestamp 1654395037
transform 1 0 62608 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _158_
timestamp 1654395037
transform 1 0 66864 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _159_
timestamp 1654395037
transform 1 0 71232 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _160_
timestamp 1654395037
transform -1 0 10304 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _161_
timestamp 1654395037
transform -1 0 195104 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _162_
timestamp 1654395037
transform -1 0 196000 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _163_
timestamp 1654395037
transform -1 0 196896 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _164_
timestamp 1654395037
transform -1 0 197008 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _165_
timestamp 1654395037
transform -1 0 197792 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _166_
timestamp 1654395037
transform 1 0 17584 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _167_
timestamp 1654395037
transform 1 0 19712 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _168_
timestamp 1654395037
transform 1 0 21728 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _169_
timestamp 1654395037
transform 1 0 25424 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _170_
timestamp 1654395037
transform 1 0 26432 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _171_
timestamp 1654395037
transform 1 0 29344 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _172_
timestamp 1654395037
transform 1 0 31360 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _173_
timestamp 1654395037
transform 1 0 33824 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _174_
timestamp 1654395037
transform 1 0 36176 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _175_
timestamp 1654395037
transform 1 0 38528 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _176_
timestamp 1654395037
transform 1 0 40544 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _177_
timestamp 1654395037
transform 1 0 42336 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _178_
timestamp 1654395037
transform 1 0 44128 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _179_
timestamp 1654395037
transform 1 0 46256 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _180_
timestamp 1654395037
transform 1 0 49280 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _181_
timestamp 1654395037
transform 1 0 44352 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _182_
timestamp 1654395037
transform 1 0 41776 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _183_
timestamp 1654395037
transform 1 0 42672 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _184_
timestamp 1654395037
transform 1 0 45024 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _185_
timestamp 1654395037
transform 1 0 47152 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _186_
timestamp 1654395037
transform 1 0 49728 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _187_
timestamp 1654395037
transform 1 0 51968 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _188_
timestamp 1654395037
transform 1 0 57232 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _189_
timestamp 1654395037
transform 1 0 61040 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _190_
timestamp 1654395037
transform 1 0 65520 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _191_
timestamp 1654395037
transform 1 0 69664 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _192_
timestamp 1654395037
transform 1 0 73920 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _193_
timestamp 1654395037
transform -1 0 167552 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _194_
timestamp 1654395037
transform -1 0 168112 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _195_
timestamp 1654395037
transform -1 0 169232 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _196_
timestamp 1654395037
transform -1 0 171920 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _197_
timestamp 1654395037
transform -1 0 10416 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _198_
timestamp 1654395037
transform -1 0 12208 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _199_
timestamp 1654395037
transform -1 0 11200 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _200_
timestamp 1654395037
transform 1 0 212576 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _201_
timestamp 1654395037
transform -1 0 11312 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  la_buf\[0\] pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform -1 0 18368 0 1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  la_buf\[1\]
timestamp 1654395037
transform -1 0 18480 0 1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  la_buf\[2\]
timestamp 1654395037
transform -1 0 17024 0 -1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  la_buf\[3\]
timestamp 1654395037
transform -1 0 17024 0 -1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  la_buf\[4\]
timestamp 1654395037
transform -1 0 12992 0 1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  la_buf\[5\]
timestamp 1654395037
transform -1 0 12992 0 1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  la_buf\[6\]
timestamp 1654395037
transform -1 0 9072 0 -1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  la_buf\[7\]
timestamp 1654395037
transform -1 0 15232 0 -1 9408
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  la_buf\[8\]
timestamp 1654395037
transform -1 0 24192 0 -1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  la_buf\[9\]
timestamp 1654395037
transform -1 0 29792 0 -1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  la_buf\[10\]
timestamp 1654395037
transform -1 0 34832 0 1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  la_buf\[11\]
timestamp 1654395037
transform -1 0 38976 0 -1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  la_buf\[12\]
timestamp 1654395037
transform -1 0 43568 0 1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  la_buf\[13\]
timestamp 1654395037
transform -1 0 48832 0 -1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  la_buf\[14\]
timestamp 1654395037
transform -1 0 56336 0 -1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  la_buf\[15\]
timestamp 1654395037
transform -1 0 65968 0 1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  la_buf\[16\]
timestamp 1654395037
transform -1 0 74368 0 1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  la_buf\[17\]
timestamp 1654395037
transform 1 0 78736 0 1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  la_buf\[18\]
timestamp 1654395037
transform 1 0 86576 0 1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  la_buf\[19\]
timestamp 1654395037
transform 1 0 92736 0 -1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  la_buf\[20\]
timestamp 1654395037
transform 1 0 98000 0 -1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  la_buf\[21\]
timestamp 1654395037
transform 1 0 102032 0 1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  la_buf\[22\]
timestamp 1654395037
transform -1 0 25200 0 1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  la_buf\[23\]
timestamp 1654395037
transform -1 0 57008 0 1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  la_buf\[24\]
timestamp 1654395037
transform -1 0 56784 0 -1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  la_buf\[25\]
timestamp 1654395037
transform -1 0 56672 0 -1 9408
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  la_buf\[26\]
timestamp 1654395037
transform -1 0 58576 0 1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  la_buf\[27\]
timestamp 1654395037
transform -1 0 65072 0 1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  la_buf\[28\]
timestamp 1654395037
transform -1 0 76608 0 1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  la_buf\[29\]
timestamp 1654395037
transform -1 0 72688 0 -1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  la_buf\[30\]
timestamp 1654395037
transform -1 0 52752 0 1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  la_buf\[31\]
timestamp 1654395037
transform -1 0 84560 0 1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  la_buf\[32\]
timestamp 1654395037
transform -1 0 100464 0 1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  la_buf\[33\]
timestamp 1654395037
transform 1 0 107632 0 -1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  la_buf\[34\]
timestamp 1654395037
transform 1 0 116816 0 1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  la_buf\[35\]
timestamp 1654395037
transform 1 0 121744 0 -1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  la_buf\[36\]
timestamp 1654395037
transform 1 0 124880 0 1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  la_buf\[37\]
timestamp 1654395037
transform 1 0 129136 0 -1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  la_buf\[38\]
timestamp 1654395037
transform 1 0 134400 0 1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  la_buf\[39\]
timestamp 1654395037
transform -1 0 144480 0 1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  la_buf\[40\]
timestamp 1654395037
transform -1 0 149744 0 -1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  la_buf\[41\]
timestamp 1654395037
transform -1 0 156128 0 1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  la_buf\[42\]
timestamp 1654395037
transform -1 0 161056 0 1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  la_buf\[43\]
timestamp 1654395037
transform -1 0 164416 0 -1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  la_buf\[44\]
timestamp 1654395037
transform -1 0 166208 0 -1 9408
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  la_buf\[45\]
timestamp 1654395037
transform -1 0 164976 0 -1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  la_buf\[46\]
timestamp 1654395037
transform -1 0 169456 0 1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  la_buf\[47\]
timestamp 1654395037
transform -1 0 172368 0 -1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  la_buf\[48\]
timestamp 1654395037
transform -1 0 174832 0 -1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  la_buf\[49\]
timestamp 1654395037
transform -1 0 176288 0 1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  la_buf\[50\]
timestamp 1654395037
transform -1 0 180320 0 -1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  la_buf\[51\]
timestamp 1654395037
transform -1 0 181440 0 -1 9408
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  la_buf\[52\]
timestamp 1654395037
transform -1 0 175168 0 -1 9408
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  la_buf\[53\]
timestamp 1654395037
transform -1 0 177744 0 1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  la_buf\[54\]
timestamp 1654395037
transform -1 0 180320 0 -1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  la_buf\[55\]
timestamp 1654395037
transform -1 0 184800 0 1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  la_buf\[56\]
timestamp 1654395037
transform 1 0 192080 0 1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  la_buf\[57\]
timestamp 1654395037
transform 1 0 196336 0 1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  la_buf\[58\]
timestamp 1654395037
transform -1 0 202720 0 1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  la_buf\[59\]
timestamp 1654395037
transform -1 0 205072 0 -1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  la_buf\[60\]
timestamp 1654395037
transform -1 0 208096 0 1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  la_buf\[61\]
timestamp 1654395037
transform -1 0 212128 0 -1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  la_buf\[62\]
timestamp 1654395037
transform -1 0 208768 0 1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  la_buf\[63\]
timestamp 1654395037
transform -1 0 207872 0 -1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_irq_buffers\[0\] pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 208992 0 1 7840
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_irq_buffers\[1\]
timestamp 1654395037
transform -1 0 208880 0 1 9408
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_irq_buffers\[2\]
timestamp 1654395037
transform -1 0 210336 0 -1 9408
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_irq_gates\[0\] pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 206080 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_irq_gates\[1\]
timestamp 1654395037
transform -1 0 210112 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_irq_gates\[2\]
timestamp 1654395037
transform -1 0 211120 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_to_mprj_in_buffers\[0\]
timestamp 1654395037
transform -1 0 20720 0 1 4704
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_to_mprj_in_buffers\[1\]
timestamp 1654395037
transform -1 0 24640 0 -1 9408
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_to_mprj_in_buffers\[2\]
timestamp 1654395037
transform -1 0 22736 0 -1 6272
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_to_mprj_in_buffers\[3\]
timestamp 1654395037
transform -1 0 24976 0 -1 6272
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_to_mprj_in_buffers\[4\]
timestamp 1654395037
transform -1 0 24640 0 1 6272
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_to_mprj_in_buffers\[5\]
timestamp 1654395037
transform -1 0 20496 0 -1 6272
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_to_mprj_in_buffers\[6\]
timestamp 1654395037
transform -1 0 24640 0 1 4704
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_to_mprj_in_buffers\[7\]
timestamp 1654395037
transform -1 0 28000 0 1 6272
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_to_mprj_in_buffers\[8\]
timestamp 1654395037
transform -1 0 28560 0 1 4704
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_to_mprj_in_buffers\[9\]
timestamp 1654395037
transform -1 0 30688 0 -1 6272
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_to_mprj_in_buffers\[10\]
timestamp 1654395037
transform -1 0 32928 0 -1 6272
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_to_mprj_in_buffers\[11\]
timestamp 1654395037
transform -1 0 35280 0 1 4704
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_to_mprj_in_buffers\[12\]
timestamp 1654395037
transform -1 0 37296 0 -1 6272
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_to_mprj_in_buffers\[13\]
timestamp 1654395037
transform 1 0 10976 0 -1 6272
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_to_mprj_in_buffers\[14\]
timestamp 1654395037
transform 1 0 10864 0 1 4704
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_to_mprj_in_buffers\[15\]
timestamp 1654395037
transform -1 0 12992 0 -1 7840
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_to_mprj_in_buffers\[16\]
timestamp 1654395037
transform -1 0 8960 0 1 4704
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_to_mprj_in_buffers\[17\]
timestamp 1654395037
transform -1 0 9072 0 -1 6272
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_to_mprj_in_buffers\[18\]
timestamp 1654395037
transform -1 0 16016 0 1 4704
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_to_mprj_in_buffers\[19\]
timestamp 1654395037
transform -1 0 20944 0 1 6272
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_to_mprj_in_buffers\[20\]
timestamp 1654395037
transform -1 0 28448 0 -1 6272
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_to_mprj_in_buffers\[21\]
timestamp 1654395037
transform -1 0 32480 0 1 4704
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_to_mprj_in_buffers\[22\]
timestamp 1654395037
transform -1 0 38864 0 1 4704
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_to_mprj_in_buffers\[23\]
timestamp 1654395037
transform -1 0 43344 0 1 4704
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_to_mprj_in_buffers\[24\]
timestamp 1654395037
transform -1 0 46816 0 -1 6272
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_to_mprj_in_buffers\[25\]
timestamp 1654395037
transform -1 0 48160 0 1 4704
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_to_mprj_in_buffers\[26\]
timestamp 1654395037
transform -1 0 51296 0 -1 6272
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_to_mprj_in_buffers\[27\]
timestamp 1654395037
transform -1 0 52080 0 1 4704
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_to_mprj_in_buffers\[28\]
timestamp 1654395037
transform -1 0 56000 0 1 4704
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_to_mprj_in_buffers\[29\]
timestamp 1654395037
transform -1 0 59920 0 1 4704
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_to_mprj_in_buffers\[30\]
timestamp 1654395037
transform -1 0 63840 0 1 4704
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_to_mprj_in_buffers\[31\]
timestamp 1654395037
transform -1 0 67648 0 1 4704
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_to_mprj_in_buffers\[32\]
timestamp 1654395037
transform 1 0 68880 0 1 4704
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_to_mprj_in_buffers\[33\]
timestamp 1654395037
transform -1 0 74144 0 1 4704
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_to_mprj_in_buffers\[34\]
timestamp 1654395037
transform -1 0 77168 0 -1 6272
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_to_mprj_in_buffers\[35\]
timestamp 1654395037
transform -1 0 79520 0 1 4704
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_to_mprj_in_buffers\[36\]
timestamp 1654395037
transform -1 0 83104 0 -1 6272
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_to_mprj_in_buffers\[37\]
timestamp 1654395037
transform -1 0 83440 0 1 4704
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_to_mprj_in_buffers\[38\]
timestamp 1654395037
transform -1 0 85568 0 -1 6272
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_to_mprj_in_buffers\[39\]
timestamp 1654395037
transform -1 0 87360 0 1 4704
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_to_mprj_in_buffers\[40\]
timestamp 1654395037
transform -1 0 90832 0 1 4704
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_to_mprj_in_buffers\[41\]
timestamp 1654395037
transform -1 0 94416 0 1 4704
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_to_mprj_in_buffers\[42\]
timestamp 1654395037
transform -1 0 97664 0 1 4704
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_to_mprj_in_buffers\[43\]
timestamp 1654395037
transform -1 0 100912 0 -1 6272
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_to_mprj_in_buffers\[44\]
timestamp 1654395037
transform -1 0 103040 0 1 4704
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_to_mprj_in_buffers\[45\]
timestamp 1654395037
transform -1 0 106960 0 1 4704
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_to_mprj_in_buffers\[46\]
timestamp 1654395037
transform -1 0 110544 0 1 4704
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_to_mprj_in_buffers\[47\]
timestamp 1654395037
transform -1 0 113792 0 1 4704
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_to_mprj_in_buffers\[48\]
timestamp 1654395037
transform -1 0 117264 0 1 4704
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_to_mprj_in_buffers\[49\]
timestamp 1654395037
transform -1 0 119504 0 -1 6272
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_to_mprj_in_buffers\[50\]
timestamp 1654395037
transform -1 0 122416 0 1 4704
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_to_mprj_in_buffers\[51\]
timestamp 1654395037
transform -1 0 125104 0 1 4704
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_to_mprj_in_buffers\[52\]
timestamp 1654395037
transform -1 0 129024 0 1 4704
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_to_mprj_in_buffers\[53\]
timestamp 1654395037
transform -1 0 130816 0 -1 6272
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_to_mprj_in_buffers\[54\]
timestamp 1654395037
transform -1 0 133056 0 1 4704
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_to_mprj_in_buffers\[55\]
timestamp 1654395037
transform 1 0 132832 0 -1 6272
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_to_mprj_in_buffers\[56\]
timestamp 1654395037
transform -1 0 136864 0 1 4704
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_to_mprj_in_buffers\[57\]
timestamp 1654395037
transform -1 0 138992 0 -1 6272
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_to_mprj_in_buffers\[58\]
timestamp 1654395037
transform -1 0 140896 0 1 4704
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_to_mprj_in_buffers\[59\]
timestamp 1654395037
transform -1 0 146160 0 1 4704
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_to_mprj_in_buffers\[60\]
timestamp 1654395037
transform -1 0 152880 0 1 4704
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_to_mprj_in_buffers\[61\]
timestamp 1654395037
transform -1 0 164304 0 1 4704
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_to_mprj_in_buffers\[62\]
timestamp 1654395037
transform -1 0 171696 0 1 6272
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_to_mprj_in_buffers\[63\]
timestamp 1654395037
transform -1 0 178528 0 1 6272
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_to_mprj_in_gates\[0\]
timestamp 1654395037
transform 1 0 47712 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_to_mprj_in_gates\[1\]
timestamp 1654395037
transform -1 0 52304 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_to_mprj_in_gates\[2\]
timestamp 1654395037
transform 1 0 53872 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_to_mprj_in_gates\[3\]
timestamp 1654395037
transform -1 0 59136 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_to_mprj_in_gates\[4\]
timestamp 1654395037
transform -1 0 63168 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_to_mprj_in_gates\[5\]
timestamp 1654395037
transform -1 0 66976 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_to_mprj_in_gates\[6\]
timestamp 1654395037
transform -1 0 70896 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_to_mprj_in_gates\[7\]
timestamp 1654395037
transform -1 0 74928 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_to_mprj_in_gates\[8\]
timestamp 1654395037
transform -1 0 78624 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_to_mprj_in_gates\[9\]
timestamp 1654395037
transform -1 0 82880 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_to_mprj_in_gates\[10\]
timestamp 1654395037
transform -1 0 85120 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_to_mprj_in_gates\[11\]
timestamp 1654395037
transform -1 0 87696 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_to_mprj_in_gates\[12\]
timestamp 1654395037
transform -1 0 90832 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_to_mprj_in_gates\[13\]
timestamp 1654395037
transform -1 0 95648 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_to_mprj_in_gates\[14\]
timestamp 1654395037
transform -1 0 97552 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_to_mprj_in_gates\[15\]
timestamp 1654395037
transform -1 0 99344 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_to_mprj_in_gates\[16\]
timestamp 1654395037
transform -1 0 100464 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_to_mprj_in_gates\[17\]
timestamp 1654395037
transform -1 0 103264 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_to_mprj_in_gates\[18\]
timestamp 1654395037
transform -1 0 104496 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_to_mprj_in_gates\[19\]
timestamp 1654395037
transform -1 0 107408 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_to_mprj_in_gates\[20\]
timestamp 1654395037
transform -1 0 110656 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_to_mprj_in_gates\[21\]
timestamp 1654395037
transform -1 0 112896 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_to_mprj_in_gates\[22\]
timestamp 1654395037
transform -1 0 115696 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_to_mprj_in_gates\[23\]
timestamp 1654395037
transform -1 0 118272 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_to_mprj_in_gates\[24\]
timestamp 1654395037
transform -1 0 120400 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_to_mprj_in_gates\[25\]
timestamp 1654395037
transform -1 0 122752 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_to_mprj_in_gates\[26\]
timestamp 1654395037
transform -1 0 126560 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_to_mprj_in_gates\[27\]
timestamp 1654395037
transform -1 0 128688 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_to_mprj_in_gates\[28\]
timestamp 1654395037
transform -1 0 131040 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_to_mprj_in_gates\[29\]
timestamp 1654395037
transform -1 0 134512 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_to_mprj_in_gates\[30\]
timestamp 1654395037
transform -1 0 136528 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_to_mprj_in_gates\[31\]
timestamp 1654395037
transform -1 0 138544 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_to_mprj_in_gates\[32\]
timestamp 1654395037
transform -1 0 140560 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_to_mprj_in_gates\[33\]
timestamp 1654395037
transform -1 0 140224 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_to_mprj_in_gates\[34\]
timestamp 1654395037
transform -1 0 141008 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_to_mprj_in_gates\[35\]
timestamp 1654395037
transform -1 0 142464 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_to_mprj_in_gates\[36\]
timestamp 1654395037
transform -1 0 142576 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_to_mprj_in_gates\[37\]
timestamp 1654395037
transform -1 0 143024 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_to_mprj_in_gates\[38\]
timestamp 1654395037
transform -1 0 144480 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_to_mprj_in_gates\[39\]
timestamp 1654395037
transform -1 0 146496 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_to_mprj_in_gates\[40\]
timestamp 1654395037
transform -1 0 146496 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_to_mprj_in_gates\[41\]
timestamp 1654395037
transform -1 0 148512 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_to_mprj_in_gates\[42\]
timestamp 1654395037
transform -1 0 150416 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_to_mprj_in_gates\[43\]
timestamp 1654395037
transform -1 0 151424 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_to_mprj_in_gates\[44\]
timestamp 1654395037
transform -1 0 154448 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_to_mprj_in_gates\[45\]
timestamp 1654395037
transform -1 0 156128 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_to_mprj_in_gates\[46\]
timestamp 1654395037
transform -1 0 157696 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_to_mprj_in_gates\[47\]
timestamp 1654395037
transform -1 0 157920 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_to_mprj_in_gates\[48\]
timestamp 1654395037
transform -1 0 154448 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_to_mprj_in_gates\[49\]
timestamp 1654395037
transform -1 0 171920 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_to_mprj_in_gates\[50\]
timestamp 1654395037
transform -1 0 179760 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_to_mprj_in_gates\[51\]
timestamp 1654395037
transform -1 0 179760 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_to_mprj_in_gates\[52\]
timestamp 1654395037
transform -1 0 182224 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_to_mprj_in_gates\[53\]
timestamp 1654395037
transform -1 0 183456 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_to_mprj_in_gates\[54\]
timestamp 1654395037
transform -1 0 184240 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_to_mprj_in_gates\[55\]
timestamp 1654395037
transform -1 0 186816 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_to_mprj_in_gates\[56\]
timestamp 1654395037
transform -1 0 186256 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_to_mprj_in_gates\[57\]
timestamp 1654395037
transform -1 0 186256 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_to_mprj_in_gates\[58\]
timestamp 1654395037
transform -1 0 188272 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_to_mprj_in_gates\[59\]
timestamp 1654395037
transform -1 0 187600 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_to_mprj_in_gates\[60\]
timestamp 1654395037
transform -1 0 188496 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_to_mprj_in_gates\[61\]
timestamp 1654395037
transform -1 0 190176 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_to_mprj_in_gates\[62\]
timestamp 1654395037
transform -1 0 190288 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_to_mprj_in_gates\[63\]
timestamp 1654395037
transform -1 0 190512 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_wb_ack_buffer
timestamp 1654395037
transform -1 0 210336 0 1 6272
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_wb_ack_gate
timestamp 1654395037
transform -1 0 212352 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_wb_dat_buffers\[0\]
timestamp 1654395037
transform 1 0 155904 0 1 4704
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_wb_dat_buffers\[1\]
timestamp 1654395037
transform 1 0 158368 0 1 4704
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_wb_dat_buffers\[2\]
timestamp 1654395037
transform 1 0 158704 0 1 6272
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_wb_dat_buffers\[3\]
timestamp 1654395037
transform 1 0 158144 0 -1 7840
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_wb_dat_buffers\[4\]
timestamp 1654395037
transform 1 0 165200 0 -1 6272
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_wb_dat_buffers\[5\]
timestamp 1654395037
transform 1 0 166208 0 1 4704
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_wb_dat_buffers\[6\]
timestamp 1654395037
transform 1 0 170128 0 1 4704
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_wb_dat_buffers\[7\]
timestamp 1654395037
transform 1 0 166432 0 1 9408
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_wb_dat_buffers\[8\]
timestamp 1654395037
transform 1 0 169008 0 1 7840
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_wb_dat_buffers\[9\]
timestamp 1654395037
transform 1 0 174048 0 1 4704
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_wb_dat_buffers\[10\]
timestamp 1654395037
transform 1 0 172592 0 -1 7840
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_wb_dat_buffers\[11\]
timestamp 1654395037
transform 1 0 177968 0 1 4704
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_wb_dat_buffers\[12\]
timestamp 1654395037
transform 1 0 174608 0 1 9408
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_wb_dat_buffers\[13\]
timestamp 1654395037
transform 1 0 180544 0 -1 6272
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_wb_dat_buffers\[14\]
timestamp 1654395037
transform 1 0 181888 0 1 4704
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_wb_dat_buffers\[15\]
timestamp 1654395037
transform 1 0 181328 0 -1 7840
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_wb_dat_buffers\[16\]
timestamp 1654395037
transform 1 0 184464 0 -1 6272
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_wb_dat_buffers\[17\]
timestamp 1654395037
transform 1 0 157920 0 -1 6272
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_wb_dat_buffers\[18\]
timestamp 1654395037
transform 1 0 160944 0 1 6272
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_wb_dat_buffers\[19\]
timestamp 1654395037
transform 1 0 161280 0 1 7840
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_wb_dat_buffers\[20\]
timestamp 1654395037
transform 1 0 164640 0 -1 7840
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_wb_dat_buffers\[21\]
timestamp 1654395037
transform 1 0 164528 0 1 7840
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_wb_dat_buffers\[22\]
timestamp 1654395037
transform 1 0 168560 0 -1 6272
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_wb_dat_buffers\[23\]
timestamp 1654395037
transform 1 0 166768 0 1 7840
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_wb_dat_buffers\[24\]
timestamp 1654395037
transform 1 0 196224 0 -1 6272
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_wb_dat_buffers\[25\]
timestamp 1654395037
transform 1 0 197568 0 1 4704
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_wb_dat_buffers\[26\]
timestamp 1654395037
transform 1 0 201488 0 1 4704
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_wb_dat_buffers\[27\]
timestamp 1654395037
transform 1 0 200368 0 -1 7840
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_wb_dat_buffers\[28\]
timestamp 1654395037
transform 1 0 205408 0 1 4704
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_wb_dat_buffers\[29\]
timestamp 1654395037
transform 1 0 205296 0 -1 6272
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_wb_dat_buffers\[30\]
timestamp 1654395037
transform 1 0 203616 0 -1 9408
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  user_wb_dat_buffers\[31\]
timestamp 1654395037
transform 1 0 209328 0 1 4704
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_wb_dat_gates\[0\]
timestamp 1654395037
transform 1 0 131712 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_wb_dat_gates\[1\]
timestamp 1654395037
transform 1 0 131936 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_wb_dat_gates\[2\]
timestamp 1654395037
transform 1 0 133728 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_wb_dat_gates\[3\]
timestamp 1654395037
transform 1 0 133168 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_wb_dat_gates\[4\]
timestamp 1654395037
transform 1 0 134848 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_wb_dat_gates\[5\]
timestamp 1654395037
transform 1 0 136752 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_wb_dat_gates\[6\]
timestamp 1654395037
transform 1 0 136752 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_wb_dat_gates\[7\]
timestamp 1654395037
transform 1 0 138768 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_wb_dat_gates\[8\]
timestamp 1654395037
transform 1 0 139664 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_wb_dat_gates\[9\]
timestamp 1654395037
transform 1 0 142240 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_wb_dat_gates\[10\]
timestamp 1654395037
transform 1 0 145040 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_wb_dat_gates\[11\]
timestamp 1654395037
transform 1 0 148624 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_wb_dat_gates\[12\]
timestamp 1654395037
transform 1 0 151536 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_wb_dat_gates\[13\]
timestamp 1654395037
transform 1 0 154672 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_wb_dat_gates\[14\]
timestamp 1654395037
transform 1 0 156688 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_wb_dat_gates\[15\]
timestamp 1654395037
transform 1 0 162288 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_wb_dat_gates\[16\]
timestamp 1654395037
transform 1 0 168560 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_wb_dat_gates\[17\]
timestamp 1654395037
transform 1 0 144928 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_wb_dat_gates\[18\]
timestamp 1654395037
transform 1 0 147952 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_wb_dat_gates\[19\]
timestamp 1654395037
transform 1 0 150304 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_wb_dat_gates\[20\]
timestamp 1654395037
transform 1 0 152768 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_wb_dat_gates\[21\]
timestamp 1654395037
transform 1 0 154784 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_wb_dat_gates\[22\]
timestamp 1654395037
transform 1 0 157136 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_wb_dat_gates\[23\]
timestamp 1654395037
transform 1 0 159264 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_wb_dat_gates\[24\]
timestamp 1654395037
transform 1 0 181888 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_wb_dat_gates\[25\]
timestamp 1654395037
transform 1 0 184464 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_wb_dat_gates\[26\]
timestamp 1654395037
transform 1 0 186480 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_wb_dat_gates\[27\]
timestamp 1654395037
transform 1 0 185808 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_wb_dat_gates\[28\]
timestamp 1654395037
transform 1 0 188496 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_wb_dat_gates\[29\]
timestamp 1654395037
transform 1 0 188384 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_wb_dat_gates\[30\]
timestamp 1654395037
transform 1 0 189728 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  user_wb_dat_gates\[31\]
timestamp 1654395037
transform 1 0 192416 0 -1 9408
box -86 -86 1878 870
<< labels >>
flabel metal4 s 28348 4644 28668 10252 0 FreeSans 1280 90 0 0 VDD
port 0 nsew power bidirectional
flabel metal4 s 82676 4644 82996 10252 0 FreeSans 1280 90 0 0 VDD
port 0 nsew power bidirectional
flabel metal4 s 137004 4644 137324 10252 0 FreeSans 1280 90 0 0 VDD
port 0 nsew power bidirectional
flabel metal4 s 191332 4644 191652 10252 0 FreeSans 1280 90 0 0 VDD
port 0 nsew power bidirectional
flabel metal5 s 1284 5243 218684 5563 0 FreeSans 2304 0 0 0 VDD
port 0 nsew power bidirectional
flabel metal5 s 1284 6641 218684 6961 0 FreeSans 2304 0 0 0 VDD
port 0 nsew power bidirectional
flabel metal5 s 1284 8039 218684 8359 0 FreeSans 2304 0 0 0 VDD
port 0 nsew power bidirectional
flabel metal5 s 1284 9437 218684 9757 0 FreeSans 2304 0 0 0 VDD
port 0 nsew power bidirectional
flabel metal4 s 55512 4644 55832 10252 0 FreeSans 1280 90 0 0 VSS
port 1 nsew ground bidirectional
flabel metal4 s 109840 4644 110160 10252 0 FreeSans 1280 90 0 0 VSS
port 1 nsew ground bidirectional
flabel metal4 s 164168 4644 164488 10252 0 FreeSans 1280 90 0 0 VSS
port 1 nsew ground bidirectional
flabel metal5 s 1284 5942 218684 6262 0 FreeSans 2304 0 0 0 VSS
port 1 nsew ground bidirectional
flabel metal5 s 1284 7340 218684 7660 0 FreeSans 2304 0 0 0 VSS
port 1 nsew ground bidirectional
flabel metal5 s 1284 8738 218684 9058 0 FreeSans 2304 0 0 0 VSS
port 1 nsew ground bidirectional
flabel metal3 s 0 2520 800 2632 0 FreeSans 448 0 0 0 caravel_clk
port 2 nsew signal input
flabel metal3 s 0 7448 800 7560 0 FreeSans 448 0 0 0 caravel_clk2
port 3 nsew signal input
flabel metal3 s 0 12376 800 12488 0 FreeSans 448 0 0 0 caravel_rstn
port 4 nsew signal input
flabel metal2 s 77448 14200 77560 15000 0 FreeSans 448 90 0 0 la_data_in_core[0]
port 5 nsew signal tristate
flabel metal2 s 99288 14200 99400 15000 0 FreeSans 448 90 0 0 la_data_in_core[10]
port 6 nsew signal tristate
flabel metal2 s 101528 14200 101640 15000 0 FreeSans 448 90 0 0 la_data_in_core[11]
port 7 nsew signal tristate
flabel metal2 s 103656 14200 103768 15000 0 FreeSans 448 90 0 0 la_data_in_core[12]
port 8 nsew signal tristate
flabel metal2 s 105896 14200 106008 15000 0 FreeSans 448 90 0 0 la_data_in_core[13]
port 9 nsew signal tristate
flabel metal2 s 108024 14200 108136 15000 0 FreeSans 448 90 0 0 la_data_in_core[14]
port 10 nsew signal tristate
flabel metal2 s 110264 14200 110376 15000 0 FreeSans 448 90 0 0 la_data_in_core[15]
port 11 nsew signal tristate
flabel metal2 s 112504 14200 112616 15000 0 FreeSans 448 90 0 0 la_data_in_core[16]
port 12 nsew signal tristate
flabel metal2 s 114632 14200 114744 15000 0 FreeSans 448 90 0 0 la_data_in_core[17]
port 13 nsew signal tristate
flabel metal2 s 116872 14200 116984 15000 0 FreeSans 448 90 0 0 la_data_in_core[18]
port 14 nsew signal tristate
flabel metal2 s 119000 14200 119112 15000 0 FreeSans 448 90 0 0 la_data_in_core[19]
port 15 nsew signal tristate
flabel metal2 s 79688 14200 79800 15000 0 FreeSans 448 90 0 0 la_data_in_core[1]
port 16 nsew signal tristate
flabel metal2 s 121240 14200 121352 15000 0 FreeSans 448 90 0 0 la_data_in_core[20]
port 17 nsew signal tristate
flabel metal2 s 123368 14200 123480 15000 0 FreeSans 448 90 0 0 la_data_in_core[21]
port 18 nsew signal tristate
flabel metal2 s 125608 14200 125720 15000 0 FreeSans 448 90 0 0 la_data_in_core[22]
port 19 nsew signal tristate
flabel metal2 s 127736 14200 127848 15000 0 FreeSans 448 90 0 0 la_data_in_core[23]
port 20 nsew signal tristate
flabel metal2 s 129976 14200 130088 15000 0 FreeSans 448 90 0 0 la_data_in_core[24]
port 21 nsew signal tristate
flabel metal2 s 132104 14200 132216 15000 0 FreeSans 448 90 0 0 la_data_in_core[25]
port 22 nsew signal tristate
flabel metal2 s 134344 14200 134456 15000 0 FreeSans 448 90 0 0 la_data_in_core[26]
port 23 nsew signal tristate
flabel metal2 s 136472 14200 136584 15000 0 FreeSans 448 90 0 0 la_data_in_core[27]
port 24 nsew signal tristate
flabel metal2 s 138712 14200 138824 15000 0 FreeSans 448 90 0 0 la_data_in_core[28]
port 25 nsew signal tristate
flabel metal2 s 140840 14200 140952 15000 0 FreeSans 448 90 0 0 la_data_in_core[29]
port 26 nsew signal tristate
flabel metal2 s 81816 14200 81928 15000 0 FreeSans 448 90 0 0 la_data_in_core[2]
port 27 nsew signal tristate
flabel metal2 s 143080 14200 143192 15000 0 FreeSans 448 90 0 0 la_data_in_core[30]
port 28 nsew signal tristate
flabel metal2 s 145208 14200 145320 15000 0 FreeSans 448 90 0 0 la_data_in_core[31]
port 29 nsew signal tristate
flabel metal2 s 147448 14200 147560 15000 0 FreeSans 448 90 0 0 la_data_in_core[32]
port 30 nsew signal tristate
flabel metal2 s 149576 14200 149688 15000 0 FreeSans 448 90 0 0 la_data_in_core[33]
port 31 nsew signal tristate
flabel metal2 s 151816 14200 151928 15000 0 FreeSans 448 90 0 0 la_data_in_core[34]
port 32 nsew signal tristate
flabel metal2 s 153944 14200 154056 15000 0 FreeSans 448 90 0 0 la_data_in_core[35]
port 33 nsew signal tristate
flabel metal2 s 156184 14200 156296 15000 0 FreeSans 448 90 0 0 la_data_in_core[36]
port 34 nsew signal tristate
flabel metal2 s 158312 14200 158424 15000 0 FreeSans 448 90 0 0 la_data_in_core[37]
port 35 nsew signal tristate
flabel metal2 s 160552 14200 160664 15000 0 FreeSans 448 90 0 0 la_data_in_core[38]
port 36 nsew signal tristate
flabel metal2 s 162680 14200 162792 15000 0 FreeSans 448 90 0 0 la_data_in_core[39]
port 37 nsew signal tristate
flabel metal2 s 84056 14200 84168 15000 0 FreeSans 448 90 0 0 la_data_in_core[3]
port 38 nsew signal tristate
flabel metal2 s 164920 14200 165032 15000 0 FreeSans 448 90 0 0 la_data_in_core[40]
port 39 nsew signal tristate
flabel metal2 s 167160 14200 167272 15000 0 FreeSans 448 90 0 0 la_data_in_core[41]
port 40 nsew signal tristate
flabel metal2 s 169288 14200 169400 15000 0 FreeSans 448 90 0 0 la_data_in_core[42]
port 41 nsew signal tristate
flabel metal2 s 171528 14200 171640 15000 0 FreeSans 448 90 0 0 la_data_in_core[43]
port 42 nsew signal tristate
flabel metal2 s 173656 14200 173768 15000 0 FreeSans 448 90 0 0 la_data_in_core[44]
port 43 nsew signal tristate
flabel metal2 s 175896 14200 176008 15000 0 FreeSans 448 90 0 0 la_data_in_core[45]
port 44 nsew signal tristate
flabel metal2 s 178024 14200 178136 15000 0 FreeSans 448 90 0 0 la_data_in_core[46]
port 45 nsew signal tristate
flabel metal2 s 180264 14200 180376 15000 0 FreeSans 448 90 0 0 la_data_in_core[47]
port 46 nsew signal tristate
flabel metal2 s 182392 14200 182504 15000 0 FreeSans 448 90 0 0 la_data_in_core[48]
port 47 nsew signal tristate
flabel metal2 s 184632 14200 184744 15000 0 FreeSans 448 90 0 0 la_data_in_core[49]
port 48 nsew signal tristate
flabel metal2 s 86184 14200 86296 15000 0 FreeSans 448 90 0 0 la_data_in_core[4]
port 49 nsew signal tristate
flabel metal2 s 186760 14200 186872 15000 0 FreeSans 448 90 0 0 la_data_in_core[50]
port 50 nsew signal tristate
flabel metal2 s 189000 14200 189112 15000 0 FreeSans 448 90 0 0 la_data_in_core[51]
port 51 nsew signal tristate
flabel metal2 s 191128 14200 191240 15000 0 FreeSans 448 90 0 0 la_data_in_core[52]
port 52 nsew signal tristate
flabel metal2 s 193368 14200 193480 15000 0 FreeSans 448 90 0 0 la_data_in_core[53]
port 53 nsew signal tristate
flabel metal2 s 195496 14200 195608 15000 0 FreeSans 448 90 0 0 la_data_in_core[54]
port 54 nsew signal tristate
flabel metal2 s 197736 14200 197848 15000 0 FreeSans 448 90 0 0 la_data_in_core[55]
port 55 nsew signal tristate
flabel metal2 s 199864 14200 199976 15000 0 FreeSans 448 90 0 0 la_data_in_core[56]
port 56 nsew signal tristate
flabel metal2 s 202104 14200 202216 15000 0 FreeSans 448 90 0 0 la_data_in_core[57]
port 57 nsew signal tristate
flabel metal2 s 204232 14200 204344 15000 0 FreeSans 448 90 0 0 la_data_in_core[58]
port 58 nsew signal tristate
flabel metal2 s 206472 14200 206584 15000 0 FreeSans 448 90 0 0 la_data_in_core[59]
port 59 nsew signal tristate
flabel metal2 s 88424 14200 88536 15000 0 FreeSans 448 90 0 0 la_data_in_core[5]
port 60 nsew signal tristate
flabel metal2 s 208600 14200 208712 15000 0 FreeSans 448 90 0 0 la_data_in_core[60]
port 61 nsew signal tristate
flabel metal2 s 210840 14200 210952 15000 0 FreeSans 448 90 0 0 la_data_in_core[61]
port 62 nsew signal tristate
flabel metal2 s 212968 14200 213080 15000 0 FreeSans 448 90 0 0 la_data_in_core[62]
port 63 nsew signal tristate
flabel metal2 s 215208 14200 215320 15000 0 FreeSans 448 90 0 0 la_data_in_core[63]
port 64 nsew signal tristate
flabel metal2 s 90552 14200 90664 15000 0 FreeSans 448 90 0 0 la_data_in_core[6]
port 65 nsew signal tristate
flabel metal2 s 92792 14200 92904 15000 0 FreeSans 448 90 0 0 la_data_in_core[7]
port 66 nsew signal tristate
flabel metal2 s 94920 14200 95032 15000 0 FreeSans 448 90 0 0 la_data_in_core[8]
port 67 nsew signal tristate
flabel metal2 s 97160 14200 97272 15000 0 FreeSans 448 90 0 0 la_data_in_core[9]
port 68 nsew signal tristate
flabel metal2 s 168 0 280 800 0 FreeSans 448 90 0 0 la_data_in_mprj[0]
port 69 nsew signal tristate
flabel metal2 s 6216 0 6328 800 0 FreeSans 448 90 0 0 la_data_in_mprj[10]
port 70 nsew signal tristate
flabel metal2 s 6776 0 6888 800 0 FreeSans 448 90 0 0 la_data_in_mprj[11]
port 71 nsew signal tristate
flabel metal2 s 7448 0 7560 800 0 FreeSans 448 90 0 0 la_data_in_mprj[12]
port 72 nsew signal tristate
flabel metal2 s 8008 0 8120 800 0 FreeSans 448 90 0 0 la_data_in_mprj[13]
port 73 nsew signal tristate
flabel metal2 s 8680 0 8792 800 0 FreeSans 448 90 0 0 la_data_in_mprj[14]
port 74 nsew signal tristate
flabel metal2 s 9240 0 9352 800 0 FreeSans 448 90 0 0 la_data_in_mprj[15]
port 75 nsew signal tristate
flabel metal2 s 9912 0 10024 800 0 FreeSans 448 90 0 0 la_data_in_mprj[16]
port 76 nsew signal tristate
flabel metal2 s 10472 0 10584 800 0 FreeSans 448 90 0 0 la_data_in_mprj[17]
port 77 nsew signal tristate
flabel metal2 s 11032 0 11144 800 0 FreeSans 448 90 0 0 la_data_in_mprj[18]
port 78 nsew signal tristate
flabel metal2 s 11704 0 11816 800 0 FreeSans 448 90 0 0 la_data_in_mprj[19]
port 79 nsew signal tristate
flabel metal2 s 728 0 840 800 0 FreeSans 448 90 0 0 la_data_in_mprj[1]
port 80 nsew signal tristate
flabel metal2 s 12264 0 12376 800 0 FreeSans 448 90 0 0 la_data_in_mprj[20]
port 81 nsew signal tristate
flabel metal2 s 12936 0 13048 800 0 FreeSans 448 90 0 0 la_data_in_mprj[21]
port 82 nsew signal tristate
flabel metal2 s 13496 0 13608 800 0 FreeSans 448 90 0 0 la_data_in_mprj[22]
port 83 nsew signal tristate
flabel metal2 s 14168 0 14280 800 0 FreeSans 448 90 0 0 la_data_in_mprj[23]
port 84 nsew signal tristate
flabel metal2 s 14728 0 14840 800 0 FreeSans 448 90 0 0 la_data_in_mprj[24]
port 85 nsew signal tristate
flabel metal2 s 15400 0 15512 800 0 FreeSans 448 90 0 0 la_data_in_mprj[25]
port 86 nsew signal tristate
flabel metal2 s 15960 0 16072 800 0 FreeSans 448 90 0 0 la_data_in_mprj[26]
port 87 nsew signal tristate
flabel metal2 s 16520 0 16632 800 0 FreeSans 448 90 0 0 la_data_in_mprj[27]
port 88 nsew signal tristate
flabel metal2 s 17192 0 17304 800 0 FreeSans 448 90 0 0 la_data_in_mprj[28]
port 89 nsew signal tristate
flabel metal2 s 17752 0 17864 800 0 FreeSans 448 90 0 0 la_data_in_mprj[29]
port 90 nsew signal tristate
flabel metal2 s 1288 0 1400 800 0 FreeSans 448 90 0 0 la_data_in_mprj[2]
port 91 nsew signal tristate
flabel metal2 s 18424 0 18536 800 0 FreeSans 448 90 0 0 la_data_in_mprj[30]
port 92 nsew signal tristate
flabel metal2 s 18984 0 19096 800 0 FreeSans 448 90 0 0 la_data_in_mprj[31]
port 93 nsew signal tristate
flabel metal2 s 19656 0 19768 800 0 FreeSans 448 90 0 0 la_data_in_mprj[32]
port 94 nsew signal tristate
flabel metal2 s 20216 0 20328 800 0 FreeSans 448 90 0 0 la_data_in_mprj[33]
port 95 nsew signal tristate
flabel metal2 s 20888 0 21000 800 0 FreeSans 448 90 0 0 la_data_in_mprj[34]
port 96 nsew signal tristate
flabel metal2 s 21448 0 21560 800 0 FreeSans 448 90 0 0 la_data_in_mprj[35]
port 97 nsew signal tristate
flabel metal2 s 22008 0 22120 800 0 FreeSans 448 90 0 0 la_data_in_mprj[36]
port 98 nsew signal tristate
flabel metal2 s 22680 0 22792 800 0 FreeSans 448 90 0 0 la_data_in_mprj[37]
port 99 nsew signal tristate
flabel metal2 s 23240 0 23352 800 0 FreeSans 448 90 0 0 la_data_in_mprj[38]
port 100 nsew signal tristate
flabel metal2 s 23912 0 24024 800 0 FreeSans 448 90 0 0 la_data_in_mprj[39]
port 101 nsew signal tristate
flabel metal2 s 1960 0 2072 800 0 FreeSans 448 90 0 0 la_data_in_mprj[3]
port 102 nsew signal tristate
flabel metal2 s 24472 0 24584 800 0 FreeSans 448 90 0 0 la_data_in_mprj[40]
port 103 nsew signal tristate
flabel metal2 s 25144 0 25256 800 0 FreeSans 448 90 0 0 la_data_in_mprj[41]
port 104 nsew signal tristate
flabel metal2 s 25704 0 25816 800 0 FreeSans 448 90 0 0 la_data_in_mprj[42]
port 105 nsew signal tristate
flabel metal2 s 26376 0 26488 800 0 FreeSans 448 90 0 0 la_data_in_mprj[43]
port 106 nsew signal tristate
flabel metal2 s 26936 0 27048 800 0 FreeSans 448 90 0 0 la_data_in_mprj[44]
port 107 nsew signal tristate
flabel metal2 s 27496 0 27608 800 0 FreeSans 448 90 0 0 la_data_in_mprj[45]
port 108 nsew signal tristate
flabel metal2 s 28168 0 28280 800 0 FreeSans 448 90 0 0 la_data_in_mprj[46]
port 109 nsew signal tristate
flabel metal2 s 28728 0 28840 800 0 FreeSans 448 90 0 0 la_data_in_mprj[47]
port 110 nsew signal tristate
flabel metal2 s 29400 0 29512 800 0 FreeSans 448 90 0 0 la_data_in_mprj[48]
port 111 nsew signal tristate
flabel metal2 s 29960 0 30072 800 0 FreeSans 448 90 0 0 la_data_in_mprj[49]
port 112 nsew signal tristate
flabel metal2 s 2520 0 2632 800 0 FreeSans 448 90 0 0 la_data_in_mprj[4]
port 113 nsew signal tristate
flabel metal2 s 30632 0 30744 800 0 FreeSans 448 90 0 0 la_data_in_mprj[50]
port 114 nsew signal tristate
flabel metal2 s 31192 0 31304 800 0 FreeSans 448 90 0 0 la_data_in_mprj[51]
port 115 nsew signal tristate
flabel metal2 s 31864 0 31976 800 0 FreeSans 448 90 0 0 la_data_in_mprj[52]
port 116 nsew signal tristate
flabel metal2 s 32424 0 32536 800 0 FreeSans 448 90 0 0 la_data_in_mprj[53]
port 117 nsew signal tristate
flabel metal2 s 32984 0 33096 800 0 FreeSans 448 90 0 0 la_data_in_mprj[54]
port 118 nsew signal tristate
flabel metal2 s 33656 0 33768 800 0 FreeSans 448 90 0 0 la_data_in_mprj[55]
port 119 nsew signal tristate
flabel metal2 s 34216 0 34328 800 0 FreeSans 448 90 0 0 la_data_in_mprj[56]
port 120 nsew signal tristate
flabel metal2 s 34888 0 35000 800 0 FreeSans 448 90 0 0 la_data_in_mprj[57]
port 121 nsew signal tristate
flabel metal2 s 35448 0 35560 800 0 FreeSans 448 90 0 0 la_data_in_mprj[58]
port 122 nsew signal tristate
flabel metal2 s 36120 0 36232 800 0 FreeSans 448 90 0 0 la_data_in_mprj[59]
port 123 nsew signal tristate
flabel metal2 s 3192 0 3304 800 0 FreeSans 448 90 0 0 la_data_in_mprj[5]
port 124 nsew signal tristate
flabel metal2 s 36680 0 36792 800 0 FreeSans 448 90 0 0 la_data_in_mprj[60]
port 125 nsew signal tristate
flabel metal2 s 37352 0 37464 800 0 FreeSans 448 90 0 0 la_data_in_mprj[61]
port 126 nsew signal tristate
flabel metal2 s 37912 0 38024 800 0 FreeSans 448 90 0 0 la_data_in_mprj[62]
port 127 nsew signal tristate
flabel metal2 s 38472 0 38584 800 0 FreeSans 448 90 0 0 la_data_in_mprj[63]
port 128 nsew signal tristate
flabel metal2 s 3752 0 3864 800 0 FreeSans 448 90 0 0 la_data_in_mprj[6]
port 129 nsew signal tristate
flabel metal2 s 4424 0 4536 800 0 FreeSans 448 90 0 0 la_data_in_mprj[7]
port 130 nsew signal tristate
flabel metal2 s 4984 0 5096 800 0 FreeSans 448 90 0 0 la_data_in_mprj[8]
port 131 nsew signal tristate
flabel metal2 s 5544 0 5656 800 0 FreeSans 448 90 0 0 la_data_in_mprj[9]
port 132 nsew signal tristate
flabel metal2 s 78232 14200 78344 15000 0 FreeSans 448 90 0 0 la_data_out_core[0]
port 133 nsew signal input
flabel metal2 s 100072 14200 100184 15000 0 FreeSans 448 90 0 0 la_data_out_core[10]
port 134 nsew signal input
flabel metal2 s 102200 14200 102312 15000 0 FreeSans 448 90 0 0 la_data_out_core[11]
port 135 nsew signal input
flabel metal2 s 104440 14200 104552 15000 0 FreeSans 448 90 0 0 la_data_out_core[12]
port 136 nsew signal input
flabel metal2 s 106568 14200 106680 15000 0 FreeSans 448 90 0 0 la_data_out_core[13]
port 137 nsew signal input
flabel metal2 s 108808 14200 108920 15000 0 FreeSans 448 90 0 0 la_data_out_core[14]
port 138 nsew signal input
flabel metal2 s 111048 14200 111160 15000 0 FreeSans 448 90 0 0 la_data_out_core[15]
port 139 nsew signal input
flabel metal2 s 113176 14200 113288 15000 0 FreeSans 448 90 0 0 la_data_out_core[16]
port 140 nsew signal input
flabel metal2 s 115416 14200 115528 15000 0 FreeSans 448 90 0 0 la_data_out_core[17]
port 141 nsew signal input
flabel metal2 s 117544 14200 117656 15000 0 FreeSans 448 90 0 0 la_data_out_core[18]
port 142 nsew signal input
flabel metal2 s 119784 14200 119896 15000 0 FreeSans 448 90 0 0 la_data_out_core[19]
port 143 nsew signal input
flabel metal2 s 80360 14200 80472 15000 0 FreeSans 448 90 0 0 la_data_out_core[1]
port 144 nsew signal input
flabel metal2 s 121912 14200 122024 15000 0 FreeSans 448 90 0 0 la_data_out_core[20]
port 145 nsew signal input
flabel metal2 s 124152 14200 124264 15000 0 FreeSans 448 90 0 0 la_data_out_core[21]
port 146 nsew signal input
flabel metal2 s 126280 14200 126392 15000 0 FreeSans 448 90 0 0 la_data_out_core[22]
port 147 nsew signal input
flabel metal2 s 128520 14200 128632 15000 0 FreeSans 448 90 0 0 la_data_out_core[23]
port 148 nsew signal input
flabel metal2 s 130648 14200 130760 15000 0 FreeSans 448 90 0 0 la_data_out_core[24]
port 149 nsew signal input
flabel metal2 s 132888 14200 133000 15000 0 FreeSans 448 90 0 0 la_data_out_core[25]
port 150 nsew signal input
flabel metal2 s 135016 14200 135128 15000 0 FreeSans 448 90 0 0 la_data_out_core[26]
port 151 nsew signal input
flabel metal2 s 137256 14200 137368 15000 0 FreeSans 448 90 0 0 la_data_out_core[27]
port 152 nsew signal input
flabel metal2 s 139384 14200 139496 15000 0 FreeSans 448 90 0 0 la_data_out_core[28]
port 153 nsew signal input
flabel metal2 s 141624 14200 141736 15000 0 FreeSans 448 90 0 0 la_data_out_core[29]
port 154 nsew signal input
flabel metal2 s 82600 14200 82712 15000 0 FreeSans 448 90 0 0 la_data_out_core[2]
port 155 nsew signal input
flabel metal2 s 143752 14200 143864 15000 0 FreeSans 448 90 0 0 la_data_out_core[30]
port 156 nsew signal input
flabel metal2 s 145992 14200 146104 15000 0 FreeSans 448 90 0 0 la_data_out_core[31]
port 157 nsew signal input
flabel metal2 s 148120 14200 148232 15000 0 FreeSans 448 90 0 0 la_data_out_core[32]
port 158 nsew signal input
flabel metal2 s 150360 14200 150472 15000 0 FreeSans 448 90 0 0 la_data_out_core[33]
port 159 nsew signal input
flabel metal2 s 152488 14200 152600 15000 0 FreeSans 448 90 0 0 la_data_out_core[34]
port 160 nsew signal input
flabel metal2 s 154728 14200 154840 15000 0 FreeSans 448 90 0 0 la_data_out_core[35]
port 161 nsew signal input
flabel metal2 s 156856 14200 156968 15000 0 FreeSans 448 90 0 0 la_data_out_core[36]
port 162 nsew signal input
flabel metal2 s 159096 14200 159208 15000 0 FreeSans 448 90 0 0 la_data_out_core[37]
port 163 nsew signal input
flabel metal2 s 161224 14200 161336 15000 0 FreeSans 448 90 0 0 la_data_out_core[38]
port 164 nsew signal input
flabel metal2 s 163464 14200 163576 15000 0 FreeSans 448 90 0 0 la_data_out_core[39]
port 165 nsew signal input
flabel metal2 s 84728 14200 84840 15000 0 FreeSans 448 90 0 0 la_data_out_core[3]
port 166 nsew signal input
flabel metal2 s 165704 14200 165816 15000 0 FreeSans 448 90 0 0 la_data_out_core[40]
port 167 nsew signal input
flabel metal2 s 167832 14200 167944 15000 0 FreeSans 448 90 0 0 la_data_out_core[41]
port 168 nsew signal input
flabel metal2 s 170072 14200 170184 15000 0 FreeSans 448 90 0 0 la_data_out_core[42]
port 169 nsew signal input
flabel metal2 s 172200 14200 172312 15000 0 FreeSans 448 90 0 0 la_data_out_core[43]
port 170 nsew signal input
flabel metal2 s 174440 14200 174552 15000 0 FreeSans 448 90 0 0 la_data_out_core[44]
port 171 nsew signal input
flabel metal2 s 176568 14200 176680 15000 0 FreeSans 448 90 0 0 la_data_out_core[45]
port 172 nsew signal input
flabel metal2 s 178808 14200 178920 15000 0 FreeSans 448 90 0 0 la_data_out_core[46]
port 173 nsew signal input
flabel metal2 s 180936 14200 181048 15000 0 FreeSans 448 90 0 0 la_data_out_core[47]
port 174 nsew signal input
flabel metal2 s 183176 14200 183288 15000 0 FreeSans 448 90 0 0 la_data_out_core[48]
port 175 nsew signal input
flabel metal2 s 185304 14200 185416 15000 0 FreeSans 448 90 0 0 la_data_out_core[49]
port 176 nsew signal input
flabel metal2 s 86968 14200 87080 15000 0 FreeSans 448 90 0 0 la_data_out_core[4]
port 177 nsew signal input
flabel metal2 s 187544 14200 187656 15000 0 FreeSans 448 90 0 0 la_data_out_core[50]
port 178 nsew signal input
flabel metal2 s 189672 14200 189784 15000 0 FreeSans 448 90 0 0 la_data_out_core[51]
port 179 nsew signal input
flabel metal2 s 191912 14200 192024 15000 0 FreeSans 448 90 0 0 la_data_out_core[52]
port 180 nsew signal input
flabel metal2 s 194040 14200 194152 15000 0 FreeSans 448 90 0 0 la_data_out_core[53]
port 181 nsew signal input
flabel metal2 s 196280 14200 196392 15000 0 FreeSans 448 90 0 0 la_data_out_core[54]
port 182 nsew signal input
flabel metal2 s 198408 14200 198520 15000 0 FreeSans 448 90 0 0 la_data_out_core[55]
port 183 nsew signal input
flabel metal2 s 200648 14200 200760 15000 0 FreeSans 448 90 0 0 la_data_out_core[56]
port 184 nsew signal input
flabel metal2 s 202776 14200 202888 15000 0 FreeSans 448 90 0 0 la_data_out_core[57]
port 185 nsew signal input
flabel metal2 s 205016 14200 205128 15000 0 FreeSans 448 90 0 0 la_data_out_core[58]
port 186 nsew signal input
flabel metal2 s 207144 14200 207256 15000 0 FreeSans 448 90 0 0 la_data_out_core[59]
port 187 nsew signal input
flabel metal2 s 89096 14200 89208 15000 0 FreeSans 448 90 0 0 la_data_out_core[5]
port 188 nsew signal input
flabel metal2 s 209384 14200 209496 15000 0 FreeSans 448 90 0 0 la_data_out_core[60]
port 189 nsew signal input
flabel metal2 s 211512 14200 211624 15000 0 FreeSans 448 90 0 0 la_data_out_core[61]
port 190 nsew signal input
flabel metal2 s 213752 14200 213864 15000 0 FreeSans 448 90 0 0 la_data_out_core[62]
port 191 nsew signal input
flabel metal2 s 215880 14200 215992 15000 0 FreeSans 448 90 0 0 la_data_out_core[63]
port 192 nsew signal input
flabel metal2 s 91336 14200 91448 15000 0 FreeSans 448 90 0 0 la_data_out_core[6]
port 193 nsew signal input
flabel metal2 s 93464 14200 93576 15000 0 FreeSans 448 90 0 0 la_data_out_core[7]
port 194 nsew signal input
flabel metal2 s 95704 14200 95816 15000 0 FreeSans 448 90 0 0 la_data_out_core[8]
port 195 nsew signal input
flabel metal2 s 97832 14200 97944 15000 0 FreeSans 448 90 0 0 la_data_out_core[9]
port 196 nsew signal input
flabel metal2 s 39144 0 39256 800 0 FreeSans 448 90 0 0 la_data_out_mprj[0]
port 197 nsew signal input
flabel metal2 s 45192 0 45304 800 0 FreeSans 448 90 0 0 la_data_out_mprj[10]
port 198 nsew signal input
flabel metal2 s 45864 0 45976 800 0 FreeSans 448 90 0 0 la_data_out_mprj[11]
port 199 nsew signal input
flabel metal2 s 46424 0 46536 800 0 FreeSans 448 90 0 0 la_data_out_mprj[12]
port 200 nsew signal input
flabel metal2 s 47096 0 47208 800 0 FreeSans 448 90 0 0 la_data_out_mprj[13]
port 201 nsew signal input
flabel metal2 s 47656 0 47768 800 0 FreeSans 448 90 0 0 la_data_out_mprj[14]
port 202 nsew signal input
flabel metal2 s 48328 0 48440 800 0 FreeSans 448 90 0 0 la_data_out_mprj[15]
port 203 nsew signal input
flabel metal2 s 48888 0 49000 800 0 FreeSans 448 90 0 0 la_data_out_mprj[16]
port 204 nsew signal input
flabel metal2 s 49448 0 49560 800 0 FreeSans 448 90 0 0 la_data_out_mprj[17]
port 205 nsew signal input
flabel metal2 s 50120 0 50232 800 0 FreeSans 448 90 0 0 la_data_out_mprj[18]
port 206 nsew signal input
flabel metal2 s 50680 0 50792 800 0 FreeSans 448 90 0 0 la_data_out_mprj[19]
port 207 nsew signal input
flabel metal2 s 39704 0 39816 800 0 FreeSans 448 90 0 0 la_data_out_mprj[1]
port 208 nsew signal input
flabel metal2 s 51352 0 51464 800 0 FreeSans 448 90 0 0 la_data_out_mprj[20]
port 209 nsew signal input
flabel metal2 s 51912 0 52024 800 0 FreeSans 448 90 0 0 la_data_out_mprj[21]
port 210 nsew signal input
flabel metal2 s 52584 0 52696 800 0 FreeSans 448 90 0 0 la_data_out_mprj[22]
port 211 nsew signal input
flabel metal2 s 53144 0 53256 800 0 FreeSans 448 90 0 0 la_data_out_mprj[23]
port 212 nsew signal input
flabel metal2 s 53816 0 53928 800 0 FreeSans 448 90 0 0 la_data_out_mprj[24]
port 213 nsew signal input
flabel metal2 s 54376 0 54488 800 0 FreeSans 448 90 0 0 la_data_out_mprj[25]
port 214 nsew signal input
flabel metal2 s 54936 0 55048 800 0 FreeSans 448 90 0 0 la_data_out_mprj[26]
port 215 nsew signal input
flabel metal2 s 55608 0 55720 800 0 FreeSans 448 90 0 0 la_data_out_mprj[27]
port 216 nsew signal input
flabel metal2 s 56168 0 56280 800 0 FreeSans 448 90 0 0 la_data_out_mprj[28]
port 217 nsew signal input
flabel metal2 s 56840 0 56952 800 0 FreeSans 448 90 0 0 la_data_out_mprj[29]
port 218 nsew signal input
flabel metal2 s 40376 0 40488 800 0 FreeSans 448 90 0 0 la_data_out_mprj[2]
port 219 nsew signal input
flabel metal2 s 57400 0 57512 800 0 FreeSans 448 90 0 0 la_data_out_mprj[30]
port 220 nsew signal input
flabel metal2 s 58072 0 58184 800 0 FreeSans 448 90 0 0 la_data_out_mprj[31]
port 221 nsew signal input
flabel metal2 s 58632 0 58744 800 0 FreeSans 448 90 0 0 la_data_out_mprj[32]
port 222 nsew signal input
flabel metal2 s 59192 0 59304 800 0 FreeSans 448 90 0 0 la_data_out_mprj[33]
port 223 nsew signal input
flabel metal2 s 59864 0 59976 800 0 FreeSans 448 90 0 0 la_data_out_mprj[34]
port 224 nsew signal input
flabel metal2 s 60424 0 60536 800 0 FreeSans 448 90 0 0 la_data_out_mprj[35]
port 225 nsew signal input
flabel metal2 s 61096 0 61208 800 0 FreeSans 448 90 0 0 la_data_out_mprj[36]
port 226 nsew signal input
flabel metal2 s 61656 0 61768 800 0 FreeSans 448 90 0 0 la_data_out_mprj[37]
port 227 nsew signal input
flabel metal2 s 62328 0 62440 800 0 FreeSans 448 90 0 0 la_data_out_mprj[38]
port 228 nsew signal input
flabel metal2 s 62888 0 63000 800 0 FreeSans 448 90 0 0 la_data_out_mprj[39]
port 229 nsew signal input
flabel metal2 s 40936 0 41048 800 0 FreeSans 448 90 0 0 la_data_out_mprj[3]
port 230 nsew signal input
flabel metal2 s 63560 0 63672 800 0 FreeSans 448 90 0 0 la_data_out_mprj[40]
port 231 nsew signal input
flabel metal2 s 64120 0 64232 800 0 FreeSans 448 90 0 0 la_data_out_mprj[41]
port 232 nsew signal input
flabel metal2 s 64680 0 64792 800 0 FreeSans 448 90 0 0 la_data_out_mprj[42]
port 233 nsew signal input
flabel metal2 s 65352 0 65464 800 0 FreeSans 448 90 0 0 la_data_out_mprj[43]
port 234 nsew signal input
flabel metal2 s 65912 0 66024 800 0 FreeSans 448 90 0 0 la_data_out_mprj[44]
port 235 nsew signal input
flabel metal2 s 66584 0 66696 800 0 FreeSans 448 90 0 0 la_data_out_mprj[45]
port 236 nsew signal input
flabel metal2 s 67144 0 67256 800 0 FreeSans 448 90 0 0 la_data_out_mprj[46]
port 237 nsew signal input
flabel metal2 s 67816 0 67928 800 0 FreeSans 448 90 0 0 la_data_out_mprj[47]
port 238 nsew signal input
flabel metal2 s 68376 0 68488 800 0 FreeSans 448 90 0 0 la_data_out_mprj[48]
port 239 nsew signal input
flabel metal2 s 69048 0 69160 800 0 FreeSans 448 90 0 0 la_data_out_mprj[49]
port 240 nsew signal input
flabel metal2 s 41608 0 41720 800 0 FreeSans 448 90 0 0 la_data_out_mprj[4]
port 241 nsew signal input
flabel metal2 s 69608 0 69720 800 0 FreeSans 448 90 0 0 la_data_out_mprj[50]
port 242 nsew signal input
flabel metal2 s 70168 0 70280 800 0 FreeSans 448 90 0 0 la_data_out_mprj[51]
port 243 nsew signal input
flabel metal2 s 70840 0 70952 800 0 FreeSans 448 90 0 0 la_data_out_mprj[52]
port 244 nsew signal input
flabel metal2 s 71400 0 71512 800 0 FreeSans 448 90 0 0 la_data_out_mprj[53]
port 245 nsew signal input
flabel metal2 s 72072 0 72184 800 0 FreeSans 448 90 0 0 la_data_out_mprj[54]
port 246 nsew signal input
flabel metal2 s 72632 0 72744 800 0 FreeSans 448 90 0 0 la_data_out_mprj[55]
port 247 nsew signal input
flabel metal2 s 73304 0 73416 800 0 FreeSans 448 90 0 0 la_data_out_mprj[56]
port 248 nsew signal input
flabel metal2 s 73864 0 73976 800 0 FreeSans 448 90 0 0 la_data_out_mprj[57]
port 249 nsew signal input
flabel metal2 s 74536 0 74648 800 0 FreeSans 448 90 0 0 la_data_out_mprj[58]
port 250 nsew signal input
flabel metal2 s 75096 0 75208 800 0 FreeSans 448 90 0 0 la_data_out_mprj[59]
port 251 nsew signal input
flabel metal2 s 42168 0 42280 800 0 FreeSans 448 90 0 0 la_data_out_mprj[5]
port 252 nsew signal input
flabel metal2 s 75656 0 75768 800 0 FreeSans 448 90 0 0 la_data_out_mprj[60]
port 253 nsew signal input
flabel metal2 s 76328 0 76440 800 0 FreeSans 448 90 0 0 la_data_out_mprj[61]
port 254 nsew signal input
flabel metal2 s 76888 0 77000 800 0 FreeSans 448 90 0 0 la_data_out_mprj[62]
port 255 nsew signal input
flabel metal2 s 77560 0 77672 800 0 FreeSans 448 90 0 0 la_data_out_mprj[63]
port 256 nsew signal input
flabel metal2 s 42840 0 42952 800 0 FreeSans 448 90 0 0 la_data_out_mprj[6]
port 257 nsew signal input
flabel metal2 s 43400 0 43512 800 0 FreeSans 448 90 0 0 la_data_out_mprj[7]
port 258 nsew signal input
flabel metal2 s 43960 0 44072 800 0 FreeSans 448 90 0 0 la_data_out_mprj[8]
port 259 nsew signal input
flabel metal2 s 44632 0 44744 800 0 FreeSans 448 90 0 0 la_data_out_mprj[9]
port 260 nsew signal input
flabel metal2 s 117208 0 117320 800 0 FreeSans 448 90 0 0 la_iena_mprj[0]
port 261 nsew signal input
flabel metal2 s 123256 0 123368 800 0 FreeSans 448 90 0 0 la_iena_mprj[10]
port 262 nsew signal input
flabel metal2 s 123816 0 123928 800 0 FreeSans 448 90 0 0 la_iena_mprj[11]
port 263 nsew signal input
flabel metal2 s 124488 0 124600 800 0 FreeSans 448 90 0 0 la_iena_mprj[12]
port 264 nsew signal input
flabel metal2 s 125048 0 125160 800 0 FreeSans 448 90 0 0 la_iena_mprj[13]
port 265 nsew signal input
flabel metal2 s 125720 0 125832 800 0 FreeSans 448 90 0 0 la_iena_mprj[14]
port 266 nsew signal input
flabel metal2 s 126280 0 126392 800 0 FreeSans 448 90 0 0 la_iena_mprj[15]
port 267 nsew signal input
flabel metal2 s 126952 0 127064 800 0 FreeSans 448 90 0 0 la_iena_mprj[16]
port 268 nsew signal input
flabel metal2 s 127512 0 127624 800 0 FreeSans 448 90 0 0 la_iena_mprj[17]
port 269 nsew signal input
flabel metal2 s 128184 0 128296 800 0 FreeSans 448 90 0 0 la_iena_mprj[18]
port 270 nsew signal input
flabel metal2 s 128744 0 128856 800 0 FreeSans 448 90 0 0 la_iena_mprj[19]
port 271 nsew signal input
flabel metal2 s 117768 0 117880 800 0 FreeSans 448 90 0 0 la_iena_mprj[1]
port 272 nsew signal input
flabel metal2 s 129304 0 129416 800 0 FreeSans 448 90 0 0 la_iena_mprj[20]
port 273 nsew signal input
flabel metal2 s 129976 0 130088 800 0 FreeSans 448 90 0 0 la_iena_mprj[21]
port 274 nsew signal input
flabel metal2 s 130536 0 130648 800 0 FreeSans 448 90 0 0 la_iena_mprj[22]
port 275 nsew signal input
flabel metal2 s 131208 0 131320 800 0 FreeSans 448 90 0 0 la_iena_mprj[23]
port 276 nsew signal input
flabel metal2 s 131768 0 131880 800 0 FreeSans 448 90 0 0 la_iena_mprj[24]
port 277 nsew signal input
flabel metal2 s 132440 0 132552 800 0 FreeSans 448 90 0 0 la_iena_mprj[25]
port 278 nsew signal input
flabel metal2 s 133000 0 133112 800 0 FreeSans 448 90 0 0 la_iena_mprj[26]
port 279 nsew signal input
flabel metal2 s 133672 0 133784 800 0 FreeSans 448 90 0 0 la_iena_mprj[27]
port 280 nsew signal input
flabel metal2 s 134232 0 134344 800 0 FreeSans 448 90 0 0 la_iena_mprj[28]
port 281 nsew signal input
flabel metal2 s 134792 0 134904 800 0 FreeSans 448 90 0 0 la_iena_mprj[29]
port 282 nsew signal input
flabel metal2 s 118328 0 118440 800 0 FreeSans 448 90 0 0 la_iena_mprj[2]
port 283 nsew signal input
flabel metal2 s 135464 0 135576 800 0 FreeSans 448 90 0 0 la_iena_mprj[30]
port 284 nsew signal input
flabel metal2 s 136024 0 136136 800 0 FreeSans 448 90 0 0 la_iena_mprj[31]
port 285 nsew signal input
flabel metal2 s 136696 0 136808 800 0 FreeSans 448 90 0 0 la_iena_mprj[32]
port 286 nsew signal input
flabel metal2 s 137256 0 137368 800 0 FreeSans 448 90 0 0 la_iena_mprj[33]
port 287 nsew signal input
flabel metal2 s 137928 0 138040 800 0 FreeSans 448 90 0 0 la_iena_mprj[34]
port 288 nsew signal input
flabel metal2 s 138488 0 138600 800 0 FreeSans 448 90 0 0 la_iena_mprj[35]
port 289 nsew signal input
flabel metal2 s 139160 0 139272 800 0 FreeSans 448 90 0 0 la_iena_mprj[36]
port 290 nsew signal input
flabel metal2 s 139720 0 139832 800 0 FreeSans 448 90 0 0 la_iena_mprj[37]
port 291 nsew signal input
flabel metal2 s 140280 0 140392 800 0 FreeSans 448 90 0 0 la_iena_mprj[38]
port 292 nsew signal input
flabel metal2 s 140952 0 141064 800 0 FreeSans 448 90 0 0 la_iena_mprj[39]
port 293 nsew signal input
flabel metal2 s 119000 0 119112 800 0 FreeSans 448 90 0 0 la_iena_mprj[3]
port 294 nsew signal input
flabel metal2 s 141512 0 141624 800 0 FreeSans 448 90 0 0 la_iena_mprj[40]
port 295 nsew signal input
flabel metal2 s 142184 0 142296 800 0 FreeSans 448 90 0 0 la_iena_mprj[41]
port 296 nsew signal input
flabel metal2 s 142744 0 142856 800 0 FreeSans 448 90 0 0 la_iena_mprj[42]
port 297 nsew signal input
flabel metal2 s 143416 0 143528 800 0 FreeSans 448 90 0 0 la_iena_mprj[43]
port 298 nsew signal input
flabel metal2 s 143976 0 144088 800 0 FreeSans 448 90 0 0 la_iena_mprj[44]
port 299 nsew signal input
flabel metal2 s 144648 0 144760 800 0 FreeSans 448 90 0 0 la_iena_mprj[45]
port 300 nsew signal input
flabel metal2 s 145208 0 145320 800 0 FreeSans 448 90 0 0 la_iena_mprj[46]
port 301 nsew signal input
flabel metal2 s 145768 0 145880 800 0 FreeSans 448 90 0 0 la_iena_mprj[47]
port 302 nsew signal input
flabel metal2 s 146440 0 146552 800 0 FreeSans 448 90 0 0 la_iena_mprj[48]
port 303 nsew signal input
flabel metal2 s 147000 0 147112 800 0 FreeSans 448 90 0 0 la_iena_mprj[49]
port 304 nsew signal input
flabel metal2 s 119560 0 119672 800 0 FreeSans 448 90 0 0 la_iena_mprj[4]
port 305 nsew signal input
flabel metal2 s 147672 0 147784 800 0 FreeSans 448 90 0 0 la_iena_mprj[50]
port 306 nsew signal input
flabel metal2 s 148232 0 148344 800 0 FreeSans 448 90 0 0 la_iena_mprj[51]
port 307 nsew signal input
flabel metal2 s 148904 0 149016 800 0 FreeSans 448 90 0 0 la_iena_mprj[52]
port 308 nsew signal input
flabel metal2 s 149464 0 149576 800 0 FreeSans 448 90 0 0 la_iena_mprj[53]
port 309 nsew signal input
flabel metal2 s 150136 0 150248 800 0 FreeSans 448 90 0 0 la_iena_mprj[54]
port 310 nsew signal input
flabel metal2 s 150696 0 150808 800 0 FreeSans 448 90 0 0 la_iena_mprj[55]
port 311 nsew signal input
flabel metal2 s 151256 0 151368 800 0 FreeSans 448 90 0 0 la_iena_mprj[56]
port 312 nsew signal input
flabel metal2 s 151928 0 152040 800 0 FreeSans 448 90 0 0 la_iena_mprj[57]
port 313 nsew signal input
flabel metal2 s 152488 0 152600 800 0 FreeSans 448 90 0 0 la_iena_mprj[58]
port 314 nsew signal input
flabel metal2 s 153160 0 153272 800 0 FreeSans 448 90 0 0 la_iena_mprj[59]
port 315 nsew signal input
flabel metal2 s 120232 0 120344 800 0 FreeSans 448 90 0 0 la_iena_mprj[5]
port 316 nsew signal input
flabel metal2 s 153720 0 153832 800 0 FreeSans 448 90 0 0 la_iena_mprj[60]
port 317 nsew signal input
flabel metal2 s 154392 0 154504 800 0 FreeSans 448 90 0 0 la_iena_mprj[61]
port 318 nsew signal input
flabel metal2 s 154952 0 155064 800 0 FreeSans 448 90 0 0 la_iena_mprj[62]
port 319 nsew signal input
flabel metal2 s 155624 0 155736 800 0 FreeSans 448 90 0 0 la_iena_mprj[63]
port 320 nsew signal input
flabel metal2 s 120792 0 120904 800 0 FreeSans 448 90 0 0 la_iena_mprj[6]
port 321 nsew signal input
flabel metal2 s 121464 0 121576 800 0 FreeSans 448 90 0 0 la_iena_mprj[7]
port 322 nsew signal input
flabel metal2 s 122024 0 122136 800 0 FreeSans 448 90 0 0 la_iena_mprj[8]
port 323 nsew signal input
flabel metal2 s 122696 0 122808 800 0 FreeSans 448 90 0 0 la_iena_mprj[9]
port 324 nsew signal input
flabel metal2 s 78904 14200 79016 15000 0 FreeSans 448 90 0 0 la_oenb_core[0]
port 325 nsew signal tristate
flabel metal2 s 100744 14200 100856 15000 0 FreeSans 448 90 0 0 la_oenb_core[10]
port 326 nsew signal tristate
flabel metal2 s 102984 14200 103096 15000 0 FreeSans 448 90 0 0 la_oenb_core[11]
port 327 nsew signal tristate
flabel metal2 s 105112 14200 105224 15000 0 FreeSans 448 90 0 0 la_oenb_core[12]
port 328 nsew signal tristate
flabel metal2 s 107352 14200 107464 15000 0 FreeSans 448 90 0 0 la_oenb_core[13]
port 329 nsew signal tristate
flabel metal2 s 109480 14200 109592 15000 0 FreeSans 448 90 0 0 la_oenb_core[14]
port 330 nsew signal tristate
flabel metal2 s 111720 14200 111832 15000 0 FreeSans 448 90 0 0 la_oenb_core[15]
port 331 nsew signal tristate
flabel metal2 s 113960 14200 114072 15000 0 FreeSans 448 90 0 0 la_oenb_core[16]
port 332 nsew signal tristate
flabel metal2 s 116088 14200 116200 15000 0 FreeSans 448 90 0 0 la_oenb_core[17]
port 333 nsew signal tristate
flabel metal2 s 118328 14200 118440 15000 0 FreeSans 448 90 0 0 la_oenb_core[18]
port 334 nsew signal tristate
flabel metal2 s 120456 14200 120568 15000 0 FreeSans 448 90 0 0 la_oenb_core[19]
port 335 nsew signal tristate
flabel metal2 s 81144 14200 81256 15000 0 FreeSans 448 90 0 0 la_oenb_core[1]
port 336 nsew signal tristate
flabel metal2 s 122696 14200 122808 15000 0 FreeSans 448 90 0 0 la_oenb_core[20]
port 337 nsew signal tristate
flabel metal2 s 124824 14200 124936 15000 0 FreeSans 448 90 0 0 la_oenb_core[21]
port 338 nsew signal tristate
flabel metal2 s 127064 14200 127176 15000 0 FreeSans 448 90 0 0 la_oenb_core[22]
port 339 nsew signal tristate
flabel metal2 s 129192 14200 129304 15000 0 FreeSans 448 90 0 0 la_oenb_core[23]
port 340 nsew signal tristate
flabel metal2 s 131432 14200 131544 15000 0 FreeSans 448 90 0 0 la_oenb_core[24]
port 341 nsew signal tristate
flabel metal2 s 133560 14200 133672 15000 0 FreeSans 448 90 0 0 la_oenb_core[25]
port 342 nsew signal tristate
flabel metal2 s 135800 14200 135912 15000 0 FreeSans 448 90 0 0 la_oenb_core[26]
port 343 nsew signal tristate
flabel metal2 s 137928 14200 138040 15000 0 FreeSans 448 90 0 0 la_oenb_core[27]
port 344 nsew signal tristate
flabel metal2 s 140168 14200 140280 15000 0 FreeSans 448 90 0 0 la_oenb_core[28]
port 345 nsew signal tristate
flabel metal2 s 142296 14200 142408 15000 0 FreeSans 448 90 0 0 la_oenb_core[29]
port 346 nsew signal tristate
flabel metal2 s 83272 14200 83384 15000 0 FreeSans 448 90 0 0 la_oenb_core[2]
port 347 nsew signal tristate
flabel metal2 s 144536 14200 144648 15000 0 FreeSans 448 90 0 0 la_oenb_core[30]
port 348 nsew signal tristate
flabel metal2 s 146664 14200 146776 15000 0 FreeSans 448 90 0 0 la_oenb_core[31]
port 349 nsew signal tristate
flabel metal2 s 148904 14200 149016 15000 0 FreeSans 448 90 0 0 la_oenb_core[32]
port 350 nsew signal tristate
flabel metal2 s 151032 14200 151144 15000 0 FreeSans 448 90 0 0 la_oenb_core[33]
port 351 nsew signal tristate
flabel metal2 s 153272 14200 153384 15000 0 FreeSans 448 90 0 0 la_oenb_core[34]
port 352 nsew signal tristate
flabel metal2 s 155400 14200 155512 15000 0 FreeSans 448 90 0 0 la_oenb_core[35]
port 353 nsew signal tristate
flabel metal2 s 157640 14200 157752 15000 0 FreeSans 448 90 0 0 la_oenb_core[36]
port 354 nsew signal tristate
flabel metal2 s 159768 14200 159880 15000 0 FreeSans 448 90 0 0 la_oenb_core[37]
port 355 nsew signal tristate
flabel metal2 s 162008 14200 162120 15000 0 FreeSans 448 90 0 0 la_oenb_core[38]
port 356 nsew signal tristate
flabel metal2 s 164136 14200 164248 15000 0 FreeSans 448 90 0 0 la_oenb_core[39]
port 357 nsew signal tristate
flabel metal2 s 85512 14200 85624 15000 0 FreeSans 448 90 0 0 la_oenb_core[3]
port 358 nsew signal tristate
flabel metal2 s 166376 14200 166488 15000 0 FreeSans 448 90 0 0 la_oenb_core[40]
port 359 nsew signal tristate
flabel metal2 s 168616 14200 168728 15000 0 FreeSans 448 90 0 0 la_oenb_core[41]
port 360 nsew signal tristate
flabel metal2 s 170744 14200 170856 15000 0 FreeSans 448 90 0 0 la_oenb_core[42]
port 361 nsew signal tristate
flabel metal2 s 172984 14200 173096 15000 0 FreeSans 448 90 0 0 la_oenb_core[43]
port 362 nsew signal tristate
flabel metal2 s 175112 14200 175224 15000 0 FreeSans 448 90 0 0 la_oenb_core[44]
port 363 nsew signal tristate
flabel metal2 s 177352 14200 177464 15000 0 FreeSans 448 90 0 0 la_oenb_core[45]
port 364 nsew signal tristate
flabel metal2 s 179480 14200 179592 15000 0 FreeSans 448 90 0 0 la_oenb_core[46]
port 365 nsew signal tristate
flabel metal2 s 181720 14200 181832 15000 0 FreeSans 448 90 0 0 la_oenb_core[47]
port 366 nsew signal tristate
flabel metal2 s 183848 14200 183960 15000 0 FreeSans 448 90 0 0 la_oenb_core[48]
port 367 nsew signal tristate
flabel metal2 s 186088 14200 186200 15000 0 FreeSans 448 90 0 0 la_oenb_core[49]
port 368 nsew signal tristate
flabel metal2 s 87640 14200 87752 15000 0 FreeSans 448 90 0 0 la_oenb_core[4]
port 369 nsew signal tristate
flabel metal2 s 188216 14200 188328 15000 0 FreeSans 448 90 0 0 la_oenb_core[50]
port 370 nsew signal tristate
flabel metal2 s 190456 14200 190568 15000 0 FreeSans 448 90 0 0 la_oenb_core[51]
port 371 nsew signal tristate
flabel metal2 s 192584 14200 192696 15000 0 FreeSans 448 90 0 0 la_oenb_core[52]
port 372 nsew signal tristate
flabel metal2 s 194824 14200 194936 15000 0 FreeSans 448 90 0 0 la_oenb_core[53]
port 373 nsew signal tristate
flabel metal2 s 196952 14200 197064 15000 0 FreeSans 448 90 0 0 la_oenb_core[54]
port 374 nsew signal tristate
flabel metal2 s 199192 14200 199304 15000 0 FreeSans 448 90 0 0 la_oenb_core[55]
port 375 nsew signal tristate
flabel metal2 s 201320 14200 201432 15000 0 FreeSans 448 90 0 0 la_oenb_core[56]
port 376 nsew signal tristate
flabel metal2 s 203560 14200 203672 15000 0 FreeSans 448 90 0 0 la_oenb_core[57]
port 377 nsew signal tristate
flabel metal2 s 205688 14200 205800 15000 0 FreeSans 448 90 0 0 la_oenb_core[58]
port 378 nsew signal tristate
flabel metal2 s 207928 14200 208040 15000 0 FreeSans 448 90 0 0 la_oenb_core[59]
port 379 nsew signal tristate
flabel metal2 s 89880 14200 89992 15000 0 FreeSans 448 90 0 0 la_oenb_core[5]
port 380 nsew signal tristate
flabel metal2 s 210056 14200 210168 15000 0 FreeSans 448 90 0 0 la_oenb_core[60]
port 381 nsew signal tristate
flabel metal2 s 212296 14200 212408 15000 0 FreeSans 448 90 0 0 la_oenb_core[61]
port 382 nsew signal tristate
flabel metal2 s 214424 14200 214536 15000 0 FreeSans 448 90 0 0 la_oenb_core[62]
port 383 nsew signal tristate
flabel metal2 s 216664 14200 216776 15000 0 FreeSans 448 90 0 0 la_oenb_core[63]
port 384 nsew signal tristate
flabel metal2 s 92008 14200 92120 15000 0 FreeSans 448 90 0 0 la_oenb_core[6]
port 385 nsew signal tristate
flabel metal2 s 94248 14200 94360 15000 0 FreeSans 448 90 0 0 la_oenb_core[7]
port 386 nsew signal tristate
flabel metal2 s 96376 14200 96488 15000 0 FreeSans 448 90 0 0 la_oenb_core[8]
port 387 nsew signal tristate
flabel metal2 s 98616 14200 98728 15000 0 FreeSans 448 90 0 0 la_oenb_core[9]
port 388 nsew signal tristate
flabel metal2 s 78120 0 78232 800 0 FreeSans 448 90 0 0 la_oenb_mprj[0]
port 389 nsew signal input
flabel metal2 s 84280 0 84392 800 0 FreeSans 448 90 0 0 la_oenb_mprj[10]
port 390 nsew signal input
flabel metal2 s 84840 0 84952 800 0 FreeSans 448 90 0 0 la_oenb_mprj[11]
port 391 nsew signal input
flabel metal2 s 85512 0 85624 800 0 FreeSans 448 90 0 0 la_oenb_mprj[12]
port 392 nsew signal input
flabel metal2 s 86072 0 86184 800 0 FreeSans 448 90 0 0 la_oenb_mprj[13]
port 393 nsew signal input
flabel metal2 s 86632 0 86744 800 0 FreeSans 448 90 0 0 la_oenb_mprj[14]
port 394 nsew signal input
flabel metal2 s 87304 0 87416 800 0 FreeSans 448 90 0 0 la_oenb_mprj[15]
port 395 nsew signal input
flabel metal2 s 87864 0 87976 800 0 FreeSans 448 90 0 0 la_oenb_mprj[16]
port 396 nsew signal input
flabel metal2 s 88536 0 88648 800 0 FreeSans 448 90 0 0 la_oenb_mprj[17]
port 397 nsew signal input
flabel metal2 s 89096 0 89208 800 0 FreeSans 448 90 0 0 la_oenb_mprj[18]
port 398 nsew signal input
flabel metal2 s 89768 0 89880 800 0 FreeSans 448 90 0 0 la_oenb_mprj[19]
port 399 nsew signal input
flabel metal2 s 78792 0 78904 800 0 FreeSans 448 90 0 0 la_oenb_mprj[1]
port 400 nsew signal input
flabel metal2 s 90328 0 90440 800 0 FreeSans 448 90 0 0 la_oenb_mprj[20]
port 401 nsew signal input
flabel metal2 s 91000 0 91112 800 0 FreeSans 448 90 0 0 la_oenb_mprj[21]
port 402 nsew signal input
flabel metal2 s 91560 0 91672 800 0 FreeSans 448 90 0 0 la_oenb_mprj[22]
port 403 nsew signal input
flabel metal2 s 92120 0 92232 800 0 FreeSans 448 90 0 0 la_oenb_mprj[23]
port 404 nsew signal input
flabel metal2 s 92792 0 92904 800 0 FreeSans 448 90 0 0 la_oenb_mprj[24]
port 405 nsew signal input
flabel metal2 s 93352 0 93464 800 0 FreeSans 448 90 0 0 la_oenb_mprj[25]
port 406 nsew signal input
flabel metal2 s 94024 0 94136 800 0 FreeSans 448 90 0 0 la_oenb_mprj[26]
port 407 nsew signal input
flabel metal2 s 94584 0 94696 800 0 FreeSans 448 90 0 0 la_oenb_mprj[27]
port 408 nsew signal input
flabel metal2 s 95256 0 95368 800 0 FreeSans 448 90 0 0 la_oenb_mprj[28]
port 409 nsew signal input
flabel metal2 s 95816 0 95928 800 0 FreeSans 448 90 0 0 la_oenb_mprj[29]
port 410 nsew signal input
flabel metal2 s 79352 0 79464 800 0 FreeSans 448 90 0 0 la_oenb_mprj[2]
port 411 nsew signal input
flabel metal2 s 96488 0 96600 800 0 FreeSans 448 90 0 0 la_oenb_mprj[30]
port 412 nsew signal input
flabel metal2 s 97048 0 97160 800 0 FreeSans 448 90 0 0 la_oenb_mprj[31]
port 413 nsew signal input
flabel metal2 s 97608 0 97720 800 0 FreeSans 448 90 0 0 la_oenb_mprj[32]
port 414 nsew signal input
flabel metal2 s 98280 0 98392 800 0 FreeSans 448 90 0 0 la_oenb_mprj[33]
port 415 nsew signal input
flabel metal2 s 98840 0 98952 800 0 FreeSans 448 90 0 0 la_oenb_mprj[34]
port 416 nsew signal input
flabel metal2 s 99512 0 99624 800 0 FreeSans 448 90 0 0 la_oenb_mprj[35]
port 417 nsew signal input
flabel metal2 s 100072 0 100184 800 0 FreeSans 448 90 0 0 la_oenb_mprj[36]
port 418 nsew signal input
flabel metal2 s 100744 0 100856 800 0 FreeSans 448 90 0 0 la_oenb_mprj[37]
port 419 nsew signal input
flabel metal2 s 101304 0 101416 800 0 FreeSans 448 90 0 0 la_oenb_mprj[38]
port 420 nsew signal input
flabel metal2 s 101976 0 102088 800 0 FreeSans 448 90 0 0 la_oenb_mprj[39]
port 421 nsew signal input
flabel metal2 s 80024 0 80136 800 0 FreeSans 448 90 0 0 la_oenb_mprj[3]
port 422 nsew signal input
flabel metal2 s 102536 0 102648 800 0 FreeSans 448 90 0 0 la_oenb_mprj[40]
port 423 nsew signal input
flabel metal2 s 103096 0 103208 800 0 FreeSans 448 90 0 0 la_oenb_mprj[41]
port 424 nsew signal input
flabel metal2 s 103768 0 103880 800 0 FreeSans 448 90 0 0 la_oenb_mprj[42]
port 425 nsew signal input
flabel metal2 s 104328 0 104440 800 0 FreeSans 448 90 0 0 la_oenb_mprj[43]
port 426 nsew signal input
flabel metal2 s 105000 0 105112 800 0 FreeSans 448 90 0 0 la_oenb_mprj[44]
port 427 nsew signal input
flabel metal2 s 105560 0 105672 800 0 FreeSans 448 90 0 0 la_oenb_mprj[45]
port 428 nsew signal input
flabel metal2 s 106232 0 106344 800 0 FreeSans 448 90 0 0 la_oenb_mprj[46]
port 429 nsew signal input
flabel metal2 s 106792 0 106904 800 0 FreeSans 448 90 0 0 la_oenb_mprj[47]
port 430 nsew signal input
flabel metal2 s 107464 0 107576 800 0 FreeSans 448 90 0 0 la_oenb_mprj[48]
port 431 nsew signal input
flabel metal2 s 108024 0 108136 800 0 FreeSans 448 90 0 0 la_oenb_mprj[49]
port 432 nsew signal input
flabel metal2 s 80584 0 80696 800 0 FreeSans 448 90 0 0 la_oenb_mprj[4]
port 433 nsew signal input
flabel metal2 s 108584 0 108696 800 0 FreeSans 448 90 0 0 la_oenb_mprj[50]
port 434 nsew signal input
flabel metal2 s 109256 0 109368 800 0 FreeSans 448 90 0 0 la_oenb_mprj[51]
port 435 nsew signal input
flabel metal2 s 109816 0 109928 800 0 FreeSans 448 90 0 0 la_oenb_mprj[52]
port 436 nsew signal input
flabel metal2 s 110488 0 110600 800 0 FreeSans 448 90 0 0 la_oenb_mprj[53]
port 437 nsew signal input
flabel metal2 s 111048 0 111160 800 0 FreeSans 448 90 0 0 la_oenb_mprj[54]
port 438 nsew signal input
flabel metal2 s 111720 0 111832 800 0 FreeSans 448 90 0 0 la_oenb_mprj[55]
port 439 nsew signal input
flabel metal2 s 112280 0 112392 800 0 FreeSans 448 90 0 0 la_oenb_mprj[56]
port 440 nsew signal input
flabel metal2 s 112840 0 112952 800 0 FreeSans 448 90 0 0 la_oenb_mprj[57]
port 441 nsew signal input
flabel metal2 s 113512 0 113624 800 0 FreeSans 448 90 0 0 la_oenb_mprj[58]
port 442 nsew signal input
flabel metal2 s 114072 0 114184 800 0 FreeSans 448 90 0 0 la_oenb_mprj[59]
port 443 nsew signal input
flabel metal2 s 81144 0 81256 800 0 FreeSans 448 90 0 0 la_oenb_mprj[5]
port 444 nsew signal input
flabel metal2 s 114744 0 114856 800 0 FreeSans 448 90 0 0 la_oenb_mprj[60]
port 445 nsew signal input
flabel metal2 s 115304 0 115416 800 0 FreeSans 448 90 0 0 la_oenb_mprj[61]
port 446 nsew signal input
flabel metal2 s 115976 0 116088 800 0 FreeSans 448 90 0 0 la_oenb_mprj[62]
port 447 nsew signal input
flabel metal2 s 116536 0 116648 800 0 FreeSans 448 90 0 0 la_oenb_mprj[63]
port 448 nsew signal input
flabel metal2 s 81816 0 81928 800 0 FreeSans 448 90 0 0 la_oenb_mprj[6]
port 449 nsew signal input
flabel metal2 s 82376 0 82488 800 0 FreeSans 448 90 0 0 la_oenb_mprj[7]
port 450 nsew signal input
flabel metal2 s 83048 0 83160 800 0 FreeSans 448 90 0 0 la_oenb_mprj[8]
port 451 nsew signal input
flabel metal2 s 83608 0 83720 800 0 FreeSans 448 90 0 0 la_oenb_mprj[9]
port 452 nsew signal input
flabel metal2 s 219016 0 219128 800 0 FreeSans 448 90 0 0 mprj_ack_i_core
port 453 nsew signal tristate
flabel metal2 s 1736 14200 1848 15000 0 FreeSans 448 90 0 0 mprj_ack_i_user
port 454 nsew signal input
flabel metal2 s 178136 0 178248 800 0 FreeSans 448 90 0 0 mprj_adr_o_core[0]
port 455 nsew signal input
flabel metal2 s 184184 0 184296 800 0 FreeSans 448 90 0 0 mprj_adr_o_core[10]
port 456 nsew signal input
flabel metal2 s 184856 0 184968 800 0 FreeSans 448 90 0 0 mprj_adr_o_core[11]
port 457 nsew signal input
flabel metal2 s 185416 0 185528 800 0 FreeSans 448 90 0 0 mprj_adr_o_core[12]
port 458 nsew signal input
flabel metal2 s 186088 0 186200 800 0 FreeSans 448 90 0 0 mprj_adr_o_core[13]
port 459 nsew signal input
flabel metal2 s 186648 0 186760 800 0 FreeSans 448 90 0 0 mprj_adr_o_core[14]
port 460 nsew signal input
flabel metal2 s 187320 0 187432 800 0 FreeSans 448 90 0 0 mprj_adr_o_core[15]
port 461 nsew signal input
flabel metal2 s 187880 0 187992 800 0 FreeSans 448 90 0 0 mprj_adr_o_core[16]
port 462 nsew signal input
flabel metal2 s 188440 0 188552 800 0 FreeSans 448 90 0 0 mprj_adr_o_core[17]
port 463 nsew signal input
flabel metal2 s 189112 0 189224 800 0 FreeSans 448 90 0 0 mprj_adr_o_core[18]
port 464 nsew signal input
flabel metal2 s 189672 0 189784 800 0 FreeSans 448 90 0 0 mprj_adr_o_core[19]
port 465 nsew signal input
flabel metal2 s 178696 0 178808 800 0 FreeSans 448 90 0 0 mprj_adr_o_core[1]
port 466 nsew signal input
flabel metal2 s 190344 0 190456 800 0 FreeSans 448 90 0 0 mprj_adr_o_core[20]
port 467 nsew signal input
flabel metal2 s 190904 0 191016 800 0 FreeSans 448 90 0 0 mprj_adr_o_core[21]
port 468 nsew signal input
flabel metal2 s 191576 0 191688 800 0 FreeSans 448 90 0 0 mprj_adr_o_core[22]
port 469 nsew signal input
flabel metal2 s 192136 0 192248 800 0 FreeSans 448 90 0 0 mprj_adr_o_core[23]
port 470 nsew signal input
flabel metal2 s 192808 0 192920 800 0 FreeSans 448 90 0 0 mprj_adr_o_core[24]
port 471 nsew signal input
flabel metal2 s 193368 0 193480 800 0 FreeSans 448 90 0 0 mprj_adr_o_core[25]
port 472 nsew signal input
flabel metal2 s 193928 0 194040 800 0 FreeSans 448 90 0 0 mprj_adr_o_core[26]
port 473 nsew signal input
flabel metal2 s 194600 0 194712 800 0 FreeSans 448 90 0 0 mprj_adr_o_core[27]
port 474 nsew signal input
flabel metal2 s 195160 0 195272 800 0 FreeSans 448 90 0 0 mprj_adr_o_core[28]
port 475 nsew signal input
flabel metal2 s 195832 0 195944 800 0 FreeSans 448 90 0 0 mprj_adr_o_core[29]
port 476 nsew signal input
flabel metal2 s 179368 0 179480 800 0 FreeSans 448 90 0 0 mprj_adr_o_core[2]
port 477 nsew signal input
flabel metal2 s 196392 0 196504 800 0 FreeSans 448 90 0 0 mprj_adr_o_core[30]
port 478 nsew signal input
flabel metal2 s 197064 0 197176 800 0 FreeSans 448 90 0 0 mprj_adr_o_core[31]
port 479 nsew signal input
flabel metal2 s 179928 0 180040 800 0 FreeSans 448 90 0 0 mprj_adr_o_core[3]
port 480 nsew signal input
flabel metal2 s 180600 0 180712 800 0 FreeSans 448 90 0 0 mprj_adr_o_core[4]
port 481 nsew signal input
flabel metal2 s 181160 0 181272 800 0 FreeSans 448 90 0 0 mprj_adr_o_core[5]
port 482 nsew signal input
flabel metal2 s 181832 0 181944 800 0 FreeSans 448 90 0 0 mprj_adr_o_core[6]
port 483 nsew signal input
flabel metal2 s 182392 0 182504 800 0 FreeSans 448 90 0 0 mprj_adr_o_core[7]
port 484 nsew signal input
flabel metal2 s 182952 0 183064 800 0 FreeSans 448 90 0 0 mprj_adr_o_core[8]
port 485 nsew signal input
flabel metal2 s 183624 0 183736 800 0 FreeSans 448 90 0 0 mprj_adr_o_core[9]
port 486 nsew signal input
flabel metal2 s 4648 14200 4760 15000 0 FreeSans 448 90 0 0 mprj_adr_o_user[0]
port 487 nsew signal tristate
flabel metal2 s 29400 14200 29512 15000 0 FreeSans 448 90 0 0 mprj_adr_o_user[10]
port 488 nsew signal tristate
flabel metal2 s 31528 14200 31640 15000 0 FreeSans 448 90 0 0 mprj_adr_o_user[11]
port 489 nsew signal tristate
flabel metal2 s 33768 14200 33880 15000 0 FreeSans 448 90 0 0 mprj_adr_o_user[12]
port 490 nsew signal tristate
flabel metal2 s 35896 14200 36008 15000 0 FreeSans 448 90 0 0 mprj_adr_o_user[13]
port 491 nsew signal tristate
flabel metal2 s 38136 14200 38248 15000 0 FreeSans 448 90 0 0 mprj_adr_o_user[14]
port 492 nsew signal tristate
flabel metal2 s 40264 14200 40376 15000 0 FreeSans 448 90 0 0 mprj_adr_o_user[15]
port 493 nsew signal tristate
flabel metal2 s 42504 14200 42616 15000 0 FreeSans 448 90 0 0 mprj_adr_o_user[16]
port 494 nsew signal tristate
flabel metal2 s 44632 14200 44744 15000 0 FreeSans 448 90 0 0 mprj_adr_o_user[17]
port 495 nsew signal tristate
flabel metal2 s 46872 14200 46984 15000 0 FreeSans 448 90 0 0 mprj_adr_o_user[18]
port 496 nsew signal tristate
flabel metal2 s 49000 14200 49112 15000 0 FreeSans 448 90 0 0 mprj_adr_o_user[19]
port 497 nsew signal tristate
flabel metal2 s 7560 14200 7672 15000 0 FreeSans 448 90 0 0 mprj_adr_o_user[1]
port 498 nsew signal tristate
flabel metal2 s 51240 14200 51352 15000 0 FreeSans 448 90 0 0 mprj_adr_o_user[20]
port 499 nsew signal tristate
flabel metal2 s 53368 14200 53480 15000 0 FreeSans 448 90 0 0 mprj_adr_o_user[21]
port 500 nsew signal tristate
flabel metal2 s 55608 14200 55720 15000 0 FreeSans 448 90 0 0 mprj_adr_o_user[22]
port 501 nsew signal tristate
flabel metal2 s 57848 14200 57960 15000 0 FreeSans 448 90 0 0 mprj_adr_o_user[23]
port 502 nsew signal tristate
flabel metal2 s 59976 14200 60088 15000 0 FreeSans 448 90 0 0 mprj_adr_o_user[24]
port 503 nsew signal tristate
flabel metal2 s 62216 14200 62328 15000 0 FreeSans 448 90 0 0 mprj_adr_o_user[25]
port 504 nsew signal tristate
flabel metal2 s 64344 14200 64456 15000 0 FreeSans 448 90 0 0 mprj_adr_o_user[26]
port 505 nsew signal tristate
flabel metal2 s 66584 14200 66696 15000 0 FreeSans 448 90 0 0 mprj_adr_o_user[27]
port 506 nsew signal tristate
flabel metal2 s 68712 14200 68824 15000 0 FreeSans 448 90 0 0 mprj_adr_o_user[28]
port 507 nsew signal tristate
flabel metal2 s 70952 14200 71064 15000 0 FreeSans 448 90 0 0 mprj_adr_o_user[29]
port 508 nsew signal tristate
flabel metal2 s 10472 14200 10584 15000 0 FreeSans 448 90 0 0 mprj_adr_o_user[2]
port 509 nsew signal tristate
flabel metal2 s 73080 14200 73192 15000 0 FreeSans 448 90 0 0 mprj_adr_o_user[30]
port 510 nsew signal tristate
flabel metal2 s 75320 14200 75432 15000 0 FreeSans 448 90 0 0 mprj_adr_o_user[31]
port 511 nsew signal tristate
flabel metal2 s 13384 14200 13496 15000 0 FreeSans 448 90 0 0 mprj_adr_o_user[3]
port 512 nsew signal tristate
flabel metal2 s 16296 14200 16408 15000 0 FreeSans 448 90 0 0 mprj_adr_o_user[4]
port 513 nsew signal tristate
flabel metal2 s 18424 14200 18536 15000 0 FreeSans 448 90 0 0 mprj_adr_o_user[5]
port 514 nsew signal tristate
flabel metal2 s 20664 14200 20776 15000 0 FreeSans 448 90 0 0 mprj_adr_o_user[6]
port 515 nsew signal tristate
flabel metal2 s 22792 14200 22904 15000 0 FreeSans 448 90 0 0 mprj_adr_o_user[7]
port 516 nsew signal tristate
flabel metal2 s 25032 14200 25144 15000 0 FreeSans 448 90 0 0 mprj_adr_o_user[8]
port 517 nsew signal tristate
flabel metal2 s 27160 14200 27272 15000 0 FreeSans 448 90 0 0 mprj_adr_o_user[9]
port 518 nsew signal tristate
flabel metal2 s 217784 0 217896 800 0 FreeSans 448 90 0 0 mprj_cyc_o_core
port 519 nsew signal input
flabel metal2 s 2408 14200 2520 15000 0 FreeSans 448 90 0 0 mprj_cyc_o_user
port 520 nsew signal tristate
flabel metal2 s 156184 0 156296 800 0 FreeSans 448 90 0 0 mprj_dat_i_core[0]
port 521 nsew signal tristate
flabel metal2 s 162232 0 162344 800 0 FreeSans 448 90 0 0 mprj_dat_i_core[10]
port 522 nsew signal tristate
flabel metal2 s 162904 0 163016 800 0 FreeSans 448 90 0 0 mprj_dat_i_core[11]
port 523 nsew signal tristate
flabel metal2 s 163464 0 163576 800 0 FreeSans 448 90 0 0 mprj_dat_i_core[12]
port 524 nsew signal tristate
flabel metal2 s 164136 0 164248 800 0 FreeSans 448 90 0 0 mprj_dat_i_core[13]
port 525 nsew signal tristate
flabel metal2 s 164696 0 164808 800 0 FreeSans 448 90 0 0 mprj_dat_i_core[14]
port 526 nsew signal tristate
flabel metal2 s 165368 0 165480 800 0 FreeSans 448 90 0 0 mprj_dat_i_core[15]
port 527 nsew signal tristate
flabel metal2 s 165928 0 166040 800 0 FreeSans 448 90 0 0 mprj_dat_i_core[16]
port 528 nsew signal tristate
flabel metal2 s 166488 0 166600 800 0 FreeSans 448 90 0 0 mprj_dat_i_core[17]
port 529 nsew signal tristate
flabel metal2 s 167160 0 167272 800 0 FreeSans 448 90 0 0 mprj_dat_i_core[18]
port 530 nsew signal tristate
flabel metal2 s 167720 0 167832 800 0 FreeSans 448 90 0 0 mprj_dat_i_core[19]
port 531 nsew signal tristate
flabel metal2 s 156744 0 156856 800 0 FreeSans 448 90 0 0 mprj_dat_i_core[1]
port 532 nsew signal tristate
flabel metal2 s 168392 0 168504 800 0 FreeSans 448 90 0 0 mprj_dat_i_core[20]
port 533 nsew signal tristate
flabel metal2 s 168952 0 169064 800 0 FreeSans 448 90 0 0 mprj_dat_i_core[21]
port 534 nsew signal tristate
flabel metal2 s 169624 0 169736 800 0 FreeSans 448 90 0 0 mprj_dat_i_core[22]
port 535 nsew signal tristate
flabel metal2 s 170184 0 170296 800 0 FreeSans 448 90 0 0 mprj_dat_i_core[23]
port 536 nsew signal tristate
flabel metal2 s 170856 0 170968 800 0 FreeSans 448 90 0 0 mprj_dat_i_core[24]
port 537 nsew signal tristate
flabel metal2 s 171416 0 171528 800 0 FreeSans 448 90 0 0 mprj_dat_i_core[25]
port 538 nsew signal tristate
flabel metal2 s 171976 0 172088 800 0 FreeSans 448 90 0 0 mprj_dat_i_core[26]
port 539 nsew signal tristate
flabel metal2 s 172648 0 172760 800 0 FreeSans 448 90 0 0 mprj_dat_i_core[27]
port 540 nsew signal tristate
flabel metal2 s 173208 0 173320 800 0 FreeSans 448 90 0 0 mprj_dat_i_core[28]
port 541 nsew signal tristate
flabel metal2 s 173880 0 173992 800 0 FreeSans 448 90 0 0 mprj_dat_i_core[29]
port 542 nsew signal tristate
flabel metal2 s 157416 0 157528 800 0 FreeSans 448 90 0 0 mprj_dat_i_core[2]
port 543 nsew signal tristate
flabel metal2 s 174440 0 174552 800 0 FreeSans 448 90 0 0 mprj_dat_i_core[30]
port 544 nsew signal tristate
flabel metal2 s 175112 0 175224 800 0 FreeSans 448 90 0 0 mprj_dat_i_core[31]
port 545 nsew signal tristate
flabel metal2 s 157976 0 158088 800 0 FreeSans 448 90 0 0 mprj_dat_i_core[3]
port 546 nsew signal tristate
flabel metal2 s 158648 0 158760 800 0 FreeSans 448 90 0 0 mprj_dat_i_core[4]
port 547 nsew signal tristate
flabel metal2 s 159208 0 159320 800 0 FreeSans 448 90 0 0 mprj_dat_i_core[5]
port 548 nsew signal tristate
flabel metal2 s 159880 0 159992 800 0 FreeSans 448 90 0 0 mprj_dat_i_core[6]
port 549 nsew signal tristate
flabel metal2 s 160440 0 160552 800 0 FreeSans 448 90 0 0 mprj_dat_i_core[7]
port 550 nsew signal tristate
flabel metal2 s 161112 0 161224 800 0 FreeSans 448 90 0 0 mprj_dat_i_core[8]
port 551 nsew signal tristate
flabel metal2 s 161672 0 161784 800 0 FreeSans 448 90 0 0 mprj_dat_i_core[9]
port 552 nsew signal tristate
flabel metal2 s 5320 14200 5432 15000 0 FreeSans 448 90 0 0 mprj_dat_i_user[0]
port 553 nsew signal input
flabel metal2 s 30072 14200 30184 15000 0 FreeSans 448 90 0 0 mprj_dat_i_user[10]
port 554 nsew signal input
flabel metal2 s 32312 14200 32424 15000 0 FreeSans 448 90 0 0 mprj_dat_i_user[11]
port 555 nsew signal input
flabel metal2 s 34440 14200 34552 15000 0 FreeSans 448 90 0 0 mprj_dat_i_user[12]
port 556 nsew signal input
flabel metal2 s 36680 14200 36792 15000 0 FreeSans 448 90 0 0 mprj_dat_i_user[13]
port 557 nsew signal input
flabel metal2 s 38808 14200 38920 15000 0 FreeSans 448 90 0 0 mprj_dat_i_user[14]
port 558 nsew signal input
flabel metal2 s 41048 14200 41160 15000 0 FreeSans 448 90 0 0 mprj_dat_i_user[15]
port 559 nsew signal input
flabel metal2 s 43176 14200 43288 15000 0 FreeSans 448 90 0 0 mprj_dat_i_user[16]
port 560 nsew signal input
flabel metal2 s 45416 14200 45528 15000 0 FreeSans 448 90 0 0 mprj_dat_i_user[17]
port 561 nsew signal input
flabel metal2 s 47544 14200 47656 15000 0 FreeSans 448 90 0 0 mprj_dat_i_user[18]
port 562 nsew signal input
flabel metal2 s 49784 14200 49896 15000 0 FreeSans 448 90 0 0 mprj_dat_i_user[19]
port 563 nsew signal input
flabel metal2 s 8232 14200 8344 15000 0 FreeSans 448 90 0 0 mprj_dat_i_user[1]
port 564 nsew signal input
flabel metal2 s 51912 14200 52024 15000 0 FreeSans 448 90 0 0 mprj_dat_i_user[20]
port 565 nsew signal input
flabel metal2 s 54152 14200 54264 15000 0 FreeSans 448 90 0 0 mprj_dat_i_user[21]
port 566 nsew signal input
flabel metal2 s 56392 14200 56504 15000 0 FreeSans 448 90 0 0 mprj_dat_i_user[22]
port 567 nsew signal input
flabel metal2 s 58520 14200 58632 15000 0 FreeSans 448 90 0 0 mprj_dat_i_user[23]
port 568 nsew signal input
flabel metal2 s 60760 14200 60872 15000 0 FreeSans 448 90 0 0 mprj_dat_i_user[24]
port 569 nsew signal input
flabel metal2 s 62888 14200 63000 15000 0 FreeSans 448 90 0 0 mprj_dat_i_user[25]
port 570 nsew signal input
flabel metal2 s 65128 14200 65240 15000 0 FreeSans 448 90 0 0 mprj_dat_i_user[26]
port 571 nsew signal input
flabel metal2 s 67256 14200 67368 15000 0 FreeSans 448 90 0 0 mprj_dat_i_user[27]
port 572 nsew signal input
flabel metal2 s 69496 14200 69608 15000 0 FreeSans 448 90 0 0 mprj_dat_i_user[28]
port 573 nsew signal input
flabel metal2 s 71624 14200 71736 15000 0 FreeSans 448 90 0 0 mprj_dat_i_user[29]
port 574 nsew signal input
flabel metal2 s 11144 14200 11256 15000 0 FreeSans 448 90 0 0 mprj_dat_i_user[2]
port 575 nsew signal input
flabel metal2 s 73864 14200 73976 15000 0 FreeSans 448 90 0 0 mprj_dat_i_user[30]
port 576 nsew signal input
flabel metal2 s 75992 14200 76104 15000 0 FreeSans 448 90 0 0 mprj_dat_i_user[31]
port 577 nsew signal input
flabel metal2 s 14056 14200 14168 15000 0 FreeSans 448 90 0 0 mprj_dat_i_user[3]
port 578 nsew signal input
flabel metal2 s 16968 14200 17080 15000 0 FreeSans 448 90 0 0 mprj_dat_i_user[4]
port 579 nsew signal input
flabel metal2 s 19208 14200 19320 15000 0 FreeSans 448 90 0 0 mprj_dat_i_user[5]
port 580 nsew signal input
flabel metal2 s 21336 14200 21448 15000 0 FreeSans 448 90 0 0 mprj_dat_i_user[6]
port 581 nsew signal input
flabel metal2 s 23576 14200 23688 15000 0 FreeSans 448 90 0 0 mprj_dat_i_user[7]
port 582 nsew signal input
flabel metal2 s 25704 14200 25816 15000 0 FreeSans 448 90 0 0 mprj_dat_i_user[8]
port 583 nsew signal input
flabel metal2 s 27944 14200 28056 15000 0 FreeSans 448 90 0 0 mprj_dat_i_user[9]
port 584 nsew signal input
flabel metal2 s 197624 0 197736 800 0 FreeSans 448 90 0 0 mprj_dat_o_core[0]
port 585 nsew signal input
flabel metal2 s 203784 0 203896 800 0 FreeSans 448 90 0 0 mprj_dat_o_core[10]
port 586 nsew signal input
flabel metal2 s 204344 0 204456 800 0 FreeSans 448 90 0 0 mprj_dat_o_core[11]
port 587 nsew signal input
flabel metal2 s 204904 0 205016 800 0 FreeSans 448 90 0 0 mprj_dat_o_core[12]
port 588 nsew signal input
flabel metal2 s 205576 0 205688 800 0 FreeSans 448 90 0 0 mprj_dat_o_core[13]
port 589 nsew signal input
flabel metal2 s 206136 0 206248 800 0 FreeSans 448 90 0 0 mprj_dat_o_core[14]
port 590 nsew signal input
flabel metal2 s 206808 0 206920 800 0 FreeSans 448 90 0 0 mprj_dat_o_core[15]
port 591 nsew signal input
flabel metal2 s 207368 0 207480 800 0 FreeSans 448 90 0 0 mprj_dat_o_core[16]
port 592 nsew signal input
flabel metal2 s 208040 0 208152 800 0 FreeSans 448 90 0 0 mprj_dat_o_core[17]
port 593 nsew signal input
flabel metal2 s 208600 0 208712 800 0 FreeSans 448 90 0 0 mprj_dat_o_core[18]
port 594 nsew signal input
flabel metal2 s 209272 0 209384 800 0 FreeSans 448 90 0 0 mprj_dat_o_core[19]
port 595 nsew signal input
flabel metal2 s 198296 0 198408 800 0 FreeSans 448 90 0 0 mprj_dat_o_core[1]
port 596 nsew signal input
flabel metal2 s 209832 0 209944 800 0 FreeSans 448 90 0 0 mprj_dat_o_core[20]
port 597 nsew signal input
flabel metal2 s 210392 0 210504 800 0 FreeSans 448 90 0 0 mprj_dat_o_core[21]
port 598 nsew signal input
flabel metal2 s 211064 0 211176 800 0 FreeSans 448 90 0 0 mprj_dat_o_core[22]
port 599 nsew signal input
flabel metal2 s 211624 0 211736 800 0 FreeSans 448 90 0 0 mprj_dat_o_core[23]
port 600 nsew signal input
flabel metal2 s 212296 0 212408 800 0 FreeSans 448 90 0 0 mprj_dat_o_core[24]
port 601 nsew signal input
flabel metal2 s 212856 0 212968 800 0 FreeSans 448 90 0 0 mprj_dat_o_core[25]
port 602 nsew signal input
flabel metal2 s 213528 0 213640 800 0 FreeSans 448 90 0 0 mprj_dat_o_core[26]
port 603 nsew signal input
flabel metal2 s 214088 0 214200 800 0 FreeSans 448 90 0 0 mprj_dat_o_core[27]
port 604 nsew signal input
flabel metal2 s 214760 0 214872 800 0 FreeSans 448 90 0 0 mprj_dat_o_core[28]
port 605 nsew signal input
flabel metal2 s 215320 0 215432 800 0 FreeSans 448 90 0 0 mprj_dat_o_core[29]
port 606 nsew signal input
flabel metal2 s 198856 0 198968 800 0 FreeSans 448 90 0 0 mprj_dat_o_core[2]
port 607 nsew signal input
flabel metal2 s 215880 0 215992 800 0 FreeSans 448 90 0 0 mprj_dat_o_core[30]
port 608 nsew signal input
flabel metal2 s 216552 0 216664 800 0 FreeSans 448 90 0 0 mprj_dat_o_core[31]
port 609 nsew signal input
flabel metal2 s 199416 0 199528 800 0 FreeSans 448 90 0 0 mprj_dat_o_core[3]
port 610 nsew signal input
flabel metal2 s 200088 0 200200 800 0 FreeSans 448 90 0 0 mprj_dat_o_core[4]
port 611 nsew signal input
flabel metal2 s 200648 0 200760 800 0 FreeSans 448 90 0 0 mprj_dat_o_core[5]
port 612 nsew signal input
flabel metal2 s 201320 0 201432 800 0 FreeSans 448 90 0 0 mprj_dat_o_core[6]
port 613 nsew signal input
flabel metal2 s 201880 0 201992 800 0 FreeSans 448 90 0 0 mprj_dat_o_core[7]
port 614 nsew signal input
flabel metal2 s 202552 0 202664 800 0 FreeSans 448 90 0 0 mprj_dat_o_core[8]
port 615 nsew signal input
flabel metal2 s 203112 0 203224 800 0 FreeSans 448 90 0 0 mprj_dat_o_core[9]
port 616 nsew signal input
flabel metal2 s 6104 14200 6216 15000 0 FreeSans 448 90 0 0 mprj_dat_o_user[0]
port 617 nsew signal tristate
flabel metal2 s 30856 14200 30968 15000 0 FreeSans 448 90 0 0 mprj_dat_o_user[10]
port 618 nsew signal tristate
flabel metal2 s 32984 14200 33096 15000 0 FreeSans 448 90 0 0 mprj_dat_o_user[11]
port 619 nsew signal tristate
flabel metal2 s 35224 14200 35336 15000 0 FreeSans 448 90 0 0 mprj_dat_o_user[12]
port 620 nsew signal tristate
flabel metal2 s 37352 14200 37464 15000 0 FreeSans 448 90 0 0 mprj_dat_o_user[13]
port 621 nsew signal tristate
flabel metal2 s 39592 14200 39704 15000 0 FreeSans 448 90 0 0 mprj_dat_o_user[14]
port 622 nsew signal tristate
flabel metal2 s 41720 14200 41832 15000 0 FreeSans 448 90 0 0 mprj_dat_o_user[15]
port 623 nsew signal tristate
flabel metal2 s 43960 14200 44072 15000 0 FreeSans 448 90 0 0 mprj_dat_o_user[16]
port 624 nsew signal tristate
flabel metal2 s 46088 14200 46200 15000 0 FreeSans 448 90 0 0 mprj_dat_o_user[17]
port 625 nsew signal tristate
flabel metal2 s 48328 14200 48440 15000 0 FreeSans 448 90 0 0 mprj_dat_o_user[18]
port 626 nsew signal tristate
flabel metal2 s 50456 14200 50568 15000 0 FreeSans 448 90 0 0 mprj_dat_o_user[19]
port 627 nsew signal tristate
flabel metal2 s 9016 14200 9128 15000 0 FreeSans 448 90 0 0 mprj_dat_o_user[1]
port 628 nsew signal tristate
flabel metal2 s 52696 14200 52808 15000 0 FreeSans 448 90 0 0 mprj_dat_o_user[20]
port 629 nsew signal tristate
flabel metal2 s 54824 14200 54936 15000 0 FreeSans 448 90 0 0 mprj_dat_o_user[21]
port 630 nsew signal tristate
flabel metal2 s 57064 14200 57176 15000 0 FreeSans 448 90 0 0 mprj_dat_o_user[22]
port 631 nsew signal tristate
flabel metal2 s 59304 14200 59416 15000 0 FreeSans 448 90 0 0 mprj_dat_o_user[23]
port 632 nsew signal tristate
flabel metal2 s 61432 14200 61544 15000 0 FreeSans 448 90 0 0 mprj_dat_o_user[24]
port 633 nsew signal tristate
flabel metal2 s 63672 14200 63784 15000 0 FreeSans 448 90 0 0 mprj_dat_o_user[25]
port 634 nsew signal tristate
flabel metal2 s 65800 14200 65912 15000 0 FreeSans 448 90 0 0 mprj_dat_o_user[26]
port 635 nsew signal tristate
flabel metal2 s 68040 14200 68152 15000 0 FreeSans 448 90 0 0 mprj_dat_o_user[27]
port 636 nsew signal tristate
flabel metal2 s 70168 14200 70280 15000 0 FreeSans 448 90 0 0 mprj_dat_o_user[28]
port 637 nsew signal tristate
flabel metal2 s 72408 14200 72520 15000 0 FreeSans 448 90 0 0 mprj_dat_o_user[29]
port 638 nsew signal tristate
flabel metal2 s 11928 14200 12040 15000 0 FreeSans 448 90 0 0 mprj_dat_o_user[2]
port 639 nsew signal tristate
flabel metal2 s 74536 14200 74648 15000 0 FreeSans 448 90 0 0 mprj_dat_o_user[30]
port 640 nsew signal tristate
flabel metal2 s 76776 14200 76888 15000 0 FreeSans 448 90 0 0 mprj_dat_o_user[31]
port 641 nsew signal tristate
flabel metal2 s 14840 14200 14952 15000 0 FreeSans 448 90 0 0 mprj_dat_o_user[3]
port 642 nsew signal tristate
flabel metal2 s 17752 14200 17864 15000 0 FreeSans 448 90 0 0 mprj_dat_o_user[4]
port 643 nsew signal tristate
flabel metal2 s 19880 14200 19992 15000 0 FreeSans 448 90 0 0 mprj_dat_o_user[5]
port 644 nsew signal tristate
flabel metal2 s 22120 14200 22232 15000 0 FreeSans 448 90 0 0 mprj_dat_o_user[6]
port 645 nsew signal tristate
flabel metal2 s 24248 14200 24360 15000 0 FreeSans 448 90 0 0 mprj_dat_o_user[7]
port 646 nsew signal tristate
flabel metal2 s 26488 14200 26600 15000 0 FreeSans 448 90 0 0 mprj_dat_o_user[8]
port 647 nsew signal tristate
flabel metal2 s 28616 14200 28728 15000 0 FreeSans 448 90 0 0 mprj_dat_o_user[9]
port 648 nsew signal tristate
flabel metal2 s 219576 0 219688 800 0 FreeSans 448 90 0 0 mprj_iena_wb
port 649 nsew signal input
flabel metal2 s 175672 0 175784 800 0 FreeSans 448 90 0 0 mprj_sel_o_core[0]
port 650 nsew signal input
flabel metal2 s 176344 0 176456 800 0 FreeSans 448 90 0 0 mprj_sel_o_core[1]
port 651 nsew signal input
flabel metal2 s 176904 0 177016 800 0 FreeSans 448 90 0 0 mprj_sel_o_core[2]
port 652 nsew signal input
flabel metal2 s 177464 0 177576 800 0 FreeSans 448 90 0 0 mprj_sel_o_core[3]
port 653 nsew signal input
flabel metal2 s 6776 14200 6888 15000 0 FreeSans 448 90 0 0 mprj_sel_o_user[0]
port 654 nsew signal tristate
flabel metal2 s 9688 14200 9800 15000 0 FreeSans 448 90 0 0 mprj_sel_o_user[1]
port 655 nsew signal tristate
flabel metal2 s 12600 14200 12712 15000 0 FreeSans 448 90 0 0 mprj_sel_o_user[2]
port 656 nsew signal tristate
flabel metal2 s 15512 14200 15624 15000 0 FreeSans 448 90 0 0 mprj_sel_o_user[3]
port 657 nsew signal tristate
flabel metal2 s 218344 0 218456 800 0 FreeSans 448 90 0 0 mprj_stb_o_core
port 658 nsew signal input
flabel metal2 s 3192 14200 3304 15000 0 FreeSans 448 90 0 0 mprj_stb_o_user
port 659 nsew signal tristate
flabel metal2 s 217112 0 217224 800 0 FreeSans 448 90 0 0 mprj_we_o_core
port 660 nsew signal input
flabel metal2 s 3864 14200 3976 15000 0 FreeSans 448 90 0 0 mprj_we_o_user
port 661 nsew signal tristate
flabel metal2 s 280 14200 392 15000 0 FreeSans 448 90 0 0 user_clock
port 662 nsew signal tristate
flabel metal2 s 217336 14200 217448 15000 0 FreeSans 448 90 0 0 user_clock2
port 663 nsew signal tristate
flabel metal3 s 219200 8680 220000 8792 0 FreeSans 448 0 0 0 user_irq[0]
port 664 nsew signal tristate
flabel metal3 s 219200 11144 220000 11256 0 FreeSans 448 0 0 0 user_irq[1]
port 665 nsew signal tristate
flabel metal3 s 219200 13608 220000 13720 0 FreeSans 448 0 0 0 user_irq[2]
port 666 nsew signal tristate
flabel metal2 s 218120 14200 218232 15000 0 FreeSans 448 90 0 0 user_irq_core[0]
port 667 nsew signal input
flabel metal2 s 218792 14200 218904 15000 0 FreeSans 448 90 0 0 user_irq_core[1]
port 668 nsew signal input
flabel metal2 s 219576 14200 219688 15000 0 FreeSans 448 90 0 0 user_irq_core[2]
port 669 nsew signal input
flabel metal3 s 219200 1288 220000 1400 0 FreeSans 448 0 0 0 user_irq_ena[0]
port 670 nsew signal input
flabel metal3 s 219200 3752 220000 3864 0 FreeSans 448 0 0 0 user_irq_ena[1]
port 671 nsew signal input
flabel metal3 s 219200 6216 220000 6328 0 FreeSans 448 0 0 0 user_irq_ena[2]
port 672 nsew signal input
flabel metal2 s 952 14200 1064 15000 0 FreeSans 448 90 0 0 user_reset
port 673 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 220000 15000
<< end >>
