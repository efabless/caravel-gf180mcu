VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO copyright_block
  CLASS BLOCK ;
  FOREIGN copyright_block ;
  ORIGIN 0.000 0.000 ;
  SIZE 93.495 BY 44.990 ;
  OBS
      LAYER Metal5 ;
        RECT 2.635 42.780 5.155 43.140 ;
        RECT 2.275 42.420 5.155 42.780 ;
        RECT 1.915 41.700 5.155 42.420 ;
        RECT 1.915 37.020 2.995 41.700 ;
        RECT 6.175 40.575 9.055 40.935 ;
        RECT 10.480 40.575 13.000 40.935 ;
        RECT 14.830 40.575 17.710 40.935 ;
        RECT 6.175 39.855 9.415 40.575 ;
        RECT 8.335 38.775 9.415 39.855 ;
        RECT 6.535 38.415 9.415 38.775 ;
        RECT 6.175 37.695 9.415 38.415 ;
        RECT 1.915 36.300 5.155 37.020 ;
        RECT 2.275 35.940 5.155 36.300 ;
        RECT 2.635 35.580 5.155 35.940 ;
        RECT 6.175 36.615 7.255 37.695 ;
        RECT 8.335 36.615 9.415 37.695 ;
        RECT 6.175 35.895 9.415 36.615 ;
        RECT 6.535 35.535 9.415 35.895 ;
        RECT 10.480 40.215 13.360 40.575 ;
        RECT 10.480 39.495 13.720 40.215 ;
        RECT 14.830 39.855 18.070 40.575 ;
        RECT 10.480 35.535 11.560 39.495 ;
        RECT 12.640 38.775 13.720 39.495 ;
        RECT 16.990 38.775 18.070 39.855 ;
        RECT 15.190 38.415 18.070 38.775 ;
        RECT 14.830 37.695 18.070 38.415 ;
        RECT 14.830 36.615 15.910 37.695 ;
        RECT 16.990 36.615 18.070 37.695 ;
        RECT 19.370 37.695 20.450 40.935 ;
        RECT 21.530 37.695 22.610 40.935 ;
        RECT 23.890 40.665 26.410 41.025 ;
        RECT 19.370 36.615 22.610 37.695 ;
        RECT 23.530 39.945 26.770 40.665 ;
        RECT 23.530 38.865 24.610 39.945 ;
        RECT 25.690 38.865 26.770 39.945 ;
        RECT 23.530 38.145 26.770 38.865 ;
        RECT 23.530 37.785 26.410 38.145 ;
        RECT 23.530 36.705 24.610 37.785 ;
        RECT 14.830 35.895 18.070 36.615 ;
        RECT 19.730 36.255 22.250 36.615 ;
        RECT 15.190 35.535 18.070 35.895 ;
        RECT 20.450 35.535 21.530 36.255 ;
        RECT 23.530 35.985 26.770 36.705 ;
        RECT 23.890 35.625 26.770 35.985 ;
        RECT 27.835 35.535 28.915 43.095 ;
        RECT 33.000 42.825 34.800 43.185 ;
        RECT 32.640 42.465 35.160 42.825 ;
        RECT 32.280 41.745 35.520 42.465 ;
        RECT 32.280 37.065 33.360 41.745 ;
        RECT 34.440 41.025 35.520 41.745 ;
        RECT 36.680 42.105 39.920 43.185 ;
        RECT 43.565 42.855 45.005 43.215 ;
        RECT 43.205 42.495 45.005 42.855 ;
        RECT 36.680 39.945 37.760 42.105 ;
        RECT 42.845 41.775 45.005 42.495 ;
        RECT 50.345 42.765 51.785 43.125 ;
        RECT 50.345 42.405 52.145 42.765 ;
        RECT 34.440 37.065 35.520 39.945 ;
        RECT 32.280 36.345 35.520 37.065 ;
        RECT 32.640 35.985 35.520 36.345 ;
        RECT 33.000 35.625 35.520 35.985 ;
        RECT 36.680 38.865 38.840 39.945 ;
        RECT 36.680 35.625 37.760 38.865 ;
        RECT 42.845 37.095 43.925 41.775 ;
        RECT 46.765 41.545 48.565 41.905 ;
        RECT 50.345 41.685 52.505 42.405 ;
        RECT 46.405 41.185 48.925 41.545 ;
        RECT 46.045 40.465 49.285 41.185 ;
        RECT 46.045 37.945 47.125 40.465 ;
        RECT 48.205 39.745 49.285 40.465 ;
        RECT 48.205 37.945 49.285 38.305 ;
        RECT 46.045 37.225 49.285 37.945 ;
        RECT 42.845 36.375 45.005 37.095 ;
        RECT 46.405 36.865 48.925 37.225 ;
        RECT 51.425 37.005 52.505 41.685 ;
        RECT 46.765 36.505 48.565 36.865 ;
        RECT 43.205 36.015 45.005 36.375 ;
        RECT 43.565 35.655 45.005 36.015 ;
        RECT 50.345 36.285 52.505 37.005 ;
        RECT 57.295 42.045 60.535 43.125 ;
        RECT 63.035 42.765 64.835 43.125 ;
        RECT 62.675 42.045 64.835 42.765 ;
        RECT 57.295 39.885 58.375 42.045 ;
        RECT 62.675 40.965 63.755 42.045 ;
        RECT 70.295 40.965 71.375 43.125 ;
        RECT 61.595 39.885 64.835 40.965 ;
        RECT 65.945 40.555 68.825 40.915 ;
        RECT 70.295 40.605 72.815 40.965 ;
        RECT 57.295 38.805 59.455 39.885 ;
        RECT 57.295 36.645 58.375 38.805 ;
        RECT 50.345 35.925 52.145 36.285 ;
        RECT 50.345 35.565 51.785 35.925 ;
        RECT 57.295 35.565 60.535 36.645 ;
        RECT 62.675 35.565 63.755 39.885 ;
        RECT 65.945 39.835 69.185 40.555 ;
        RECT 68.105 38.755 69.185 39.835 ;
        RECT 66.305 38.395 69.185 38.755 ;
        RECT 65.945 37.675 69.185 38.395 ;
        RECT 65.945 36.595 67.025 37.675 ;
        RECT 68.105 36.595 69.185 37.675 ;
        RECT 65.945 35.875 69.185 36.595 ;
        RECT 66.305 35.515 69.185 35.875 ;
        RECT 70.295 40.245 73.175 40.605 ;
        RECT 70.295 39.525 73.535 40.245 ;
        RECT 70.295 37.005 71.375 39.525 ;
        RECT 72.455 37.005 73.535 39.525 ;
        RECT 70.295 36.285 73.535 37.005 ;
        RECT 70.295 35.925 73.175 36.285 ;
        RECT 70.295 35.565 72.815 35.925 ;
        RECT 74.645 35.565 75.725 43.125 ;
        RECT 77.155 40.605 79.675 40.965 ;
        RECT 81.865 40.645 84.385 41.005 ;
        RECT 86.165 40.645 88.685 41.005 ;
        RECT 76.795 39.885 80.035 40.605 ;
        RECT 81.505 40.285 84.385 40.645 ;
        RECT 85.805 40.285 88.685 40.645 ;
        RECT 76.795 38.805 77.875 39.885 ;
        RECT 78.955 38.805 80.035 39.885 ;
        RECT 76.795 38.085 80.035 38.805 ;
        RECT 81.145 39.925 84.385 40.285 ;
        RECT 85.445 39.925 88.685 40.285 ;
        RECT 81.145 38.845 82.585 39.925 ;
        RECT 85.445 38.845 86.885 39.925 ;
        RECT 81.145 38.485 83.665 38.845 ;
        RECT 85.445 38.485 87.965 38.845 ;
        RECT 81.505 38.125 84.025 38.485 ;
        RECT 85.805 38.125 88.325 38.485 ;
        RECT 76.795 37.725 79.675 38.085 ;
        RECT 81.865 37.765 84.385 38.125 ;
        RECT 86.165 37.765 88.685 38.125 ;
        RECT 76.795 36.645 77.875 37.725 ;
        RECT 82.945 36.685 84.385 37.765 ;
        RECT 87.245 36.685 88.685 37.765 ;
        RECT 76.795 35.925 80.035 36.645 ;
        RECT 77.155 35.565 80.035 35.925 ;
        RECT 81.145 36.325 84.385 36.685 ;
        RECT 85.445 36.325 88.685 36.685 ;
        RECT 81.145 35.965 84.025 36.325 ;
        RECT 85.445 35.965 88.325 36.325 ;
        RECT 81.145 35.605 83.665 35.965 ;
        RECT 85.445 35.605 87.965 35.965 ;
        RECT 3.060 32.205 4.860 32.565 ;
        RECT 2.700 31.845 5.220 32.205 ;
        RECT 2.340 31.125 5.580 31.845 ;
        RECT 2.340 26.445 3.420 31.125 ;
        RECT 4.500 30.405 5.580 31.125 ;
        RECT 7.260 30.130 9.060 30.490 ;
        RECT 6.900 29.770 9.420 30.130 ;
        RECT 11.515 30.080 13.315 30.440 ;
        RECT 4.500 26.445 5.580 29.325 ;
        RECT 2.340 25.725 5.580 26.445 ;
        RECT 6.540 29.050 9.780 29.770 ;
        RECT 11.155 29.720 13.675 30.080 ;
        RECT 15.910 30.035 17.710 30.395 ;
        RECT 6.540 26.530 7.620 29.050 ;
        RECT 8.700 26.530 9.780 29.050 ;
        RECT 6.540 25.810 9.780 26.530 ;
        RECT 10.795 29.000 14.035 29.720 ;
        RECT 15.550 29.675 18.070 30.035 ;
        RECT 10.795 26.480 11.875 29.000 ;
        RECT 12.955 26.480 14.035 29.000 ;
        RECT 2.700 25.365 5.580 25.725 ;
        RECT 6.900 25.450 9.420 25.810 ;
        RECT 10.795 25.760 14.035 26.480 ;
        RECT 15.190 28.955 18.430 29.675 ;
        RECT 15.190 26.435 16.270 28.955 ;
        RECT 17.350 26.435 18.430 28.955 ;
        RECT 3.060 25.005 5.580 25.365 ;
        RECT 7.260 25.090 9.060 25.450 ;
        RECT 11.155 25.400 13.675 25.760 ;
        RECT 15.190 25.715 18.430 26.435 ;
        RECT 11.515 25.040 13.315 25.400 ;
        RECT 15.550 25.355 18.430 25.715 ;
        RECT 15.910 24.995 18.430 25.355 ;
        RECT 16.990 23.915 18.430 24.995 ;
        RECT 19.535 24.950 20.615 32.510 ;
        RECT 32.020 32.205 33.820 32.565 ;
        RECT 31.660 31.845 34.180 32.205 ;
        RECT 31.300 31.125 34.540 31.845 ;
        RECT 22.095 29.990 24.615 30.350 ;
        RECT 21.735 29.270 24.975 29.990 ;
        RECT 21.735 28.190 22.815 29.270 ;
        RECT 23.895 28.190 24.975 29.270 ;
        RECT 21.735 27.470 24.975 28.190 ;
        RECT 25.985 28.140 30.305 29.220 ;
        RECT 21.735 27.110 24.615 27.470 ;
        RECT 21.735 26.030 22.815 27.110 ;
        RECT 31.300 26.445 32.380 31.125 ;
        RECT 33.460 30.405 34.540 31.125 ;
        RECT 33.460 26.445 34.540 29.325 ;
        RECT 21.735 25.310 24.975 26.030 ;
        RECT 31.300 25.725 34.540 26.445 ;
        RECT 31.660 25.365 34.540 25.725 ;
        RECT 22.095 24.950 24.975 25.310 ;
        RECT 32.020 25.005 34.540 25.365 ;
        RECT 35.600 24.875 36.680 32.435 ;
        RECT 42.105 30.320 43.185 32.480 ;
        RECT 38.520 29.865 40.320 30.225 ;
        RECT 42.105 29.960 44.625 30.320 ;
        RECT 46.410 29.960 49.290 30.320 ;
        RECT 38.160 29.505 40.680 29.865 ;
        RECT 42.105 29.600 44.985 29.960 ;
        RECT 37.800 28.785 41.040 29.505 ;
        RECT 37.800 26.265 38.880 28.785 ;
        RECT 39.960 26.265 41.040 28.785 ;
        RECT 37.800 25.545 41.040 26.265 ;
        RECT 42.105 28.880 45.345 29.600 ;
        RECT 46.410 29.240 49.650 29.960 ;
        RECT 42.105 26.360 43.185 28.880 ;
        RECT 44.265 26.360 45.345 28.880 ;
        RECT 48.570 28.160 49.650 29.240 ;
        RECT 46.770 27.800 49.650 28.160 ;
        RECT 42.105 25.640 45.345 26.360 ;
        RECT 46.410 27.080 49.650 27.800 ;
        RECT 46.410 26.000 47.490 27.080 ;
        RECT 48.570 26.000 49.650 27.080 ;
        RECT 38.160 25.185 40.680 25.545 ;
        RECT 42.105 25.280 44.985 25.640 ;
        RECT 46.410 25.280 49.650 26.000 ;
        RECT 38.520 24.825 40.320 25.185 ;
        RECT 42.105 24.920 44.625 25.280 ;
        RECT 46.770 24.920 49.650 25.280 ;
        RECT 50.760 24.825 51.840 32.385 ;
        RECT 55.250 31.260 58.490 32.340 ;
        RECT 55.250 29.100 56.330 31.260 ;
        RECT 74.580 30.405 75.660 32.565 ;
        RECT 81.030 30.405 83.190 32.565 ;
        RECT 60.230 30.000 62.030 30.360 ;
        RECT 59.870 29.640 62.390 30.000 ;
        RECT 55.250 28.020 57.410 29.100 ;
        RECT 59.510 28.920 62.750 29.640 ;
        RECT 55.250 24.780 56.330 28.020 ;
        RECT 59.510 26.400 60.590 28.920 ;
        RECT 61.670 26.400 62.750 28.920 ;
        RECT 59.510 25.680 62.750 26.400 ;
        RECT 63.815 26.445 64.895 30.405 ;
        RECT 65.975 26.445 67.055 30.405 ;
        RECT 63.815 25.725 67.055 26.445 ;
        RECT 59.870 25.320 62.390 25.680 ;
        RECT 64.175 25.365 67.055 25.725 ;
        RECT 60.230 24.960 62.030 25.320 ;
        RECT 64.535 25.005 67.055 25.365 ;
        RECT 68.025 29.955 70.545 30.315 ;
        RECT 73.140 30.045 75.660 30.405 ;
        RECT 68.025 29.595 70.905 29.955 ;
        RECT 72.780 29.685 75.660 30.045 ;
        RECT 68.025 28.875 71.265 29.595 ;
        RECT 68.025 24.915 69.105 28.875 ;
        RECT 70.185 24.915 71.265 28.875 ;
        RECT 72.420 28.965 75.660 29.685 ;
        RECT 72.420 26.445 73.500 28.965 ;
        RECT 74.580 26.445 75.660 28.965 ;
        RECT 72.420 25.725 75.660 26.445 ;
        RECT 72.780 25.365 75.660 25.725 ;
        RECT 73.140 25.005 75.660 25.365 ;
        RECT 76.725 30.000 79.245 30.360 ;
        RECT 84.665 30.000 87.185 30.360 ;
        RECT 89.375 30.045 91.895 30.405 ;
        RECT 76.725 29.640 79.605 30.000 ;
        RECT 76.725 28.920 79.965 29.640 ;
        RECT 76.725 24.960 77.805 28.920 ;
        RECT 78.885 28.200 79.965 28.920 ;
        RECT 81.030 28.245 83.190 29.325 ;
        RECT 82.110 26.085 83.190 28.245 ;
        RECT 81.030 25.005 83.190 26.085 ;
        RECT 84.305 29.280 87.545 30.000 ;
        RECT 89.015 29.685 91.895 30.045 ;
        RECT 84.305 28.200 85.385 29.280 ;
        RECT 86.465 28.200 87.545 29.280 ;
        RECT 84.305 27.480 87.545 28.200 ;
        RECT 88.655 29.325 91.895 29.685 ;
        RECT 88.655 28.245 90.095 29.325 ;
        RECT 88.655 27.885 91.175 28.245 ;
        RECT 89.015 27.525 91.535 27.885 ;
        RECT 84.305 27.120 87.185 27.480 ;
        RECT 89.375 27.165 91.895 27.525 ;
        RECT 84.305 26.040 85.385 27.120 ;
        RECT 90.455 26.085 91.895 27.165 ;
        RECT 84.305 25.320 87.545 26.040 ;
        RECT 84.665 24.960 87.545 25.320 ;
        RECT 88.655 25.725 91.895 26.085 ;
        RECT 88.655 25.365 91.535 25.725 ;
        RECT 88.655 25.005 91.175 25.365 ;
        RECT 15.190 23.555 18.430 23.915 ;
        RECT 15.190 23.195 18.070 23.555 ;
        RECT 15.190 22.835 17.710 23.195 ;
        RECT 23.065 20.985 25.585 21.345 ;
        RECT 23.065 20.625 25.945 20.985 ;
        RECT 27.370 20.895 29.890 21.255 ;
        RECT 23.065 19.905 26.305 20.625 ;
        RECT 2.590 18.920 4.390 19.280 ;
        RECT 6.895 18.965 8.695 19.325 ;
        RECT 2.230 18.560 4.750 18.920 ;
        RECT 6.535 18.605 9.055 18.965 ;
        RECT 10.885 18.875 13.405 19.235 ;
        RECT 1.870 17.840 5.110 18.560 ;
        RECT 1.870 15.320 2.950 17.840 ;
        RECT 4.030 15.320 5.110 17.840 ;
        RECT 1.870 14.600 5.110 15.320 ;
        RECT 6.175 17.885 9.415 18.605 ;
        RECT 6.175 15.365 7.255 17.885 ;
        RECT 8.335 15.365 9.415 17.885 ;
        RECT 6.175 14.645 9.415 15.365 ;
        RECT 10.525 18.155 13.765 18.875 ;
        RECT 10.525 17.075 11.605 18.155 ;
        RECT 12.685 17.075 13.765 18.155 ;
        RECT 10.525 16.355 13.765 17.075 ;
        RECT 14.785 18.780 17.305 19.140 ;
        RECT 14.785 18.420 17.665 18.780 ;
        RECT 14.785 17.700 18.025 18.420 ;
        RECT 10.525 15.995 13.405 16.355 ;
        RECT 10.525 14.915 11.605 15.995 ;
        RECT 2.230 14.240 4.750 14.600 ;
        RECT 6.175 14.285 9.055 14.645 ;
        RECT 2.590 13.880 4.390 14.240 ;
        RECT 6.175 13.925 8.695 14.285 ;
        RECT 10.525 14.195 13.765 14.915 ;
        RECT 6.175 11.765 7.255 13.925 ;
        RECT 10.885 13.835 13.765 14.195 ;
        RECT 14.785 13.740 15.865 17.700 ;
        RECT 16.945 13.740 18.025 17.700 ;
        RECT 23.065 17.385 24.145 19.905 ;
        RECT 25.225 17.385 26.305 19.905 ;
        RECT 23.065 16.665 26.305 17.385 ;
        RECT 27.370 20.535 30.250 20.895 ;
        RECT 27.370 19.815 30.610 20.535 ;
        RECT 23.065 16.305 25.945 16.665 ;
        RECT 23.065 15.945 25.585 16.305 ;
        RECT 23.065 13.785 24.145 15.945 ;
        RECT 27.370 15.135 28.450 19.815 ;
        RECT 29.530 15.135 30.610 19.815 ;
        RECT 27.370 14.415 30.610 15.135 ;
        RECT 31.670 19.455 32.750 21.255 ;
        RECT 33.830 19.455 34.910 21.255 ;
        RECT 31.670 18.735 34.910 19.455 ;
        RECT 31.670 18.015 34.550 18.735 ;
        RECT 31.670 16.935 34.190 18.015 ;
        RECT 31.670 16.215 34.550 16.935 ;
        RECT 31.670 15.495 34.910 16.215 ;
        RECT 27.370 14.055 30.250 14.415 ;
        RECT 27.370 13.695 29.890 14.055 ;
        RECT 31.670 13.695 32.750 15.495 ;
        RECT 33.830 13.695 34.910 15.495 ;
        RECT 1.355 8.820 3.875 9.180 ;
        RECT 1.355 8.460 4.235 8.820 ;
        RECT 1.355 7.740 4.595 8.460 ;
        RECT 22.410 8.095 25.650 9.175 ;
        RECT 1.355 3.060 2.435 7.740 ;
        RECT 3.515 3.060 4.595 7.740 ;
        RECT 24.570 7.015 25.650 8.095 ;
        RECT 6.020 6.615 8.540 6.975 ;
        RECT 10.685 6.615 12.485 6.975 ;
        RECT 1.355 2.340 4.595 3.060 ;
        RECT 5.660 5.895 8.900 6.615 ;
        RECT 10.325 6.255 12.845 6.615 ;
        RECT 5.660 4.815 6.740 5.895 ;
        RECT 7.820 4.815 8.900 5.895 ;
        RECT 5.660 4.095 8.900 4.815 ;
        RECT 9.965 5.535 13.205 6.255 ;
        RECT 5.660 3.735 8.540 4.095 ;
        RECT 5.660 2.655 6.740 3.735 ;
        RECT 9.965 3.015 11.045 5.535 ;
        RECT 12.125 4.815 13.205 5.535 ;
        RECT 22.410 5.935 25.650 7.015 ;
        RECT 26.760 8.140 30.000 9.220 ;
        RECT 12.125 3.015 13.205 3.375 ;
        RECT 1.355 1.980 4.235 2.340 ;
        RECT 1.355 1.620 3.875 1.980 ;
        RECT 5.660 1.935 8.900 2.655 ;
        RECT 9.965 2.295 13.205 3.015 ;
        RECT 22.410 2.695 23.490 5.935 ;
        RECT 26.760 2.740 27.840 8.140 ;
        RECT 28.920 2.740 30.000 8.140 ;
        RECT 31.160 8.100 34.400 9.180 ;
        RECT 35.600 8.140 38.840 9.220 ;
        RECT 33.320 7.020 34.400 8.100 ;
        RECT 37.760 7.060 38.840 8.140 ;
        RECT 10.325 1.935 12.845 2.295 ;
        RECT 6.020 1.575 8.900 1.935 ;
        RECT 10.685 1.575 12.485 1.935 ;
        RECT 22.410 1.615 25.650 2.695 ;
        RECT 26.760 1.660 30.000 2.740 ;
        RECT 31.160 5.940 34.400 7.020 ;
        RECT 35.600 5.980 38.840 7.060 ;
        RECT 31.160 2.700 32.240 5.940 ;
        RECT 35.600 2.740 36.680 5.980 ;
        RECT 31.160 1.620 34.400 2.700 ;
        RECT 35.600 1.660 38.840 2.740 ;
  END
END copyright_block
END LIBRARY

