magic
tech gf180mcuC
magscale 1 5
timestamp 1668623937
<< checkpaint >>
rect 931130 41485 991195 50375
rect 928530 38430 991195 41485
rect 928530 36340 990930 38430
rect 931330 35955 990930 36340
rect 931340 35880 990930 35955
rect 942275 35785 990930 35880
<< fillblock >>
rect 933525 37510 943030 39210
use font_6C  font_6C_0 alpha
timestamp 1654634570
transform 1 0 935855 0 1 37855
box 0 0 108 756
use font_6E  font_6E_0 alpha
timestamp 1654634570
transform 1 0 936585 0 1 37855
box 0 0 324 540
use font_22  font_22_0 alpha
timestamp 1654634570
transform 1 0 933765 0 1 38225
box 0 324 324 756
use font_22  font_22_1
timestamp 1654634570
transform 1 0 942425 0 1 38225
box 0 324 324 756
use font_43  font_43_0 alpha
timestamp 1654634570
transform 1 0 941275 0 1 37850
box 0 0 324 756
use font_49  font_49_0 alpha
timestamp 1654634570
transform 1 0 940680 0 1 37860
box 0 0 324 756
use font_53  font_53_0 alpha
timestamp 1654634570
transform 1 0 934370 0 1 37865
box 0 0 324 756
use font_54  font_54_0 alpha
timestamp 1654634570
transform 1 0 938340 0 1 37855
box 0 0 324 756
use font_61  font_61_0 alpha
timestamp 1654634570
transform 1 0 934910 0 1 37860
box 0 0 324 540
use font_65  font_65_0 alpha
timestamp 1654634570
transform 1 0 939395 0 1 37855
box 0 0 324 540
use font_67  font_67_0 alpha
timestamp 1654634570
transform 1 0 937085 0 1 37855
box 0 -216 324 540
use font_68  font_68_0 alpha
timestamp 1654634570
transform 1 0 938865 0 1 37855
box 0 0 324 756
use font_69  font_69_0 alpha
timestamp 1654634570
transform 1 0 935440 0 1 37860
box 0 0 216 756
use font_69  font_69_1
timestamp 1654634570
transform 1 0 936190 0 1 37855
box 0 0 216 756
use font_73  font_73_0 alpha
timestamp 1654634570
transform 1 0 941865 0 1 37855
box 0 0 324 540
<< end >>
