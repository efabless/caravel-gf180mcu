magic
tech gf180mcuC
magscale 1 10
timestamp 1655304105
<< error_p >>
rect -730 -255 -719 -209
rect -516 -255 -505 -209
rect -302 -255 -291 -209
rect -88 -255 -77 -209
rect 126 -255 137 -209
rect 340 -255 351 -209
rect 554 -255 565 -209
<< nwell >>
rect -1050 -486 980 486
<< mvpmos >>
rect -732 -176 -622 224
rect -518 -176 -408 224
rect -304 -176 -194 224
rect -90 -176 20 224
rect 124 -176 234 224
rect 338 -176 448 224
rect 552 -176 662 224
<< mvpdiff >>
rect -820 211 -732 224
rect -820 -163 -807 211
rect -761 -163 -732 211
rect -820 -176 -732 -163
rect -622 211 -518 224
rect -622 -163 -593 211
rect -547 -163 -518 211
rect -622 -176 -518 -163
rect -408 211 -304 224
rect -408 -163 -379 211
rect -333 -163 -304 211
rect -408 -176 -304 -163
rect -194 211 -90 224
rect -194 -163 -165 211
rect -119 -163 -90 211
rect -194 -176 -90 -163
rect 20 211 124 224
rect 20 -163 49 211
rect 95 -163 124 211
rect 20 -176 124 -163
rect 234 211 338 224
rect 234 -163 263 211
rect 309 -163 338 211
rect 234 -176 338 -163
rect 448 211 552 224
rect 448 -163 477 211
rect 523 -163 552 211
rect 448 -176 552 -163
rect 662 211 750 224
rect 662 -163 691 211
rect 737 -163 750 211
rect 662 -176 750 -163
<< mvpdiffc >>
rect -807 -163 -761 211
rect -593 -163 -547 211
rect -379 -163 -333 211
rect -165 -163 -119 211
rect 49 -163 95 211
rect 263 -163 309 211
rect 477 -163 523 211
rect 691 -163 737 211
<< mvnsubdiff >>
rect -964 387 894 400
rect -964 341 -848 387
rect 778 341 894 387
rect -964 328 894 341
rect -964 284 -892 328
rect -964 -284 -951 284
rect -905 -284 -892 284
rect 822 284 894 328
rect -964 -328 -892 -284
rect 822 -284 835 284
rect 881 -284 894 284
rect 822 -328 894 -284
rect -964 -400 894 -328
<< mvnsubdiffcont >>
rect -848 341 778 387
rect -951 -284 -905 284
rect 835 -284 881 284
<< polysilicon >>
rect -732 224 -622 268
rect -518 224 -408 268
rect -304 224 -194 268
rect -90 224 20 268
rect 124 224 234 268
rect 338 224 448 268
rect 552 224 662 268
rect -732 -209 -622 -176
rect -732 -255 -719 -209
rect -635 -255 -622 -209
rect -732 -268 -622 -255
rect -518 -209 -408 -176
rect -518 -255 -505 -209
rect -421 -255 -408 -209
rect -518 -268 -408 -255
rect -304 -209 -194 -176
rect -304 -255 -291 -209
rect -207 -255 -194 -209
rect -304 -268 -194 -255
rect -90 -209 20 -176
rect -90 -255 -77 -209
rect 7 -255 20 -209
rect -90 -268 20 -255
rect 124 -209 234 -176
rect 124 -255 137 -209
rect 221 -255 234 -209
rect 124 -268 234 -255
rect 338 -209 448 -176
rect 338 -255 351 -209
rect 435 -255 448 -209
rect 338 -268 448 -255
rect 552 -209 662 -176
rect 552 -255 565 -209
rect 649 -255 662 -209
rect 552 -268 662 -255
<< polycontact >>
rect -719 -255 -635 -209
rect -505 -255 -421 -209
rect -291 -255 -207 -209
rect -77 -255 7 -209
rect 137 -255 221 -209
rect 351 -255 435 -209
rect 565 -255 649 -209
<< metal1 >>
rect -951 341 -848 387
rect 778 341 881 387
rect -951 284 -905 341
rect 835 284 881 341
rect -807 211 -761 222
rect -807 -174 -761 -163
rect -593 211 -547 222
rect -593 -174 -547 -163
rect -379 211 -333 222
rect -379 -174 -333 -163
rect -165 211 -119 222
rect -165 -174 -119 -163
rect 49 211 95 222
rect 49 -174 95 -163
rect 263 211 309 222
rect 263 -174 309 -163
rect 477 211 523 222
rect 477 -174 523 -163
rect 691 211 737 222
rect 691 -174 737 -163
rect -730 -255 -719 -209
rect -635 -255 -624 -209
rect -516 -255 -505 -209
rect -421 -255 -410 -209
rect -302 -255 -291 -209
rect -207 -255 -196 -209
rect -88 -255 -77 -209
rect 7 -255 18 -209
rect 126 -255 137 -209
rect 221 -255 232 -209
rect 340 -255 351 -209
rect 435 -255 446 -209
rect 554 -255 565 -209
rect 649 -255 660 -209
rect -951 -341 -905 -284
rect 835 -341 881 -284
rect -951 -387 881 -341
<< properties >>
string FIXED_BBOX -858 -364 858 364
string gencell pmos_6p0
string library gf180mcu
string parameters w 2 l 0.5 m 1 nf 7 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 0 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.5 wmin 0.3 full_metal 1 compatible {pmos_3p3 pmos_6p0}
<< end >>
