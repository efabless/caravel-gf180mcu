VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_id_programming
  CLASS BLOCK ;
  FOREIGN user_id_programming ;
  ORIGIN 0.000 0.000 ;
  SIZE 108.360 BY 11.565 ;
  PIN mask_rev[0]
    PORT
      LAYER Metal2 ;
        RECT 0.000 0.000 0.280 5.380 ;
    END
  END mask_rev[0]
  PIN mask_rev[10]
    PORT
      LAYER Metal2 ;
        RECT 34.720 0.000 35.000 9.545 ;
    END
  END mask_rev[10]
  PIN mask_rev[11]
    PORT
      LAYER Metal2 ;
        RECT 38.640 0.000 38.920 4.500 ;
    END
  END mask_rev[11]
  PIN mask_rev[12]
    PORT
      LAYER Metal2 ;
        RECT 42.000 0.000 42.280 9.545 ;
    END
  END mask_rev[12]
  PIN mask_rev[13]
    PORT
      LAYER Metal2 ;
        RECT 45.360 0.000 45.640 4.495 ;
    END
  END mask_rev[13]
  PIN mask_rev[14]
    PORT
      LAYER Metal2 ;
        RECT 48.720 0.000 49.000 9.545 ;
    END
  END mask_rev[14]
  PIN mask_rev[15]
    PORT
      LAYER Metal2 ;
        RECT 52.080 0.000 52.360 4.495 ;
    END
  END mask_rev[15]
  PIN mask_rev[16]
    PORT
      LAYER Metal2 ;
        RECT 56.000 0.000 56.280 9.545 ;
    END
  END mask_rev[16]
  PIN mask_rev[17]
    PORT
      LAYER Metal2 ;
        RECT 59.360 0.000 59.640 4.495 ;
    END
  END mask_rev[17]
  PIN mask_rev[18]
    PORT
      LAYER Metal2 ;
        RECT 62.720 0.000 63.000 9.545 ;
    END
  END mask_rev[18]
  PIN mask_rev[19]
    PORT
      LAYER Metal2 ;
        RECT 66.080 0.000 66.360 4.390 ;
    END
  END mask_rev[19]
  PIN mask_rev[1]
    PORT
      LAYER Metal2 ;
        RECT 3.360 0.000 3.640 4.495 ;
    END
  END mask_rev[1]
  PIN mask_rev[20]
    PORT
      LAYER Metal2 ;
        RECT 70.000 0.000 70.280 3.045 ;
    END
  END mask_rev[20]
  PIN mask_rev[21]
    PORT
      LAYER Metal2 ;
        RECT 73.360 0.000 73.640 4.495 ;
    END
  END mask_rev[21]
  PIN mask_rev[22]
    PORT
      LAYER Metal2 ;
        RECT 76.720 0.000 77.000 3.545 ;
    END
  END mask_rev[22]
  PIN mask_rev[23]
    PORT
      LAYER Metal2 ;
        RECT 80.080 0.000 80.360 4.495 ;
    END
  END mask_rev[23]
  PIN mask_rev[24]
    PORT
      LAYER Metal2 ;
        RECT 83.440 0.000 83.720 3.585 ;
    END
  END mask_rev[24]
  PIN mask_rev[25]
    PORT
      LAYER Metal2 ;
        RECT 87.360 0.000 87.640 4.495 ;
    END
  END mask_rev[25]
  PIN mask_rev[26]
    PORT
      LAYER Metal2 ;
        RECT 90.720 0.000 91.000 3.870 ;
    END
  END mask_rev[26]
  PIN mask_rev[27]
    PORT
      LAYER Metal2 ;
        RECT 94.080 0.000 94.360 3.655 ;
    END
  END mask_rev[27]
  PIN mask_rev[28]
    PORT
      LAYER Metal2 ;
        RECT 97.440 0.000 97.720 3.895 ;
    END
  END mask_rev[28]
  PIN mask_rev[29]
    PORT
      LAYER Metal2 ;
        RECT 101.360 0.000 101.640 3.835 ;
    END
  END mask_rev[29]
  PIN mask_rev[2]
    PORT
      LAYER Metal2 ;
        RECT 7.280 0.000 7.560 3.830 ;
    END
  END mask_rev[2]
  PIN mask_rev[30]
    PORT
      LAYER Metal2 ;
        RECT 104.720 0.000 105.000 3.845 ;
    END
  END mask_rev[30]
  PIN mask_rev[31]
    PORT
      LAYER Metal2 ;
        RECT 108.080 0.000 108.360 4.495 ;
    END
  END mask_rev[31]
  PIN mask_rev[3]
    PORT
      LAYER Metal2 ;
        RECT 10.640 0.000 10.920 3.040 ;
    END
  END mask_rev[3]
  PIN mask_rev[4]
    PORT
      LAYER Metal2 ;
        RECT 14.000 0.000 14.280 3.090 ;
    END
  END mask_rev[4]
  PIN mask_rev[5]
    PORT
      LAYER Metal2 ;
        RECT 17.360 0.000 17.640 4.495 ;
    END
  END mask_rev[5]
  PIN mask_rev[6]
    PORT
      LAYER Metal2 ;
        RECT 20.720 0.000 21.000 3.610 ;
    END
  END mask_rev[6]
  PIN mask_rev[7]
    PORT
      LAYER Metal2 ;
        RECT 24.640 0.000 24.920 4.495 ;
    END
  END mask_rev[7]
  PIN mask_rev[8]
    PORT
      LAYER Metal2 ;
        RECT 28.000 0.000 28.280 3.295 ;
    END
  END mask_rev[8]
  PIN mask_rev[9]
    PORT
      LAYER Metal2 ;
        RECT 31.360 0.000 31.640 4.495 ;
    END
  END mask_rev[9]
  PIN VDD
    USE POWER ;
    PORT
      LAYER Metal5 ;
        RECT 3.705 6.125 31.045 7.725 ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    PORT
      LAYER Metal5 ;
        RECT 3.705 2.125 8.545 3.725 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 4.445 2.640 104.125 11.080 ;
      LAYER Metal2 ;
        RECT 0.280 9.845 108.080 11.565 ;
        RECT 0.280 5.680 34.420 9.845 ;
        RECT 0.580 4.795 34.420 5.680 ;
        RECT 0.580 2.125 3.060 4.795 ;
        RECT 3.940 4.130 17.060 4.795 ;
        RECT 3.940 2.125 6.980 4.130 ;
        RECT 7.860 3.390 17.060 4.130 ;
        RECT 7.860 3.340 13.700 3.390 ;
        RECT 7.860 2.125 10.340 3.340 ;
        RECT 11.220 2.125 13.700 3.340 ;
        RECT 14.580 2.125 17.060 3.390 ;
        RECT 17.940 3.910 24.340 4.795 ;
        RECT 17.940 2.125 20.420 3.910 ;
        RECT 21.300 2.125 24.340 3.910 ;
        RECT 25.220 3.595 31.060 4.795 ;
        RECT 25.220 2.125 27.700 3.595 ;
        RECT 28.580 2.125 31.060 3.595 ;
        RECT 31.940 2.125 34.420 4.795 ;
        RECT 35.300 4.800 41.700 9.845 ;
        RECT 35.300 2.125 38.340 4.800 ;
        RECT 39.220 2.125 41.700 4.800 ;
        RECT 42.580 4.795 48.420 9.845 ;
        RECT 42.580 2.125 45.060 4.795 ;
        RECT 45.940 2.125 48.420 4.795 ;
        RECT 49.300 4.795 55.700 9.845 ;
        RECT 49.300 2.125 51.780 4.795 ;
        RECT 52.660 2.125 55.700 4.795 ;
        RECT 56.580 4.795 62.420 9.845 ;
        RECT 56.580 2.125 59.060 4.795 ;
        RECT 59.940 2.125 62.420 4.795 ;
        RECT 63.300 4.795 108.080 9.845 ;
        RECT 63.300 4.690 73.060 4.795 ;
        RECT 63.300 2.125 65.780 4.690 ;
        RECT 66.660 3.345 73.060 4.690 ;
        RECT 66.660 2.125 69.700 3.345 ;
        RECT 70.580 2.125 73.060 3.345 ;
        RECT 73.940 3.845 79.780 4.795 ;
        RECT 73.940 2.125 76.420 3.845 ;
        RECT 77.300 2.125 79.780 3.845 ;
        RECT 80.660 3.885 87.060 4.795 ;
        RECT 80.660 2.125 83.140 3.885 ;
        RECT 84.020 2.125 87.060 3.885 ;
        RECT 87.940 4.195 107.780 4.795 ;
        RECT 87.940 4.170 97.140 4.195 ;
        RECT 87.940 2.125 90.420 4.170 ;
        RECT 91.300 3.955 97.140 4.170 ;
        RECT 91.300 2.125 93.780 3.955 ;
        RECT 94.660 2.125 97.140 3.955 ;
        RECT 98.020 4.145 107.780 4.195 ;
        RECT 98.020 4.135 104.420 4.145 ;
        RECT 98.020 2.125 101.060 4.135 ;
        RECT 101.940 2.125 104.420 4.135 ;
        RECT 105.300 2.125 107.780 4.145 ;
      LAYER Metal3 ;
        RECT 8.480 2.125 100.070 11.565 ;
      LAYER Metal4 ;
        RECT 8.480 2.125 100.065 11.565 ;
      LAYER Metal5 ;
        RECT 3.705 8.225 104.580 11.565 ;
        RECT 31.545 5.625 104.580 8.225 ;
        RECT 3.705 4.225 104.580 5.625 ;
        RECT 9.045 2.125 104.580 4.225 ;
  END
END user_id_programming
END LIBRARY

