VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO copyright_block
  CLASS BLOCK ;
  FOREIGN copyright_block ;
  ORIGIN 0.000 0.000 ;
  SIZE 40.000 BY 25.000 ;
END copyright_block
END LIBRARY