* Simple Schmitt trigger inverter testbench (No. 1:  Using hand-written netlist)

.include /usr/share/pdk/gf180mcuC/libs.tech/ngspice/design.ngspice
.lib /usr/share/pdk/gf180mcuC/libs.tech/ngspice/sm141064.ngspice typical
.lib /usr/share/pdk/gf180mcuC/libs.tech/ngspice/sm141064.ngspice res_typical
.include simple_por.spice

V0 VDD 0 5
V1 In 0 PWL(0 0 100u 5 200u 5 300u 0)

X0 VDD 0 In Out schmitt_inverter

.control
tran 500n 350u
plot V(In) V(Out)
.endc
