magic
tech gf180mcuC
magscale 1 5
timestamp 1654634570
<< metal5 >>
rect 72 504 252 540
rect 36 468 288 504
rect 0 396 324 468
rect 0 144 108 396
rect 216 144 324 396
rect 0 72 324 144
rect 36 36 324 72
rect 72 0 324 36
rect 180 -108 324 0
rect 0 -144 324 -108
rect 0 -180 288 -144
rect 0 -216 252 -180
<< properties >>
string FIXED_BBOX 0 -216 432 756
<< end >>
