magic
tech gf180mcuC
magscale 1 10
timestamp 1668701476
<< metal1 >>
rect 598 2766 673 3020
rect 916 2887 991 3030
rect 916 2827 923 2887
rect 983 2827 991 2887
rect 916 2806 991 2827
rect 468 2694 673 2766
rect 468 2675 540 2694
rect 468 2010 540 2029
rect 1812 2010 1884 2029
rect 2932 2010 3004 2029
rect 468 1938 673 2010
rect 1812 1938 2017 2010
rect 2932 1938 3137 2010
rect 598 1877 673 1938
rect 598 1817 605 1877
rect 665 1817 673 1877
rect 598 1684 673 1817
rect 916 1674 991 1898
rect 1942 1684 2017 1938
rect 2260 1877 2335 1898
rect 2260 1817 2267 1877
rect 2327 1817 2335 1877
rect 2260 1674 2335 1817
rect 3062 1877 3137 1938
rect 3062 1817 3069 1877
rect 3129 1817 3137 1877
rect 3062 1684 3137 1817
rect 3380 1674 3455 1898
rect 598 1319 673 1452
rect 598 1259 605 1319
rect 665 1259 673 1319
rect 598 1198 673 1259
rect 916 1238 991 1462
rect 1942 1198 2017 1452
rect 2260 1319 2335 1462
rect 2260 1259 2267 1319
rect 2327 1259 2335 1319
rect 2260 1238 2335 1259
rect 3062 1198 3137 1452
rect 3380 1319 3455 1462
rect 3380 1259 3387 1319
rect 3447 1259 3455 1319
rect 3380 1238 3455 1259
rect 468 1126 673 1198
rect 1812 1126 2017 1198
rect 2932 1126 3137 1198
rect 468 1107 540 1126
rect 1812 1107 1884 1126
rect 2932 1107 3004 1126
rect 468 442 540 461
rect 1812 442 1884 461
rect 2932 442 3004 461
rect 468 370 673 442
rect 1812 370 2017 442
rect 2932 370 3137 442
rect 598 309 673 370
rect 598 249 605 309
rect 665 249 673 309
rect 598 116 673 249
rect 916 106 991 330
rect 1942 116 2017 370
rect 2260 309 2335 330
rect 2260 249 2267 309
rect 2327 249 2335 309
rect 2260 106 2335 249
rect 3062 116 3137 370
rect 3380 309 3455 330
rect 3380 249 3387 309
rect 3447 249 3455 309
rect 3380 106 3455 249
<< via1 >>
rect 83 3110 652 3170
rect 923 2827 983 2887
rect 1793 2330 2362 2390
rect 605 1817 665 1877
rect 2267 1817 2327 1877
rect 3069 1817 3129 1877
rect 83 1540 652 1600
rect 605 1259 665 1319
rect 2267 1259 2327 1319
rect 3387 1259 3447 1319
rect 1793 750 2362 810
rect 605 249 665 309
rect 2267 249 2327 309
rect 3387 249 3447 309
rect 92 -29 621 31
<< metal2 >>
rect 70 3170 666 3181
rect 70 3110 83 3170
rect 652 3110 666 3170
rect 70 3098 666 3110
rect 576 2887 1699 2889
rect 576 2827 923 2887
rect 983 2827 1699 2887
rect 576 2825 1699 2827
rect 585 1877 1428 1879
rect 585 1817 605 1877
rect 665 1817 1428 1877
rect 585 1815 1428 1817
rect 70 1600 666 1611
rect 70 1540 83 1600
rect 652 1540 666 1600
rect 70 1528 666 1540
rect 585 1319 1132 1321
rect 585 1259 605 1319
rect 665 1259 1132 1319
rect 585 1257 1132 1259
rect 572 309 1004 311
rect 572 249 605 309
rect 665 249 1004 309
rect 572 247 1004 249
rect 80 31 633 43
rect 80 -29 92 31
rect 621 -29 633 31
rect 80 -40 633 -29
rect 700 -84 756 247
rect 1076 157 1132 1257
rect 1036 97 1132 157
rect 1036 -84 1092 97
rect 1372 -84 1428 1815
rect 1643 496 1699 2825
rect 1780 2390 2376 2401
rect 1780 2330 1793 2390
rect 2362 2330 2376 2390
rect 1780 2318 2376 2330
rect 1929 1877 2772 1879
rect 1929 1817 2267 1877
rect 2327 1817 2772 1877
rect 1929 1815 2772 1817
rect 1929 1319 2496 1321
rect 1929 1259 2267 1319
rect 2327 1259 2496 1319
rect 1929 1257 2496 1259
rect 1780 810 2376 821
rect 1780 750 1793 810
rect 2362 750 2376 810
rect 1780 738 2376 750
rect 1643 440 1764 496
rect 1708 -84 1764 440
rect 1915 309 2348 311
rect 1915 249 2267 309
rect 2327 249 2348 309
rect 1915 247 2348 249
rect 2044 -84 2100 247
rect 2440 174 2496 1257
rect 2380 118 2496 174
rect 2380 -84 2436 118
rect 2716 -84 2772 1815
rect 2921 1877 3468 1879
rect 2921 1817 3069 1877
rect 3129 1817 3468 1877
rect 2921 1815 3468 1817
rect 2921 177 2977 1815
rect 3041 1319 3780 1321
rect 3041 1259 3387 1319
rect 3447 1259 3780 1319
rect 3041 1257 3780 1259
rect 3043 309 3462 311
rect 3043 249 3387 309
rect 3447 249 3462 309
rect 3043 247 3462 249
rect 2921 121 3108 177
rect 3052 -84 3108 121
rect 3388 -84 3444 247
rect 3724 -84 3780 1257
<< via2 >>
rect 83 3110 652 3170
rect 83 1540 652 1600
rect 92 -29 621 31
rect 1793 2330 2362 2390
rect 1793 750 2362 810
<< metal3 >>
rect 66 3170 672 3192
rect 66 3110 83 3170
rect 652 3110 672 3170
rect 66 1600 672 3110
rect 66 1540 83 1600
rect 652 1540 672 1600
rect 66 31 672 1540
rect 66 -29 92 31
rect 621 -29 672 31
rect 66 -53 672 -29
rect 1773 2390 2379 3192
rect 1773 2330 1793 2390
rect 2362 2330 2379 2390
rect 1773 810 2379 2330
rect 1773 750 1793 810
rect 2362 750 2379 810
rect 1773 -53 2379 750
use gf180mcu_fd_sc_mcu7t5v0__endcap  gf180mcu_fd_sc_mcu7t5v0__endcap_0 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1664373539
transform 1 0 0 0 1 0
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  gf180mcu_fd_sc_mcu7t5v0__endcap_1
timestamp 1664373539
transform 1 0 2464 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  gf180mcu_fd_sc_mcu7t5v0__endcap_2
timestamp 1664373539
transform 1 0 3584 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  gf180mcu_fd_sc_mcu7t5v0__endcap_3
timestamp 1664373539
transform 1 0 0 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  gf180mcu_fd_sc_mcu7t5v0__endcap_4
timestamp 1664373539
transform 1 0 0 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  gf180mcu_fd_sc_mcu7t5v0__endcap_5
timestamp 1664373539
transform 1 0 2464 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  gf180mcu_fd_sc_mcu7t5v0__endcap_6
timestamp 1664373539
transform 1 0 3584 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  gf180mcu_fd_sc_mcu7t5v0__fillcap_4_0 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1664373539
transform 1 0 1120 0 1 0
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  gf180mcu_fd_sc_mcu7t5v0__fillcap_4_1
timestamp 1664373539
transform 1 0 1120 0 -1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  gf180mcu_fd_sc_mcu7t5v0__fillcap_4_2
timestamp 1664373539
transform 1 0 2016 0 -1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  gf180mcu_fd_sc_mcu7t5v0__fillcap_4_3
timestamp 1664373539
transform 1 0 1120 0 -1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  gf180mcu_fd_sc_mcu7t5v0__fillcap_4_4
timestamp 1664373539
transform 1 0 3136 0 -1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  gf180mcu_fd_sc_mcu7t5v0__fillcap_4_5
timestamp 1664373539
transform 1 0 1568 0 -1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  gf180mcu_fd_sc_mcu7t5v0__fillcap_4_6
timestamp 1664373539
transform 1 0 1120 0 1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  gf180mcu_fd_sc_mcu7t5v0__fillcap_4_7
timestamp 1664373539
transform 1 0 2688 0 -1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  gf180mcu_fd_sc_mcu7t5v0__filltie_0 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1664373539
transform 1 0 2464 0 1 0
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  gf180mcu_fd_sc_mcu7t5v0__filltie_1
timestamp 1664373539
transform 1 0 3584 0 1 0
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  gf180mcu_fd_sc_mcu7t5v0__filltie_2
timestamp 1664373539
transform 1 0 3584 0 -1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  gf180mcu_fd_sc_mcu7t5v0__filltie_4
timestamp 1664373539
transform 1 0 0 0 -1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  gf180mcu_fd_sc_mcu7t5v0__filltie_5
timestamp 1664373539
transform 1 0 2464 0 -1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  gf180mcu_fd_sc_mcu7t5v0__tieh_0 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1664373539
transform 1 0 224 0 1 0
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  gf180mcu_fd_sc_mcu7t5v0__tieh_1
timestamp 1664373539
transform 1 0 1568 0 1 0
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  gf180mcu_fd_sc_mcu7t5v0__tieh_2
timestamp 1664373539
transform 1 0 2688 0 1 0
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  gf180mcu_fd_sc_mcu7t5v0__tieh_4
timestamp 1664373539
transform 1 0 2688 0 -1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  gf180mcu_fd_sc_mcu7t5v0__tieh_7
timestamp 1664373539
transform 1 0 224 0 -1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  gf180mcu_fd_sc_mcu7t5v0__tieh_8
timestamp 1664373539
transform 1 0 224 0 1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  gf180mcu_fd_sc_mcu7t5v0__tieh_9
timestamp 1664373539
transform 1 0 1568 0 1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  gf180mcu_fd_sc_mcu7t5v0__tieh_11
timestamp 1664373539
transform 1 0 2688 0 1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  gf180mcu_fd_sc_mcu7t5v0__tieh_12
timestamp 1664373539
transform 1 0 1568 0 -1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  gf180mcu_fd_sc_mcu7t5v0__tieh_13
timestamp 1664373539
transform 1 0 224 0 -1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  gf180mcu_fd_sc_mcu7t5v0__tiel_0 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1664373539
transform 1 0 672 0 1 0
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  gf180mcu_fd_sc_mcu7t5v0__tiel_1
timestamp 1664373539
transform 1 0 2016 0 1 0
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  gf180mcu_fd_sc_mcu7t5v0__tiel_2
timestamp 1664373539
transform 1 0 3136 0 1 0
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  gf180mcu_fd_sc_mcu7t5v0__tiel_4
timestamp 1664373539
transform 1 0 3136 0 -1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  gf180mcu_fd_sc_mcu7t5v0__tiel_7
timestamp 1664373539
transform 1 0 672 0 -1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  gf180mcu_fd_sc_mcu7t5v0__tiel_8
timestamp 1664373539
transform 1 0 672 0 1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  gf180mcu_fd_sc_mcu7t5v0__tiel_9
timestamp 1664373539
transform 1 0 2016 0 1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  gf180mcu_fd_sc_mcu7t5v0__tiel_11
timestamp 1664373539
transform 1 0 3136 0 1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  gf180mcu_fd_sc_mcu7t5v0__tiel_12
timestamp 1664373539
transform 1 0 2016 0 -1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  gf180mcu_fd_sc_mcu7t5v0__tiel_13
timestamp 1664373539
transform 1 0 672 0 -1 1568
box -86 -86 534 870
<< labels >>
flabel metal3 1773 -53 2379 750 0 FreeSans 1600 0 0 0 VDD
port 11 nsew
flabel metal3 66 55 672 858 0 FreeSans 1600 0 0 0 VSS
port 12 nsew
flabel metal2 700 -84 756 150 0 FreeSans 400 90 0 0 gpio_defaults[0]
port 1 nsew
flabel metal2 1036 -84 1092 150 0 FreeSans 400 90 0 0 gpio_defaults[1]
port 5 nsew
flabel metal2 1372 -84 1428 150 0 FreeSans 400 90 0 0 gpio_defaults[2]
port 9 nsew
flabel metal2 1708 -84 1764 150 0 FreeSans 400 90 0 0 gpio_defaults[3]
port 8 nsew
flabel metal2 2044 -84 2100 150 0 FreeSans 400 90 0 0 gpio_defaults[4]
port 2 nsew
flabel metal2 2380 -84 2436 150 0 FreeSans 400 90 0 0 gpio_defaults[5]
port 6 nsew
flabel metal2 2716 -84 2772 150 0 FreeSans 400 90 0 0 gpio_defaults[6]
port 10 nsew
flabel metal2 3052 -84 3108 150 0 FreeSans 400 90 0 0 gpio_defaults[7]
port 4 nsew
flabel metal2 3388 -84 3444 150 0 FreeSans 400 90 0 0 gpio_defaults[8]
port 3 nsew
flabel metal2 3724 -84 3780 150 0 FreeSans 400 90 0 0 gpio_defaults[9]
port 7 nsew
<< end >>
