magic
tech gf180mcuC
magscale 1 5
timestamp 1654634570
<< metal5 >>
rect 0 324 432 432
<< properties >>
string FIXED_BBOX 0 -216 540 756
<< end >>
