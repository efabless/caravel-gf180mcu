magic
tech gf180mcuC
magscale 1 10
timestamp 1483923398
<< checkpaint >>
rect 67800 67800 710200 952200
<< metal2 >>
rect 381272 949926 383172 950200
rect 381272 949870 381342 949926
rect 381398 949870 381466 949926
rect 381522 949870 381590 949926
rect 381646 949870 381714 949926
rect 381770 949870 381838 949926
rect 381894 949870 381962 949926
rect 382018 949870 382086 949926
rect 382142 949870 382210 949926
rect 382266 949870 382334 949926
rect 382390 949870 382458 949926
rect 382514 949870 382582 949926
rect 382638 949870 382706 949926
rect 382762 949870 382830 949926
rect 382886 949870 382954 949926
rect 383010 949870 383078 949926
rect 383134 949870 383172 949926
rect 381272 949800 383172 949870
rect 383752 949926 385802 950200
rect 383752 949870 383822 949926
rect 383878 949870 383946 949926
rect 384002 949870 384070 949926
rect 384126 949870 384194 949926
rect 384250 949870 384318 949926
rect 384374 949870 384442 949926
rect 384498 949870 384566 949926
rect 384622 949870 384690 949926
rect 384746 949870 384814 949926
rect 384870 949870 384938 949926
rect 384994 949870 385062 949926
rect 385118 949870 385186 949926
rect 385242 949870 385310 949926
rect 385366 949870 385434 949926
rect 385490 949870 385558 949926
rect 385614 949870 385682 949926
rect 385738 949870 385802 949926
rect 383752 949800 385802 949870
rect 386122 949926 388172 950200
rect 386122 949870 386192 949926
rect 386248 949870 386316 949926
rect 386372 949870 386440 949926
rect 386496 949870 386564 949926
rect 386620 949870 386688 949926
rect 386744 949870 386812 949926
rect 386868 949870 386936 949926
rect 386992 949870 387060 949926
rect 387116 949870 387184 949926
rect 387240 949870 387308 949926
rect 387364 949870 387432 949926
rect 387488 949870 387556 949926
rect 387612 949870 387680 949926
rect 387736 949870 387804 949926
rect 387860 949870 387928 949926
rect 387984 949870 388052 949926
rect 388108 949870 388172 949926
rect 386122 949800 388172 949870
rect 388828 949926 390878 950200
rect 388828 949870 388892 949926
rect 388948 949870 389016 949926
rect 389072 949870 389140 949926
rect 389196 949870 389264 949926
rect 389320 949870 389388 949926
rect 389444 949870 389512 949926
rect 389568 949870 389636 949926
rect 389692 949870 389760 949926
rect 389816 949870 389884 949926
rect 389940 949870 390008 949926
rect 390064 949870 390132 949926
rect 390188 949870 390256 949926
rect 390312 949870 390380 949926
rect 390436 949870 390504 949926
rect 390560 949870 390628 949926
rect 390684 949870 390752 949926
rect 390808 949870 390878 949926
rect 388828 949800 390878 949870
rect 391198 949926 393248 950200
rect 391198 949870 391262 949926
rect 391318 949870 391386 949926
rect 391442 949870 391510 949926
rect 391566 949870 391634 949926
rect 391690 949870 391758 949926
rect 391814 949870 391882 949926
rect 391938 949870 392006 949926
rect 392062 949870 392130 949926
rect 392186 949870 392254 949926
rect 392310 949870 392378 949926
rect 392434 949870 392502 949926
rect 392558 949870 392626 949926
rect 392682 949870 392750 949926
rect 392806 949870 392874 949926
rect 392930 949870 392998 949926
rect 393054 949870 393122 949926
rect 393178 949870 393248 949926
rect 391198 949800 393248 949870
rect 393828 949926 395728 950200
rect 393828 949870 393866 949926
rect 393922 949870 393990 949926
rect 394046 949870 394114 949926
rect 394170 949870 394238 949926
rect 394294 949870 394362 949926
rect 394418 949870 394486 949926
rect 394542 949870 394610 949926
rect 394666 949870 394734 949926
rect 394790 949870 394858 949926
rect 394914 949870 394982 949926
rect 395038 949870 395106 949926
rect 395162 949870 395230 949926
rect 395286 949870 395354 949926
rect 395410 949870 395478 949926
rect 395534 949870 395602 949926
rect 395658 949870 395728 949926
rect 393828 949800 395728 949870
rect 601272 949926 603172 950200
rect 601272 949870 601342 949926
rect 601398 949870 601466 949926
rect 601522 949870 601590 949926
rect 601646 949870 601714 949926
rect 601770 949870 601838 949926
rect 601894 949870 601962 949926
rect 602018 949870 602086 949926
rect 602142 949870 602210 949926
rect 602266 949870 602334 949926
rect 602390 949870 602458 949926
rect 602514 949870 602582 949926
rect 602638 949870 602706 949926
rect 602762 949870 602830 949926
rect 602886 949870 602954 949926
rect 603010 949870 603078 949926
rect 603134 949870 603172 949926
rect 601272 949800 603172 949870
rect 603752 949926 605802 950200
rect 603752 949870 603822 949926
rect 603878 949870 603946 949926
rect 604002 949870 604070 949926
rect 604126 949870 604194 949926
rect 604250 949870 604318 949926
rect 604374 949870 604442 949926
rect 604498 949870 604566 949926
rect 604622 949870 604690 949926
rect 604746 949870 604814 949926
rect 604870 949870 604938 949926
rect 604994 949870 605062 949926
rect 605118 949870 605186 949926
rect 605242 949870 605310 949926
rect 605366 949870 605434 949926
rect 605490 949870 605558 949926
rect 605614 949870 605682 949926
rect 605738 949870 605802 949926
rect 603752 949800 605802 949870
rect 606122 949926 608172 950200
rect 606122 949870 606192 949926
rect 606248 949870 606316 949926
rect 606372 949870 606440 949926
rect 606496 949870 606564 949926
rect 606620 949870 606688 949926
rect 606744 949870 606812 949926
rect 606868 949870 606936 949926
rect 606992 949870 607060 949926
rect 607116 949870 607184 949926
rect 607240 949870 607308 949926
rect 607364 949870 607432 949926
rect 607488 949870 607556 949926
rect 607612 949870 607680 949926
rect 607736 949870 607804 949926
rect 607860 949870 607928 949926
rect 607984 949870 608052 949926
rect 608108 949870 608172 949926
rect 606122 949800 608172 949870
rect 608828 949926 610878 950200
rect 608828 949870 608892 949926
rect 608948 949870 609016 949926
rect 609072 949870 609140 949926
rect 609196 949870 609264 949926
rect 609320 949870 609388 949926
rect 609444 949870 609512 949926
rect 609568 949870 609636 949926
rect 609692 949870 609760 949926
rect 609816 949870 609884 949926
rect 609940 949870 610008 949926
rect 610064 949870 610132 949926
rect 610188 949870 610256 949926
rect 610312 949870 610380 949926
rect 610436 949870 610504 949926
rect 610560 949870 610628 949926
rect 610684 949870 610752 949926
rect 610808 949870 610878 949926
rect 608828 949800 610878 949870
rect 611198 949926 613248 950200
rect 611198 949870 611262 949926
rect 611318 949870 611386 949926
rect 611442 949870 611510 949926
rect 611566 949870 611634 949926
rect 611690 949870 611758 949926
rect 611814 949870 611882 949926
rect 611938 949870 612006 949926
rect 612062 949870 612130 949926
rect 612186 949870 612254 949926
rect 612310 949870 612378 949926
rect 612434 949870 612502 949926
rect 612558 949870 612626 949926
rect 612682 949870 612750 949926
rect 612806 949870 612874 949926
rect 612930 949870 612998 949926
rect 613054 949870 613122 949926
rect 613178 949870 613248 949926
rect 611198 949800 613248 949870
rect 613828 949926 615728 950200
rect 613828 949870 613866 949926
rect 613922 949870 613990 949926
rect 614046 949870 614114 949926
rect 614170 949870 614238 949926
rect 614294 949870 614362 949926
rect 614418 949870 614486 949926
rect 614542 949870 614610 949926
rect 614666 949870 614734 949926
rect 614790 949870 614858 949926
rect 614914 949870 614982 949926
rect 615038 949870 615106 949926
rect 615162 949870 615230 949926
rect 615286 949870 615354 949926
rect 615410 949870 615478 949926
rect 615534 949870 615602 949926
rect 615658 949870 615728 949926
rect 613828 949800 615728 949870
rect 69800 884658 70200 884728
rect 69800 884602 70074 884658
rect 70130 884602 70200 884658
rect 69800 884534 70200 884602
rect 69800 884478 70074 884534
rect 70130 884478 70200 884534
rect 69800 884410 70200 884478
rect 69800 884354 70074 884410
rect 70130 884354 70200 884410
rect 69800 884286 70200 884354
rect 69800 884230 70074 884286
rect 70130 884230 70200 884286
rect 69800 884162 70200 884230
rect 69800 884106 70074 884162
rect 70130 884106 70200 884162
rect 69800 884038 70200 884106
rect 69800 883982 70074 884038
rect 70130 883982 70200 884038
rect 69800 883914 70200 883982
rect 69800 883858 70074 883914
rect 70130 883858 70200 883914
rect 69800 883790 70200 883858
rect 69800 883734 70074 883790
rect 70130 883734 70200 883790
rect 69800 883666 70200 883734
rect 69800 883610 70074 883666
rect 70130 883610 70200 883666
rect 69800 883542 70200 883610
rect 69800 883486 70074 883542
rect 70130 883486 70200 883542
rect 69800 883418 70200 883486
rect 69800 883362 70074 883418
rect 70130 883362 70200 883418
rect 69800 883294 70200 883362
rect 69800 883238 70074 883294
rect 70130 883238 70200 883294
rect 69800 883170 70200 883238
rect 69800 883114 70074 883170
rect 70130 883114 70200 883170
rect 69800 883046 70200 883114
rect 69800 882990 70074 883046
rect 70130 882990 70200 883046
rect 69800 882922 70200 882990
rect 69800 882866 70074 882922
rect 70130 882866 70200 882922
rect 69800 882828 70200 882866
rect 707800 883658 708200 883728
rect 707800 883602 707870 883658
rect 707926 883602 708200 883658
rect 707800 883534 708200 883602
rect 707800 883478 707870 883534
rect 707926 883478 708200 883534
rect 707800 883410 708200 883478
rect 707800 883354 707870 883410
rect 707926 883354 708200 883410
rect 707800 883286 708200 883354
rect 707800 883230 707870 883286
rect 707926 883230 708200 883286
rect 707800 883162 708200 883230
rect 707800 883106 707870 883162
rect 707926 883106 708200 883162
rect 707800 883038 708200 883106
rect 707800 882982 707870 883038
rect 707926 882982 708200 883038
rect 707800 882914 708200 882982
rect 707800 882858 707870 882914
rect 707926 882858 708200 882914
rect 707800 882790 708200 882858
rect 707800 882734 707870 882790
rect 707926 882734 708200 882790
rect 707800 882666 708200 882734
rect 707800 882610 707870 882666
rect 707926 882610 708200 882666
rect 707800 882542 708200 882610
rect 707800 882486 707870 882542
rect 707926 882486 708200 882542
rect 707800 882418 708200 882486
rect 707800 882362 707870 882418
rect 707926 882362 708200 882418
rect 707800 882294 708200 882362
rect 69800 882184 70200 882248
rect 69800 882128 70074 882184
rect 70130 882128 70200 882184
rect 69800 882060 70200 882128
rect 69800 882004 70074 882060
rect 70130 882004 70200 882060
rect 69800 881936 70200 882004
rect 69800 881880 70074 881936
rect 70130 881880 70200 881936
rect 69800 881812 70200 881880
rect 707800 882238 707870 882294
rect 707926 882238 708200 882294
rect 707800 882170 708200 882238
rect 707800 882114 707870 882170
rect 707926 882114 708200 882170
rect 707800 882046 708200 882114
rect 707800 881990 707870 882046
rect 707926 881990 708200 882046
rect 707800 881922 708200 881990
rect 707800 881866 707870 881922
rect 707926 881866 708200 881922
rect 707800 881828 708200 881866
rect 69800 881756 70074 881812
rect 70130 881756 70200 881812
rect 69800 881688 70200 881756
rect 69800 881632 70074 881688
rect 70130 881632 70200 881688
rect 69800 881564 70200 881632
rect 69800 881508 70074 881564
rect 70130 881508 70200 881564
rect 69800 881440 70200 881508
rect 69800 881384 70074 881440
rect 70130 881384 70200 881440
rect 69800 881316 70200 881384
rect 69800 881260 70074 881316
rect 70130 881260 70200 881316
rect 69800 881192 70200 881260
rect 69800 881136 70074 881192
rect 70130 881136 70200 881192
rect 69800 881068 70200 881136
rect 69800 881012 70074 881068
rect 70130 881012 70200 881068
rect 69800 880944 70200 881012
rect 69800 880888 70074 880944
rect 70130 880888 70200 880944
rect 69800 880820 70200 880888
rect 69800 880764 70074 880820
rect 70130 880764 70200 880820
rect 69800 880696 70200 880764
rect 69800 880640 70074 880696
rect 70130 880640 70200 880696
rect 69800 880572 70200 880640
rect 69800 880516 70074 880572
rect 70130 880516 70200 880572
rect 69800 880448 70200 880516
rect 69800 880392 70074 880448
rect 70130 880392 70200 880448
rect 69800 880324 70200 880392
rect 69800 880268 70074 880324
rect 70130 880268 70200 880324
rect 69800 880198 70200 880268
rect 707800 881178 708200 881248
rect 707800 881122 707870 881178
rect 707926 881122 708200 881178
rect 707800 881054 708200 881122
rect 707800 880998 707870 881054
rect 707926 880998 708200 881054
rect 707800 880930 708200 880998
rect 707800 880874 707870 880930
rect 707926 880874 708200 880930
rect 707800 880806 708200 880874
rect 707800 880750 707870 880806
rect 707926 880750 708200 880806
rect 707800 880682 708200 880750
rect 707800 880626 707870 880682
rect 707926 880626 708200 880682
rect 707800 880558 708200 880626
rect 707800 880502 707870 880558
rect 707926 880502 708200 880558
rect 707800 880434 708200 880502
rect 707800 880378 707870 880434
rect 707926 880378 708200 880434
rect 707800 880310 708200 880378
rect 707800 880254 707870 880310
rect 707926 880254 708200 880310
rect 707800 880186 708200 880254
rect 707800 880130 707870 880186
rect 707926 880130 708200 880186
rect 707800 880062 708200 880130
rect 707800 880006 707870 880062
rect 707926 880006 708200 880062
rect 707800 879938 708200 880006
rect 707800 879882 707870 879938
rect 707926 879882 708200 879938
rect 69800 879814 70200 879878
rect 69800 879758 70074 879814
rect 70130 879758 70200 879814
rect 69800 879690 70200 879758
rect 69800 879634 70074 879690
rect 70130 879634 70200 879690
rect 69800 879566 70200 879634
rect 69800 879510 70074 879566
rect 70130 879510 70200 879566
rect 69800 879442 70200 879510
rect 69800 879386 70074 879442
rect 70130 879386 70200 879442
rect 69800 879318 70200 879386
rect 69800 879262 70074 879318
rect 70130 879262 70200 879318
rect 69800 879194 70200 879262
rect 707800 879814 708200 879882
rect 707800 879758 707870 879814
rect 707926 879758 708200 879814
rect 707800 879690 708200 879758
rect 707800 879634 707870 879690
rect 707926 879634 708200 879690
rect 707800 879566 708200 879634
rect 707800 879510 707870 879566
rect 707926 879510 708200 879566
rect 707800 879442 708200 879510
rect 707800 879386 707870 879442
rect 707926 879386 708200 879442
rect 707800 879318 708200 879386
rect 707800 879262 707870 879318
rect 707926 879262 708200 879318
rect 707800 879198 708200 879262
rect 69800 879138 70074 879194
rect 70130 879138 70200 879194
rect 69800 879070 70200 879138
rect 69800 879014 70074 879070
rect 70130 879014 70200 879070
rect 69800 878946 70200 879014
rect 69800 878890 70074 878946
rect 70130 878890 70200 878946
rect 69800 878822 70200 878890
rect 69800 878766 70074 878822
rect 70130 878766 70200 878822
rect 69800 878698 70200 878766
rect 69800 878642 70074 878698
rect 70130 878642 70200 878698
rect 69800 878574 70200 878642
rect 69800 878518 70074 878574
rect 70130 878518 70200 878574
rect 69800 878450 70200 878518
rect 69800 878394 70074 878450
rect 70130 878394 70200 878450
rect 69800 878326 70200 878394
rect 69800 878270 70074 878326
rect 70130 878270 70200 878326
rect 69800 878202 70200 878270
rect 69800 878146 70074 878202
rect 70130 878146 70200 878202
rect 69800 878078 70200 878146
rect 69800 878022 70074 878078
rect 70130 878022 70200 878078
rect 69800 877954 70200 878022
rect 69800 877898 70074 877954
rect 70130 877898 70200 877954
rect 69800 877828 70200 877898
rect 707800 878808 708200 878878
rect 707800 878752 707870 878808
rect 707926 878752 708200 878808
rect 707800 878684 708200 878752
rect 707800 878628 707870 878684
rect 707926 878628 708200 878684
rect 707800 878560 708200 878628
rect 707800 878504 707870 878560
rect 707926 878504 708200 878560
rect 707800 878436 708200 878504
rect 707800 878380 707870 878436
rect 707926 878380 708200 878436
rect 707800 878312 708200 878380
rect 707800 878256 707870 878312
rect 707926 878256 708200 878312
rect 707800 878188 708200 878256
rect 707800 878132 707870 878188
rect 707926 878132 708200 878188
rect 707800 878064 708200 878132
rect 707800 878008 707870 878064
rect 707926 878008 708200 878064
rect 707800 877940 708200 878008
rect 707800 877884 707870 877940
rect 707926 877884 708200 877940
rect 707800 877816 708200 877884
rect 707800 877760 707870 877816
rect 707926 877760 708200 877816
rect 707800 877692 708200 877760
rect 707800 877636 707870 877692
rect 707926 877636 708200 877692
rect 707800 877568 708200 877636
rect 707800 877512 707870 877568
rect 707926 877512 708200 877568
rect 707800 877444 708200 877512
rect 707800 877388 707870 877444
rect 707926 877388 708200 877444
rect 707800 877320 708200 877388
rect 707800 877264 707870 877320
rect 707926 877264 708200 877320
rect 707800 877196 708200 877264
rect 69800 877108 70200 877172
rect 69800 877052 70074 877108
rect 70130 877052 70200 877108
rect 69800 876984 70200 877052
rect 69800 876928 70074 876984
rect 70130 876928 70200 876984
rect 69800 876860 70200 876928
rect 69800 876804 70074 876860
rect 70130 876804 70200 876860
rect 707800 877140 707870 877196
rect 707926 877140 708200 877196
rect 707800 877072 708200 877140
rect 707800 877016 707870 877072
rect 707926 877016 708200 877072
rect 707800 876948 708200 877016
rect 707800 876892 707870 876948
rect 707926 876892 708200 876948
rect 707800 876828 708200 876892
rect 69800 876736 70200 876804
rect 69800 876680 70074 876736
rect 70130 876680 70200 876736
rect 69800 876612 70200 876680
rect 69800 876556 70074 876612
rect 70130 876556 70200 876612
rect 69800 876488 70200 876556
rect 69800 876432 70074 876488
rect 70130 876432 70200 876488
rect 69800 876364 70200 876432
rect 69800 876308 70074 876364
rect 70130 876308 70200 876364
rect 69800 876240 70200 876308
rect 69800 876184 70074 876240
rect 70130 876184 70200 876240
rect 69800 876116 70200 876184
rect 69800 876060 70074 876116
rect 70130 876060 70200 876116
rect 69800 875992 70200 876060
rect 69800 875936 70074 875992
rect 70130 875936 70200 875992
rect 69800 875868 70200 875936
rect 69800 875812 70074 875868
rect 70130 875812 70200 875868
rect 69800 875744 70200 875812
rect 69800 875688 70074 875744
rect 70130 875688 70200 875744
rect 69800 875620 70200 875688
rect 69800 875564 70074 875620
rect 70130 875564 70200 875620
rect 69800 875496 70200 875564
rect 69800 875440 70074 875496
rect 70130 875440 70200 875496
rect 69800 875372 70200 875440
rect 69800 875316 70074 875372
rect 70130 875316 70200 875372
rect 69800 875248 70200 875316
rect 69800 875192 70074 875248
rect 70130 875192 70200 875248
rect 69800 875122 70200 875192
rect 707800 876102 708200 876172
rect 707800 876046 707870 876102
rect 707926 876046 708200 876102
rect 707800 875978 708200 876046
rect 707800 875922 707870 875978
rect 707926 875922 708200 875978
rect 707800 875854 708200 875922
rect 707800 875798 707870 875854
rect 707926 875798 708200 875854
rect 707800 875730 708200 875798
rect 707800 875674 707870 875730
rect 707926 875674 708200 875730
rect 707800 875606 708200 875674
rect 707800 875550 707870 875606
rect 707926 875550 708200 875606
rect 707800 875482 708200 875550
rect 707800 875426 707870 875482
rect 707926 875426 708200 875482
rect 707800 875358 708200 875426
rect 707800 875302 707870 875358
rect 707926 875302 708200 875358
rect 707800 875234 708200 875302
rect 707800 875178 707870 875234
rect 707926 875178 708200 875234
rect 707800 875110 708200 875178
rect 707800 875054 707870 875110
rect 707926 875054 708200 875110
rect 707800 874986 708200 875054
rect 707800 874930 707870 874986
rect 707926 874930 708200 874986
rect 707800 874862 708200 874930
rect 707800 874806 707870 874862
rect 707926 874806 708200 874862
rect 69800 874738 70200 874802
rect 69800 874682 70074 874738
rect 70130 874682 70200 874738
rect 69800 874614 70200 874682
rect 69800 874558 70074 874614
rect 70130 874558 70200 874614
rect 69800 874490 70200 874558
rect 69800 874434 70074 874490
rect 70130 874434 70200 874490
rect 69800 874366 70200 874434
rect 69800 874310 70074 874366
rect 70130 874310 70200 874366
rect 69800 874242 70200 874310
rect 69800 874186 70074 874242
rect 70130 874186 70200 874242
rect 69800 874118 70200 874186
rect 707800 874738 708200 874806
rect 707800 874682 707870 874738
rect 707926 874682 708200 874738
rect 707800 874614 708200 874682
rect 707800 874558 707870 874614
rect 707926 874558 708200 874614
rect 707800 874490 708200 874558
rect 707800 874434 707870 874490
rect 707926 874434 708200 874490
rect 707800 874366 708200 874434
rect 707800 874310 707870 874366
rect 707926 874310 708200 874366
rect 707800 874242 708200 874310
rect 707800 874186 707870 874242
rect 707926 874186 708200 874242
rect 707800 874122 708200 874186
rect 69800 874062 70074 874118
rect 70130 874062 70200 874118
rect 69800 873994 70200 874062
rect 69800 873938 70074 873994
rect 70130 873938 70200 873994
rect 69800 873870 70200 873938
rect 69800 873814 70074 873870
rect 70130 873814 70200 873870
rect 69800 873746 70200 873814
rect 69800 873690 70074 873746
rect 70130 873690 70200 873746
rect 69800 873622 70200 873690
rect 69800 873566 70074 873622
rect 70130 873566 70200 873622
rect 69800 873498 70200 873566
rect 69800 873442 70074 873498
rect 70130 873442 70200 873498
rect 69800 873374 70200 873442
rect 69800 873318 70074 873374
rect 70130 873318 70200 873374
rect 69800 873250 70200 873318
rect 69800 873194 70074 873250
rect 70130 873194 70200 873250
rect 69800 873126 70200 873194
rect 69800 873070 70074 873126
rect 70130 873070 70200 873126
rect 69800 873002 70200 873070
rect 69800 872946 70074 873002
rect 70130 872946 70200 873002
rect 69800 872878 70200 872946
rect 69800 872822 70074 872878
rect 70130 872822 70200 872878
rect 69800 872752 70200 872822
rect 707800 873732 708200 873802
rect 707800 873676 707870 873732
rect 707926 873676 708200 873732
rect 707800 873608 708200 873676
rect 707800 873552 707870 873608
rect 707926 873552 708200 873608
rect 707800 873484 708200 873552
rect 707800 873428 707870 873484
rect 707926 873428 708200 873484
rect 707800 873360 708200 873428
rect 707800 873304 707870 873360
rect 707926 873304 708200 873360
rect 707800 873236 708200 873304
rect 707800 873180 707870 873236
rect 707926 873180 708200 873236
rect 707800 873112 708200 873180
rect 707800 873056 707870 873112
rect 707926 873056 708200 873112
rect 707800 872988 708200 873056
rect 707800 872932 707870 872988
rect 707926 872932 708200 872988
rect 707800 872864 708200 872932
rect 707800 872808 707870 872864
rect 707926 872808 708200 872864
rect 707800 872740 708200 872808
rect 707800 872684 707870 872740
rect 707926 872684 708200 872740
rect 707800 872616 708200 872684
rect 707800 872560 707870 872616
rect 707926 872560 708200 872616
rect 707800 872492 708200 872560
rect 707800 872436 707870 872492
rect 707926 872436 708200 872492
rect 707800 872368 708200 872436
rect 707800 872312 707870 872368
rect 707926 872312 708200 872368
rect 707800 872244 708200 872312
rect 707800 872188 707870 872244
rect 707926 872188 708200 872244
rect 69800 872134 70200 872172
rect 69800 872078 70074 872134
rect 70130 872078 70200 872134
rect 69800 872010 70200 872078
rect 69800 871954 70074 872010
rect 70130 871954 70200 872010
rect 69800 871886 70200 871954
rect 69800 871830 70074 871886
rect 70130 871830 70200 871886
rect 69800 871762 70200 871830
rect 69800 871706 70074 871762
rect 70130 871706 70200 871762
rect 707800 872120 708200 872188
rect 707800 872064 707870 872120
rect 707926 872064 708200 872120
rect 707800 871996 708200 872064
rect 707800 871940 707870 871996
rect 707926 871940 708200 871996
rect 707800 871872 708200 871940
rect 707800 871816 707870 871872
rect 707926 871816 708200 871872
rect 707800 871752 708200 871816
rect 69800 871638 70200 871706
rect 69800 871582 70074 871638
rect 70130 871582 70200 871638
rect 69800 871514 70200 871582
rect 69800 871458 70074 871514
rect 70130 871458 70200 871514
rect 69800 871390 70200 871458
rect 69800 871334 70074 871390
rect 70130 871334 70200 871390
rect 69800 871266 70200 871334
rect 69800 871210 70074 871266
rect 70130 871210 70200 871266
rect 69800 871142 70200 871210
rect 69800 871086 70074 871142
rect 70130 871086 70200 871142
rect 69800 871018 70200 871086
rect 69800 870962 70074 871018
rect 70130 870962 70200 871018
rect 69800 870894 70200 870962
rect 69800 870838 70074 870894
rect 70130 870838 70200 870894
rect 69800 870770 70200 870838
rect 69800 870714 70074 870770
rect 70130 870714 70200 870770
rect 69800 870646 70200 870714
rect 69800 870590 70074 870646
rect 70130 870590 70200 870646
rect 69800 870522 70200 870590
rect 69800 870466 70074 870522
rect 70130 870466 70200 870522
rect 69800 870398 70200 870466
rect 69800 870342 70074 870398
rect 70130 870342 70200 870398
rect 69800 870272 70200 870342
rect 707800 871134 708200 871172
rect 707800 871078 707870 871134
rect 707926 871078 708200 871134
rect 707800 871010 708200 871078
rect 707800 870954 707870 871010
rect 707926 870954 708200 871010
rect 707800 870886 708200 870954
rect 707800 870830 707870 870886
rect 707926 870830 708200 870886
rect 707800 870762 708200 870830
rect 707800 870706 707870 870762
rect 707926 870706 708200 870762
rect 707800 870638 708200 870706
rect 707800 870582 707870 870638
rect 707926 870582 708200 870638
rect 707800 870514 708200 870582
rect 707800 870458 707870 870514
rect 707926 870458 708200 870514
rect 707800 870390 708200 870458
rect 707800 870334 707870 870390
rect 707926 870334 708200 870390
rect 707800 870266 708200 870334
rect 707800 870210 707870 870266
rect 707926 870210 708200 870266
rect 707800 870142 708200 870210
rect 707800 870086 707870 870142
rect 707926 870086 708200 870142
rect 707800 870018 708200 870086
rect 707800 869962 707870 870018
rect 707926 869962 708200 870018
rect 707800 869894 708200 869962
rect 707800 869838 707870 869894
rect 707926 869838 708200 869894
rect 707800 869770 708200 869838
rect 707800 869714 707870 869770
rect 707926 869714 708200 869770
rect 707800 869646 708200 869714
rect 707800 869590 707870 869646
rect 707926 869590 708200 869646
rect 707800 869522 708200 869590
rect 707800 869466 707870 869522
rect 707926 869466 708200 869522
rect 707800 869398 708200 869466
rect 707800 869342 707870 869398
rect 707926 869342 708200 869398
rect 707800 869272 708200 869342
rect 69800 843658 70200 843728
rect 69800 843602 70074 843658
rect 70130 843602 70200 843658
rect 69800 843534 70200 843602
rect 69800 843478 70074 843534
rect 70130 843478 70200 843534
rect 69800 843410 70200 843478
rect 69800 843354 70074 843410
rect 70130 843354 70200 843410
rect 69800 843286 70200 843354
rect 69800 843230 70074 843286
rect 70130 843230 70200 843286
rect 69800 843162 70200 843230
rect 69800 843106 70074 843162
rect 70130 843106 70200 843162
rect 69800 843038 70200 843106
rect 69800 842982 70074 843038
rect 70130 842982 70200 843038
rect 69800 842914 70200 842982
rect 69800 842858 70074 842914
rect 70130 842858 70200 842914
rect 69800 842790 70200 842858
rect 69800 842734 70074 842790
rect 70130 842734 70200 842790
rect 69800 842666 70200 842734
rect 69800 842610 70074 842666
rect 70130 842610 70200 842666
rect 69800 842542 70200 842610
rect 69800 842486 70074 842542
rect 70130 842486 70200 842542
rect 69800 842418 70200 842486
rect 69800 842362 70074 842418
rect 70130 842362 70200 842418
rect 69800 842294 70200 842362
rect 69800 842238 70074 842294
rect 70130 842238 70200 842294
rect 69800 842170 70200 842238
rect 69800 842114 70074 842170
rect 70130 842114 70200 842170
rect 69800 842046 70200 842114
rect 69800 841990 70074 842046
rect 70130 841990 70200 842046
rect 69800 841922 70200 841990
rect 69800 841866 70074 841922
rect 70130 841866 70200 841922
rect 69800 841828 70200 841866
rect 69800 841184 70200 841248
rect 69800 841128 70074 841184
rect 70130 841128 70200 841184
rect 69800 841060 70200 841128
rect 69800 841004 70074 841060
rect 70130 841004 70200 841060
rect 69800 840936 70200 841004
rect 69800 840880 70074 840936
rect 70130 840880 70200 840936
rect 69800 840812 70200 840880
rect 69800 840756 70074 840812
rect 70130 840756 70200 840812
rect 69800 840688 70200 840756
rect 69800 840632 70074 840688
rect 70130 840632 70200 840688
rect 69800 840564 70200 840632
rect 69800 840508 70074 840564
rect 70130 840508 70200 840564
rect 69800 840440 70200 840508
rect 69800 840384 70074 840440
rect 70130 840384 70200 840440
rect 69800 840316 70200 840384
rect 69800 840260 70074 840316
rect 70130 840260 70200 840316
rect 69800 840192 70200 840260
rect 69800 840136 70074 840192
rect 70130 840136 70200 840192
rect 69800 840068 70200 840136
rect 69800 840012 70074 840068
rect 70130 840012 70200 840068
rect 69800 839944 70200 840012
rect 69800 839888 70074 839944
rect 70130 839888 70200 839944
rect 69800 839820 70200 839888
rect 69800 839764 70074 839820
rect 70130 839764 70200 839820
rect 69800 839696 70200 839764
rect 69800 839640 70074 839696
rect 70130 839640 70200 839696
rect 69800 839572 70200 839640
rect 69800 839516 70074 839572
rect 70130 839516 70200 839572
rect 69800 839448 70200 839516
rect 69800 839392 70074 839448
rect 70130 839392 70200 839448
rect 69800 839324 70200 839392
rect 69800 839268 70074 839324
rect 70130 839268 70200 839324
rect 69800 839198 70200 839268
rect 69800 838814 70200 838878
rect 69800 838758 70074 838814
rect 70130 838758 70200 838814
rect 69800 838690 70200 838758
rect 69800 838634 70074 838690
rect 70130 838634 70200 838690
rect 69800 838566 70200 838634
rect 69800 838510 70074 838566
rect 70130 838510 70200 838566
rect 69800 838442 70200 838510
rect 69800 838386 70074 838442
rect 70130 838386 70200 838442
rect 69800 838318 70200 838386
rect 69800 838262 70074 838318
rect 70130 838262 70200 838318
rect 69800 838194 70200 838262
rect 69800 838138 70074 838194
rect 70130 838138 70200 838194
rect 69800 838070 70200 838138
rect 69800 838014 70074 838070
rect 70130 838014 70200 838070
rect 69800 837946 70200 838014
rect 69800 837890 70074 837946
rect 70130 837890 70200 837946
rect 69800 837822 70200 837890
rect 69800 837766 70074 837822
rect 70130 837766 70200 837822
rect 69800 837698 70200 837766
rect 69800 837642 70074 837698
rect 70130 837642 70200 837698
rect 69800 837574 70200 837642
rect 69800 837518 70074 837574
rect 70130 837518 70200 837574
rect 69800 837450 70200 837518
rect 69800 837394 70074 837450
rect 70130 837394 70200 837450
rect 69800 837326 70200 837394
rect 69800 837270 70074 837326
rect 70130 837270 70200 837326
rect 69800 837202 70200 837270
rect 69800 837146 70074 837202
rect 70130 837146 70200 837202
rect 69800 837078 70200 837146
rect 69800 837022 70074 837078
rect 70130 837022 70200 837078
rect 69800 836954 70200 837022
rect 69800 836898 70074 836954
rect 70130 836898 70200 836954
rect 69800 836828 70200 836898
rect 69800 836108 70200 836172
rect 69800 836052 70074 836108
rect 70130 836052 70200 836108
rect 69800 835984 70200 836052
rect 69800 835928 70074 835984
rect 70130 835928 70200 835984
rect 69800 835860 70200 835928
rect 69800 835804 70074 835860
rect 70130 835804 70200 835860
rect 69800 835736 70200 835804
rect 69800 835680 70074 835736
rect 70130 835680 70200 835736
rect 69800 835612 70200 835680
rect 69800 835556 70074 835612
rect 70130 835556 70200 835612
rect 69800 835488 70200 835556
rect 69800 835432 70074 835488
rect 70130 835432 70200 835488
rect 69800 835364 70200 835432
rect 69800 835308 70074 835364
rect 70130 835308 70200 835364
rect 69800 835240 70200 835308
rect 69800 835184 70074 835240
rect 70130 835184 70200 835240
rect 69800 835116 70200 835184
rect 69800 835060 70074 835116
rect 70130 835060 70200 835116
rect 69800 834992 70200 835060
rect 69800 834936 70074 834992
rect 70130 834936 70200 834992
rect 69800 834868 70200 834936
rect 69800 834812 70074 834868
rect 70130 834812 70200 834868
rect 69800 834744 70200 834812
rect 69800 834688 70074 834744
rect 70130 834688 70200 834744
rect 69800 834620 70200 834688
rect 69800 834564 70074 834620
rect 70130 834564 70200 834620
rect 69800 834496 70200 834564
rect 69800 834440 70074 834496
rect 70130 834440 70200 834496
rect 69800 834372 70200 834440
rect 69800 834316 70074 834372
rect 70130 834316 70200 834372
rect 69800 834248 70200 834316
rect 69800 834192 70074 834248
rect 70130 834192 70200 834248
rect 69800 834122 70200 834192
rect 69800 833738 70200 833802
rect 69800 833682 70074 833738
rect 70130 833682 70200 833738
rect 69800 833614 70200 833682
rect 69800 833558 70074 833614
rect 70130 833558 70200 833614
rect 69800 833490 70200 833558
rect 69800 833434 70074 833490
rect 70130 833434 70200 833490
rect 69800 833366 70200 833434
rect 69800 833310 70074 833366
rect 70130 833310 70200 833366
rect 69800 833242 70200 833310
rect 69800 833186 70074 833242
rect 70130 833186 70200 833242
rect 69800 833118 70200 833186
rect 69800 833062 70074 833118
rect 70130 833062 70200 833118
rect 69800 832994 70200 833062
rect 69800 832938 70074 832994
rect 70130 832938 70200 832994
rect 69800 832870 70200 832938
rect 69800 832814 70074 832870
rect 70130 832814 70200 832870
rect 69800 832746 70200 832814
rect 69800 832690 70074 832746
rect 70130 832690 70200 832746
rect 69800 832622 70200 832690
rect 69800 832566 70074 832622
rect 70130 832566 70200 832622
rect 69800 832498 70200 832566
rect 69800 832442 70074 832498
rect 70130 832442 70200 832498
rect 69800 832374 70200 832442
rect 69800 832318 70074 832374
rect 70130 832318 70200 832374
rect 69800 832250 70200 832318
rect 69800 832194 70074 832250
rect 70130 832194 70200 832250
rect 69800 832126 70200 832194
rect 69800 832070 70074 832126
rect 70130 832070 70200 832126
rect 69800 832002 70200 832070
rect 69800 831946 70074 832002
rect 70130 831946 70200 832002
rect 69800 831878 70200 831946
rect 69800 831822 70074 831878
rect 70130 831822 70200 831878
rect 69800 831752 70200 831822
rect 69800 831134 70200 831172
rect 69800 831078 70074 831134
rect 70130 831078 70200 831134
rect 69800 831010 70200 831078
rect 69800 830954 70074 831010
rect 70130 830954 70200 831010
rect 69800 830886 70200 830954
rect 69800 830830 70074 830886
rect 70130 830830 70200 830886
rect 69800 830762 70200 830830
rect 69800 830706 70074 830762
rect 70130 830706 70200 830762
rect 69800 830638 70200 830706
rect 69800 830582 70074 830638
rect 70130 830582 70200 830638
rect 69800 830514 70200 830582
rect 69800 830458 70074 830514
rect 70130 830458 70200 830514
rect 69800 830390 70200 830458
rect 69800 830334 70074 830390
rect 70130 830334 70200 830390
rect 69800 830266 70200 830334
rect 69800 830210 70074 830266
rect 70130 830210 70200 830266
rect 69800 830142 70200 830210
rect 69800 830086 70074 830142
rect 70130 830086 70200 830142
rect 69800 830018 70200 830086
rect 69800 829962 70074 830018
rect 70130 829962 70200 830018
rect 69800 829894 70200 829962
rect 69800 829838 70074 829894
rect 70130 829838 70200 829894
rect 69800 829770 70200 829838
rect 69800 829714 70074 829770
rect 70130 829714 70200 829770
rect 69800 829646 70200 829714
rect 69800 829590 70074 829646
rect 70130 829590 70200 829646
rect 69800 829522 70200 829590
rect 69800 829466 70074 829522
rect 70130 829466 70200 829522
rect 69800 829398 70200 829466
rect 69800 829342 70074 829398
rect 70130 829342 70200 829398
rect 69800 829272 70200 829342
rect 69800 802658 70200 802728
rect 69800 802602 70074 802658
rect 70130 802602 70200 802658
rect 69800 802534 70200 802602
rect 69800 802478 70074 802534
rect 70130 802478 70200 802534
rect 69800 802410 70200 802478
rect 69800 802354 70074 802410
rect 70130 802354 70200 802410
rect 69800 802286 70200 802354
rect 69800 802230 70074 802286
rect 70130 802230 70200 802286
rect 69800 802162 70200 802230
rect 69800 802106 70074 802162
rect 70130 802106 70200 802162
rect 69800 802038 70200 802106
rect 69800 801982 70074 802038
rect 70130 801982 70200 802038
rect 69800 801914 70200 801982
rect 69800 801858 70074 801914
rect 70130 801858 70200 801914
rect 69800 801790 70200 801858
rect 69800 801734 70074 801790
rect 70130 801734 70200 801790
rect 69800 801666 70200 801734
rect 69800 801610 70074 801666
rect 70130 801610 70200 801666
rect 69800 801542 70200 801610
rect 69800 801486 70074 801542
rect 70130 801486 70200 801542
rect 69800 801418 70200 801486
rect 69800 801362 70074 801418
rect 70130 801362 70200 801418
rect 69800 801294 70200 801362
rect 69800 801238 70074 801294
rect 70130 801238 70200 801294
rect 69800 801170 70200 801238
rect 69800 801114 70074 801170
rect 70130 801114 70200 801170
rect 69800 801046 70200 801114
rect 69800 800990 70074 801046
rect 70130 800990 70200 801046
rect 69800 800922 70200 800990
rect 69800 800866 70074 800922
rect 70130 800866 70200 800922
rect 69800 800828 70200 800866
rect 69800 800184 70200 800248
rect 69800 800128 70074 800184
rect 70130 800128 70200 800184
rect 69800 800060 70200 800128
rect 69800 800004 70074 800060
rect 70130 800004 70200 800060
rect 69800 799936 70200 800004
rect 69800 799880 70074 799936
rect 70130 799880 70200 799936
rect 69800 799812 70200 799880
rect 69800 799756 70074 799812
rect 70130 799756 70200 799812
rect 69800 799688 70200 799756
rect 69800 799632 70074 799688
rect 70130 799632 70200 799688
rect 69800 799564 70200 799632
rect 69800 799508 70074 799564
rect 70130 799508 70200 799564
rect 69800 799440 70200 799508
rect 69800 799384 70074 799440
rect 70130 799384 70200 799440
rect 69800 799316 70200 799384
rect 69800 799260 70074 799316
rect 70130 799260 70200 799316
rect 69800 799192 70200 799260
rect 69800 799136 70074 799192
rect 70130 799136 70200 799192
rect 69800 799068 70200 799136
rect 69800 799012 70074 799068
rect 70130 799012 70200 799068
rect 69800 798944 70200 799012
rect 69800 798888 70074 798944
rect 70130 798888 70200 798944
rect 69800 798820 70200 798888
rect 69800 798764 70074 798820
rect 70130 798764 70200 798820
rect 69800 798696 70200 798764
rect 69800 798640 70074 798696
rect 70130 798640 70200 798696
rect 69800 798572 70200 798640
rect 69800 798516 70074 798572
rect 70130 798516 70200 798572
rect 69800 798448 70200 798516
rect 69800 798392 70074 798448
rect 70130 798392 70200 798448
rect 69800 798324 70200 798392
rect 69800 798268 70074 798324
rect 70130 798268 70200 798324
rect 69800 798198 70200 798268
rect 69800 797814 70200 797878
rect 69800 797758 70074 797814
rect 70130 797758 70200 797814
rect 69800 797690 70200 797758
rect 69800 797634 70074 797690
rect 70130 797634 70200 797690
rect 69800 797566 70200 797634
rect 69800 797510 70074 797566
rect 70130 797510 70200 797566
rect 69800 797442 70200 797510
rect 69800 797386 70074 797442
rect 70130 797386 70200 797442
rect 69800 797318 70200 797386
rect 69800 797262 70074 797318
rect 70130 797262 70200 797318
rect 69800 797194 70200 797262
rect 69800 797138 70074 797194
rect 70130 797138 70200 797194
rect 69800 797070 70200 797138
rect 69800 797014 70074 797070
rect 70130 797014 70200 797070
rect 69800 796946 70200 797014
rect 69800 796890 70074 796946
rect 70130 796890 70200 796946
rect 69800 796822 70200 796890
rect 69800 796766 70074 796822
rect 70130 796766 70200 796822
rect 69800 796698 70200 796766
rect 69800 796642 70074 796698
rect 70130 796642 70200 796698
rect 69800 796574 70200 796642
rect 69800 796518 70074 796574
rect 70130 796518 70200 796574
rect 69800 796450 70200 796518
rect 69800 796394 70074 796450
rect 70130 796394 70200 796450
rect 69800 796326 70200 796394
rect 69800 796270 70074 796326
rect 70130 796270 70200 796326
rect 69800 796202 70200 796270
rect 69800 796146 70074 796202
rect 70130 796146 70200 796202
rect 69800 796078 70200 796146
rect 69800 796022 70074 796078
rect 70130 796022 70200 796078
rect 69800 795954 70200 796022
rect 69800 795898 70074 795954
rect 70130 795898 70200 795954
rect 69800 795828 70200 795898
rect 707800 797658 708200 797728
rect 707800 797602 707870 797658
rect 707926 797602 708200 797658
rect 707800 797534 708200 797602
rect 707800 797478 707870 797534
rect 707926 797478 708200 797534
rect 707800 797410 708200 797478
rect 707800 797354 707870 797410
rect 707926 797354 708200 797410
rect 707800 797286 708200 797354
rect 707800 797230 707870 797286
rect 707926 797230 708200 797286
rect 707800 797162 708200 797230
rect 707800 797106 707870 797162
rect 707926 797106 708200 797162
rect 707800 797038 708200 797106
rect 707800 796982 707870 797038
rect 707926 796982 708200 797038
rect 707800 796914 708200 796982
rect 707800 796858 707870 796914
rect 707926 796858 708200 796914
rect 707800 796790 708200 796858
rect 707800 796734 707870 796790
rect 707926 796734 708200 796790
rect 707800 796666 708200 796734
rect 707800 796610 707870 796666
rect 707926 796610 708200 796666
rect 707800 796542 708200 796610
rect 707800 796486 707870 796542
rect 707926 796486 708200 796542
rect 707800 796418 708200 796486
rect 707800 796362 707870 796418
rect 707926 796362 708200 796418
rect 707800 796294 708200 796362
rect 707800 796238 707870 796294
rect 707926 796238 708200 796294
rect 707800 796170 708200 796238
rect 707800 796114 707870 796170
rect 707926 796114 708200 796170
rect 707800 796046 708200 796114
rect 707800 795990 707870 796046
rect 707926 795990 708200 796046
rect 707800 795922 708200 795990
rect 707800 795866 707870 795922
rect 707926 795866 708200 795922
rect 707800 795828 708200 795866
rect 707800 795178 708200 795248
rect 69800 795108 70200 795172
rect 69800 795052 70074 795108
rect 70130 795052 70200 795108
rect 69800 794984 70200 795052
rect 69800 794928 70074 794984
rect 70130 794928 70200 794984
rect 69800 794860 70200 794928
rect 69800 794804 70074 794860
rect 70130 794804 70200 794860
rect 69800 794736 70200 794804
rect 69800 794680 70074 794736
rect 70130 794680 70200 794736
rect 69800 794612 70200 794680
rect 69800 794556 70074 794612
rect 70130 794556 70200 794612
rect 69800 794488 70200 794556
rect 69800 794432 70074 794488
rect 70130 794432 70200 794488
rect 69800 794364 70200 794432
rect 69800 794308 70074 794364
rect 70130 794308 70200 794364
rect 69800 794240 70200 794308
rect 69800 794184 70074 794240
rect 70130 794184 70200 794240
rect 69800 794116 70200 794184
rect 69800 794060 70074 794116
rect 70130 794060 70200 794116
rect 69800 793992 70200 794060
rect 69800 793936 70074 793992
rect 70130 793936 70200 793992
rect 69800 793868 70200 793936
rect 69800 793812 70074 793868
rect 70130 793812 70200 793868
rect 69800 793744 70200 793812
rect 69800 793688 70074 793744
rect 70130 793688 70200 793744
rect 69800 793620 70200 793688
rect 69800 793564 70074 793620
rect 70130 793564 70200 793620
rect 69800 793496 70200 793564
rect 69800 793440 70074 793496
rect 70130 793440 70200 793496
rect 69800 793372 70200 793440
rect 69800 793316 70074 793372
rect 70130 793316 70200 793372
rect 69800 793248 70200 793316
rect 69800 793192 70074 793248
rect 70130 793192 70200 793248
rect 707800 795122 707870 795178
rect 707926 795122 708200 795178
rect 707800 795054 708200 795122
rect 707800 794998 707870 795054
rect 707926 794998 708200 795054
rect 707800 794930 708200 794998
rect 707800 794874 707870 794930
rect 707926 794874 708200 794930
rect 707800 794806 708200 794874
rect 707800 794750 707870 794806
rect 707926 794750 708200 794806
rect 707800 794682 708200 794750
rect 707800 794626 707870 794682
rect 707926 794626 708200 794682
rect 707800 794558 708200 794626
rect 707800 794502 707870 794558
rect 707926 794502 708200 794558
rect 707800 794434 708200 794502
rect 707800 794378 707870 794434
rect 707926 794378 708200 794434
rect 707800 794310 708200 794378
rect 707800 794254 707870 794310
rect 707926 794254 708200 794310
rect 707800 794186 708200 794254
rect 707800 794130 707870 794186
rect 707926 794130 708200 794186
rect 707800 794062 708200 794130
rect 707800 794006 707870 794062
rect 707926 794006 708200 794062
rect 707800 793938 708200 794006
rect 707800 793882 707870 793938
rect 707926 793882 708200 793938
rect 707800 793814 708200 793882
rect 707800 793758 707870 793814
rect 707926 793758 708200 793814
rect 707800 793690 708200 793758
rect 707800 793634 707870 793690
rect 707926 793634 708200 793690
rect 707800 793566 708200 793634
rect 707800 793510 707870 793566
rect 707926 793510 708200 793566
rect 707800 793442 708200 793510
rect 707800 793386 707870 793442
rect 707926 793386 708200 793442
rect 707800 793318 708200 793386
rect 707800 793262 707870 793318
rect 707926 793262 708200 793318
rect 707800 793198 708200 793262
rect 69800 793122 70200 793192
rect 707800 792808 708200 792878
rect 69800 792738 70200 792802
rect 69800 792682 70074 792738
rect 70130 792682 70200 792738
rect 69800 792614 70200 792682
rect 69800 792558 70074 792614
rect 70130 792558 70200 792614
rect 69800 792490 70200 792558
rect 69800 792434 70074 792490
rect 70130 792434 70200 792490
rect 69800 792366 70200 792434
rect 69800 792310 70074 792366
rect 70130 792310 70200 792366
rect 69800 792242 70200 792310
rect 69800 792186 70074 792242
rect 70130 792186 70200 792242
rect 69800 792118 70200 792186
rect 69800 792062 70074 792118
rect 70130 792062 70200 792118
rect 69800 791994 70200 792062
rect 69800 791938 70074 791994
rect 70130 791938 70200 791994
rect 69800 791870 70200 791938
rect 69800 791814 70074 791870
rect 70130 791814 70200 791870
rect 69800 791746 70200 791814
rect 69800 791690 70074 791746
rect 70130 791690 70200 791746
rect 69800 791622 70200 791690
rect 69800 791566 70074 791622
rect 70130 791566 70200 791622
rect 69800 791498 70200 791566
rect 69800 791442 70074 791498
rect 70130 791442 70200 791498
rect 69800 791374 70200 791442
rect 69800 791318 70074 791374
rect 70130 791318 70200 791374
rect 69800 791250 70200 791318
rect 69800 791194 70074 791250
rect 70130 791194 70200 791250
rect 69800 791126 70200 791194
rect 69800 791070 70074 791126
rect 70130 791070 70200 791126
rect 69800 791002 70200 791070
rect 69800 790946 70074 791002
rect 70130 790946 70200 791002
rect 69800 790878 70200 790946
rect 69800 790822 70074 790878
rect 70130 790822 70200 790878
rect 707800 792752 707870 792808
rect 707926 792752 708200 792808
rect 707800 792684 708200 792752
rect 707800 792628 707870 792684
rect 707926 792628 708200 792684
rect 707800 792560 708200 792628
rect 707800 792504 707870 792560
rect 707926 792504 708200 792560
rect 707800 792436 708200 792504
rect 707800 792380 707870 792436
rect 707926 792380 708200 792436
rect 707800 792312 708200 792380
rect 707800 792256 707870 792312
rect 707926 792256 708200 792312
rect 707800 792188 708200 792256
rect 707800 792132 707870 792188
rect 707926 792132 708200 792188
rect 707800 792064 708200 792132
rect 707800 792008 707870 792064
rect 707926 792008 708200 792064
rect 707800 791940 708200 792008
rect 707800 791884 707870 791940
rect 707926 791884 708200 791940
rect 707800 791816 708200 791884
rect 707800 791760 707870 791816
rect 707926 791760 708200 791816
rect 707800 791692 708200 791760
rect 707800 791636 707870 791692
rect 707926 791636 708200 791692
rect 707800 791568 708200 791636
rect 707800 791512 707870 791568
rect 707926 791512 708200 791568
rect 707800 791444 708200 791512
rect 707800 791388 707870 791444
rect 707926 791388 708200 791444
rect 707800 791320 708200 791388
rect 707800 791264 707870 791320
rect 707926 791264 708200 791320
rect 707800 791196 708200 791264
rect 707800 791140 707870 791196
rect 707926 791140 708200 791196
rect 707800 791072 708200 791140
rect 707800 791016 707870 791072
rect 707926 791016 708200 791072
rect 707800 790948 708200 791016
rect 707800 790892 707870 790948
rect 707926 790892 708200 790948
rect 707800 790828 708200 790892
rect 69800 790752 70200 790822
rect 69800 790134 70200 790172
rect 69800 790078 70074 790134
rect 70130 790078 70200 790134
rect 69800 790010 70200 790078
rect 69800 789954 70074 790010
rect 70130 789954 70200 790010
rect 69800 789886 70200 789954
rect 69800 789830 70074 789886
rect 70130 789830 70200 789886
rect 69800 789762 70200 789830
rect 69800 789706 70074 789762
rect 70130 789706 70200 789762
rect 69800 789638 70200 789706
rect 69800 789582 70074 789638
rect 70130 789582 70200 789638
rect 69800 789514 70200 789582
rect 69800 789458 70074 789514
rect 70130 789458 70200 789514
rect 69800 789390 70200 789458
rect 69800 789334 70074 789390
rect 70130 789334 70200 789390
rect 69800 789266 70200 789334
rect 69800 789210 70074 789266
rect 70130 789210 70200 789266
rect 69800 789142 70200 789210
rect 69800 789086 70074 789142
rect 70130 789086 70200 789142
rect 69800 789018 70200 789086
rect 69800 788962 70074 789018
rect 70130 788962 70200 789018
rect 69800 788894 70200 788962
rect 69800 788838 70074 788894
rect 70130 788838 70200 788894
rect 69800 788770 70200 788838
rect 69800 788714 70074 788770
rect 70130 788714 70200 788770
rect 69800 788646 70200 788714
rect 69800 788590 70074 788646
rect 70130 788590 70200 788646
rect 69800 788522 70200 788590
rect 69800 788466 70074 788522
rect 70130 788466 70200 788522
rect 69800 788398 70200 788466
rect 69800 788342 70074 788398
rect 70130 788342 70200 788398
rect 69800 788272 70200 788342
rect 707800 790102 708200 790172
rect 707800 790046 707870 790102
rect 707926 790046 708200 790102
rect 707800 789978 708200 790046
rect 707800 789922 707870 789978
rect 707926 789922 708200 789978
rect 707800 789854 708200 789922
rect 707800 789798 707870 789854
rect 707926 789798 708200 789854
rect 707800 789730 708200 789798
rect 707800 789674 707870 789730
rect 707926 789674 708200 789730
rect 707800 789606 708200 789674
rect 707800 789550 707870 789606
rect 707926 789550 708200 789606
rect 707800 789482 708200 789550
rect 707800 789426 707870 789482
rect 707926 789426 708200 789482
rect 707800 789358 708200 789426
rect 707800 789302 707870 789358
rect 707926 789302 708200 789358
rect 707800 789234 708200 789302
rect 707800 789178 707870 789234
rect 707926 789178 708200 789234
rect 707800 789110 708200 789178
rect 707800 789054 707870 789110
rect 707926 789054 708200 789110
rect 707800 788986 708200 789054
rect 707800 788930 707870 788986
rect 707926 788930 708200 788986
rect 707800 788862 708200 788930
rect 707800 788806 707870 788862
rect 707926 788806 708200 788862
rect 707800 788738 708200 788806
rect 707800 788682 707870 788738
rect 707926 788682 708200 788738
rect 707800 788614 708200 788682
rect 707800 788558 707870 788614
rect 707926 788558 708200 788614
rect 707800 788490 708200 788558
rect 707800 788434 707870 788490
rect 707926 788434 708200 788490
rect 707800 788366 708200 788434
rect 707800 788310 707870 788366
rect 707926 788310 708200 788366
rect 707800 788242 708200 788310
rect 707800 788186 707870 788242
rect 707926 788186 708200 788242
rect 707800 788122 708200 788186
rect 707800 787732 708200 787802
rect 707800 787676 707870 787732
rect 707926 787676 708200 787732
rect 707800 787608 708200 787676
rect 707800 787552 707870 787608
rect 707926 787552 708200 787608
rect 707800 787484 708200 787552
rect 707800 787428 707870 787484
rect 707926 787428 708200 787484
rect 707800 787360 708200 787428
rect 707800 787304 707870 787360
rect 707926 787304 708200 787360
rect 707800 787236 708200 787304
rect 707800 787180 707870 787236
rect 707926 787180 708200 787236
rect 707800 787112 708200 787180
rect 707800 787056 707870 787112
rect 707926 787056 708200 787112
rect 707800 786988 708200 787056
rect 707800 786932 707870 786988
rect 707926 786932 708200 786988
rect 707800 786864 708200 786932
rect 707800 786808 707870 786864
rect 707926 786808 708200 786864
rect 707800 786740 708200 786808
rect 707800 786684 707870 786740
rect 707926 786684 708200 786740
rect 707800 786616 708200 786684
rect 707800 786560 707870 786616
rect 707926 786560 708200 786616
rect 707800 786492 708200 786560
rect 707800 786436 707870 786492
rect 707926 786436 708200 786492
rect 707800 786368 708200 786436
rect 707800 786312 707870 786368
rect 707926 786312 708200 786368
rect 707800 786244 708200 786312
rect 707800 786188 707870 786244
rect 707926 786188 708200 786244
rect 707800 786120 708200 786188
rect 707800 786064 707870 786120
rect 707926 786064 708200 786120
rect 707800 785996 708200 786064
rect 707800 785940 707870 785996
rect 707926 785940 708200 785996
rect 707800 785872 708200 785940
rect 707800 785816 707870 785872
rect 707926 785816 708200 785872
rect 707800 785752 708200 785816
rect 707800 785134 708200 785172
rect 707800 785078 707870 785134
rect 707926 785078 708200 785134
rect 707800 785010 708200 785078
rect 707800 784954 707870 785010
rect 707926 784954 708200 785010
rect 707800 784886 708200 784954
rect 707800 784830 707870 784886
rect 707926 784830 708200 784886
rect 707800 784762 708200 784830
rect 707800 784706 707870 784762
rect 707926 784706 708200 784762
rect 707800 784638 708200 784706
rect 707800 784582 707870 784638
rect 707926 784582 708200 784638
rect 707800 784514 708200 784582
rect 707800 784458 707870 784514
rect 707926 784458 708200 784514
rect 707800 784390 708200 784458
rect 707800 784334 707870 784390
rect 707926 784334 708200 784390
rect 707800 784266 708200 784334
rect 707800 784210 707870 784266
rect 707926 784210 708200 784266
rect 707800 784142 708200 784210
rect 707800 784086 707870 784142
rect 707926 784086 708200 784142
rect 707800 784018 708200 784086
rect 707800 783962 707870 784018
rect 707926 783962 708200 784018
rect 707800 783894 708200 783962
rect 707800 783838 707870 783894
rect 707926 783838 708200 783894
rect 707800 783770 708200 783838
rect 707800 783714 707870 783770
rect 707926 783714 708200 783770
rect 707800 783646 708200 783714
rect 707800 783590 707870 783646
rect 707926 783590 708200 783646
rect 707800 783522 708200 783590
rect 707800 783466 707870 783522
rect 707926 783466 708200 783522
rect 707800 783398 708200 783466
rect 707800 783342 707870 783398
rect 707926 783342 708200 783398
rect 707800 783272 708200 783342
rect 707800 496658 708200 496728
rect 707800 496602 707870 496658
rect 707926 496602 708200 496658
rect 707800 496534 708200 496602
rect 707800 496478 707870 496534
rect 707926 496478 708200 496534
rect 707800 496410 708200 496478
rect 707800 496354 707870 496410
rect 707926 496354 708200 496410
rect 707800 496286 708200 496354
rect 707800 496230 707870 496286
rect 707926 496230 708200 496286
rect 707800 496162 708200 496230
rect 707800 496106 707870 496162
rect 707926 496106 708200 496162
rect 707800 496038 708200 496106
rect 707800 495982 707870 496038
rect 707926 495982 708200 496038
rect 707800 495914 708200 495982
rect 707800 495858 707870 495914
rect 707926 495858 708200 495914
rect 707800 495790 708200 495858
rect 707800 495734 707870 495790
rect 707926 495734 708200 495790
rect 707800 495666 708200 495734
rect 707800 495610 707870 495666
rect 707926 495610 708200 495666
rect 707800 495542 708200 495610
rect 707800 495486 707870 495542
rect 707926 495486 708200 495542
rect 707800 495418 708200 495486
rect 707800 495362 707870 495418
rect 707926 495362 708200 495418
rect 707800 495294 708200 495362
rect 707800 495238 707870 495294
rect 707926 495238 708200 495294
rect 707800 495170 708200 495238
rect 707800 495114 707870 495170
rect 707926 495114 708200 495170
rect 707800 495046 708200 495114
rect 707800 494990 707870 495046
rect 707926 494990 708200 495046
rect 707800 494922 708200 494990
rect 707800 494866 707870 494922
rect 707926 494866 708200 494922
rect 707800 494828 708200 494866
rect 707800 494178 708200 494248
rect 707800 494122 707870 494178
rect 707926 494122 708200 494178
rect 707800 494054 708200 494122
rect 707800 493998 707870 494054
rect 707926 493998 708200 494054
rect 707800 493930 708200 493998
rect 707800 493874 707870 493930
rect 707926 493874 708200 493930
rect 707800 493806 708200 493874
rect 707800 493750 707870 493806
rect 707926 493750 708200 493806
rect 707800 493682 708200 493750
rect 707800 493626 707870 493682
rect 707926 493626 708200 493682
rect 707800 493558 708200 493626
rect 707800 493502 707870 493558
rect 707926 493502 708200 493558
rect 707800 493434 708200 493502
rect 707800 493378 707870 493434
rect 707926 493378 708200 493434
rect 707800 493310 708200 493378
rect 707800 493254 707870 493310
rect 707926 493254 708200 493310
rect 707800 493186 708200 493254
rect 707800 493130 707870 493186
rect 707926 493130 708200 493186
rect 707800 493062 708200 493130
rect 707800 493006 707870 493062
rect 707926 493006 708200 493062
rect 707800 492938 708200 493006
rect 707800 492882 707870 492938
rect 707926 492882 708200 492938
rect 707800 492814 708200 492882
rect 707800 492758 707870 492814
rect 707926 492758 708200 492814
rect 707800 492690 708200 492758
rect 707800 492634 707870 492690
rect 707926 492634 708200 492690
rect 707800 492566 708200 492634
rect 707800 492510 707870 492566
rect 707926 492510 708200 492566
rect 707800 492442 708200 492510
rect 707800 492386 707870 492442
rect 707926 492386 708200 492442
rect 707800 492318 708200 492386
rect 707800 492262 707870 492318
rect 707926 492262 708200 492318
rect 707800 492198 708200 492262
rect 707800 491808 708200 491878
rect 707800 491752 707870 491808
rect 707926 491752 708200 491808
rect 707800 491684 708200 491752
rect 707800 491628 707870 491684
rect 707926 491628 708200 491684
rect 707800 491560 708200 491628
rect 707800 491504 707870 491560
rect 707926 491504 708200 491560
rect 707800 491436 708200 491504
rect 707800 491380 707870 491436
rect 707926 491380 708200 491436
rect 707800 491312 708200 491380
rect 707800 491256 707870 491312
rect 707926 491256 708200 491312
rect 707800 491188 708200 491256
rect 707800 491132 707870 491188
rect 707926 491132 708200 491188
rect 707800 491064 708200 491132
rect 707800 491008 707870 491064
rect 707926 491008 708200 491064
rect 707800 490940 708200 491008
rect 707800 490884 707870 490940
rect 707926 490884 708200 490940
rect 707800 490816 708200 490884
rect 707800 490760 707870 490816
rect 707926 490760 708200 490816
rect 707800 490692 708200 490760
rect 707800 490636 707870 490692
rect 707926 490636 708200 490692
rect 707800 490568 708200 490636
rect 707800 490512 707870 490568
rect 707926 490512 708200 490568
rect 707800 490444 708200 490512
rect 707800 490388 707870 490444
rect 707926 490388 708200 490444
rect 707800 490320 708200 490388
rect 707800 490264 707870 490320
rect 707926 490264 708200 490320
rect 707800 490196 708200 490264
rect 707800 490140 707870 490196
rect 707926 490140 708200 490196
rect 707800 490072 708200 490140
rect 707800 490016 707870 490072
rect 707926 490016 708200 490072
rect 707800 489948 708200 490016
rect 707800 489892 707870 489948
rect 707926 489892 708200 489948
rect 707800 489828 708200 489892
rect 707800 489102 708200 489172
rect 707800 489046 707870 489102
rect 707926 489046 708200 489102
rect 707800 488978 708200 489046
rect 707800 488922 707870 488978
rect 707926 488922 708200 488978
rect 707800 488854 708200 488922
rect 707800 488798 707870 488854
rect 707926 488798 708200 488854
rect 707800 488730 708200 488798
rect 707800 488674 707870 488730
rect 707926 488674 708200 488730
rect 707800 488606 708200 488674
rect 707800 488550 707870 488606
rect 707926 488550 708200 488606
rect 707800 488482 708200 488550
rect 707800 488426 707870 488482
rect 707926 488426 708200 488482
rect 707800 488358 708200 488426
rect 707800 488302 707870 488358
rect 707926 488302 708200 488358
rect 707800 488234 708200 488302
rect 707800 488178 707870 488234
rect 707926 488178 708200 488234
rect 707800 488110 708200 488178
rect 707800 488054 707870 488110
rect 707926 488054 708200 488110
rect 707800 487986 708200 488054
rect 707800 487930 707870 487986
rect 707926 487930 708200 487986
rect 707800 487862 708200 487930
rect 707800 487806 707870 487862
rect 707926 487806 708200 487862
rect 707800 487738 708200 487806
rect 707800 487682 707870 487738
rect 707926 487682 708200 487738
rect 707800 487614 708200 487682
rect 707800 487558 707870 487614
rect 707926 487558 708200 487614
rect 707800 487490 708200 487558
rect 707800 487434 707870 487490
rect 707926 487434 708200 487490
rect 707800 487366 708200 487434
rect 707800 487310 707870 487366
rect 707926 487310 708200 487366
rect 707800 487242 708200 487310
rect 707800 487186 707870 487242
rect 707926 487186 708200 487242
rect 707800 487122 708200 487186
rect 707800 486732 708200 486802
rect 707800 486676 707870 486732
rect 707926 486676 708200 486732
rect 707800 486608 708200 486676
rect 707800 486552 707870 486608
rect 707926 486552 708200 486608
rect 707800 486484 708200 486552
rect 707800 486428 707870 486484
rect 707926 486428 708200 486484
rect 707800 486360 708200 486428
rect 707800 486304 707870 486360
rect 707926 486304 708200 486360
rect 707800 486236 708200 486304
rect 707800 486180 707870 486236
rect 707926 486180 708200 486236
rect 707800 486112 708200 486180
rect 707800 486056 707870 486112
rect 707926 486056 708200 486112
rect 707800 485988 708200 486056
rect 707800 485932 707870 485988
rect 707926 485932 708200 485988
rect 707800 485864 708200 485932
rect 707800 485808 707870 485864
rect 707926 485808 708200 485864
rect 707800 485740 708200 485808
rect 707800 485684 707870 485740
rect 707926 485684 708200 485740
rect 707800 485616 708200 485684
rect 707800 485560 707870 485616
rect 707926 485560 708200 485616
rect 707800 485492 708200 485560
rect 707800 485436 707870 485492
rect 707926 485436 708200 485492
rect 707800 485368 708200 485436
rect 707800 485312 707870 485368
rect 707926 485312 708200 485368
rect 707800 485244 708200 485312
rect 707800 485188 707870 485244
rect 707926 485188 708200 485244
rect 707800 485120 708200 485188
rect 707800 485064 707870 485120
rect 707926 485064 708200 485120
rect 707800 484996 708200 485064
rect 707800 484940 707870 484996
rect 707926 484940 708200 484996
rect 707800 484872 708200 484940
rect 707800 484816 707870 484872
rect 707926 484816 708200 484872
rect 707800 484752 708200 484816
rect 707800 484134 708200 484172
rect 707800 484078 707870 484134
rect 707926 484078 708200 484134
rect 707800 484010 708200 484078
rect 707800 483954 707870 484010
rect 707926 483954 708200 484010
rect 707800 483886 708200 483954
rect 707800 483830 707870 483886
rect 707926 483830 708200 483886
rect 707800 483762 708200 483830
rect 707800 483706 707870 483762
rect 707926 483706 708200 483762
rect 707800 483638 708200 483706
rect 707800 483582 707870 483638
rect 707926 483582 708200 483638
rect 707800 483514 708200 483582
rect 707800 483458 707870 483514
rect 707926 483458 708200 483514
rect 707800 483390 708200 483458
rect 707800 483334 707870 483390
rect 707926 483334 708200 483390
rect 707800 483266 708200 483334
rect 707800 483210 707870 483266
rect 707926 483210 708200 483266
rect 707800 483142 708200 483210
rect 707800 483086 707870 483142
rect 707926 483086 708200 483142
rect 707800 483018 708200 483086
rect 707800 482962 707870 483018
rect 707926 482962 708200 483018
rect 707800 482894 708200 482962
rect 707800 482838 707870 482894
rect 707926 482838 708200 482894
rect 707800 482770 708200 482838
rect 707800 482714 707870 482770
rect 707926 482714 708200 482770
rect 707800 482646 708200 482714
rect 707800 482590 707870 482646
rect 707926 482590 708200 482646
rect 707800 482522 708200 482590
rect 707800 482466 707870 482522
rect 707926 482466 708200 482522
rect 707800 482398 708200 482466
rect 707800 482342 707870 482398
rect 707926 482342 708200 482398
rect 707800 482272 708200 482342
rect 69800 474658 70200 474728
rect 69800 474602 70074 474658
rect 70130 474602 70200 474658
rect 69800 474534 70200 474602
rect 69800 474478 70074 474534
rect 70130 474478 70200 474534
rect 69800 474410 70200 474478
rect 69800 474354 70074 474410
rect 70130 474354 70200 474410
rect 69800 474286 70200 474354
rect 69800 474230 70074 474286
rect 70130 474230 70200 474286
rect 69800 474162 70200 474230
rect 69800 474106 70074 474162
rect 70130 474106 70200 474162
rect 69800 474038 70200 474106
rect 69800 473982 70074 474038
rect 70130 473982 70200 474038
rect 69800 473914 70200 473982
rect 69800 473858 70074 473914
rect 70130 473858 70200 473914
rect 69800 473790 70200 473858
rect 69800 473734 70074 473790
rect 70130 473734 70200 473790
rect 69800 473666 70200 473734
rect 69800 473610 70074 473666
rect 70130 473610 70200 473666
rect 69800 473542 70200 473610
rect 69800 473486 70074 473542
rect 70130 473486 70200 473542
rect 69800 473418 70200 473486
rect 69800 473362 70074 473418
rect 70130 473362 70200 473418
rect 69800 473294 70200 473362
rect 69800 473238 70074 473294
rect 70130 473238 70200 473294
rect 69800 473170 70200 473238
rect 69800 473114 70074 473170
rect 70130 473114 70200 473170
rect 69800 473046 70200 473114
rect 69800 472990 70074 473046
rect 70130 472990 70200 473046
rect 69800 472922 70200 472990
rect 69800 472866 70074 472922
rect 70130 472866 70200 472922
rect 69800 472828 70200 472866
rect 69800 472184 70200 472248
rect 69800 472128 70074 472184
rect 70130 472128 70200 472184
rect 69800 472060 70200 472128
rect 69800 472004 70074 472060
rect 70130 472004 70200 472060
rect 69800 471936 70200 472004
rect 69800 471880 70074 471936
rect 70130 471880 70200 471936
rect 69800 471812 70200 471880
rect 69800 471756 70074 471812
rect 70130 471756 70200 471812
rect 69800 471688 70200 471756
rect 69800 471632 70074 471688
rect 70130 471632 70200 471688
rect 69800 471564 70200 471632
rect 69800 471508 70074 471564
rect 70130 471508 70200 471564
rect 69800 471440 70200 471508
rect 69800 471384 70074 471440
rect 70130 471384 70200 471440
rect 69800 471316 70200 471384
rect 69800 471260 70074 471316
rect 70130 471260 70200 471316
rect 69800 471192 70200 471260
rect 69800 471136 70074 471192
rect 70130 471136 70200 471192
rect 69800 471068 70200 471136
rect 69800 471012 70074 471068
rect 70130 471012 70200 471068
rect 69800 470944 70200 471012
rect 69800 470888 70074 470944
rect 70130 470888 70200 470944
rect 69800 470820 70200 470888
rect 69800 470764 70074 470820
rect 70130 470764 70200 470820
rect 69800 470696 70200 470764
rect 69800 470640 70074 470696
rect 70130 470640 70200 470696
rect 69800 470572 70200 470640
rect 69800 470516 70074 470572
rect 70130 470516 70200 470572
rect 69800 470448 70200 470516
rect 69800 470392 70074 470448
rect 70130 470392 70200 470448
rect 69800 470324 70200 470392
rect 69800 470268 70074 470324
rect 70130 470268 70200 470324
rect 69800 470198 70200 470268
rect 69800 469814 70200 469878
rect 69800 469758 70074 469814
rect 70130 469758 70200 469814
rect 69800 469690 70200 469758
rect 69800 469634 70074 469690
rect 70130 469634 70200 469690
rect 69800 469566 70200 469634
rect 69800 469510 70074 469566
rect 70130 469510 70200 469566
rect 69800 469442 70200 469510
rect 69800 469386 70074 469442
rect 70130 469386 70200 469442
rect 69800 469318 70200 469386
rect 69800 469262 70074 469318
rect 70130 469262 70200 469318
rect 69800 469194 70200 469262
rect 69800 469138 70074 469194
rect 70130 469138 70200 469194
rect 69800 469070 70200 469138
rect 69800 469014 70074 469070
rect 70130 469014 70200 469070
rect 69800 468946 70200 469014
rect 69800 468890 70074 468946
rect 70130 468890 70200 468946
rect 69800 468822 70200 468890
rect 69800 468766 70074 468822
rect 70130 468766 70200 468822
rect 69800 468698 70200 468766
rect 69800 468642 70074 468698
rect 70130 468642 70200 468698
rect 69800 468574 70200 468642
rect 69800 468518 70074 468574
rect 70130 468518 70200 468574
rect 69800 468450 70200 468518
rect 69800 468394 70074 468450
rect 70130 468394 70200 468450
rect 69800 468326 70200 468394
rect 69800 468270 70074 468326
rect 70130 468270 70200 468326
rect 69800 468202 70200 468270
rect 69800 468146 70074 468202
rect 70130 468146 70200 468202
rect 69800 468078 70200 468146
rect 69800 468022 70074 468078
rect 70130 468022 70200 468078
rect 69800 467954 70200 468022
rect 69800 467898 70074 467954
rect 70130 467898 70200 467954
rect 69800 467828 70200 467898
rect 69800 467108 70200 467172
rect 69800 467052 70074 467108
rect 70130 467052 70200 467108
rect 69800 466984 70200 467052
rect 69800 466928 70074 466984
rect 70130 466928 70200 466984
rect 69800 466860 70200 466928
rect 69800 466804 70074 466860
rect 70130 466804 70200 466860
rect 69800 466736 70200 466804
rect 69800 466680 70074 466736
rect 70130 466680 70200 466736
rect 69800 466612 70200 466680
rect 69800 466556 70074 466612
rect 70130 466556 70200 466612
rect 69800 466488 70200 466556
rect 69800 466432 70074 466488
rect 70130 466432 70200 466488
rect 69800 466364 70200 466432
rect 69800 466308 70074 466364
rect 70130 466308 70200 466364
rect 69800 466240 70200 466308
rect 69800 466184 70074 466240
rect 70130 466184 70200 466240
rect 69800 466116 70200 466184
rect 69800 466060 70074 466116
rect 70130 466060 70200 466116
rect 69800 465992 70200 466060
rect 69800 465936 70074 465992
rect 70130 465936 70200 465992
rect 69800 465868 70200 465936
rect 69800 465812 70074 465868
rect 70130 465812 70200 465868
rect 69800 465744 70200 465812
rect 69800 465688 70074 465744
rect 70130 465688 70200 465744
rect 69800 465620 70200 465688
rect 69800 465564 70074 465620
rect 70130 465564 70200 465620
rect 69800 465496 70200 465564
rect 69800 465440 70074 465496
rect 70130 465440 70200 465496
rect 69800 465372 70200 465440
rect 69800 465316 70074 465372
rect 70130 465316 70200 465372
rect 69800 465248 70200 465316
rect 69800 465192 70074 465248
rect 70130 465192 70200 465248
rect 69800 465122 70200 465192
rect 69800 464738 70200 464802
rect 69800 464682 70074 464738
rect 70130 464682 70200 464738
rect 69800 464614 70200 464682
rect 69800 464558 70074 464614
rect 70130 464558 70200 464614
rect 69800 464490 70200 464558
rect 69800 464434 70074 464490
rect 70130 464434 70200 464490
rect 69800 464366 70200 464434
rect 69800 464310 70074 464366
rect 70130 464310 70200 464366
rect 69800 464242 70200 464310
rect 69800 464186 70074 464242
rect 70130 464186 70200 464242
rect 69800 464118 70200 464186
rect 69800 464062 70074 464118
rect 70130 464062 70200 464118
rect 69800 463994 70200 464062
rect 69800 463938 70074 463994
rect 70130 463938 70200 463994
rect 69800 463870 70200 463938
rect 69800 463814 70074 463870
rect 70130 463814 70200 463870
rect 69800 463746 70200 463814
rect 69800 463690 70074 463746
rect 70130 463690 70200 463746
rect 69800 463622 70200 463690
rect 69800 463566 70074 463622
rect 70130 463566 70200 463622
rect 69800 463498 70200 463566
rect 69800 463442 70074 463498
rect 70130 463442 70200 463498
rect 69800 463374 70200 463442
rect 69800 463318 70074 463374
rect 70130 463318 70200 463374
rect 69800 463250 70200 463318
rect 69800 463194 70074 463250
rect 70130 463194 70200 463250
rect 69800 463126 70200 463194
rect 69800 463070 70074 463126
rect 70130 463070 70200 463126
rect 69800 463002 70200 463070
rect 69800 462946 70074 463002
rect 70130 462946 70200 463002
rect 69800 462878 70200 462946
rect 69800 462822 70074 462878
rect 70130 462822 70200 462878
rect 69800 462752 70200 462822
rect 69800 462134 70200 462172
rect 69800 462078 70074 462134
rect 70130 462078 70200 462134
rect 69800 462010 70200 462078
rect 69800 461954 70074 462010
rect 70130 461954 70200 462010
rect 69800 461886 70200 461954
rect 69800 461830 70074 461886
rect 70130 461830 70200 461886
rect 69800 461762 70200 461830
rect 69800 461706 70074 461762
rect 70130 461706 70200 461762
rect 69800 461638 70200 461706
rect 69800 461582 70074 461638
rect 70130 461582 70200 461638
rect 69800 461514 70200 461582
rect 69800 461458 70074 461514
rect 70130 461458 70200 461514
rect 69800 461390 70200 461458
rect 69800 461334 70074 461390
rect 70130 461334 70200 461390
rect 69800 461266 70200 461334
rect 69800 461210 70074 461266
rect 70130 461210 70200 461266
rect 69800 461142 70200 461210
rect 69800 461086 70074 461142
rect 70130 461086 70200 461142
rect 69800 461018 70200 461086
rect 69800 460962 70074 461018
rect 70130 460962 70200 461018
rect 69800 460894 70200 460962
rect 69800 460838 70074 460894
rect 70130 460838 70200 460894
rect 69800 460770 70200 460838
rect 69800 460714 70074 460770
rect 70130 460714 70200 460770
rect 69800 460646 70200 460714
rect 69800 460590 70074 460646
rect 70130 460590 70200 460646
rect 69800 460522 70200 460590
rect 69800 460466 70074 460522
rect 70130 460466 70200 460522
rect 69800 460398 70200 460466
rect 69800 460342 70074 460398
rect 70130 460342 70200 460398
rect 69800 460272 70200 460342
rect 707800 453658 708200 453728
rect 707800 453602 707870 453658
rect 707926 453602 708200 453658
rect 707800 453534 708200 453602
rect 707800 453478 707870 453534
rect 707926 453478 708200 453534
rect 707800 453410 708200 453478
rect 707800 453354 707870 453410
rect 707926 453354 708200 453410
rect 707800 453286 708200 453354
rect 707800 453230 707870 453286
rect 707926 453230 708200 453286
rect 707800 453162 708200 453230
rect 707800 453106 707870 453162
rect 707926 453106 708200 453162
rect 707800 453038 708200 453106
rect 707800 452982 707870 453038
rect 707926 452982 708200 453038
rect 707800 452914 708200 452982
rect 707800 452858 707870 452914
rect 707926 452858 708200 452914
rect 707800 452790 708200 452858
rect 707800 452734 707870 452790
rect 707926 452734 708200 452790
rect 707800 452666 708200 452734
rect 707800 452610 707870 452666
rect 707926 452610 708200 452666
rect 707800 452542 708200 452610
rect 707800 452486 707870 452542
rect 707926 452486 708200 452542
rect 707800 452418 708200 452486
rect 707800 452362 707870 452418
rect 707926 452362 708200 452418
rect 707800 452294 708200 452362
rect 707800 452238 707870 452294
rect 707926 452238 708200 452294
rect 707800 452170 708200 452238
rect 707800 452114 707870 452170
rect 707926 452114 708200 452170
rect 707800 452046 708200 452114
rect 707800 451990 707870 452046
rect 707926 451990 708200 452046
rect 707800 451922 708200 451990
rect 707800 451866 707870 451922
rect 707926 451866 708200 451922
rect 707800 451828 708200 451866
rect 707800 451178 708200 451248
rect 707800 451122 707870 451178
rect 707926 451122 708200 451178
rect 707800 451054 708200 451122
rect 707800 450998 707870 451054
rect 707926 450998 708200 451054
rect 707800 450930 708200 450998
rect 707800 450874 707870 450930
rect 707926 450874 708200 450930
rect 707800 450806 708200 450874
rect 707800 450750 707870 450806
rect 707926 450750 708200 450806
rect 707800 450682 708200 450750
rect 707800 450626 707870 450682
rect 707926 450626 708200 450682
rect 707800 450558 708200 450626
rect 707800 450502 707870 450558
rect 707926 450502 708200 450558
rect 707800 450434 708200 450502
rect 707800 450378 707870 450434
rect 707926 450378 708200 450434
rect 707800 450310 708200 450378
rect 707800 450254 707870 450310
rect 707926 450254 708200 450310
rect 707800 450186 708200 450254
rect 707800 450130 707870 450186
rect 707926 450130 708200 450186
rect 707800 450062 708200 450130
rect 707800 450006 707870 450062
rect 707926 450006 708200 450062
rect 707800 449938 708200 450006
rect 707800 449882 707870 449938
rect 707926 449882 708200 449938
rect 707800 449814 708200 449882
rect 707800 449758 707870 449814
rect 707926 449758 708200 449814
rect 707800 449690 708200 449758
rect 707800 449634 707870 449690
rect 707926 449634 708200 449690
rect 707800 449566 708200 449634
rect 707800 449510 707870 449566
rect 707926 449510 708200 449566
rect 707800 449442 708200 449510
rect 707800 449386 707870 449442
rect 707926 449386 708200 449442
rect 707800 449318 708200 449386
rect 707800 449262 707870 449318
rect 707926 449262 708200 449318
rect 707800 449198 708200 449262
rect 707800 448808 708200 448878
rect 707800 448752 707870 448808
rect 707926 448752 708200 448808
rect 707800 448684 708200 448752
rect 707800 448628 707870 448684
rect 707926 448628 708200 448684
rect 707800 448560 708200 448628
rect 707800 448504 707870 448560
rect 707926 448504 708200 448560
rect 707800 448436 708200 448504
rect 707800 448380 707870 448436
rect 707926 448380 708200 448436
rect 707800 448312 708200 448380
rect 707800 448256 707870 448312
rect 707926 448256 708200 448312
rect 707800 448188 708200 448256
rect 707800 448132 707870 448188
rect 707926 448132 708200 448188
rect 707800 448064 708200 448132
rect 707800 448008 707870 448064
rect 707926 448008 708200 448064
rect 707800 447940 708200 448008
rect 707800 447884 707870 447940
rect 707926 447884 708200 447940
rect 707800 447816 708200 447884
rect 707800 447760 707870 447816
rect 707926 447760 708200 447816
rect 707800 447692 708200 447760
rect 707800 447636 707870 447692
rect 707926 447636 708200 447692
rect 707800 447568 708200 447636
rect 707800 447512 707870 447568
rect 707926 447512 708200 447568
rect 707800 447444 708200 447512
rect 707800 447388 707870 447444
rect 707926 447388 708200 447444
rect 707800 447320 708200 447388
rect 707800 447264 707870 447320
rect 707926 447264 708200 447320
rect 707800 447196 708200 447264
rect 707800 447140 707870 447196
rect 707926 447140 708200 447196
rect 707800 447072 708200 447140
rect 707800 447016 707870 447072
rect 707926 447016 708200 447072
rect 707800 446948 708200 447016
rect 707800 446892 707870 446948
rect 707926 446892 708200 446948
rect 707800 446828 708200 446892
rect 707800 446102 708200 446172
rect 707800 446046 707870 446102
rect 707926 446046 708200 446102
rect 707800 445978 708200 446046
rect 707800 445922 707870 445978
rect 707926 445922 708200 445978
rect 707800 445854 708200 445922
rect 707800 445798 707870 445854
rect 707926 445798 708200 445854
rect 707800 445730 708200 445798
rect 707800 445674 707870 445730
rect 707926 445674 708200 445730
rect 707800 445606 708200 445674
rect 707800 445550 707870 445606
rect 707926 445550 708200 445606
rect 707800 445482 708200 445550
rect 707800 445426 707870 445482
rect 707926 445426 708200 445482
rect 707800 445358 708200 445426
rect 707800 445302 707870 445358
rect 707926 445302 708200 445358
rect 707800 445234 708200 445302
rect 707800 445178 707870 445234
rect 707926 445178 708200 445234
rect 707800 445110 708200 445178
rect 707800 445054 707870 445110
rect 707926 445054 708200 445110
rect 707800 444986 708200 445054
rect 707800 444930 707870 444986
rect 707926 444930 708200 444986
rect 707800 444862 708200 444930
rect 707800 444806 707870 444862
rect 707926 444806 708200 444862
rect 707800 444738 708200 444806
rect 707800 444682 707870 444738
rect 707926 444682 708200 444738
rect 707800 444614 708200 444682
rect 707800 444558 707870 444614
rect 707926 444558 708200 444614
rect 707800 444490 708200 444558
rect 707800 444434 707870 444490
rect 707926 444434 708200 444490
rect 707800 444366 708200 444434
rect 707800 444310 707870 444366
rect 707926 444310 708200 444366
rect 707800 444242 708200 444310
rect 707800 444186 707870 444242
rect 707926 444186 708200 444242
rect 707800 444122 708200 444186
rect 707800 443732 708200 443802
rect 707800 443676 707870 443732
rect 707926 443676 708200 443732
rect 707800 443608 708200 443676
rect 707800 443552 707870 443608
rect 707926 443552 708200 443608
rect 707800 443484 708200 443552
rect 707800 443428 707870 443484
rect 707926 443428 708200 443484
rect 707800 443360 708200 443428
rect 707800 443304 707870 443360
rect 707926 443304 708200 443360
rect 707800 443236 708200 443304
rect 707800 443180 707870 443236
rect 707926 443180 708200 443236
rect 707800 443112 708200 443180
rect 707800 443056 707870 443112
rect 707926 443056 708200 443112
rect 707800 442988 708200 443056
rect 707800 442932 707870 442988
rect 707926 442932 708200 442988
rect 707800 442864 708200 442932
rect 707800 442808 707870 442864
rect 707926 442808 708200 442864
rect 707800 442740 708200 442808
rect 707800 442684 707870 442740
rect 707926 442684 708200 442740
rect 707800 442616 708200 442684
rect 707800 442560 707870 442616
rect 707926 442560 708200 442616
rect 707800 442492 708200 442560
rect 707800 442436 707870 442492
rect 707926 442436 708200 442492
rect 707800 442368 708200 442436
rect 707800 442312 707870 442368
rect 707926 442312 708200 442368
rect 707800 442244 708200 442312
rect 707800 442188 707870 442244
rect 707926 442188 708200 442244
rect 707800 442120 708200 442188
rect 707800 442064 707870 442120
rect 707926 442064 708200 442120
rect 707800 441996 708200 442064
rect 707800 441940 707870 441996
rect 707926 441940 708200 441996
rect 707800 441872 708200 441940
rect 707800 441816 707870 441872
rect 707926 441816 708200 441872
rect 707800 441752 708200 441816
rect 707800 441134 708200 441172
rect 707800 441078 707870 441134
rect 707926 441078 708200 441134
rect 707800 441010 708200 441078
rect 707800 440954 707870 441010
rect 707926 440954 708200 441010
rect 707800 440886 708200 440954
rect 707800 440830 707870 440886
rect 707926 440830 708200 440886
rect 707800 440762 708200 440830
rect 707800 440706 707870 440762
rect 707926 440706 708200 440762
rect 707800 440638 708200 440706
rect 707800 440582 707870 440638
rect 707926 440582 708200 440638
rect 707800 440514 708200 440582
rect 707800 440458 707870 440514
rect 707926 440458 708200 440514
rect 707800 440390 708200 440458
rect 707800 440334 707870 440390
rect 707926 440334 708200 440390
rect 707800 440266 708200 440334
rect 707800 440210 707870 440266
rect 707926 440210 708200 440266
rect 707800 440142 708200 440210
rect 707800 440086 707870 440142
rect 707926 440086 708200 440142
rect 707800 440018 708200 440086
rect 707800 439962 707870 440018
rect 707926 439962 708200 440018
rect 707800 439894 708200 439962
rect 707800 439838 707870 439894
rect 707926 439838 708200 439894
rect 707800 439770 708200 439838
rect 707800 439714 707870 439770
rect 707926 439714 708200 439770
rect 707800 439646 708200 439714
rect 707800 439590 707870 439646
rect 707926 439590 708200 439646
rect 707800 439522 708200 439590
rect 707800 439466 707870 439522
rect 707926 439466 708200 439522
rect 707800 439398 708200 439466
rect 707800 439342 707870 439398
rect 707926 439342 708200 439398
rect 707800 439272 708200 439342
rect 69800 433658 70200 433728
rect 69800 433602 70074 433658
rect 70130 433602 70200 433658
rect 69800 433534 70200 433602
rect 69800 433478 70074 433534
rect 70130 433478 70200 433534
rect 69800 433410 70200 433478
rect 69800 433354 70074 433410
rect 70130 433354 70200 433410
rect 69800 433286 70200 433354
rect 69800 433230 70074 433286
rect 70130 433230 70200 433286
rect 69800 433162 70200 433230
rect 69800 433106 70074 433162
rect 70130 433106 70200 433162
rect 69800 433038 70200 433106
rect 69800 432982 70074 433038
rect 70130 432982 70200 433038
rect 69800 432914 70200 432982
rect 69800 432858 70074 432914
rect 70130 432858 70200 432914
rect 69800 432790 70200 432858
rect 69800 432734 70074 432790
rect 70130 432734 70200 432790
rect 69800 432666 70200 432734
rect 69800 432610 70074 432666
rect 70130 432610 70200 432666
rect 69800 432542 70200 432610
rect 69800 432486 70074 432542
rect 70130 432486 70200 432542
rect 69800 432418 70200 432486
rect 69800 432362 70074 432418
rect 70130 432362 70200 432418
rect 69800 432294 70200 432362
rect 69800 432238 70074 432294
rect 70130 432238 70200 432294
rect 69800 432170 70200 432238
rect 69800 432114 70074 432170
rect 70130 432114 70200 432170
rect 69800 432046 70200 432114
rect 69800 431990 70074 432046
rect 70130 431990 70200 432046
rect 69800 431922 70200 431990
rect 69800 431866 70074 431922
rect 70130 431866 70200 431922
rect 69800 431828 70200 431866
rect 69800 431184 70200 431248
rect 69800 431128 70074 431184
rect 70130 431128 70200 431184
rect 69800 431060 70200 431128
rect 69800 431004 70074 431060
rect 70130 431004 70200 431060
rect 69800 430936 70200 431004
rect 69800 430880 70074 430936
rect 70130 430880 70200 430936
rect 69800 430812 70200 430880
rect 69800 430756 70074 430812
rect 70130 430756 70200 430812
rect 69800 430688 70200 430756
rect 69800 430632 70074 430688
rect 70130 430632 70200 430688
rect 69800 430564 70200 430632
rect 69800 430508 70074 430564
rect 70130 430508 70200 430564
rect 69800 430440 70200 430508
rect 69800 430384 70074 430440
rect 70130 430384 70200 430440
rect 69800 430316 70200 430384
rect 69800 430260 70074 430316
rect 70130 430260 70200 430316
rect 69800 430192 70200 430260
rect 69800 430136 70074 430192
rect 70130 430136 70200 430192
rect 69800 430068 70200 430136
rect 69800 430012 70074 430068
rect 70130 430012 70200 430068
rect 69800 429944 70200 430012
rect 69800 429888 70074 429944
rect 70130 429888 70200 429944
rect 69800 429820 70200 429888
rect 69800 429764 70074 429820
rect 70130 429764 70200 429820
rect 69800 429696 70200 429764
rect 69800 429640 70074 429696
rect 70130 429640 70200 429696
rect 69800 429572 70200 429640
rect 69800 429516 70074 429572
rect 70130 429516 70200 429572
rect 69800 429448 70200 429516
rect 69800 429392 70074 429448
rect 70130 429392 70200 429448
rect 69800 429324 70200 429392
rect 69800 429268 70074 429324
rect 70130 429268 70200 429324
rect 69800 429198 70200 429268
rect 69800 428814 70200 428878
rect 69800 428758 70074 428814
rect 70130 428758 70200 428814
rect 69800 428690 70200 428758
rect 69800 428634 70074 428690
rect 70130 428634 70200 428690
rect 69800 428566 70200 428634
rect 69800 428510 70074 428566
rect 70130 428510 70200 428566
rect 69800 428442 70200 428510
rect 69800 428386 70074 428442
rect 70130 428386 70200 428442
rect 69800 428318 70200 428386
rect 69800 428262 70074 428318
rect 70130 428262 70200 428318
rect 69800 428194 70200 428262
rect 69800 428138 70074 428194
rect 70130 428138 70200 428194
rect 69800 428070 70200 428138
rect 69800 428014 70074 428070
rect 70130 428014 70200 428070
rect 69800 427946 70200 428014
rect 69800 427890 70074 427946
rect 70130 427890 70200 427946
rect 69800 427822 70200 427890
rect 69800 427766 70074 427822
rect 70130 427766 70200 427822
rect 69800 427698 70200 427766
rect 69800 427642 70074 427698
rect 70130 427642 70200 427698
rect 69800 427574 70200 427642
rect 69800 427518 70074 427574
rect 70130 427518 70200 427574
rect 69800 427450 70200 427518
rect 69800 427394 70074 427450
rect 70130 427394 70200 427450
rect 69800 427326 70200 427394
rect 69800 427270 70074 427326
rect 70130 427270 70200 427326
rect 69800 427202 70200 427270
rect 69800 427146 70074 427202
rect 70130 427146 70200 427202
rect 69800 427078 70200 427146
rect 69800 427022 70074 427078
rect 70130 427022 70200 427078
rect 69800 426954 70200 427022
rect 69800 426898 70074 426954
rect 70130 426898 70200 426954
rect 69800 426828 70200 426898
rect 69800 426108 70200 426172
rect 69800 426052 70074 426108
rect 70130 426052 70200 426108
rect 69800 425984 70200 426052
rect 69800 425928 70074 425984
rect 70130 425928 70200 425984
rect 69800 425860 70200 425928
rect 69800 425804 70074 425860
rect 70130 425804 70200 425860
rect 69800 425736 70200 425804
rect 69800 425680 70074 425736
rect 70130 425680 70200 425736
rect 69800 425612 70200 425680
rect 69800 425556 70074 425612
rect 70130 425556 70200 425612
rect 69800 425488 70200 425556
rect 69800 425432 70074 425488
rect 70130 425432 70200 425488
rect 69800 425364 70200 425432
rect 69800 425308 70074 425364
rect 70130 425308 70200 425364
rect 69800 425240 70200 425308
rect 69800 425184 70074 425240
rect 70130 425184 70200 425240
rect 69800 425116 70200 425184
rect 69800 425060 70074 425116
rect 70130 425060 70200 425116
rect 69800 424992 70200 425060
rect 69800 424936 70074 424992
rect 70130 424936 70200 424992
rect 69800 424868 70200 424936
rect 69800 424812 70074 424868
rect 70130 424812 70200 424868
rect 69800 424744 70200 424812
rect 69800 424688 70074 424744
rect 70130 424688 70200 424744
rect 69800 424620 70200 424688
rect 69800 424564 70074 424620
rect 70130 424564 70200 424620
rect 69800 424496 70200 424564
rect 69800 424440 70074 424496
rect 70130 424440 70200 424496
rect 69800 424372 70200 424440
rect 69800 424316 70074 424372
rect 70130 424316 70200 424372
rect 69800 424248 70200 424316
rect 69800 424192 70074 424248
rect 70130 424192 70200 424248
rect 69800 424122 70200 424192
rect 69800 423738 70200 423802
rect 69800 423682 70074 423738
rect 70130 423682 70200 423738
rect 69800 423614 70200 423682
rect 69800 423558 70074 423614
rect 70130 423558 70200 423614
rect 69800 423490 70200 423558
rect 69800 423434 70074 423490
rect 70130 423434 70200 423490
rect 69800 423366 70200 423434
rect 69800 423310 70074 423366
rect 70130 423310 70200 423366
rect 69800 423242 70200 423310
rect 69800 423186 70074 423242
rect 70130 423186 70200 423242
rect 69800 423118 70200 423186
rect 69800 423062 70074 423118
rect 70130 423062 70200 423118
rect 69800 422994 70200 423062
rect 69800 422938 70074 422994
rect 70130 422938 70200 422994
rect 69800 422870 70200 422938
rect 69800 422814 70074 422870
rect 70130 422814 70200 422870
rect 69800 422746 70200 422814
rect 69800 422690 70074 422746
rect 70130 422690 70200 422746
rect 69800 422622 70200 422690
rect 69800 422566 70074 422622
rect 70130 422566 70200 422622
rect 69800 422498 70200 422566
rect 69800 422442 70074 422498
rect 70130 422442 70200 422498
rect 69800 422374 70200 422442
rect 69800 422318 70074 422374
rect 70130 422318 70200 422374
rect 69800 422250 70200 422318
rect 69800 422194 70074 422250
rect 70130 422194 70200 422250
rect 69800 422126 70200 422194
rect 69800 422070 70074 422126
rect 70130 422070 70200 422126
rect 69800 422002 70200 422070
rect 69800 421946 70074 422002
rect 70130 421946 70200 422002
rect 69800 421878 70200 421946
rect 69800 421822 70074 421878
rect 70130 421822 70200 421878
rect 69800 421752 70200 421822
rect 69800 421134 70200 421172
rect 69800 421078 70074 421134
rect 70130 421078 70200 421134
rect 69800 421010 70200 421078
rect 69800 420954 70074 421010
rect 70130 420954 70200 421010
rect 69800 420886 70200 420954
rect 69800 420830 70074 420886
rect 70130 420830 70200 420886
rect 69800 420762 70200 420830
rect 69800 420706 70074 420762
rect 70130 420706 70200 420762
rect 69800 420638 70200 420706
rect 69800 420582 70074 420638
rect 70130 420582 70200 420638
rect 69800 420514 70200 420582
rect 69800 420458 70074 420514
rect 70130 420458 70200 420514
rect 69800 420390 70200 420458
rect 69800 420334 70074 420390
rect 70130 420334 70200 420390
rect 69800 420266 70200 420334
rect 69800 420210 70074 420266
rect 70130 420210 70200 420266
rect 69800 420142 70200 420210
rect 69800 420086 70074 420142
rect 70130 420086 70200 420142
rect 69800 420018 70200 420086
rect 69800 419962 70074 420018
rect 70130 419962 70200 420018
rect 69800 419894 70200 419962
rect 69800 419838 70074 419894
rect 70130 419838 70200 419894
rect 69800 419770 70200 419838
rect 69800 419714 70074 419770
rect 70130 419714 70200 419770
rect 69800 419646 70200 419714
rect 69800 419590 70074 419646
rect 70130 419590 70200 419646
rect 69800 419522 70200 419590
rect 69800 419466 70074 419522
rect 70130 419466 70200 419522
rect 69800 419398 70200 419466
rect 69800 419342 70074 419398
rect 70130 419342 70200 419398
rect 69800 419272 70200 419342
rect 707800 410658 708200 410728
rect 707800 410602 707870 410658
rect 707926 410602 708200 410658
rect 707800 410534 708200 410602
rect 707800 410478 707870 410534
rect 707926 410478 708200 410534
rect 707800 410410 708200 410478
rect 707800 410354 707870 410410
rect 707926 410354 708200 410410
rect 707800 410286 708200 410354
rect 707800 410230 707870 410286
rect 707926 410230 708200 410286
rect 707800 410162 708200 410230
rect 707800 410106 707870 410162
rect 707926 410106 708200 410162
rect 707800 410038 708200 410106
rect 707800 409982 707870 410038
rect 707926 409982 708200 410038
rect 707800 409914 708200 409982
rect 707800 409858 707870 409914
rect 707926 409858 708200 409914
rect 707800 409790 708200 409858
rect 707800 409734 707870 409790
rect 707926 409734 708200 409790
rect 707800 409666 708200 409734
rect 707800 409610 707870 409666
rect 707926 409610 708200 409666
rect 707800 409542 708200 409610
rect 707800 409486 707870 409542
rect 707926 409486 708200 409542
rect 707800 409418 708200 409486
rect 707800 409362 707870 409418
rect 707926 409362 708200 409418
rect 707800 409294 708200 409362
rect 707800 409238 707870 409294
rect 707926 409238 708200 409294
rect 707800 409170 708200 409238
rect 707800 409114 707870 409170
rect 707926 409114 708200 409170
rect 707800 409046 708200 409114
rect 707800 408990 707870 409046
rect 707926 408990 708200 409046
rect 707800 408922 708200 408990
rect 707800 408866 707870 408922
rect 707926 408866 708200 408922
rect 707800 408828 708200 408866
rect 707800 408178 708200 408248
rect 707800 408122 707870 408178
rect 707926 408122 708200 408178
rect 707800 408054 708200 408122
rect 707800 407998 707870 408054
rect 707926 407998 708200 408054
rect 707800 407930 708200 407998
rect 707800 407874 707870 407930
rect 707926 407874 708200 407930
rect 707800 407806 708200 407874
rect 707800 407750 707870 407806
rect 707926 407750 708200 407806
rect 707800 407682 708200 407750
rect 707800 407626 707870 407682
rect 707926 407626 708200 407682
rect 707800 407558 708200 407626
rect 707800 407502 707870 407558
rect 707926 407502 708200 407558
rect 707800 407434 708200 407502
rect 707800 407378 707870 407434
rect 707926 407378 708200 407434
rect 707800 407310 708200 407378
rect 707800 407254 707870 407310
rect 707926 407254 708200 407310
rect 707800 407186 708200 407254
rect 707800 407130 707870 407186
rect 707926 407130 708200 407186
rect 707800 407062 708200 407130
rect 707800 407006 707870 407062
rect 707926 407006 708200 407062
rect 707800 406938 708200 407006
rect 707800 406882 707870 406938
rect 707926 406882 708200 406938
rect 707800 406814 708200 406882
rect 707800 406758 707870 406814
rect 707926 406758 708200 406814
rect 707800 406690 708200 406758
rect 707800 406634 707870 406690
rect 707926 406634 708200 406690
rect 707800 406566 708200 406634
rect 707800 406510 707870 406566
rect 707926 406510 708200 406566
rect 707800 406442 708200 406510
rect 707800 406386 707870 406442
rect 707926 406386 708200 406442
rect 707800 406318 708200 406386
rect 707800 406262 707870 406318
rect 707926 406262 708200 406318
rect 707800 406198 708200 406262
rect 707800 405808 708200 405878
rect 707800 405752 707870 405808
rect 707926 405752 708200 405808
rect 707800 405684 708200 405752
rect 707800 405628 707870 405684
rect 707926 405628 708200 405684
rect 707800 405560 708200 405628
rect 707800 405504 707870 405560
rect 707926 405504 708200 405560
rect 707800 405436 708200 405504
rect 707800 405380 707870 405436
rect 707926 405380 708200 405436
rect 707800 405312 708200 405380
rect 707800 405256 707870 405312
rect 707926 405256 708200 405312
rect 707800 405188 708200 405256
rect 707800 405132 707870 405188
rect 707926 405132 708200 405188
rect 707800 405064 708200 405132
rect 707800 405008 707870 405064
rect 707926 405008 708200 405064
rect 707800 404940 708200 405008
rect 707800 404884 707870 404940
rect 707926 404884 708200 404940
rect 707800 404816 708200 404884
rect 707800 404760 707870 404816
rect 707926 404760 708200 404816
rect 707800 404692 708200 404760
rect 707800 404636 707870 404692
rect 707926 404636 708200 404692
rect 707800 404568 708200 404636
rect 707800 404512 707870 404568
rect 707926 404512 708200 404568
rect 707800 404444 708200 404512
rect 707800 404388 707870 404444
rect 707926 404388 708200 404444
rect 707800 404320 708200 404388
rect 707800 404264 707870 404320
rect 707926 404264 708200 404320
rect 707800 404196 708200 404264
rect 707800 404140 707870 404196
rect 707926 404140 708200 404196
rect 707800 404072 708200 404140
rect 707800 404016 707870 404072
rect 707926 404016 708200 404072
rect 707800 403948 708200 404016
rect 707800 403892 707870 403948
rect 707926 403892 708200 403948
rect 707800 403828 708200 403892
rect 707800 403102 708200 403172
rect 707800 403046 707870 403102
rect 707926 403046 708200 403102
rect 707800 402978 708200 403046
rect 707800 402922 707870 402978
rect 707926 402922 708200 402978
rect 707800 402854 708200 402922
rect 707800 402798 707870 402854
rect 707926 402798 708200 402854
rect 707800 402730 708200 402798
rect 707800 402674 707870 402730
rect 707926 402674 708200 402730
rect 707800 402606 708200 402674
rect 707800 402550 707870 402606
rect 707926 402550 708200 402606
rect 707800 402482 708200 402550
rect 707800 402426 707870 402482
rect 707926 402426 708200 402482
rect 707800 402358 708200 402426
rect 707800 402302 707870 402358
rect 707926 402302 708200 402358
rect 707800 402234 708200 402302
rect 707800 402178 707870 402234
rect 707926 402178 708200 402234
rect 707800 402110 708200 402178
rect 707800 402054 707870 402110
rect 707926 402054 708200 402110
rect 707800 401986 708200 402054
rect 707800 401930 707870 401986
rect 707926 401930 708200 401986
rect 707800 401862 708200 401930
rect 707800 401806 707870 401862
rect 707926 401806 708200 401862
rect 707800 401738 708200 401806
rect 707800 401682 707870 401738
rect 707926 401682 708200 401738
rect 707800 401614 708200 401682
rect 707800 401558 707870 401614
rect 707926 401558 708200 401614
rect 707800 401490 708200 401558
rect 707800 401434 707870 401490
rect 707926 401434 708200 401490
rect 707800 401366 708200 401434
rect 707800 401310 707870 401366
rect 707926 401310 708200 401366
rect 707800 401242 708200 401310
rect 707800 401186 707870 401242
rect 707926 401186 708200 401242
rect 707800 401122 708200 401186
rect 707800 400732 708200 400802
rect 707800 400676 707870 400732
rect 707926 400676 708200 400732
rect 707800 400608 708200 400676
rect 707800 400552 707870 400608
rect 707926 400552 708200 400608
rect 707800 400484 708200 400552
rect 707800 400428 707870 400484
rect 707926 400428 708200 400484
rect 707800 400360 708200 400428
rect 707800 400304 707870 400360
rect 707926 400304 708200 400360
rect 707800 400236 708200 400304
rect 707800 400180 707870 400236
rect 707926 400180 708200 400236
rect 707800 400112 708200 400180
rect 707800 400056 707870 400112
rect 707926 400056 708200 400112
rect 707800 399988 708200 400056
rect 707800 399932 707870 399988
rect 707926 399932 708200 399988
rect 707800 399864 708200 399932
rect 707800 399808 707870 399864
rect 707926 399808 708200 399864
rect 707800 399740 708200 399808
rect 707800 399684 707870 399740
rect 707926 399684 708200 399740
rect 707800 399616 708200 399684
rect 707800 399560 707870 399616
rect 707926 399560 708200 399616
rect 707800 399492 708200 399560
rect 707800 399436 707870 399492
rect 707926 399436 708200 399492
rect 707800 399368 708200 399436
rect 707800 399312 707870 399368
rect 707926 399312 708200 399368
rect 707800 399244 708200 399312
rect 707800 399188 707870 399244
rect 707926 399188 708200 399244
rect 707800 399120 708200 399188
rect 707800 399064 707870 399120
rect 707926 399064 708200 399120
rect 707800 398996 708200 399064
rect 707800 398940 707870 398996
rect 707926 398940 708200 398996
rect 707800 398872 708200 398940
rect 707800 398816 707870 398872
rect 707926 398816 708200 398872
rect 707800 398752 708200 398816
rect 707800 398134 708200 398172
rect 707800 398078 707870 398134
rect 707926 398078 708200 398134
rect 707800 398010 708200 398078
rect 707800 397954 707870 398010
rect 707926 397954 708200 398010
rect 707800 397886 708200 397954
rect 707800 397830 707870 397886
rect 707926 397830 708200 397886
rect 707800 397762 708200 397830
rect 707800 397706 707870 397762
rect 707926 397706 708200 397762
rect 707800 397638 708200 397706
rect 707800 397582 707870 397638
rect 707926 397582 708200 397638
rect 707800 397514 708200 397582
rect 707800 397458 707870 397514
rect 707926 397458 708200 397514
rect 707800 397390 708200 397458
rect 707800 397334 707870 397390
rect 707926 397334 708200 397390
rect 707800 397266 708200 397334
rect 707800 397210 707870 397266
rect 707926 397210 708200 397266
rect 707800 397142 708200 397210
rect 707800 397086 707870 397142
rect 707926 397086 708200 397142
rect 707800 397018 708200 397086
rect 707800 396962 707870 397018
rect 707926 396962 708200 397018
rect 707800 396894 708200 396962
rect 707800 396838 707870 396894
rect 707926 396838 708200 396894
rect 707800 396770 708200 396838
rect 707800 396714 707870 396770
rect 707926 396714 708200 396770
rect 707800 396646 708200 396714
rect 707800 396590 707870 396646
rect 707926 396590 708200 396646
rect 707800 396522 708200 396590
rect 707800 396466 707870 396522
rect 707926 396466 708200 396522
rect 707800 396398 708200 396466
rect 707800 396342 707870 396398
rect 707926 396342 708200 396398
rect 707800 396272 708200 396342
rect 69800 146658 70200 146728
rect 69800 146602 70074 146658
rect 70130 146602 70200 146658
rect 69800 146534 70200 146602
rect 69800 146478 70074 146534
rect 70130 146478 70200 146534
rect 69800 146410 70200 146478
rect 69800 146354 70074 146410
rect 70130 146354 70200 146410
rect 69800 146286 70200 146354
rect 69800 146230 70074 146286
rect 70130 146230 70200 146286
rect 69800 146162 70200 146230
rect 69800 146106 70074 146162
rect 70130 146106 70200 146162
rect 69800 146038 70200 146106
rect 69800 145982 70074 146038
rect 70130 145982 70200 146038
rect 69800 145914 70200 145982
rect 69800 145858 70074 145914
rect 70130 145858 70200 145914
rect 69800 145790 70200 145858
rect 69800 145734 70074 145790
rect 70130 145734 70200 145790
rect 69800 145666 70200 145734
rect 69800 145610 70074 145666
rect 70130 145610 70200 145666
rect 69800 145542 70200 145610
rect 69800 145486 70074 145542
rect 70130 145486 70200 145542
rect 69800 145418 70200 145486
rect 69800 145362 70074 145418
rect 70130 145362 70200 145418
rect 69800 145294 70200 145362
rect 69800 145238 70074 145294
rect 70130 145238 70200 145294
rect 69800 145170 70200 145238
rect 69800 145114 70074 145170
rect 70130 145114 70200 145170
rect 69800 145046 70200 145114
rect 69800 144990 70074 145046
rect 70130 144990 70200 145046
rect 69800 144922 70200 144990
rect 69800 144866 70074 144922
rect 70130 144866 70200 144922
rect 69800 144828 70200 144866
rect 69800 144184 70200 144248
rect 69800 144128 70074 144184
rect 70130 144128 70200 144184
rect 69800 144060 70200 144128
rect 69800 144004 70074 144060
rect 70130 144004 70200 144060
rect 69800 143936 70200 144004
rect 69800 143880 70074 143936
rect 70130 143880 70200 143936
rect 69800 143812 70200 143880
rect 69800 143756 70074 143812
rect 70130 143756 70200 143812
rect 69800 143688 70200 143756
rect 69800 143632 70074 143688
rect 70130 143632 70200 143688
rect 69800 143564 70200 143632
rect 69800 143508 70074 143564
rect 70130 143508 70200 143564
rect 69800 143440 70200 143508
rect 69800 143384 70074 143440
rect 70130 143384 70200 143440
rect 69800 143316 70200 143384
rect 69800 143260 70074 143316
rect 70130 143260 70200 143316
rect 69800 143192 70200 143260
rect 69800 143136 70074 143192
rect 70130 143136 70200 143192
rect 69800 143068 70200 143136
rect 69800 143012 70074 143068
rect 70130 143012 70200 143068
rect 69800 142944 70200 143012
rect 69800 142888 70074 142944
rect 70130 142888 70200 142944
rect 69800 142820 70200 142888
rect 69800 142764 70074 142820
rect 70130 142764 70200 142820
rect 69800 142696 70200 142764
rect 69800 142640 70074 142696
rect 70130 142640 70200 142696
rect 69800 142572 70200 142640
rect 69800 142516 70074 142572
rect 70130 142516 70200 142572
rect 69800 142448 70200 142516
rect 69800 142392 70074 142448
rect 70130 142392 70200 142448
rect 69800 142324 70200 142392
rect 69800 142268 70074 142324
rect 70130 142268 70200 142324
rect 69800 142198 70200 142268
rect 69800 141814 70200 141878
rect 69800 141758 70074 141814
rect 70130 141758 70200 141814
rect 69800 141690 70200 141758
rect 69800 141634 70074 141690
rect 70130 141634 70200 141690
rect 69800 141566 70200 141634
rect 69800 141510 70074 141566
rect 70130 141510 70200 141566
rect 69800 141442 70200 141510
rect 69800 141386 70074 141442
rect 70130 141386 70200 141442
rect 69800 141318 70200 141386
rect 69800 141262 70074 141318
rect 70130 141262 70200 141318
rect 69800 141194 70200 141262
rect 69800 141138 70074 141194
rect 70130 141138 70200 141194
rect 69800 141070 70200 141138
rect 69800 141014 70074 141070
rect 70130 141014 70200 141070
rect 69800 140946 70200 141014
rect 69800 140890 70074 140946
rect 70130 140890 70200 140946
rect 69800 140822 70200 140890
rect 69800 140766 70074 140822
rect 70130 140766 70200 140822
rect 69800 140698 70200 140766
rect 69800 140642 70074 140698
rect 70130 140642 70200 140698
rect 69800 140574 70200 140642
rect 69800 140518 70074 140574
rect 70130 140518 70200 140574
rect 69800 140450 70200 140518
rect 69800 140394 70074 140450
rect 70130 140394 70200 140450
rect 69800 140326 70200 140394
rect 69800 140270 70074 140326
rect 70130 140270 70200 140326
rect 69800 140202 70200 140270
rect 69800 140146 70074 140202
rect 70130 140146 70200 140202
rect 69800 140078 70200 140146
rect 69800 140022 70074 140078
rect 70130 140022 70200 140078
rect 69800 139954 70200 140022
rect 69800 139898 70074 139954
rect 70130 139898 70200 139954
rect 69800 139828 70200 139898
rect 69800 139108 70200 139172
rect 69800 139052 70074 139108
rect 70130 139052 70200 139108
rect 69800 138984 70200 139052
rect 69800 138928 70074 138984
rect 70130 138928 70200 138984
rect 69800 138860 70200 138928
rect 69800 138804 70074 138860
rect 70130 138804 70200 138860
rect 69800 138736 70200 138804
rect 69800 138680 70074 138736
rect 70130 138680 70200 138736
rect 69800 138612 70200 138680
rect 69800 138556 70074 138612
rect 70130 138556 70200 138612
rect 69800 138488 70200 138556
rect 69800 138432 70074 138488
rect 70130 138432 70200 138488
rect 69800 138364 70200 138432
rect 69800 138308 70074 138364
rect 70130 138308 70200 138364
rect 69800 138240 70200 138308
rect 69800 138184 70074 138240
rect 70130 138184 70200 138240
rect 69800 138116 70200 138184
rect 69800 138060 70074 138116
rect 70130 138060 70200 138116
rect 69800 137992 70200 138060
rect 69800 137936 70074 137992
rect 70130 137936 70200 137992
rect 69800 137868 70200 137936
rect 69800 137812 70074 137868
rect 70130 137812 70200 137868
rect 69800 137744 70200 137812
rect 69800 137688 70074 137744
rect 70130 137688 70200 137744
rect 69800 137620 70200 137688
rect 69800 137564 70074 137620
rect 70130 137564 70200 137620
rect 69800 137496 70200 137564
rect 69800 137440 70074 137496
rect 70130 137440 70200 137496
rect 69800 137372 70200 137440
rect 69800 137316 70074 137372
rect 70130 137316 70200 137372
rect 69800 137248 70200 137316
rect 69800 137192 70074 137248
rect 70130 137192 70200 137248
rect 69800 137122 70200 137192
rect 69800 136738 70200 136802
rect 69800 136682 70074 136738
rect 70130 136682 70200 136738
rect 69800 136614 70200 136682
rect 69800 136558 70074 136614
rect 70130 136558 70200 136614
rect 69800 136490 70200 136558
rect 69800 136434 70074 136490
rect 70130 136434 70200 136490
rect 69800 136366 70200 136434
rect 69800 136310 70074 136366
rect 70130 136310 70200 136366
rect 69800 136242 70200 136310
rect 69800 136186 70074 136242
rect 70130 136186 70200 136242
rect 69800 136118 70200 136186
rect 69800 136062 70074 136118
rect 70130 136062 70200 136118
rect 69800 135994 70200 136062
rect 69800 135938 70074 135994
rect 70130 135938 70200 135994
rect 69800 135870 70200 135938
rect 69800 135814 70074 135870
rect 70130 135814 70200 135870
rect 69800 135746 70200 135814
rect 69800 135690 70074 135746
rect 70130 135690 70200 135746
rect 69800 135622 70200 135690
rect 69800 135566 70074 135622
rect 70130 135566 70200 135622
rect 69800 135498 70200 135566
rect 69800 135442 70074 135498
rect 70130 135442 70200 135498
rect 69800 135374 70200 135442
rect 69800 135318 70074 135374
rect 70130 135318 70200 135374
rect 69800 135250 70200 135318
rect 69800 135194 70074 135250
rect 70130 135194 70200 135250
rect 69800 135126 70200 135194
rect 69800 135070 70074 135126
rect 70130 135070 70200 135126
rect 69800 135002 70200 135070
rect 69800 134946 70074 135002
rect 70130 134946 70200 135002
rect 69800 134878 70200 134946
rect 69800 134822 70074 134878
rect 70130 134822 70200 134878
rect 69800 134752 70200 134822
rect 69800 134134 70200 134172
rect 69800 134078 70074 134134
rect 70130 134078 70200 134134
rect 69800 134010 70200 134078
rect 69800 133954 70074 134010
rect 70130 133954 70200 134010
rect 69800 133886 70200 133954
rect 69800 133830 70074 133886
rect 70130 133830 70200 133886
rect 69800 133762 70200 133830
rect 69800 133706 70074 133762
rect 70130 133706 70200 133762
rect 69800 133638 70200 133706
rect 69800 133582 70074 133638
rect 70130 133582 70200 133638
rect 69800 133514 70200 133582
rect 69800 133458 70074 133514
rect 70130 133458 70200 133514
rect 69800 133390 70200 133458
rect 69800 133334 70074 133390
rect 70130 133334 70200 133390
rect 69800 133266 70200 133334
rect 69800 133210 70074 133266
rect 70130 133210 70200 133266
rect 69800 133142 70200 133210
rect 69800 133086 70074 133142
rect 70130 133086 70200 133142
rect 69800 133018 70200 133086
rect 69800 132962 70074 133018
rect 70130 132962 70200 133018
rect 69800 132894 70200 132962
rect 69800 132838 70074 132894
rect 70130 132838 70200 132894
rect 69800 132770 70200 132838
rect 69800 132714 70074 132770
rect 70130 132714 70200 132770
rect 69800 132646 70200 132714
rect 69800 132590 70074 132646
rect 70130 132590 70200 132646
rect 69800 132522 70200 132590
rect 69800 132466 70074 132522
rect 70130 132466 70200 132522
rect 69800 132398 70200 132466
rect 69800 132342 70074 132398
rect 70130 132342 70200 132398
rect 69800 132272 70200 132342
rect 69800 105658 70200 105728
rect 69800 105602 70074 105658
rect 70130 105602 70200 105658
rect 69800 105534 70200 105602
rect 69800 105478 70074 105534
rect 70130 105478 70200 105534
rect 69800 105410 70200 105478
rect 69800 105354 70074 105410
rect 70130 105354 70200 105410
rect 69800 105286 70200 105354
rect 69800 105230 70074 105286
rect 70130 105230 70200 105286
rect 69800 105162 70200 105230
rect 69800 105106 70074 105162
rect 70130 105106 70200 105162
rect 69800 105038 70200 105106
rect 69800 104982 70074 105038
rect 70130 104982 70200 105038
rect 69800 104914 70200 104982
rect 69800 104858 70074 104914
rect 70130 104858 70200 104914
rect 69800 104790 70200 104858
rect 69800 104734 70074 104790
rect 70130 104734 70200 104790
rect 69800 104666 70200 104734
rect 69800 104610 70074 104666
rect 70130 104610 70200 104666
rect 69800 104542 70200 104610
rect 69800 104486 70074 104542
rect 70130 104486 70200 104542
rect 69800 104418 70200 104486
rect 69800 104362 70074 104418
rect 70130 104362 70200 104418
rect 69800 104294 70200 104362
rect 69800 104238 70074 104294
rect 70130 104238 70200 104294
rect 69800 104170 70200 104238
rect 69800 104114 70074 104170
rect 70130 104114 70200 104170
rect 69800 104046 70200 104114
rect 69800 103990 70074 104046
rect 70130 103990 70200 104046
rect 69800 103922 70200 103990
rect 69800 103866 70074 103922
rect 70130 103866 70200 103922
rect 69800 103828 70200 103866
rect 69800 103184 70200 103248
rect 69800 103128 70074 103184
rect 70130 103128 70200 103184
rect 69800 103060 70200 103128
rect 69800 103004 70074 103060
rect 70130 103004 70200 103060
rect 69800 102936 70200 103004
rect 69800 102880 70074 102936
rect 70130 102880 70200 102936
rect 69800 102812 70200 102880
rect 69800 102756 70074 102812
rect 70130 102756 70200 102812
rect 69800 102688 70200 102756
rect 69800 102632 70074 102688
rect 70130 102632 70200 102688
rect 69800 102564 70200 102632
rect 69800 102508 70074 102564
rect 70130 102508 70200 102564
rect 69800 102440 70200 102508
rect 69800 102384 70074 102440
rect 70130 102384 70200 102440
rect 69800 102316 70200 102384
rect 69800 102260 70074 102316
rect 70130 102260 70200 102316
rect 69800 102192 70200 102260
rect 69800 102136 70074 102192
rect 70130 102136 70200 102192
rect 69800 102068 70200 102136
rect 69800 102012 70074 102068
rect 70130 102012 70200 102068
rect 69800 101944 70200 102012
rect 69800 101888 70074 101944
rect 70130 101888 70200 101944
rect 69800 101820 70200 101888
rect 69800 101764 70074 101820
rect 70130 101764 70200 101820
rect 69800 101696 70200 101764
rect 69800 101640 70074 101696
rect 70130 101640 70200 101696
rect 69800 101572 70200 101640
rect 69800 101516 70074 101572
rect 70130 101516 70200 101572
rect 69800 101448 70200 101516
rect 69800 101392 70074 101448
rect 70130 101392 70200 101448
rect 69800 101324 70200 101392
rect 69800 101268 70074 101324
rect 70130 101268 70200 101324
rect 69800 101198 70200 101268
rect 69800 100814 70200 100878
rect 69800 100758 70074 100814
rect 70130 100758 70200 100814
rect 69800 100690 70200 100758
rect 69800 100634 70074 100690
rect 70130 100634 70200 100690
rect 69800 100566 70200 100634
rect 69800 100510 70074 100566
rect 70130 100510 70200 100566
rect 69800 100442 70200 100510
rect 69800 100386 70074 100442
rect 70130 100386 70200 100442
rect 69800 100318 70200 100386
rect 69800 100262 70074 100318
rect 70130 100262 70200 100318
rect 69800 100194 70200 100262
rect 69800 100138 70074 100194
rect 70130 100138 70200 100194
rect 69800 100070 70200 100138
rect 69800 100014 70074 100070
rect 70130 100014 70200 100070
rect 69800 99946 70200 100014
rect 69800 99890 70074 99946
rect 70130 99890 70200 99946
rect 69800 99822 70200 99890
rect 69800 99766 70074 99822
rect 70130 99766 70200 99822
rect 69800 99698 70200 99766
rect 69800 99642 70074 99698
rect 70130 99642 70200 99698
rect 69800 99574 70200 99642
rect 69800 99518 70074 99574
rect 70130 99518 70200 99574
rect 69800 99450 70200 99518
rect 69800 99394 70074 99450
rect 70130 99394 70200 99450
rect 69800 99326 70200 99394
rect 69800 99270 70074 99326
rect 70130 99270 70200 99326
rect 69800 99202 70200 99270
rect 69800 99146 70074 99202
rect 70130 99146 70200 99202
rect 69800 99078 70200 99146
rect 69800 99022 70074 99078
rect 70130 99022 70200 99078
rect 69800 98954 70200 99022
rect 69800 98898 70074 98954
rect 70130 98898 70200 98954
rect 69800 98828 70200 98898
rect 69800 98108 70200 98172
rect 69800 98052 70074 98108
rect 70130 98052 70200 98108
rect 69800 97984 70200 98052
rect 69800 97928 70074 97984
rect 70130 97928 70200 97984
rect 69800 97860 70200 97928
rect 69800 97804 70074 97860
rect 70130 97804 70200 97860
rect 69800 97736 70200 97804
rect 69800 97680 70074 97736
rect 70130 97680 70200 97736
rect 69800 97612 70200 97680
rect 69800 97556 70074 97612
rect 70130 97556 70200 97612
rect 69800 97488 70200 97556
rect 69800 97432 70074 97488
rect 70130 97432 70200 97488
rect 69800 97364 70200 97432
rect 69800 97308 70074 97364
rect 70130 97308 70200 97364
rect 69800 97240 70200 97308
rect 69800 97184 70074 97240
rect 70130 97184 70200 97240
rect 69800 97116 70200 97184
rect 69800 97060 70074 97116
rect 70130 97060 70200 97116
rect 69800 96992 70200 97060
rect 69800 96936 70074 96992
rect 70130 96936 70200 96992
rect 69800 96868 70200 96936
rect 69800 96812 70074 96868
rect 70130 96812 70200 96868
rect 69800 96744 70200 96812
rect 69800 96688 70074 96744
rect 70130 96688 70200 96744
rect 69800 96620 70200 96688
rect 69800 96564 70074 96620
rect 70130 96564 70200 96620
rect 69800 96496 70200 96564
rect 69800 96440 70074 96496
rect 70130 96440 70200 96496
rect 69800 96372 70200 96440
rect 69800 96316 70074 96372
rect 70130 96316 70200 96372
rect 69800 96248 70200 96316
rect 69800 96192 70074 96248
rect 70130 96192 70200 96248
rect 69800 96122 70200 96192
rect 69800 95738 70200 95802
rect 69800 95682 70074 95738
rect 70130 95682 70200 95738
rect 69800 95614 70200 95682
rect 69800 95558 70074 95614
rect 70130 95558 70200 95614
rect 69800 95490 70200 95558
rect 69800 95434 70074 95490
rect 70130 95434 70200 95490
rect 69800 95366 70200 95434
rect 69800 95310 70074 95366
rect 70130 95310 70200 95366
rect 69800 95242 70200 95310
rect 69800 95186 70074 95242
rect 70130 95186 70200 95242
rect 69800 95118 70200 95186
rect 69800 95062 70074 95118
rect 70130 95062 70200 95118
rect 69800 94994 70200 95062
rect 69800 94938 70074 94994
rect 70130 94938 70200 94994
rect 69800 94870 70200 94938
rect 69800 94814 70074 94870
rect 70130 94814 70200 94870
rect 69800 94746 70200 94814
rect 69800 94690 70074 94746
rect 70130 94690 70200 94746
rect 69800 94622 70200 94690
rect 69800 94566 70074 94622
rect 70130 94566 70200 94622
rect 69800 94498 70200 94566
rect 69800 94442 70074 94498
rect 70130 94442 70200 94498
rect 69800 94374 70200 94442
rect 69800 94318 70074 94374
rect 70130 94318 70200 94374
rect 69800 94250 70200 94318
rect 69800 94194 70074 94250
rect 70130 94194 70200 94250
rect 69800 94126 70200 94194
rect 69800 94070 70074 94126
rect 70130 94070 70200 94126
rect 69800 94002 70200 94070
rect 69800 93946 70074 94002
rect 70130 93946 70200 94002
rect 69800 93878 70200 93946
rect 69800 93822 70074 93878
rect 70130 93822 70200 93878
rect 69800 93752 70200 93822
rect 69800 93134 70200 93172
rect 69800 93078 70074 93134
rect 70130 93078 70200 93134
rect 69800 93010 70200 93078
rect 69800 92954 70074 93010
rect 70130 92954 70200 93010
rect 69800 92886 70200 92954
rect 69800 92830 70074 92886
rect 70130 92830 70200 92886
rect 69800 92762 70200 92830
rect 69800 92706 70074 92762
rect 70130 92706 70200 92762
rect 69800 92638 70200 92706
rect 69800 92582 70074 92638
rect 70130 92582 70200 92638
rect 69800 92514 70200 92582
rect 69800 92458 70074 92514
rect 70130 92458 70200 92514
rect 69800 92390 70200 92458
rect 69800 92334 70074 92390
rect 70130 92334 70200 92390
rect 69800 92266 70200 92334
rect 69800 92210 70074 92266
rect 70130 92210 70200 92266
rect 69800 92142 70200 92210
rect 69800 92086 70074 92142
rect 70130 92086 70200 92142
rect 69800 92018 70200 92086
rect 69800 91962 70074 92018
rect 70130 91962 70200 92018
rect 69800 91894 70200 91962
rect 69800 91838 70074 91894
rect 70130 91838 70200 91894
rect 69800 91770 70200 91838
rect 69800 91714 70074 91770
rect 70130 91714 70200 91770
rect 69800 91646 70200 91714
rect 69800 91590 70074 91646
rect 70130 91590 70200 91646
rect 69800 91522 70200 91590
rect 69800 91466 70074 91522
rect 70130 91466 70200 91522
rect 69800 91398 70200 91466
rect 69800 91342 70074 91398
rect 70130 91342 70200 91398
rect 69800 91272 70200 91342
rect 107272 70130 109172 70200
rect 107272 70074 107342 70130
rect 107398 70074 107466 70130
rect 107522 70074 107590 70130
rect 107646 70074 107714 70130
rect 107770 70074 107838 70130
rect 107894 70074 107962 70130
rect 108018 70074 108086 70130
rect 108142 70074 108210 70130
rect 108266 70074 108334 70130
rect 108390 70074 108458 70130
rect 108514 70074 108582 70130
rect 108638 70074 108706 70130
rect 108762 70074 108830 70130
rect 108886 70074 108954 70130
rect 109010 70074 109078 70130
rect 109134 70074 109172 70130
rect 107272 69800 109172 70074
rect 109752 70130 111802 70200
rect 109752 70074 109822 70130
rect 109878 70074 109946 70130
rect 110002 70074 110070 70130
rect 110126 70074 110194 70130
rect 110250 70074 110318 70130
rect 110374 70074 110442 70130
rect 110498 70074 110566 70130
rect 110622 70074 110690 70130
rect 110746 70074 110814 70130
rect 110870 70074 110938 70130
rect 110994 70074 111062 70130
rect 111118 70074 111186 70130
rect 111242 70074 111310 70130
rect 111366 70074 111434 70130
rect 111490 70074 111558 70130
rect 111614 70074 111682 70130
rect 111738 70074 111802 70130
rect 109752 69800 111802 70074
rect 112122 70130 114172 70200
rect 112122 70074 112192 70130
rect 112248 70074 112316 70130
rect 112372 70074 112440 70130
rect 112496 70074 112564 70130
rect 112620 70074 112688 70130
rect 112744 70074 112812 70130
rect 112868 70074 112936 70130
rect 112992 70074 113060 70130
rect 113116 70074 113184 70130
rect 113240 70074 113308 70130
rect 113364 70074 113432 70130
rect 113488 70074 113556 70130
rect 113612 70074 113680 70130
rect 113736 70074 113804 70130
rect 113860 70074 113928 70130
rect 113984 70074 114052 70130
rect 114108 70074 114172 70130
rect 112122 69800 114172 70074
rect 114828 70130 116878 70200
rect 114828 70074 114892 70130
rect 114948 70074 115016 70130
rect 115072 70074 115140 70130
rect 115196 70074 115264 70130
rect 115320 70074 115388 70130
rect 115444 70074 115512 70130
rect 115568 70074 115636 70130
rect 115692 70074 115760 70130
rect 115816 70074 115884 70130
rect 115940 70074 116008 70130
rect 116064 70074 116132 70130
rect 116188 70074 116256 70130
rect 116312 70074 116380 70130
rect 116436 70074 116504 70130
rect 116560 70074 116628 70130
rect 116684 70074 116752 70130
rect 116808 70074 116878 70130
rect 114828 69800 116878 70074
rect 117198 70130 119248 70200
rect 117198 70074 117262 70130
rect 117318 70074 117386 70130
rect 117442 70074 117510 70130
rect 117566 70074 117634 70130
rect 117690 70074 117758 70130
rect 117814 70074 117882 70130
rect 117938 70074 118006 70130
rect 118062 70074 118130 70130
rect 118186 70074 118254 70130
rect 118310 70074 118378 70130
rect 118434 70074 118502 70130
rect 118558 70074 118626 70130
rect 118682 70074 118750 70130
rect 118806 70074 118874 70130
rect 118930 70074 118998 70130
rect 119054 70074 119122 70130
rect 119178 70074 119248 70130
rect 117198 69800 119248 70074
rect 119828 70130 121728 70200
rect 119828 70074 119866 70130
rect 119922 70074 119990 70130
rect 120046 70074 120114 70130
rect 120170 70074 120238 70130
rect 120294 70074 120362 70130
rect 120418 70074 120486 70130
rect 120542 70074 120610 70130
rect 120666 70074 120734 70130
rect 120790 70074 120858 70130
rect 120914 70074 120982 70130
rect 121038 70074 121106 70130
rect 121162 70074 121230 70130
rect 121286 70074 121354 70130
rect 121410 70074 121478 70130
rect 121534 70074 121602 70130
rect 121658 70074 121728 70130
rect 119828 69800 121728 70074
rect 272272 70130 274172 70200
rect 272272 70074 272342 70130
rect 272398 70074 272466 70130
rect 272522 70074 272590 70130
rect 272646 70074 272714 70130
rect 272770 70074 272838 70130
rect 272894 70074 272962 70130
rect 273018 70074 273086 70130
rect 273142 70074 273210 70130
rect 273266 70074 273334 70130
rect 273390 70074 273458 70130
rect 273514 70074 273582 70130
rect 273638 70074 273706 70130
rect 273762 70074 273830 70130
rect 273886 70074 273954 70130
rect 274010 70074 274078 70130
rect 274134 70074 274172 70130
rect 272272 69800 274172 70074
rect 274752 70130 276802 70200
rect 274752 70074 274822 70130
rect 274878 70074 274946 70130
rect 275002 70074 275070 70130
rect 275126 70074 275194 70130
rect 275250 70074 275318 70130
rect 275374 70074 275442 70130
rect 275498 70074 275566 70130
rect 275622 70074 275690 70130
rect 275746 70074 275814 70130
rect 275870 70074 275938 70130
rect 275994 70074 276062 70130
rect 276118 70074 276186 70130
rect 276242 70074 276310 70130
rect 276366 70074 276434 70130
rect 276490 70074 276558 70130
rect 276614 70074 276682 70130
rect 276738 70074 276802 70130
rect 274752 69800 276802 70074
rect 277122 70130 279172 70200
rect 277122 70074 277192 70130
rect 277248 70074 277316 70130
rect 277372 70074 277440 70130
rect 277496 70074 277564 70130
rect 277620 70074 277688 70130
rect 277744 70074 277812 70130
rect 277868 70074 277936 70130
rect 277992 70074 278060 70130
rect 278116 70074 278184 70130
rect 278240 70074 278308 70130
rect 278364 70074 278432 70130
rect 278488 70074 278556 70130
rect 278612 70074 278680 70130
rect 278736 70074 278804 70130
rect 278860 70074 278928 70130
rect 278984 70074 279052 70130
rect 279108 70074 279172 70130
rect 277122 69800 279172 70074
rect 279828 70130 281878 70200
rect 279828 70074 279892 70130
rect 279948 70074 280016 70130
rect 280072 70074 280140 70130
rect 280196 70074 280264 70130
rect 280320 70074 280388 70130
rect 280444 70074 280512 70130
rect 280568 70074 280636 70130
rect 280692 70074 280760 70130
rect 280816 70074 280884 70130
rect 280940 70074 281008 70130
rect 281064 70074 281132 70130
rect 281188 70074 281256 70130
rect 281312 70074 281380 70130
rect 281436 70074 281504 70130
rect 281560 70074 281628 70130
rect 281684 70074 281752 70130
rect 281808 70074 281878 70130
rect 279828 69800 281878 70074
rect 282198 70130 284248 70200
rect 282198 70074 282262 70130
rect 282318 70074 282386 70130
rect 282442 70074 282510 70130
rect 282566 70074 282634 70130
rect 282690 70074 282758 70130
rect 282814 70074 282882 70130
rect 282938 70074 283006 70130
rect 283062 70074 283130 70130
rect 283186 70074 283254 70130
rect 283310 70074 283378 70130
rect 283434 70074 283502 70130
rect 283558 70074 283626 70130
rect 283682 70074 283750 70130
rect 283806 70074 283874 70130
rect 283930 70074 283998 70130
rect 284054 70074 284122 70130
rect 284178 70074 284248 70130
rect 282198 69800 284248 70074
rect 284828 70130 286728 70200
rect 284828 70074 284866 70130
rect 284922 70074 284990 70130
rect 285046 70074 285114 70130
rect 285170 70074 285238 70130
rect 285294 70074 285362 70130
rect 285418 70074 285486 70130
rect 285542 70074 285610 70130
rect 285666 70074 285734 70130
rect 285790 70074 285858 70130
rect 285914 70074 285982 70130
rect 286038 70074 286106 70130
rect 286162 70074 286230 70130
rect 286286 70074 286354 70130
rect 286410 70074 286478 70130
rect 286534 70074 286602 70130
rect 286658 70074 286728 70130
rect 284828 69800 286728 70074
rect 602272 70130 604172 70200
rect 602272 70074 602342 70130
rect 602398 70074 602466 70130
rect 602522 70074 602590 70130
rect 602646 70074 602714 70130
rect 602770 70074 602838 70130
rect 602894 70074 602962 70130
rect 603018 70074 603086 70130
rect 603142 70074 603210 70130
rect 603266 70074 603334 70130
rect 603390 70074 603458 70130
rect 603514 70074 603582 70130
rect 603638 70074 603706 70130
rect 603762 70074 603830 70130
rect 603886 70074 603954 70130
rect 604010 70074 604078 70130
rect 604134 70074 604172 70130
rect 602272 69800 604172 70074
rect 604752 70130 606802 70200
rect 604752 70074 604822 70130
rect 604878 70074 604946 70130
rect 605002 70074 605070 70130
rect 605126 70074 605194 70130
rect 605250 70074 605318 70130
rect 605374 70074 605442 70130
rect 605498 70074 605566 70130
rect 605622 70074 605690 70130
rect 605746 70074 605814 70130
rect 605870 70074 605938 70130
rect 605994 70074 606062 70130
rect 606118 70074 606186 70130
rect 606242 70074 606310 70130
rect 606366 70074 606434 70130
rect 606490 70074 606558 70130
rect 606614 70074 606682 70130
rect 606738 70074 606802 70130
rect 604752 69800 606802 70074
rect 607122 70130 609172 70200
rect 607122 70074 607192 70130
rect 607248 70074 607316 70130
rect 607372 70074 607440 70130
rect 607496 70074 607564 70130
rect 607620 70074 607688 70130
rect 607744 70074 607812 70130
rect 607868 70074 607936 70130
rect 607992 70074 608060 70130
rect 608116 70074 608184 70130
rect 608240 70074 608308 70130
rect 608364 70074 608432 70130
rect 608488 70074 608556 70130
rect 608612 70074 608680 70130
rect 608736 70074 608804 70130
rect 608860 70074 608928 70130
rect 608984 70074 609052 70130
rect 609108 70074 609172 70130
rect 607122 69800 609172 70074
rect 609828 70130 611878 70200
rect 609828 70074 609892 70130
rect 609948 70074 610016 70130
rect 610072 70074 610140 70130
rect 610196 70074 610264 70130
rect 610320 70074 610388 70130
rect 610444 70074 610512 70130
rect 610568 70074 610636 70130
rect 610692 70074 610760 70130
rect 610816 70074 610884 70130
rect 610940 70074 611008 70130
rect 611064 70074 611132 70130
rect 611188 70074 611256 70130
rect 611312 70074 611380 70130
rect 611436 70074 611504 70130
rect 611560 70074 611628 70130
rect 611684 70074 611752 70130
rect 611808 70074 611878 70130
rect 609828 69800 611878 70074
rect 612198 70130 614248 70200
rect 612198 70074 612262 70130
rect 612318 70074 612386 70130
rect 612442 70074 612510 70130
rect 612566 70074 612634 70130
rect 612690 70074 612758 70130
rect 612814 70074 612882 70130
rect 612938 70074 613006 70130
rect 613062 70074 613130 70130
rect 613186 70074 613254 70130
rect 613310 70074 613378 70130
rect 613434 70074 613502 70130
rect 613558 70074 613626 70130
rect 613682 70074 613750 70130
rect 613806 70074 613874 70130
rect 613930 70074 613998 70130
rect 614054 70074 614122 70130
rect 614178 70074 614248 70130
rect 612198 69800 614248 70074
rect 614828 70130 616728 70200
rect 614828 70074 614866 70130
rect 614922 70074 614990 70130
rect 615046 70074 615114 70130
rect 615170 70074 615238 70130
rect 615294 70074 615362 70130
rect 615418 70074 615486 70130
rect 615542 70074 615610 70130
rect 615666 70074 615734 70130
rect 615790 70074 615858 70130
rect 615914 70074 615982 70130
rect 616038 70074 616106 70130
rect 616162 70074 616230 70130
rect 616286 70074 616354 70130
rect 616410 70074 616478 70130
rect 616534 70074 616602 70130
rect 616658 70074 616728 70130
rect 614828 69800 616728 70074
rect 657272 70130 659172 70200
rect 657272 70074 657342 70130
rect 657398 70074 657466 70130
rect 657522 70074 657590 70130
rect 657646 70074 657714 70130
rect 657770 70074 657838 70130
rect 657894 70074 657962 70130
rect 658018 70074 658086 70130
rect 658142 70074 658210 70130
rect 658266 70074 658334 70130
rect 658390 70074 658458 70130
rect 658514 70074 658582 70130
rect 658638 70074 658706 70130
rect 658762 70074 658830 70130
rect 658886 70074 658954 70130
rect 659010 70074 659078 70130
rect 659134 70074 659172 70130
rect 657272 69800 659172 70074
rect 659752 70130 661802 70200
rect 659752 70074 659822 70130
rect 659878 70074 659946 70130
rect 660002 70074 660070 70130
rect 660126 70074 660194 70130
rect 660250 70074 660318 70130
rect 660374 70074 660442 70130
rect 660498 70074 660566 70130
rect 660622 70074 660690 70130
rect 660746 70074 660814 70130
rect 660870 70074 660938 70130
rect 660994 70074 661062 70130
rect 661118 70074 661186 70130
rect 661242 70074 661310 70130
rect 661366 70074 661434 70130
rect 661490 70074 661558 70130
rect 661614 70074 661682 70130
rect 661738 70074 661802 70130
rect 659752 69800 661802 70074
rect 662122 70130 664172 70200
rect 662122 70074 662192 70130
rect 662248 70074 662316 70130
rect 662372 70074 662440 70130
rect 662496 70074 662564 70130
rect 662620 70074 662688 70130
rect 662744 70074 662812 70130
rect 662868 70074 662936 70130
rect 662992 70074 663060 70130
rect 663116 70074 663184 70130
rect 663240 70074 663308 70130
rect 663364 70074 663432 70130
rect 663488 70074 663556 70130
rect 663612 70074 663680 70130
rect 663736 70074 663804 70130
rect 663860 70074 663928 70130
rect 663984 70074 664052 70130
rect 664108 70074 664172 70130
rect 662122 69800 664172 70074
rect 664828 70130 666878 70200
rect 664828 70074 664892 70130
rect 664948 70074 665016 70130
rect 665072 70074 665140 70130
rect 665196 70074 665264 70130
rect 665320 70074 665388 70130
rect 665444 70074 665512 70130
rect 665568 70074 665636 70130
rect 665692 70074 665760 70130
rect 665816 70074 665884 70130
rect 665940 70074 666008 70130
rect 666064 70074 666132 70130
rect 666188 70074 666256 70130
rect 666312 70074 666380 70130
rect 666436 70074 666504 70130
rect 666560 70074 666628 70130
rect 666684 70074 666752 70130
rect 666808 70074 666878 70130
rect 664828 69800 666878 70074
rect 667198 70130 669248 70200
rect 667198 70074 667262 70130
rect 667318 70074 667386 70130
rect 667442 70074 667510 70130
rect 667566 70074 667634 70130
rect 667690 70074 667758 70130
rect 667814 70074 667882 70130
rect 667938 70074 668006 70130
rect 668062 70074 668130 70130
rect 668186 70074 668254 70130
rect 668310 70074 668378 70130
rect 668434 70074 668502 70130
rect 668558 70074 668626 70130
rect 668682 70074 668750 70130
rect 668806 70074 668874 70130
rect 668930 70074 668998 70130
rect 669054 70074 669122 70130
rect 669178 70074 669248 70130
rect 667198 69800 669248 70074
rect 669828 70130 671728 70200
rect 669828 70074 669866 70130
rect 669922 70074 669990 70130
rect 670046 70074 670114 70130
rect 670170 70074 670238 70130
rect 670294 70074 670362 70130
rect 670418 70074 670486 70130
rect 670542 70074 670610 70130
rect 670666 70074 670734 70130
rect 670790 70074 670858 70130
rect 670914 70074 670982 70130
rect 671038 70074 671106 70130
rect 671162 70074 671230 70130
rect 671286 70074 671354 70130
rect 671410 70074 671478 70130
rect 671534 70074 671602 70130
rect 671658 70074 671728 70130
rect 669828 69800 671728 70074
<< via2 >>
rect 381342 949870 381398 949926
rect 381466 949870 381522 949926
rect 381590 949870 381646 949926
rect 381714 949870 381770 949926
rect 381838 949870 381894 949926
rect 381962 949870 382018 949926
rect 382086 949870 382142 949926
rect 382210 949870 382266 949926
rect 382334 949870 382390 949926
rect 382458 949870 382514 949926
rect 382582 949870 382638 949926
rect 382706 949870 382762 949926
rect 382830 949870 382886 949926
rect 382954 949870 383010 949926
rect 383078 949870 383134 949926
rect 383822 949870 383878 949926
rect 383946 949870 384002 949926
rect 384070 949870 384126 949926
rect 384194 949870 384250 949926
rect 384318 949870 384374 949926
rect 384442 949870 384498 949926
rect 384566 949870 384622 949926
rect 384690 949870 384746 949926
rect 384814 949870 384870 949926
rect 384938 949870 384994 949926
rect 385062 949870 385118 949926
rect 385186 949870 385242 949926
rect 385310 949870 385366 949926
rect 385434 949870 385490 949926
rect 385558 949870 385614 949926
rect 385682 949870 385738 949926
rect 386192 949870 386248 949926
rect 386316 949870 386372 949926
rect 386440 949870 386496 949926
rect 386564 949870 386620 949926
rect 386688 949870 386744 949926
rect 386812 949870 386868 949926
rect 386936 949870 386992 949926
rect 387060 949870 387116 949926
rect 387184 949870 387240 949926
rect 387308 949870 387364 949926
rect 387432 949870 387488 949926
rect 387556 949870 387612 949926
rect 387680 949870 387736 949926
rect 387804 949870 387860 949926
rect 387928 949870 387984 949926
rect 388052 949870 388108 949926
rect 388892 949870 388948 949926
rect 389016 949870 389072 949926
rect 389140 949870 389196 949926
rect 389264 949870 389320 949926
rect 389388 949870 389444 949926
rect 389512 949870 389568 949926
rect 389636 949870 389692 949926
rect 389760 949870 389816 949926
rect 389884 949870 389940 949926
rect 390008 949870 390064 949926
rect 390132 949870 390188 949926
rect 390256 949870 390312 949926
rect 390380 949870 390436 949926
rect 390504 949870 390560 949926
rect 390628 949870 390684 949926
rect 390752 949870 390808 949926
rect 391262 949870 391318 949926
rect 391386 949870 391442 949926
rect 391510 949870 391566 949926
rect 391634 949870 391690 949926
rect 391758 949870 391814 949926
rect 391882 949870 391938 949926
rect 392006 949870 392062 949926
rect 392130 949870 392186 949926
rect 392254 949870 392310 949926
rect 392378 949870 392434 949926
rect 392502 949870 392558 949926
rect 392626 949870 392682 949926
rect 392750 949870 392806 949926
rect 392874 949870 392930 949926
rect 392998 949870 393054 949926
rect 393122 949870 393178 949926
rect 393866 949870 393922 949926
rect 393990 949870 394046 949926
rect 394114 949870 394170 949926
rect 394238 949870 394294 949926
rect 394362 949870 394418 949926
rect 394486 949870 394542 949926
rect 394610 949870 394666 949926
rect 394734 949870 394790 949926
rect 394858 949870 394914 949926
rect 394982 949870 395038 949926
rect 395106 949870 395162 949926
rect 395230 949870 395286 949926
rect 395354 949870 395410 949926
rect 395478 949870 395534 949926
rect 395602 949870 395658 949926
rect 601342 949870 601398 949926
rect 601466 949870 601522 949926
rect 601590 949870 601646 949926
rect 601714 949870 601770 949926
rect 601838 949870 601894 949926
rect 601962 949870 602018 949926
rect 602086 949870 602142 949926
rect 602210 949870 602266 949926
rect 602334 949870 602390 949926
rect 602458 949870 602514 949926
rect 602582 949870 602638 949926
rect 602706 949870 602762 949926
rect 602830 949870 602886 949926
rect 602954 949870 603010 949926
rect 603078 949870 603134 949926
rect 603822 949870 603878 949926
rect 603946 949870 604002 949926
rect 604070 949870 604126 949926
rect 604194 949870 604250 949926
rect 604318 949870 604374 949926
rect 604442 949870 604498 949926
rect 604566 949870 604622 949926
rect 604690 949870 604746 949926
rect 604814 949870 604870 949926
rect 604938 949870 604994 949926
rect 605062 949870 605118 949926
rect 605186 949870 605242 949926
rect 605310 949870 605366 949926
rect 605434 949870 605490 949926
rect 605558 949870 605614 949926
rect 605682 949870 605738 949926
rect 606192 949870 606248 949926
rect 606316 949870 606372 949926
rect 606440 949870 606496 949926
rect 606564 949870 606620 949926
rect 606688 949870 606744 949926
rect 606812 949870 606868 949926
rect 606936 949870 606992 949926
rect 607060 949870 607116 949926
rect 607184 949870 607240 949926
rect 607308 949870 607364 949926
rect 607432 949870 607488 949926
rect 607556 949870 607612 949926
rect 607680 949870 607736 949926
rect 607804 949870 607860 949926
rect 607928 949870 607984 949926
rect 608052 949870 608108 949926
rect 608892 949870 608948 949926
rect 609016 949870 609072 949926
rect 609140 949870 609196 949926
rect 609264 949870 609320 949926
rect 609388 949870 609444 949926
rect 609512 949870 609568 949926
rect 609636 949870 609692 949926
rect 609760 949870 609816 949926
rect 609884 949870 609940 949926
rect 610008 949870 610064 949926
rect 610132 949870 610188 949926
rect 610256 949870 610312 949926
rect 610380 949870 610436 949926
rect 610504 949870 610560 949926
rect 610628 949870 610684 949926
rect 610752 949870 610808 949926
rect 611262 949870 611318 949926
rect 611386 949870 611442 949926
rect 611510 949870 611566 949926
rect 611634 949870 611690 949926
rect 611758 949870 611814 949926
rect 611882 949870 611938 949926
rect 612006 949870 612062 949926
rect 612130 949870 612186 949926
rect 612254 949870 612310 949926
rect 612378 949870 612434 949926
rect 612502 949870 612558 949926
rect 612626 949870 612682 949926
rect 612750 949870 612806 949926
rect 612874 949870 612930 949926
rect 612998 949870 613054 949926
rect 613122 949870 613178 949926
rect 613866 949870 613922 949926
rect 613990 949870 614046 949926
rect 614114 949870 614170 949926
rect 614238 949870 614294 949926
rect 614362 949870 614418 949926
rect 614486 949870 614542 949926
rect 614610 949870 614666 949926
rect 614734 949870 614790 949926
rect 614858 949870 614914 949926
rect 614982 949870 615038 949926
rect 615106 949870 615162 949926
rect 615230 949870 615286 949926
rect 615354 949870 615410 949926
rect 615478 949870 615534 949926
rect 615602 949870 615658 949926
rect 70074 884602 70130 884658
rect 70074 884478 70130 884534
rect 70074 884354 70130 884410
rect 70074 884230 70130 884286
rect 70074 884106 70130 884162
rect 70074 883982 70130 884038
rect 70074 883858 70130 883914
rect 70074 883734 70130 883790
rect 70074 883610 70130 883666
rect 70074 883486 70130 883542
rect 70074 883362 70130 883418
rect 70074 883238 70130 883294
rect 70074 883114 70130 883170
rect 70074 882990 70130 883046
rect 70074 882866 70130 882922
rect 707870 883602 707926 883658
rect 707870 883478 707926 883534
rect 707870 883354 707926 883410
rect 707870 883230 707926 883286
rect 707870 883106 707926 883162
rect 707870 882982 707926 883038
rect 707870 882858 707926 882914
rect 707870 882734 707926 882790
rect 707870 882610 707926 882666
rect 707870 882486 707926 882542
rect 707870 882362 707926 882418
rect 70074 882128 70130 882184
rect 70074 882004 70130 882060
rect 70074 881880 70130 881936
rect 707870 882238 707926 882294
rect 707870 882114 707926 882170
rect 707870 881990 707926 882046
rect 707870 881866 707926 881922
rect 70074 881756 70130 881812
rect 70074 881632 70130 881688
rect 70074 881508 70130 881564
rect 70074 881384 70130 881440
rect 70074 881260 70130 881316
rect 70074 881136 70130 881192
rect 70074 881012 70130 881068
rect 70074 880888 70130 880944
rect 70074 880764 70130 880820
rect 70074 880640 70130 880696
rect 70074 880516 70130 880572
rect 70074 880392 70130 880448
rect 70074 880268 70130 880324
rect 707870 881122 707926 881178
rect 707870 880998 707926 881054
rect 707870 880874 707926 880930
rect 707870 880750 707926 880806
rect 707870 880626 707926 880682
rect 707870 880502 707926 880558
rect 707870 880378 707926 880434
rect 707870 880254 707926 880310
rect 707870 880130 707926 880186
rect 707870 880006 707926 880062
rect 707870 879882 707926 879938
rect 70074 879758 70130 879814
rect 70074 879634 70130 879690
rect 70074 879510 70130 879566
rect 70074 879386 70130 879442
rect 70074 879262 70130 879318
rect 707870 879758 707926 879814
rect 707870 879634 707926 879690
rect 707870 879510 707926 879566
rect 707870 879386 707926 879442
rect 707870 879262 707926 879318
rect 70074 879138 70130 879194
rect 70074 879014 70130 879070
rect 70074 878890 70130 878946
rect 70074 878766 70130 878822
rect 70074 878642 70130 878698
rect 70074 878518 70130 878574
rect 70074 878394 70130 878450
rect 70074 878270 70130 878326
rect 70074 878146 70130 878202
rect 70074 878022 70130 878078
rect 70074 877898 70130 877954
rect 707870 878752 707926 878808
rect 707870 878628 707926 878684
rect 707870 878504 707926 878560
rect 707870 878380 707926 878436
rect 707870 878256 707926 878312
rect 707870 878132 707926 878188
rect 707870 878008 707926 878064
rect 707870 877884 707926 877940
rect 707870 877760 707926 877816
rect 707870 877636 707926 877692
rect 707870 877512 707926 877568
rect 707870 877388 707926 877444
rect 707870 877264 707926 877320
rect 70074 877052 70130 877108
rect 70074 876928 70130 876984
rect 70074 876804 70130 876860
rect 707870 877140 707926 877196
rect 707870 877016 707926 877072
rect 707870 876892 707926 876948
rect 70074 876680 70130 876736
rect 70074 876556 70130 876612
rect 70074 876432 70130 876488
rect 70074 876308 70130 876364
rect 70074 876184 70130 876240
rect 70074 876060 70130 876116
rect 70074 875936 70130 875992
rect 70074 875812 70130 875868
rect 70074 875688 70130 875744
rect 70074 875564 70130 875620
rect 70074 875440 70130 875496
rect 70074 875316 70130 875372
rect 70074 875192 70130 875248
rect 707870 876046 707926 876102
rect 707870 875922 707926 875978
rect 707870 875798 707926 875854
rect 707870 875674 707926 875730
rect 707870 875550 707926 875606
rect 707870 875426 707926 875482
rect 707870 875302 707926 875358
rect 707870 875178 707926 875234
rect 707870 875054 707926 875110
rect 707870 874930 707926 874986
rect 707870 874806 707926 874862
rect 70074 874682 70130 874738
rect 70074 874558 70130 874614
rect 70074 874434 70130 874490
rect 70074 874310 70130 874366
rect 70074 874186 70130 874242
rect 707870 874682 707926 874738
rect 707870 874558 707926 874614
rect 707870 874434 707926 874490
rect 707870 874310 707926 874366
rect 707870 874186 707926 874242
rect 70074 874062 70130 874118
rect 70074 873938 70130 873994
rect 70074 873814 70130 873870
rect 70074 873690 70130 873746
rect 70074 873566 70130 873622
rect 70074 873442 70130 873498
rect 70074 873318 70130 873374
rect 70074 873194 70130 873250
rect 70074 873070 70130 873126
rect 70074 872946 70130 873002
rect 70074 872822 70130 872878
rect 707870 873676 707926 873732
rect 707870 873552 707926 873608
rect 707870 873428 707926 873484
rect 707870 873304 707926 873360
rect 707870 873180 707926 873236
rect 707870 873056 707926 873112
rect 707870 872932 707926 872988
rect 707870 872808 707926 872864
rect 707870 872684 707926 872740
rect 707870 872560 707926 872616
rect 707870 872436 707926 872492
rect 707870 872312 707926 872368
rect 707870 872188 707926 872244
rect 70074 872078 70130 872134
rect 70074 871954 70130 872010
rect 70074 871830 70130 871886
rect 70074 871706 70130 871762
rect 707870 872064 707926 872120
rect 707870 871940 707926 871996
rect 707870 871816 707926 871872
rect 70074 871582 70130 871638
rect 70074 871458 70130 871514
rect 70074 871334 70130 871390
rect 70074 871210 70130 871266
rect 70074 871086 70130 871142
rect 70074 870962 70130 871018
rect 70074 870838 70130 870894
rect 70074 870714 70130 870770
rect 70074 870590 70130 870646
rect 70074 870466 70130 870522
rect 70074 870342 70130 870398
rect 707870 871078 707926 871134
rect 707870 870954 707926 871010
rect 707870 870830 707926 870886
rect 707870 870706 707926 870762
rect 707870 870582 707926 870638
rect 707870 870458 707926 870514
rect 707870 870334 707926 870390
rect 707870 870210 707926 870266
rect 707870 870086 707926 870142
rect 707870 869962 707926 870018
rect 707870 869838 707926 869894
rect 707870 869714 707926 869770
rect 707870 869590 707926 869646
rect 707870 869466 707926 869522
rect 707870 869342 707926 869398
rect 70074 843602 70130 843658
rect 70074 843478 70130 843534
rect 70074 843354 70130 843410
rect 70074 843230 70130 843286
rect 70074 843106 70130 843162
rect 70074 842982 70130 843038
rect 70074 842858 70130 842914
rect 70074 842734 70130 842790
rect 70074 842610 70130 842666
rect 70074 842486 70130 842542
rect 70074 842362 70130 842418
rect 70074 842238 70130 842294
rect 70074 842114 70130 842170
rect 70074 841990 70130 842046
rect 70074 841866 70130 841922
rect 70074 841128 70130 841184
rect 70074 841004 70130 841060
rect 70074 840880 70130 840936
rect 70074 840756 70130 840812
rect 70074 840632 70130 840688
rect 70074 840508 70130 840564
rect 70074 840384 70130 840440
rect 70074 840260 70130 840316
rect 70074 840136 70130 840192
rect 70074 840012 70130 840068
rect 70074 839888 70130 839944
rect 70074 839764 70130 839820
rect 70074 839640 70130 839696
rect 70074 839516 70130 839572
rect 70074 839392 70130 839448
rect 70074 839268 70130 839324
rect 70074 838758 70130 838814
rect 70074 838634 70130 838690
rect 70074 838510 70130 838566
rect 70074 838386 70130 838442
rect 70074 838262 70130 838318
rect 70074 838138 70130 838194
rect 70074 838014 70130 838070
rect 70074 837890 70130 837946
rect 70074 837766 70130 837822
rect 70074 837642 70130 837698
rect 70074 837518 70130 837574
rect 70074 837394 70130 837450
rect 70074 837270 70130 837326
rect 70074 837146 70130 837202
rect 70074 837022 70130 837078
rect 70074 836898 70130 836954
rect 70074 836052 70130 836108
rect 70074 835928 70130 835984
rect 70074 835804 70130 835860
rect 70074 835680 70130 835736
rect 70074 835556 70130 835612
rect 70074 835432 70130 835488
rect 70074 835308 70130 835364
rect 70074 835184 70130 835240
rect 70074 835060 70130 835116
rect 70074 834936 70130 834992
rect 70074 834812 70130 834868
rect 70074 834688 70130 834744
rect 70074 834564 70130 834620
rect 70074 834440 70130 834496
rect 70074 834316 70130 834372
rect 70074 834192 70130 834248
rect 70074 833682 70130 833738
rect 70074 833558 70130 833614
rect 70074 833434 70130 833490
rect 70074 833310 70130 833366
rect 70074 833186 70130 833242
rect 70074 833062 70130 833118
rect 70074 832938 70130 832994
rect 70074 832814 70130 832870
rect 70074 832690 70130 832746
rect 70074 832566 70130 832622
rect 70074 832442 70130 832498
rect 70074 832318 70130 832374
rect 70074 832194 70130 832250
rect 70074 832070 70130 832126
rect 70074 831946 70130 832002
rect 70074 831822 70130 831878
rect 70074 831078 70130 831134
rect 70074 830954 70130 831010
rect 70074 830830 70130 830886
rect 70074 830706 70130 830762
rect 70074 830582 70130 830638
rect 70074 830458 70130 830514
rect 70074 830334 70130 830390
rect 70074 830210 70130 830266
rect 70074 830086 70130 830142
rect 70074 829962 70130 830018
rect 70074 829838 70130 829894
rect 70074 829714 70130 829770
rect 70074 829590 70130 829646
rect 70074 829466 70130 829522
rect 70074 829342 70130 829398
rect 70074 802602 70130 802658
rect 70074 802478 70130 802534
rect 70074 802354 70130 802410
rect 70074 802230 70130 802286
rect 70074 802106 70130 802162
rect 70074 801982 70130 802038
rect 70074 801858 70130 801914
rect 70074 801734 70130 801790
rect 70074 801610 70130 801666
rect 70074 801486 70130 801542
rect 70074 801362 70130 801418
rect 70074 801238 70130 801294
rect 70074 801114 70130 801170
rect 70074 800990 70130 801046
rect 70074 800866 70130 800922
rect 70074 800128 70130 800184
rect 70074 800004 70130 800060
rect 70074 799880 70130 799936
rect 70074 799756 70130 799812
rect 70074 799632 70130 799688
rect 70074 799508 70130 799564
rect 70074 799384 70130 799440
rect 70074 799260 70130 799316
rect 70074 799136 70130 799192
rect 70074 799012 70130 799068
rect 70074 798888 70130 798944
rect 70074 798764 70130 798820
rect 70074 798640 70130 798696
rect 70074 798516 70130 798572
rect 70074 798392 70130 798448
rect 70074 798268 70130 798324
rect 70074 797758 70130 797814
rect 70074 797634 70130 797690
rect 70074 797510 70130 797566
rect 70074 797386 70130 797442
rect 70074 797262 70130 797318
rect 70074 797138 70130 797194
rect 70074 797014 70130 797070
rect 70074 796890 70130 796946
rect 70074 796766 70130 796822
rect 70074 796642 70130 796698
rect 70074 796518 70130 796574
rect 70074 796394 70130 796450
rect 70074 796270 70130 796326
rect 70074 796146 70130 796202
rect 70074 796022 70130 796078
rect 70074 795898 70130 795954
rect 707870 797602 707926 797658
rect 707870 797478 707926 797534
rect 707870 797354 707926 797410
rect 707870 797230 707926 797286
rect 707870 797106 707926 797162
rect 707870 796982 707926 797038
rect 707870 796858 707926 796914
rect 707870 796734 707926 796790
rect 707870 796610 707926 796666
rect 707870 796486 707926 796542
rect 707870 796362 707926 796418
rect 707870 796238 707926 796294
rect 707870 796114 707926 796170
rect 707870 795990 707926 796046
rect 707870 795866 707926 795922
rect 70074 795052 70130 795108
rect 70074 794928 70130 794984
rect 70074 794804 70130 794860
rect 70074 794680 70130 794736
rect 70074 794556 70130 794612
rect 70074 794432 70130 794488
rect 70074 794308 70130 794364
rect 70074 794184 70130 794240
rect 70074 794060 70130 794116
rect 70074 793936 70130 793992
rect 70074 793812 70130 793868
rect 70074 793688 70130 793744
rect 70074 793564 70130 793620
rect 70074 793440 70130 793496
rect 70074 793316 70130 793372
rect 70074 793192 70130 793248
rect 707870 795122 707926 795178
rect 707870 794998 707926 795054
rect 707870 794874 707926 794930
rect 707870 794750 707926 794806
rect 707870 794626 707926 794682
rect 707870 794502 707926 794558
rect 707870 794378 707926 794434
rect 707870 794254 707926 794310
rect 707870 794130 707926 794186
rect 707870 794006 707926 794062
rect 707870 793882 707926 793938
rect 707870 793758 707926 793814
rect 707870 793634 707926 793690
rect 707870 793510 707926 793566
rect 707870 793386 707926 793442
rect 707870 793262 707926 793318
rect 70074 792682 70130 792738
rect 70074 792558 70130 792614
rect 70074 792434 70130 792490
rect 70074 792310 70130 792366
rect 70074 792186 70130 792242
rect 70074 792062 70130 792118
rect 70074 791938 70130 791994
rect 70074 791814 70130 791870
rect 70074 791690 70130 791746
rect 70074 791566 70130 791622
rect 70074 791442 70130 791498
rect 70074 791318 70130 791374
rect 70074 791194 70130 791250
rect 70074 791070 70130 791126
rect 70074 790946 70130 791002
rect 70074 790822 70130 790878
rect 707870 792752 707926 792808
rect 707870 792628 707926 792684
rect 707870 792504 707926 792560
rect 707870 792380 707926 792436
rect 707870 792256 707926 792312
rect 707870 792132 707926 792188
rect 707870 792008 707926 792064
rect 707870 791884 707926 791940
rect 707870 791760 707926 791816
rect 707870 791636 707926 791692
rect 707870 791512 707926 791568
rect 707870 791388 707926 791444
rect 707870 791264 707926 791320
rect 707870 791140 707926 791196
rect 707870 791016 707926 791072
rect 707870 790892 707926 790948
rect 70074 790078 70130 790134
rect 70074 789954 70130 790010
rect 70074 789830 70130 789886
rect 70074 789706 70130 789762
rect 70074 789582 70130 789638
rect 70074 789458 70130 789514
rect 70074 789334 70130 789390
rect 70074 789210 70130 789266
rect 70074 789086 70130 789142
rect 70074 788962 70130 789018
rect 70074 788838 70130 788894
rect 70074 788714 70130 788770
rect 70074 788590 70130 788646
rect 70074 788466 70130 788522
rect 70074 788342 70130 788398
rect 707870 790046 707926 790102
rect 707870 789922 707926 789978
rect 707870 789798 707926 789854
rect 707870 789674 707926 789730
rect 707870 789550 707926 789606
rect 707870 789426 707926 789482
rect 707870 789302 707926 789358
rect 707870 789178 707926 789234
rect 707870 789054 707926 789110
rect 707870 788930 707926 788986
rect 707870 788806 707926 788862
rect 707870 788682 707926 788738
rect 707870 788558 707926 788614
rect 707870 788434 707926 788490
rect 707870 788310 707926 788366
rect 707870 788186 707926 788242
rect 707870 787676 707926 787732
rect 707870 787552 707926 787608
rect 707870 787428 707926 787484
rect 707870 787304 707926 787360
rect 707870 787180 707926 787236
rect 707870 787056 707926 787112
rect 707870 786932 707926 786988
rect 707870 786808 707926 786864
rect 707870 786684 707926 786740
rect 707870 786560 707926 786616
rect 707870 786436 707926 786492
rect 707870 786312 707926 786368
rect 707870 786188 707926 786244
rect 707870 786064 707926 786120
rect 707870 785940 707926 785996
rect 707870 785816 707926 785872
rect 707870 785078 707926 785134
rect 707870 784954 707926 785010
rect 707870 784830 707926 784886
rect 707870 784706 707926 784762
rect 707870 784582 707926 784638
rect 707870 784458 707926 784514
rect 707870 784334 707926 784390
rect 707870 784210 707926 784266
rect 707870 784086 707926 784142
rect 707870 783962 707926 784018
rect 707870 783838 707926 783894
rect 707870 783714 707926 783770
rect 707870 783590 707926 783646
rect 707870 783466 707926 783522
rect 707870 783342 707926 783398
rect 707870 496602 707926 496658
rect 707870 496478 707926 496534
rect 707870 496354 707926 496410
rect 707870 496230 707926 496286
rect 707870 496106 707926 496162
rect 707870 495982 707926 496038
rect 707870 495858 707926 495914
rect 707870 495734 707926 495790
rect 707870 495610 707926 495666
rect 707870 495486 707926 495542
rect 707870 495362 707926 495418
rect 707870 495238 707926 495294
rect 707870 495114 707926 495170
rect 707870 494990 707926 495046
rect 707870 494866 707926 494922
rect 707870 494122 707926 494178
rect 707870 493998 707926 494054
rect 707870 493874 707926 493930
rect 707870 493750 707926 493806
rect 707870 493626 707926 493682
rect 707870 493502 707926 493558
rect 707870 493378 707926 493434
rect 707870 493254 707926 493310
rect 707870 493130 707926 493186
rect 707870 493006 707926 493062
rect 707870 492882 707926 492938
rect 707870 492758 707926 492814
rect 707870 492634 707926 492690
rect 707870 492510 707926 492566
rect 707870 492386 707926 492442
rect 707870 492262 707926 492318
rect 707870 491752 707926 491808
rect 707870 491628 707926 491684
rect 707870 491504 707926 491560
rect 707870 491380 707926 491436
rect 707870 491256 707926 491312
rect 707870 491132 707926 491188
rect 707870 491008 707926 491064
rect 707870 490884 707926 490940
rect 707870 490760 707926 490816
rect 707870 490636 707926 490692
rect 707870 490512 707926 490568
rect 707870 490388 707926 490444
rect 707870 490264 707926 490320
rect 707870 490140 707926 490196
rect 707870 490016 707926 490072
rect 707870 489892 707926 489948
rect 707870 489046 707926 489102
rect 707870 488922 707926 488978
rect 707870 488798 707926 488854
rect 707870 488674 707926 488730
rect 707870 488550 707926 488606
rect 707870 488426 707926 488482
rect 707870 488302 707926 488358
rect 707870 488178 707926 488234
rect 707870 488054 707926 488110
rect 707870 487930 707926 487986
rect 707870 487806 707926 487862
rect 707870 487682 707926 487738
rect 707870 487558 707926 487614
rect 707870 487434 707926 487490
rect 707870 487310 707926 487366
rect 707870 487186 707926 487242
rect 707870 486676 707926 486732
rect 707870 486552 707926 486608
rect 707870 486428 707926 486484
rect 707870 486304 707926 486360
rect 707870 486180 707926 486236
rect 707870 486056 707926 486112
rect 707870 485932 707926 485988
rect 707870 485808 707926 485864
rect 707870 485684 707926 485740
rect 707870 485560 707926 485616
rect 707870 485436 707926 485492
rect 707870 485312 707926 485368
rect 707870 485188 707926 485244
rect 707870 485064 707926 485120
rect 707870 484940 707926 484996
rect 707870 484816 707926 484872
rect 707870 484078 707926 484134
rect 707870 483954 707926 484010
rect 707870 483830 707926 483886
rect 707870 483706 707926 483762
rect 707870 483582 707926 483638
rect 707870 483458 707926 483514
rect 707870 483334 707926 483390
rect 707870 483210 707926 483266
rect 707870 483086 707926 483142
rect 707870 482962 707926 483018
rect 707870 482838 707926 482894
rect 707870 482714 707926 482770
rect 707870 482590 707926 482646
rect 707870 482466 707926 482522
rect 707870 482342 707926 482398
rect 70074 474602 70130 474658
rect 70074 474478 70130 474534
rect 70074 474354 70130 474410
rect 70074 474230 70130 474286
rect 70074 474106 70130 474162
rect 70074 473982 70130 474038
rect 70074 473858 70130 473914
rect 70074 473734 70130 473790
rect 70074 473610 70130 473666
rect 70074 473486 70130 473542
rect 70074 473362 70130 473418
rect 70074 473238 70130 473294
rect 70074 473114 70130 473170
rect 70074 472990 70130 473046
rect 70074 472866 70130 472922
rect 70074 472128 70130 472184
rect 70074 472004 70130 472060
rect 70074 471880 70130 471936
rect 70074 471756 70130 471812
rect 70074 471632 70130 471688
rect 70074 471508 70130 471564
rect 70074 471384 70130 471440
rect 70074 471260 70130 471316
rect 70074 471136 70130 471192
rect 70074 471012 70130 471068
rect 70074 470888 70130 470944
rect 70074 470764 70130 470820
rect 70074 470640 70130 470696
rect 70074 470516 70130 470572
rect 70074 470392 70130 470448
rect 70074 470268 70130 470324
rect 70074 469758 70130 469814
rect 70074 469634 70130 469690
rect 70074 469510 70130 469566
rect 70074 469386 70130 469442
rect 70074 469262 70130 469318
rect 70074 469138 70130 469194
rect 70074 469014 70130 469070
rect 70074 468890 70130 468946
rect 70074 468766 70130 468822
rect 70074 468642 70130 468698
rect 70074 468518 70130 468574
rect 70074 468394 70130 468450
rect 70074 468270 70130 468326
rect 70074 468146 70130 468202
rect 70074 468022 70130 468078
rect 70074 467898 70130 467954
rect 70074 467052 70130 467108
rect 70074 466928 70130 466984
rect 70074 466804 70130 466860
rect 70074 466680 70130 466736
rect 70074 466556 70130 466612
rect 70074 466432 70130 466488
rect 70074 466308 70130 466364
rect 70074 466184 70130 466240
rect 70074 466060 70130 466116
rect 70074 465936 70130 465992
rect 70074 465812 70130 465868
rect 70074 465688 70130 465744
rect 70074 465564 70130 465620
rect 70074 465440 70130 465496
rect 70074 465316 70130 465372
rect 70074 465192 70130 465248
rect 70074 464682 70130 464738
rect 70074 464558 70130 464614
rect 70074 464434 70130 464490
rect 70074 464310 70130 464366
rect 70074 464186 70130 464242
rect 70074 464062 70130 464118
rect 70074 463938 70130 463994
rect 70074 463814 70130 463870
rect 70074 463690 70130 463746
rect 70074 463566 70130 463622
rect 70074 463442 70130 463498
rect 70074 463318 70130 463374
rect 70074 463194 70130 463250
rect 70074 463070 70130 463126
rect 70074 462946 70130 463002
rect 70074 462822 70130 462878
rect 70074 462078 70130 462134
rect 70074 461954 70130 462010
rect 70074 461830 70130 461886
rect 70074 461706 70130 461762
rect 70074 461582 70130 461638
rect 70074 461458 70130 461514
rect 70074 461334 70130 461390
rect 70074 461210 70130 461266
rect 70074 461086 70130 461142
rect 70074 460962 70130 461018
rect 70074 460838 70130 460894
rect 70074 460714 70130 460770
rect 70074 460590 70130 460646
rect 70074 460466 70130 460522
rect 70074 460342 70130 460398
rect 707870 453602 707926 453658
rect 707870 453478 707926 453534
rect 707870 453354 707926 453410
rect 707870 453230 707926 453286
rect 707870 453106 707926 453162
rect 707870 452982 707926 453038
rect 707870 452858 707926 452914
rect 707870 452734 707926 452790
rect 707870 452610 707926 452666
rect 707870 452486 707926 452542
rect 707870 452362 707926 452418
rect 707870 452238 707926 452294
rect 707870 452114 707926 452170
rect 707870 451990 707926 452046
rect 707870 451866 707926 451922
rect 707870 451122 707926 451178
rect 707870 450998 707926 451054
rect 707870 450874 707926 450930
rect 707870 450750 707926 450806
rect 707870 450626 707926 450682
rect 707870 450502 707926 450558
rect 707870 450378 707926 450434
rect 707870 450254 707926 450310
rect 707870 450130 707926 450186
rect 707870 450006 707926 450062
rect 707870 449882 707926 449938
rect 707870 449758 707926 449814
rect 707870 449634 707926 449690
rect 707870 449510 707926 449566
rect 707870 449386 707926 449442
rect 707870 449262 707926 449318
rect 707870 448752 707926 448808
rect 707870 448628 707926 448684
rect 707870 448504 707926 448560
rect 707870 448380 707926 448436
rect 707870 448256 707926 448312
rect 707870 448132 707926 448188
rect 707870 448008 707926 448064
rect 707870 447884 707926 447940
rect 707870 447760 707926 447816
rect 707870 447636 707926 447692
rect 707870 447512 707926 447568
rect 707870 447388 707926 447444
rect 707870 447264 707926 447320
rect 707870 447140 707926 447196
rect 707870 447016 707926 447072
rect 707870 446892 707926 446948
rect 707870 446046 707926 446102
rect 707870 445922 707926 445978
rect 707870 445798 707926 445854
rect 707870 445674 707926 445730
rect 707870 445550 707926 445606
rect 707870 445426 707926 445482
rect 707870 445302 707926 445358
rect 707870 445178 707926 445234
rect 707870 445054 707926 445110
rect 707870 444930 707926 444986
rect 707870 444806 707926 444862
rect 707870 444682 707926 444738
rect 707870 444558 707926 444614
rect 707870 444434 707926 444490
rect 707870 444310 707926 444366
rect 707870 444186 707926 444242
rect 707870 443676 707926 443732
rect 707870 443552 707926 443608
rect 707870 443428 707926 443484
rect 707870 443304 707926 443360
rect 707870 443180 707926 443236
rect 707870 443056 707926 443112
rect 707870 442932 707926 442988
rect 707870 442808 707926 442864
rect 707870 442684 707926 442740
rect 707870 442560 707926 442616
rect 707870 442436 707926 442492
rect 707870 442312 707926 442368
rect 707870 442188 707926 442244
rect 707870 442064 707926 442120
rect 707870 441940 707926 441996
rect 707870 441816 707926 441872
rect 707870 441078 707926 441134
rect 707870 440954 707926 441010
rect 707870 440830 707926 440886
rect 707870 440706 707926 440762
rect 707870 440582 707926 440638
rect 707870 440458 707926 440514
rect 707870 440334 707926 440390
rect 707870 440210 707926 440266
rect 707870 440086 707926 440142
rect 707870 439962 707926 440018
rect 707870 439838 707926 439894
rect 707870 439714 707926 439770
rect 707870 439590 707926 439646
rect 707870 439466 707926 439522
rect 707870 439342 707926 439398
rect 70074 433602 70130 433658
rect 70074 433478 70130 433534
rect 70074 433354 70130 433410
rect 70074 433230 70130 433286
rect 70074 433106 70130 433162
rect 70074 432982 70130 433038
rect 70074 432858 70130 432914
rect 70074 432734 70130 432790
rect 70074 432610 70130 432666
rect 70074 432486 70130 432542
rect 70074 432362 70130 432418
rect 70074 432238 70130 432294
rect 70074 432114 70130 432170
rect 70074 431990 70130 432046
rect 70074 431866 70130 431922
rect 70074 431128 70130 431184
rect 70074 431004 70130 431060
rect 70074 430880 70130 430936
rect 70074 430756 70130 430812
rect 70074 430632 70130 430688
rect 70074 430508 70130 430564
rect 70074 430384 70130 430440
rect 70074 430260 70130 430316
rect 70074 430136 70130 430192
rect 70074 430012 70130 430068
rect 70074 429888 70130 429944
rect 70074 429764 70130 429820
rect 70074 429640 70130 429696
rect 70074 429516 70130 429572
rect 70074 429392 70130 429448
rect 70074 429268 70130 429324
rect 70074 428758 70130 428814
rect 70074 428634 70130 428690
rect 70074 428510 70130 428566
rect 70074 428386 70130 428442
rect 70074 428262 70130 428318
rect 70074 428138 70130 428194
rect 70074 428014 70130 428070
rect 70074 427890 70130 427946
rect 70074 427766 70130 427822
rect 70074 427642 70130 427698
rect 70074 427518 70130 427574
rect 70074 427394 70130 427450
rect 70074 427270 70130 427326
rect 70074 427146 70130 427202
rect 70074 427022 70130 427078
rect 70074 426898 70130 426954
rect 70074 426052 70130 426108
rect 70074 425928 70130 425984
rect 70074 425804 70130 425860
rect 70074 425680 70130 425736
rect 70074 425556 70130 425612
rect 70074 425432 70130 425488
rect 70074 425308 70130 425364
rect 70074 425184 70130 425240
rect 70074 425060 70130 425116
rect 70074 424936 70130 424992
rect 70074 424812 70130 424868
rect 70074 424688 70130 424744
rect 70074 424564 70130 424620
rect 70074 424440 70130 424496
rect 70074 424316 70130 424372
rect 70074 424192 70130 424248
rect 70074 423682 70130 423738
rect 70074 423558 70130 423614
rect 70074 423434 70130 423490
rect 70074 423310 70130 423366
rect 70074 423186 70130 423242
rect 70074 423062 70130 423118
rect 70074 422938 70130 422994
rect 70074 422814 70130 422870
rect 70074 422690 70130 422746
rect 70074 422566 70130 422622
rect 70074 422442 70130 422498
rect 70074 422318 70130 422374
rect 70074 422194 70130 422250
rect 70074 422070 70130 422126
rect 70074 421946 70130 422002
rect 70074 421822 70130 421878
rect 70074 421078 70130 421134
rect 70074 420954 70130 421010
rect 70074 420830 70130 420886
rect 70074 420706 70130 420762
rect 70074 420582 70130 420638
rect 70074 420458 70130 420514
rect 70074 420334 70130 420390
rect 70074 420210 70130 420266
rect 70074 420086 70130 420142
rect 70074 419962 70130 420018
rect 70074 419838 70130 419894
rect 70074 419714 70130 419770
rect 70074 419590 70130 419646
rect 70074 419466 70130 419522
rect 70074 419342 70130 419398
rect 707870 410602 707926 410658
rect 707870 410478 707926 410534
rect 707870 410354 707926 410410
rect 707870 410230 707926 410286
rect 707870 410106 707926 410162
rect 707870 409982 707926 410038
rect 707870 409858 707926 409914
rect 707870 409734 707926 409790
rect 707870 409610 707926 409666
rect 707870 409486 707926 409542
rect 707870 409362 707926 409418
rect 707870 409238 707926 409294
rect 707870 409114 707926 409170
rect 707870 408990 707926 409046
rect 707870 408866 707926 408922
rect 707870 408122 707926 408178
rect 707870 407998 707926 408054
rect 707870 407874 707926 407930
rect 707870 407750 707926 407806
rect 707870 407626 707926 407682
rect 707870 407502 707926 407558
rect 707870 407378 707926 407434
rect 707870 407254 707926 407310
rect 707870 407130 707926 407186
rect 707870 407006 707926 407062
rect 707870 406882 707926 406938
rect 707870 406758 707926 406814
rect 707870 406634 707926 406690
rect 707870 406510 707926 406566
rect 707870 406386 707926 406442
rect 707870 406262 707926 406318
rect 707870 405752 707926 405808
rect 707870 405628 707926 405684
rect 707870 405504 707926 405560
rect 707870 405380 707926 405436
rect 707870 405256 707926 405312
rect 707870 405132 707926 405188
rect 707870 405008 707926 405064
rect 707870 404884 707926 404940
rect 707870 404760 707926 404816
rect 707870 404636 707926 404692
rect 707870 404512 707926 404568
rect 707870 404388 707926 404444
rect 707870 404264 707926 404320
rect 707870 404140 707926 404196
rect 707870 404016 707926 404072
rect 707870 403892 707926 403948
rect 707870 403046 707926 403102
rect 707870 402922 707926 402978
rect 707870 402798 707926 402854
rect 707870 402674 707926 402730
rect 707870 402550 707926 402606
rect 707870 402426 707926 402482
rect 707870 402302 707926 402358
rect 707870 402178 707926 402234
rect 707870 402054 707926 402110
rect 707870 401930 707926 401986
rect 707870 401806 707926 401862
rect 707870 401682 707926 401738
rect 707870 401558 707926 401614
rect 707870 401434 707926 401490
rect 707870 401310 707926 401366
rect 707870 401186 707926 401242
rect 707870 400676 707926 400732
rect 707870 400552 707926 400608
rect 707870 400428 707926 400484
rect 707870 400304 707926 400360
rect 707870 400180 707926 400236
rect 707870 400056 707926 400112
rect 707870 399932 707926 399988
rect 707870 399808 707926 399864
rect 707870 399684 707926 399740
rect 707870 399560 707926 399616
rect 707870 399436 707926 399492
rect 707870 399312 707926 399368
rect 707870 399188 707926 399244
rect 707870 399064 707926 399120
rect 707870 398940 707926 398996
rect 707870 398816 707926 398872
rect 707870 398078 707926 398134
rect 707870 397954 707926 398010
rect 707870 397830 707926 397886
rect 707870 397706 707926 397762
rect 707870 397582 707926 397638
rect 707870 397458 707926 397514
rect 707870 397334 707926 397390
rect 707870 397210 707926 397266
rect 707870 397086 707926 397142
rect 707870 396962 707926 397018
rect 707870 396838 707926 396894
rect 707870 396714 707926 396770
rect 707870 396590 707926 396646
rect 707870 396466 707926 396522
rect 707870 396342 707926 396398
rect 70074 146602 70130 146658
rect 70074 146478 70130 146534
rect 70074 146354 70130 146410
rect 70074 146230 70130 146286
rect 70074 146106 70130 146162
rect 70074 145982 70130 146038
rect 70074 145858 70130 145914
rect 70074 145734 70130 145790
rect 70074 145610 70130 145666
rect 70074 145486 70130 145542
rect 70074 145362 70130 145418
rect 70074 145238 70130 145294
rect 70074 145114 70130 145170
rect 70074 144990 70130 145046
rect 70074 144866 70130 144922
rect 70074 144128 70130 144184
rect 70074 144004 70130 144060
rect 70074 143880 70130 143936
rect 70074 143756 70130 143812
rect 70074 143632 70130 143688
rect 70074 143508 70130 143564
rect 70074 143384 70130 143440
rect 70074 143260 70130 143316
rect 70074 143136 70130 143192
rect 70074 143012 70130 143068
rect 70074 142888 70130 142944
rect 70074 142764 70130 142820
rect 70074 142640 70130 142696
rect 70074 142516 70130 142572
rect 70074 142392 70130 142448
rect 70074 142268 70130 142324
rect 70074 141758 70130 141814
rect 70074 141634 70130 141690
rect 70074 141510 70130 141566
rect 70074 141386 70130 141442
rect 70074 141262 70130 141318
rect 70074 141138 70130 141194
rect 70074 141014 70130 141070
rect 70074 140890 70130 140946
rect 70074 140766 70130 140822
rect 70074 140642 70130 140698
rect 70074 140518 70130 140574
rect 70074 140394 70130 140450
rect 70074 140270 70130 140326
rect 70074 140146 70130 140202
rect 70074 140022 70130 140078
rect 70074 139898 70130 139954
rect 70074 139052 70130 139108
rect 70074 138928 70130 138984
rect 70074 138804 70130 138860
rect 70074 138680 70130 138736
rect 70074 138556 70130 138612
rect 70074 138432 70130 138488
rect 70074 138308 70130 138364
rect 70074 138184 70130 138240
rect 70074 138060 70130 138116
rect 70074 137936 70130 137992
rect 70074 137812 70130 137868
rect 70074 137688 70130 137744
rect 70074 137564 70130 137620
rect 70074 137440 70130 137496
rect 70074 137316 70130 137372
rect 70074 137192 70130 137248
rect 70074 136682 70130 136738
rect 70074 136558 70130 136614
rect 70074 136434 70130 136490
rect 70074 136310 70130 136366
rect 70074 136186 70130 136242
rect 70074 136062 70130 136118
rect 70074 135938 70130 135994
rect 70074 135814 70130 135870
rect 70074 135690 70130 135746
rect 70074 135566 70130 135622
rect 70074 135442 70130 135498
rect 70074 135318 70130 135374
rect 70074 135194 70130 135250
rect 70074 135070 70130 135126
rect 70074 134946 70130 135002
rect 70074 134822 70130 134878
rect 70074 134078 70130 134134
rect 70074 133954 70130 134010
rect 70074 133830 70130 133886
rect 70074 133706 70130 133762
rect 70074 133582 70130 133638
rect 70074 133458 70130 133514
rect 70074 133334 70130 133390
rect 70074 133210 70130 133266
rect 70074 133086 70130 133142
rect 70074 132962 70130 133018
rect 70074 132838 70130 132894
rect 70074 132714 70130 132770
rect 70074 132590 70130 132646
rect 70074 132466 70130 132522
rect 70074 132342 70130 132398
rect 70074 105602 70130 105658
rect 70074 105478 70130 105534
rect 70074 105354 70130 105410
rect 70074 105230 70130 105286
rect 70074 105106 70130 105162
rect 70074 104982 70130 105038
rect 70074 104858 70130 104914
rect 70074 104734 70130 104790
rect 70074 104610 70130 104666
rect 70074 104486 70130 104542
rect 70074 104362 70130 104418
rect 70074 104238 70130 104294
rect 70074 104114 70130 104170
rect 70074 103990 70130 104046
rect 70074 103866 70130 103922
rect 70074 103128 70130 103184
rect 70074 103004 70130 103060
rect 70074 102880 70130 102936
rect 70074 102756 70130 102812
rect 70074 102632 70130 102688
rect 70074 102508 70130 102564
rect 70074 102384 70130 102440
rect 70074 102260 70130 102316
rect 70074 102136 70130 102192
rect 70074 102012 70130 102068
rect 70074 101888 70130 101944
rect 70074 101764 70130 101820
rect 70074 101640 70130 101696
rect 70074 101516 70130 101572
rect 70074 101392 70130 101448
rect 70074 101268 70130 101324
rect 70074 100758 70130 100814
rect 70074 100634 70130 100690
rect 70074 100510 70130 100566
rect 70074 100386 70130 100442
rect 70074 100262 70130 100318
rect 70074 100138 70130 100194
rect 70074 100014 70130 100070
rect 70074 99890 70130 99946
rect 70074 99766 70130 99822
rect 70074 99642 70130 99698
rect 70074 99518 70130 99574
rect 70074 99394 70130 99450
rect 70074 99270 70130 99326
rect 70074 99146 70130 99202
rect 70074 99022 70130 99078
rect 70074 98898 70130 98954
rect 70074 98052 70130 98108
rect 70074 97928 70130 97984
rect 70074 97804 70130 97860
rect 70074 97680 70130 97736
rect 70074 97556 70130 97612
rect 70074 97432 70130 97488
rect 70074 97308 70130 97364
rect 70074 97184 70130 97240
rect 70074 97060 70130 97116
rect 70074 96936 70130 96992
rect 70074 96812 70130 96868
rect 70074 96688 70130 96744
rect 70074 96564 70130 96620
rect 70074 96440 70130 96496
rect 70074 96316 70130 96372
rect 70074 96192 70130 96248
rect 70074 95682 70130 95738
rect 70074 95558 70130 95614
rect 70074 95434 70130 95490
rect 70074 95310 70130 95366
rect 70074 95186 70130 95242
rect 70074 95062 70130 95118
rect 70074 94938 70130 94994
rect 70074 94814 70130 94870
rect 70074 94690 70130 94746
rect 70074 94566 70130 94622
rect 70074 94442 70130 94498
rect 70074 94318 70130 94374
rect 70074 94194 70130 94250
rect 70074 94070 70130 94126
rect 70074 93946 70130 94002
rect 70074 93822 70130 93878
rect 70074 93078 70130 93134
rect 70074 92954 70130 93010
rect 70074 92830 70130 92886
rect 70074 92706 70130 92762
rect 70074 92582 70130 92638
rect 70074 92458 70130 92514
rect 70074 92334 70130 92390
rect 70074 92210 70130 92266
rect 70074 92086 70130 92142
rect 70074 91962 70130 92018
rect 70074 91838 70130 91894
rect 70074 91714 70130 91770
rect 70074 91590 70130 91646
rect 70074 91466 70130 91522
rect 70074 91342 70130 91398
rect 107342 70074 107398 70130
rect 107466 70074 107522 70130
rect 107590 70074 107646 70130
rect 107714 70074 107770 70130
rect 107838 70074 107894 70130
rect 107962 70074 108018 70130
rect 108086 70074 108142 70130
rect 108210 70074 108266 70130
rect 108334 70074 108390 70130
rect 108458 70074 108514 70130
rect 108582 70074 108638 70130
rect 108706 70074 108762 70130
rect 108830 70074 108886 70130
rect 108954 70074 109010 70130
rect 109078 70074 109134 70130
rect 109822 70074 109878 70130
rect 109946 70074 110002 70130
rect 110070 70074 110126 70130
rect 110194 70074 110250 70130
rect 110318 70074 110374 70130
rect 110442 70074 110498 70130
rect 110566 70074 110622 70130
rect 110690 70074 110746 70130
rect 110814 70074 110870 70130
rect 110938 70074 110994 70130
rect 111062 70074 111118 70130
rect 111186 70074 111242 70130
rect 111310 70074 111366 70130
rect 111434 70074 111490 70130
rect 111558 70074 111614 70130
rect 111682 70074 111738 70130
rect 112192 70074 112248 70130
rect 112316 70074 112372 70130
rect 112440 70074 112496 70130
rect 112564 70074 112620 70130
rect 112688 70074 112744 70130
rect 112812 70074 112868 70130
rect 112936 70074 112992 70130
rect 113060 70074 113116 70130
rect 113184 70074 113240 70130
rect 113308 70074 113364 70130
rect 113432 70074 113488 70130
rect 113556 70074 113612 70130
rect 113680 70074 113736 70130
rect 113804 70074 113860 70130
rect 113928 70074 113984 70130
rect 114052 70074 114108 70130
rect 114892 70074 114948 70130
rect 115016 70074 115072 70130
rect 115140 70074 115196 70130
rect 115264 70074 115320 70130
rect 115388 70074 115444 70130
rect 115512 70074 115568 70130
rect 115636 70074 115692 70130
rect 115760 70074 115816 70130
rect 115884 70074 115940 70130
rect 116008 70074 116064 70130
rect 116132 70074 116188 70130
rect 116256 70074 116312 70130
rect 116380 70074 116436 70130
rect 116504 70074 116560 70130
rect 116628 70074 116684 70130
rect 116752 70074 116808 70130
rect 117262 70074 117318 70130
rect 117386 70074 117442 70130
rect 117510 70074 117566 70130
rect 117634 70074 117690 70130
rect 117758 70074 117814 70130
rect 117882 70074 117938 70130
rect 118006 70074 118062 70130
rect 118130 70074 118186 70130
rect 118254 70074 118310 70130
rect 118378 70074 118434 70130
rect 118502 70074 118558 70130
rect 118626 70074 118682 70130
rect 118750 70074 118806 70130
rect 118874 70074 118930 70130
rect 118998 70074 119054 70130
rect 119122 70074 119178 70130
rect 119866 70074 119922 70130
rect 119990 70074 120046 70130
rect 120114 70074 120170 70130
rect 120238 70074 120294 70130
rect 120362 70074 120418 70130
rect 120486 70074 120542 70130
rect 120610 70074 120666 70130
rect 120734 70074 120790 70130
rect 120858 70074 120914 70130
rect 120982 70074 121038 70130
rect 121106 70074 121162 70130
rect 121230 70074 121286 70130
rect 121354 70074 121410 70130
rect 121478 70074 121534 70130
rect 121602 70074 121658 70130
rect 272342 70074 272398 70130
rect 272466 70074 272522 70130
rect 272590 70074 272646 70130
rect 272714 70074 272770 70130
rect 272838 70074 272894 70130
rect 272962 70074 273018 70130
rect 273086 70074 273142 70130
rect 273210 70074 273266 70130
rect 273334 70074 273390 70130
rect 273458 70074 273514 70130
rect 273582 70074 273638 70130
rect 273706 70074 273762 70130
rect 273830 70074 273886 70130
rect 273954 70074 274010 70130
rect 274078 70074 274134 70130
rect 274822 70074 274878 70130
rect 274946 70074 275002 70130
rect 275070 70074 275126 70130
rect 275194 70074 275250 70130
rect 275318 70074 275374 70130
rect 275442 70074 275498 70130
rect 275566 70074 275622 70130
rect 275690 70074 275746 70130
rect 275814 70074 275870 70130
rect 275938 70074 275994 70130
rect 276062 70074 276118 70130
rect 276186 70074 276242 70130
rect 276310 70074 276366 70130
rect 276434 70074 276490 70130
rect 276558 70074 276614 70130
rect 276682 70074 276738 70130
rect 277192 70074 277248 70130
rect 277316 70074 277372 70130
rect 277440 70074 277496 70130
rect 277564 70074 277620 70130
rect 277688 70074 277744 70130
rect 277812 70074 277868 70130
rect 277936 70074 277992 70130
rect 278060 70074 278116 70130
rect 278184 70074 278240 70130
rect 278308 70074 278364 70130
rect 278432 70074 278488 70130
rect 278556 70074 278612 70130
rect 278680 70074 278736 70130
rect 278804 70074 278860 70130
rect 278928 70074 278984 70130
rect 279052 70074 279108 70130
rect 279892 70074 279948 70130
rect 280016 70074 280072 70130
rect 280140 70074 280196 70130
rect 280264 70074 280320 70130
rect 280388 70074 280444 70130
rect 280512 70074 280568 70130
rect 280636 70074 280692 70130
rect 280760 70074 280816 70130
rect 280884 70074 280940 70130
rect 281008 70074 281064 70130
rect 281132 70074 281188 70130
rect 281256 70074 281312 70130
rect 281380 70074 281436 70130
rect 281504 70074 281560 70130
rect 281628 70074 281684 70130
rect 281752 70074 281808 70130
rect 282262 70074 282318 70130
rect 282386 70074 282442 70130
rect 282510 70074 282566 70130
rect 282634 70074 282690 70130
rect 282758 70074 282814 70130
rect 282882 70074 282938 70130
rect 283006 70074 283062 70130
rect 283130 70074 283186 70130
rect 283254 70074 283310 70130
rect 283378 70074 283434 70130
rect 283502 70074 283558 70130
rect 283626 70074 283682 70130
rect 283750 70074 283806 70130
rect 283874 70074 283930 70130
rect 283998 70074 284054 70130
rect 284122 70074 284178 70130
rect 284866 70074 284922 70130
rect 284990 70074 285046 70130
rect 285114 70074 285170 70130
rect 285238 70074 285294 70130
rect 285362 70074 285418 70130
rect 285486 70074 285542 70130
rect 285610 70074 285666 70130
rect 285734 70074 285790 70130
rect 285858 70074 285914 70130
rect 285982 70074 286038 70130
rect 286106 70074 286162 70130
rect 286230 70074 286286 70130
rect 286354 70074 286410 70130
rect 286478 70074 286534 70130
rect 286602 70074 286658 70130
rect 602342 70074 602398 70130
rect 602466 70074 602522 70130
rect 602590 70074 602646 70130
rect 602714 70074 602770 70130
rect 602838 70074 602894 70130
rect 602962 70074 603018 70130
rect 603086 70074 603142 70130
rect 603210 70074 603266 70130
rect 603334 70074 603390 70130
rect 603458 70074 603514 70130
rect 603582 70074 603638 70130
rect 603706 70074 603762 70130
rect 603830 70074 603886 70130
rect 603954 70074 604010 70130
rect 604078 70074 604134 70130
rect 604822 70074 604878 70130
rect 604946 70074 605002 70130
rect 605070 70074 605126 70130
rect 605194 70074 605250 70130
rect 605318 70074 605374 70130
rect 605442 70074 605498 70130
rect 605566 70074 605622 70130
rect 605690 70074 605746 70130
rect 605814 70074 605870 70130
rect 605938 70074 605994 70130
rect 606062 70074 606118 70130
rect 606186 70074 606242 70130
rect 606310 70074 606366 70130
rect 606434 70074 606490 70130
rect 606558 70074 606614 70130
rect 606682 70074 606738 70130
rect 607192 70074 607248 70130
rect 607316 70074 607372 70130
rect 607440 70074 607496 70130
rect 607564 70074 607620 70130
rect 607688 70074 607744 70130
rect 607812 70074 607868 70130
rect 607936 70074 607992 70130
rect 608060 70074 608116 70130
rect 608184 70074 608240 70130
rect 608308 70074 608364 70130
rect 608432 70074 608488 70130
rect 608556 70074 608612 70130
rect 608680 70074 608736 70130
rect 608804 70074 608860 70130
rect 608928 70074 608984 70130
rect 609052 70074 609108 70130
rect 609892 70074 609948 70130
rect 610016 70074 610072 70130
rect 610140 70074 610196 70130
rect 610264 70074 610320 70130
rect 610388 70074 610444 70130
rect 610512 70074 610568 70130
rect 610636 70074 610692 70130
rect 610760 70074 610816 70130
rect 610884 70074 610940 70130
rect 611008 70074 611064 70130
rect 611132 70074 611188 70130
rect 611256 70074 611312 70130
rect 611380 70074 611436 70130
rect 611504 70074 611560 70130
rect 611628 70074 611684 70130
rect 611752 70074 611808 70130
rect 612262 70074 612318 70130
rect 612386 70074 612442 70130
rect 612510 70074 612566 70130
rect 612634 70074 612690 70130
rect 612758 70074 612814 70130
rect 612882 70074 612938 70130
rect 613006 70074 613062 70130
rect 613130 70074 613186 70130
rect 613254 70074 613310 70130
rect 613378 70074 613434 70130
rect 613502 70074 613558 70130
rect 613626 70074 613682 70130
rect 613750 70074 613806 70130
rect 613874 70074 613930 70130
rect 613998 70074 614054 70130
rect 614122 70074 614178 70130
rect 614866 70074 614922 70130
rect 614990 70074 615046 70130
rect 615114 70074 615170 70130
rect 615238 70074 615294 70130
rect 615362 70074 615418 70130
rect 615486 70074 615542 70130
rect 615610 70074 615666 70130
rect 615734 70074 615790 70130
rect 615858 70074 615914 70130
rect 615982 70074 616038 70130
rect 616106 70074 616162 70130
rect 616230 70074 616286 70130
rect 616354 70074 616410 70130
rect 616478 70074 616534 70130
rect 616602 70074 616658 70130
rect 657342 70074 657398 70130
rect 657466 70074 657522 70130
rect 657590 70074 657646 70130
rect 657714 70074 657770 70130
rect 657838 70074 657894 70130
rect 657962 70074 658018 70130
rect 658086 70074 658142 70130
rect 658210 70074 658266 70130
rect 658334 70074 658390 70130
rect 658458 70074 658514 70130
rect 658582 70074 658638 70130
rect 658706 70074 658762 70130
rect 658830 70074 658886 70130
rect 658954 70074 659010 70130
rect 659078 70074 659134 70130
rect 659822 70074 659878 70130
rect 659946 70074 660002 70130
rect 660070 70074 660126 70130
rect 660194 70074 660250 70130
rect 660318 70074 660374 70130
rect 660442 70074 660498 70130
rect 660566 70074 660622 70130
rect 660690 70074 660746 70130
rect 660814 70074 660870 70130
rect 660938 70074 660994 70130
rect 661062 70074 661118 70130
rect 661186 70074 661242 70130
rect 661310 70074 661366 70130
rect 661434 70074 661490 70130
rect 661558 70074 661614 70130
rect 661682 70074 661738 70130
rect 662192 70074 662248 70130
rect 662316 70074 662372 70130
rect 662440 70074 662496 70130
rect 662564 70074 662620 70130
rect 662688 70074 662744 70130
rect 662812 70074 662868 70130
rect 662936 70074 662992 70130
rect 663060 70074 663116 70130
rect 663184 70074 663240 70130
rect 663308 70074 663364 70130
rect 663432 70074 663488 70130
rect 663556 70074 663612 70130
rect 663680 70074 663736 70130
rect 663804 70074 663860 70130
rect 663928 70074 663984 70130
rect 664052 70074 664108 70130
rect 664892 70074 664948 70130
rect 665016 70074 665072 70130
rect 665140 70074 665196 70130
rect 665264 70074 665320 70130
rect 665388 70074 665444 70130
rect 665512 70074 665568 70130
rect 665636 70074 665692 70130
rect 665760 70074 665816 70130
rect 665884 70074 665940 70130
rect 666008 70074 666064 70130
rect 666132 70074 666188 70130
rect 666256 70074 666312 70130
rect 666380 70074 666436 70130
rect 666504 70074 666560 70130
rect 666628 70074 666684 70130
rect 666752 70074 666808 70130
rect 667262 70074 667318 70130
rect 667386 70074 667442 70130
rect 667510 70074 667566 70130
rect 667634 70074 667690 70130
rect 667758 70074 667814 70130
rect 667882 70074 667938 70130
rect 668006 70074 668062 70130
rect 668130 70074 668186 70130
rect 668254 70074 668310 70130
rect 668378 70074 668434 70130
rect 668502 70074 668558 70130
rect 668626 70074 668682 70130
rect 668750 70074 668806 70130
rect 668874 70074 668930 70130
rect 668998 70074 669054 70130
rect 669122 70074 669178 70130
rect 669866 70074 669922 70130
rect 669990 70074 670046 70130
rect 670114 70074 670170 70130
rect 670238 70074 670294 70130
rect 670362 70074 670418 70130
rect 670486 70074 670542 70130
rect 670610 70074 670666 70130
rect 670734 70074 670790 70130
rect 670858 70074 670914 70130
rect 670982 70074 671038 70130
rect 671106 70074 671162 70130
rect 671230 70074 671286 70130
rect 671354 70074 671410 70130
rect 671478 70074 671534 70130
rect 671602 70074 671658 70130
<< metal3 >>
rect 381272 949926 383172 950000
rect 381272 949870 381342 949926
rect 381398 949870 381466 949926
rect 381522 949870 381590 949926
rect 381646 949870 381714 949926
rect 381770 949870 381838 949926
rect 381894 949870 381962 949926
rect 382018 949870 382086 949926
rect 382142 949870 382210 949926
rect 382266 949870 382334 949926
rect 382390 949870 382458 949926
rect 382514 949870 382582 949926
rect 382638 949870 382706 949926
rect 382762 949870 382830 949926
rect 382886 949870 382954 949926
rect 383010 949870 383078 949926
rect 383134 949870 383172 949926
rect 381272 949800 383172 949870
rect 383752 949926 385802 950000
rect 383752 949870 383822 949926
rect 383878 949870 383946 949926
rect 384002 949870 384070 949926
rect 384126 949870 384194 949926
rect 384250 949870 384318 949926
rect 384374 949870 384442 949926
rect 384498 949870 384566 949926
rect 384622 949870 384690 949926
rect 384746 949870 384814 949926
rect 384870 949870 384938 949926
rect 384994 949870 385062 949926
rect 385118 949870 385186 949926
rect 385242 949870 385310 949926
rect 385366 949870 385434 949926
rect 385490 949870 385558 949926
rect 385614 949870 385682 949926
rect 385738 949870 385802 949926
rect 383752 949800 385802 949870
rect 386122 949926 388172 950000
rect 386122 949870 386192 949926
rect 386248 949870 386316 949926
rect 386372 949870 386440 949926
rect 386496 949870 386564 949926
rect 386620 949870 386688 949926
rect 386744 949870 386812 949926
rect 386868 949870 386936 949926
rect 386992 949870 387060 949926
rect 387116 949870 387184 949926
rect 387240 949870 387308 949926
rect 387364 949870 387432 949926
rect 387488 949870 387556 949926
rect 387612 949870 387680 949926
rect 387736 949870 387804 949926
rect 387860 949870 387928 949926
rect 387984 949870 388052 949926
rect 388108 949870 388172 949926
rect 386122 949800 388172 949870
rect 388828 949926 390878 950000
rect 388828 949870 388892 949926
rect 388948 949870 389016 949926
rect 389072 949870 389140 949926
rect 389196 949870 389264 949926
rect 389320 949870 389388 949926
rect 389444 949870 389512 949926
rect 389568 949870 389636 949926
rect 389692 949870 389760 949926
rect 389816 949870 389884 949926
rect 389940 949870 390008 949926
rect 390064 949870 390132 949926
rect 390188 949870 390256 949926
rect 390312 949870 390380 949926
rect 390436 949870 390504 949926
rect 390560 949870 390628 949926
rect 390684 949870 390752 949926
rect 390808 949870 390878 949926
rect 388828 949800 390878 949870
rect 391198 949926 393248 950000
rect 391198 949870 391262 949926
rect 391318 949870 391386 949926
rect 391442 949870 391510 949926
rect 391566 949870 391634 949926
rect 391690 949870 391758 949926
rect 391814 949870 391882 949926
rect 391938 949870 392006 949926
rect 392062 949870 392130 949926
rect 392186 949870 392254 949926
rect 392310 949870 392378 949926
rect 392434 949870 392502 949926
rect 392558 949870 392626 949926
rect 392682 949870 392750 949926
rect 392806 949870 392874 949926
rect 392930 949870 392998 949926
rect 393054 949870 393122 949926
rect 393178 949870 393248 949926
rect 391198 949800 393248 949870
rect 393828 949926 395728 950000
rect 393828 949870 393866 949926
rect 393922 949870 393990 949926
rect 394046 949870 394114 949926
rect 394170 949870 394238 949926
rect 394294 949870 394362 949926
rect 394418 949870 394486 949926
rect 394542 949870 394610 949926
rect 394666 949870 394734 949926
rect 394790 949870 394858 949926
rect 394914 949870 394982 949926
rect 395038 949870 395106 949926
rect 395162 949870 395230 949926
rect 395286 949870 395354 949926
rect 395410 949870 395478 949926
rect 395534 949870 395602 949926
rect 395658 949870 395728 949926
rect 393828 949800 395728 949870
rect 601272 949926 603172 950000
rect 601272 949870 601342 949926
rect 601398 949870 601466 949926
rect 601522 949870 601590 949926
rect 601646 949870 601714 949926
rect 601770 949870 601838 949926
rect 601894 949870 601962 949926
rect 602018 949870 602086 949926
rect 602142 949870 602210 949926
rect 602266 949870 602334 949926
rect 602390 949870 602458 949926
rect 602514 949870 602582 949926
rect 602638 949870 602706 949926
rect 602762 949870 602830 949926
rect 602886 949870 602954 949926
rect 603010 949870 603078 949926
rect 603134 949870 603172 949926
rect 601272 949800 603172 949870
rect 603752 949926 605802 950000
rect 603752 949870 603822 949926
rect 603878 949870 603946 949926
rect 604002 949870 604070 949926
rect 604126 949870 604194 949926
rect 604250 949870 604318 949926
rect 604374 949870 604442 949926
rect 604498 949870 604566 949926
rect 604622 949870 604690 949926
rect 604746 949870 604814 949926
rect 604870 949870 604938 949926
rect 604994 949870 605062 949926
rect 605118 949870 605186 949926
rect 605242 949870 605310 949926
rect 605366 949870 605434 949926
rect 605490 949870 605558 949926
rect 605614 949870 605682 949926
rect 605738 949870 605802 949926
rect 603752 949800 605802 949870
rect 606122 949926 608172 950000
rect 606122 949870 606192 949926
rect 606248 949870 606316 949926
rect 606372 949870 606440 949926
rect 606496 949870 606564 949926
rect 606620 949870 606688 949926
rect 606744 949870 606812 949926
rect 606868 949870 606936 949926
rect 606992 949870 607060 949926
rect 607116 949870 607184 949926
rect 607240 949870 607308 949926
rect 607364 949870 607432 949926
rect 607488 949870 607556 949926
rect 607612 949870 607680 949926
rect 607736 949870 607804 949926
rect 607860 949870 607928 949926
rect 607984 949870 608052 949926
rect 608108 949870 608172 949926
rect 606122 949800 608172 949870
rect 608828 949926 610878 950000
rect 608828 949870 608892 949926
rect 608948 949870 609016 949926
rect 609072 949870 609140 949926
rect 609196 949870 609264 949926
rect 609320 949870 609388 949926
rect 609444 949870 609512 949926
rect 609568 949870 609636 949926
rect 609692 949870 609760 949926
rect 609816 949870 609884 949926
rect 609940 949870 610008 949926
rect 610064 949870 610132 949926
rect 610188 949870 610256 949926
rect 610312 949870 610380 949926
rect 610436 949870 610504 949926
rect 610560 949870 610628 949926
rect 610684 949870 610752 949926
rect 610808 949870 610878 949926
rect 608828 949800 610878 949870
rect 611198 949926 613248 950000
rect 611198 949870 611262 949926
rect 611318 949870 611386 949926
rect 611442 949870 611510 949926
rect 611566 949870 611634 949926
rect 611690 949870 611758 949926
rect 611814 949870 611882 949926
rect 611938 949870 612006 949926
rect 612062 949870 612130 949926
rect 612186 949870 612254 949926
rect 612310 949870 612378 949926
rect 612434 949870 612502 949926
rect 612558 949870 612626 949926
rect 612682 949870 612750 949926
rect 612806 949870 612874 949926
rect 612930 949870 612998 949926
rect 613054 949870 613122 949926
rect 613178 949870 613248 949926
rect 611198 949800 613248 949870
rect 613828 949926 615728 950000
rect 613828 949870 613866 949926
rect 613922 949870 613990 949926
rect 614046 949870 614114 949926
rect 614170 949870 614238 949926
rect 614294 949870 614362 949926
rect 614418 949870 614486 949926
rect 614542 949870 614610 949926
rect 614666 949870 614734 949926
rect 614790 949870 614858 949926
rect 614914 949870 614982 949926
rect 615038 949870 615106 949926
rect 615162 949870 615230 949926
rect 615286 949870 615354 949926
rect 615410 949870 615478 949926
rect 615534 949870 615602 949926
rect 615658 949870 615728 949926
rect 613828 949800 615728 949870
rect 70000 884658 70200 884728
rect 70000 884602 70074 884658
rect 70130 884602 70200 884658
rect 70000 884534 70200 884602
rect 70000 884478 70074 884534
rect 70130 884478 70200 884534
rect 70000 884410 70200 884478
rect 70000 884354 70074 884410
rect 70130 884354 70200 884410
rect 70000 884286 70200 884354
rect 70000 884230 70074 884286
rect 70130 884230 70200 884286
rect 70000 884162 70200 884230
rect 70000 884106 70074 884162
rect 70130 884106 70200 884162
rect 70000 884038 70200 884106
rect 70000 883982 70074 884038
rect 70130 883982 70200 884038
rect 70000 883914 70200 883982
rect 70000 883858 70074 883914
rect 70130 883858 70200 883914
rect 70000 883790 70200 883858
rect 70000 883734 70074 883790
rect 70130 883734 70200 883790
rect 70000 883666 70200 883734
rect 70000 883610 70074 883666
rect 70130 883610 70200 883666
rect 70000 883542 70200 883610
rect 70000 883486 70074 883542
rect 70130 883486 70200 883542
rect 70000 883418 70200 883486
rect 70000 883362 70074 883418
rect 70130 883362 70200 883418
rect 70000 883294 70200 883362
rect 70000 883238 70074 883294
rect 70130 883238 70200 883294
rect 70000 883170 70200 883238
rect 70000 883114 70074 883170
rect 70130 883114 70200 883170
rect 70000 883046 70200 883114
rect 70000 882990 70074 883046
rect 70130 882990 70200 883046
rect 70000 882922 70200 882990
rect 70000 882866 70074 882922
rect 70130 882866 70200 882922
rect 70000 882828 70200 882866
rect 707800 883658 708000 883728
rect 707800 883602 707870 883658
rect 707926 883602 708000 883658
rect 707800 883534 708000 883602
rect 707800 883478 707870 883534
rect 707926 883478 708000 883534
rect 707800 883410 708000 883478
rect 707800 883354 707870 883410
rect 707926 883354 708000 883410
rect 707800 883286 708000 883354
rect 707800 883230 707870 883286
rect 707926 883230 708000 883286
rect 707800 883162 708000 883230
rect 707800 883106 707870 883162
rect 707926 883106 708000 883162
rect 707800 883038 708000 883106
rect 707800 882982 707870 883038
rect 707926 882982 708000 883038
rect 707800 882914 708000 882982
rect 707800 882858 707870 882914
rect 707926 882858 708000 882914
rect 707800 882790 708000 882858
rect 707800 882734 707870 882790
rect 707926 882734 708000 882790
rect 707800 882666 708000 882734
rect 707800 882610 707870 882666
rect 707926 882610 708000 882666
rect 707800 882542 708000 882610
rect 707800 882486 707870 882542
rect 707926 882486 708000 882542
rect 707800 882418 708000 882486
rect 707800 882362 707870 882418
rect 707926 882362 708000 882418
rect 707800 882294 708000 882362
rect 70000 882184 70200 882248
rect 70000 882128 70074 882184
rect 70130 882128 70200 882184
rect 70000 882060 70200 882128
rect 70000 882004 70074 882060
rect 70130 882004 70200 882060
rect 70000 881936 70200 882004
rect 70000 881880 70074 881936
rect 70130 881880 70200 881936
rect 70000 881812 70200 881880
rect 707800 882238 707870 882294
rect 707926 882238 708000 882294
rect 707800 882170 708000 882238
rect 707800 882114 707870 882170
rect 707926 882114 708000 882170
rect 707800 882046 708000 882114
rect 707800 881990 707870 882046
rect 707926 881990 708000 882046
rect 707800 881922 708000 881990
rect 707800 881866 707870 881922
rect 707926 881866 708000 881922
rect 707800 881828 708000 881866
rect 70000 881756 70074 881812
rect 70130 881756 70200 881812
rect 70000 881688 70200 881756
rect 70000 881632 70074 881688
rect 70130 881632 70200 881688
rect 70000 881564 70200 881632
rect 70000 881508 70074 881564
rect 70130 881508 70200 881564
rect 70000 881440 70200 881508
rect 70000 881384 70074 881440
rect 70130 881384 70200 881440
rect 70000 881316 70200 881384
rect 70000 881260 70074 881316
rect 70130 881260 70200 881316
rect 70000 881192 70200 881260
rect 70000 881136 70074 881192
rect 70130 881136 70200 881192
rect 70000 881068 70200 881136
rect 70000 881012 70074 881068
rect 70130 881012 70200 881068
rect 70000 880944 70200 881012
rect 70000 880888 70074 880944
rect 70130 880888 70200 880944
rect 70000 880820 70200 880888
rect 70000 880764 70074 880820
rect 70130 880764 70200 880820
rect 70000 880696 70200 880764
rect 70000 880640 70074 880696
rect 70130 880640 70200 880696
rect 70000 880572 70200 880640
rect 70000 880516 70074 880572
rect 70130 880516 70200 880572
rect 70000 880448 70200 880516
rect 70000 880392 70074 880448
rect 70130 880392 70200 880448
rect 70000 880324 70200 880392
rect 70000 880268 70074 880324
rect 70130 880268 70200 880324
rect 70000 880198 70200 880268
rect 707800 881178 708000 881248
rect 707800 881122 707870 881178
rect 707926 881122 708000 881178
rect 707800 881054 708000 881122
rect 707800 880998 707870 881054
rect 707926 880998 708000 881054
rect 707800 880930 708000 880998
rect 707800 880874 707870 880930
rect 707926 880874 708000 880930
rect 707800 880806 708000 880874
rect 707800 880750 707870 880806
rect 707926 880750 708000 880806
rect 707800 880682 708000 880750
rect 707800 880626 707870 880682
rect 707926 880626 708000 880682
rect 707800 880558 708000 880626
rect 707800 880502 707870 880558
rect 707926 880502 708000 880558
rect 707800 880434 708000 880502
rect 707800 880378 707870 880434
rect 707926 880378 708000 880434
rect 707800 880310 708000 880378
rect 707800 880254 707870 880310
rect 707926 880254 708000 880310
rect 707800 880186 708000 880254
rect 707800 880130 707870 880186
rect 707926 880130 708000 880186
rect 707800 880062 708000 880130
rect 707800 880006 707870 880062
rect 707926 880006 708000 880062
rect 707800 879938 708000 880006
rect 707800 879882 707870 879938
rect 707926 879882 708000 879938
rect 70000 879814 70200 879878
rect 70000 879758 70074 879814
rect 70130 879758 70200 879814
rect 70000 879690 70200 879758
rect 70000 879634 70074 879690
rect 70130 879634 70200 879690
rect 70000 879566 70200 879634
rect 70000 879510 70074 879566
rect 70130 879510 70200 879566
rect 70000 879442 70200 879510
rect 70000 879386 70074 879442
rect 70130 879386 70200 879442
rect 70000 879318 70200 879386
rect 70000 879262 70074 879318
rect 70130 879262 70200 879318
rect 70000 879194 70200 879262
rect 707800 879814 708000 879882
rect 707800 879758 707870 879814
rect 707926 879758 708000 879814
rect 707800 879690 708000 879758
rect 707800 879634 707870 879690
rect 707926 879634 708000 879690
rect 707800 879566 708000 879634
rect 707800 879510 707870 879566
rect 707926 879510 708000 879566
rect 707800 879442 708000 879510
rect 707800 879386 707870 879442
rect 707926 879386 708000 879442
rect 707800 879318 708000 879386
rect 707800 879262 707870 879318
rect 707926 879262 708000 879318
rect 707800 879198 708000 879262
rect 70000 879138 70074 879194
rect 70130 879138 70200 879194
rect 70000 879070 70200 879138
rect 70000 879014 70074 879070
rect 70130 879014 70200 879070
rect 70000 878946 70200 879014
rect 70000 878890 70074 878946
rect 70130 878890 70200 878946
rect 70000 878822 70200 878890
rect 70000 878766 70074 878822
rect 70130 878766 70200 878822
rect 70000 878698 70200 878766
rect 70000 878642 70074 878698
rect 70130 878642 70200 878698
rect 70000 878574 70200 878642
rect 70000 878518 70074 878574
rect 70130 878518 70200 878574
rect 70000 878450 70200 878518
rect 70000 878394 70074 878450
rect 70130 878394 70200 878450
rect 70000 878326 70200 878394
rect 70000 878270 70074 878326
rect 70130 878270 70200 878326
rect 70000 878202 70200 878270
rect 70000 878146 70074 878202
rect 70130 878146 70200 878202
rect 70000 878078 70200 878146
rect 70000 878022 70074 878078
rect 70130 878022 70200 878078
rect 70000 877954 70200 878022
rect 70000 877898 70074 877954
rect 70130 877898 70200 877954
rect 70000 877828 70200 877898
rect 707800 878808 708000 878878
rect 707800 878752 707870 878808
rect 707926 878752 708000 878808
rect 707800 878684 708000 878752
rect 707800 878628 707870 878684
rect 707926 878628 708000 878684
rect 707800 878560 708000 878628
rect 707800 878504 707870 878560
rect 707926 878504 708000 878560
rect 707800 878436 708000 878504
rect 707800 878380 707870 878436
rect 707926 878380 708000 878436
rect 707800 878312 708000 878380
rect 707800 878256 707870 878312
rect 707926 878256 708000 878312
rect 707800 878188 708000 878256
rect 707800 878132 707870 878188
rect 707926 878132 708000 878188
rect 707800 878064 708000 878132
rect 707800 878008 707870 878064
rect 707926 878008 708000 878064
rect 707800 877940 708000 878008
rect 707800 877884 707870 877940
rect 707926 877884 708000 877940
rect 707800 877816 708000 877884
rect 707800 877760 707870 877816
rect 707926 877760 708000 877816
rect 707800 877692 708000 877760
rect 707800 877636 707870 877692
rect 707926 877636 708000 877692
rect 707800 877568 708000 877636
rect 707800 877512 707870 877568
rect 707926 877512 708000 877568
rect 707800 877444 708000 877512
rect 707800 877388 707870 877444
rect 707926 877388 708000 877444
rect 707800 877320 708000 877388
rect 707800 877264 707870 877320
rect 707926 877264 708000 877320
rect 707800 877196 708000 877264
rect 70000 877108 70200 877172
rect 70000 877052 70074 877108
rect 70130 877052 70200 877108
rect 70000 876984 70200 877052
rect 70000 876928 70074 876984
rect 70130 876928 70200 876984
rect 70000 876860 70200 876928
rect 70000 876804 70074 876860
rect 70130 876804 70200 876860
rect 707800 877140 707870 877196
rect 707926 877140 708000 877196
rect 707800 877072 708000 877140
rect 707800 877016 707870 877072
rect 707926 877016 708000 877072
rect 707800 876948 708000 877016
rect 707800 876892 707870 876948
rect 707926 876892 708000 876948
rect 707800 876828 708000 876892
rect 70000 876736 70200 876804
rect 70000 876680 70074 876736
rect 70130 876680 70200 876736
rect 70000 876612 70200 876680
rect 70000 876556 70074 876612
rect 70130 876556 70200 876612
rect 70000 876488 70200 876556
rect 70000 876432 70074 876488
rect 70130 876432 70200 876488
rect 70000 876364 70200 876432
rect 70000 876308 70074 876364
rect 70130 876308 70200 876364
rect 70000 876240 70200 876308
rect 70000 876184 70074 876240
rect 70130 876184 70200 876240
rect 70000 876116 70200 876184
rect 70000 876060 70074 876116
rect 70130 876060 70200 876116
rect 70000 875992 70200 876060
rect 70000 875936 70074 875992
rect 70130 875936 70200 875992
rect 70000 875868 70200 875936
rect 70000 875812 70074 875868
rect 70130 875812 70200 875868
rect 70000 875744 70200 875812
rect 70000 875688 70074 875744
rect 70130 875688 70200 875744
rect 70000 875620 70200 875688
rect 70000 875564 70074 875620
rect 70130 875564 70200 875620
rect 70000 875496 70200 875564
rect 70000 875440 70074 875496
rect 70130 875440 70200 875496
rect 70000 875372 70200 875440
rect 70000 875316 70074 875372
rect 70130 875316 70200 875372
rect 70000 875248 70200 875316
rect 70000 875192 70074 875248
rect 70130 875192 70200 875248
rect 70000 875122 70200 875192
rect 707800 876102 708000 876172
rect 707800 876046 707870 876102
rect 707926 876046 708000 876102
rect 707800 875978 708000 876046
rect 707800 875922 707870 875978
rect 707926 875922 708000 875978
rect 707800 875854 708000 875922
rect 707800 875798 707870 875854
rect 707926 875798 708000 875854
rect 707800 875730 708000 875798
rect 707800 875674 707870 875730
rect 707926 875674 708000 875730
rect 707800 875606 708000 875674
rect 707800 875550 707870 875606
rect 707926 875550 708000 875606
rect 707800 875482 708000 875550
rect 707800 875426 707870 875482
rect 707926 875426 708000 875482
rect 707800 875358 708000 875426
rect 707800 875302 707870 875358
rect 707926 875302 708000 875358
rect 707800 875234 708000 875302
rect 707800 875178 707870 875234
rect 707926 875178 708000 875234
rect 707800 875110 708000 875178
rect 707800 875054 707870 875110
rect 707926 875054 708000 875110
rect 707800 874986 708000 875054
rect 707800 874930 707870 874986
rect 707926 874930 708000 874986
rect 707800 874862 708000 874930
rect 707800 874806 707870 874862
rect 707926 874806 708000 874862
rect 70000 874738 70200 874802
rect 70000 874682 70074 874738
rect 70130 874682 70200 874738
rect 70000 874614 70200 874682
rect 70000 874558 70074 874614
rect 70130 874558 70200 874614
rect 70000 874490 70200 874558
rect 70000 874434 70074 874490
rect 70130 874434 70200 874490
rect 70000 874366 70200 874434
rect 70000 874310 70074 874366
rect 70130 874310 70200 874366
rect 70000 874242 70200 874310
rect 70000 874186 70074 874242
rect 70130 874186 70200 874242
rect 70000 874118 70200 874186
rect 707800 874738 708000 874806
rect 707800 874682 707870 874738
rect 707926 874682 708000 874738
rect 707800 874614 708000 874682
rect 707800 874558 707870 874614
rect 707926 874558 708000 874614
rect 707800 874490 708000 874558
rect 707800 874434 707870 874490
rect 707926 874434 708000 874490
rect 707800 874366 708000 874434
rect 707800 874310 707870 874366
rect 707926 874310 708000 874366
rect 707800 874242 708000 874310
rect 707800 874186 707870 874242
rect 707926 874186 708000 874242
rect 707800 874122 708000 874186
rect 70000 874062 70074 874118
rect 70130 874062 70200 874118
rect 70000 873994 70200 874062
rect 70000 873938 70074 873994
rect 70130 873938 70200 873994
rect 70000 873870 70200 873938
rect 70000 873814 70074 873870
rect 70130 873814 70200 873870
rect 70000 873746 70200 873814
rect 70000 873690 70074 873746
rect 70130 873690 70200 873746
rect 70000 873622 70200 873690
rect 70000 873566 70074 873622
rect 70130 873566 70200 873622
rect 70000 873498 70200 873566
rect 70000 873442 70074 873498
rect 70130 873442 70200 873498
rect 70000 873374 70200 873442
rect 70000 873318 70074 873374
rect 70130 873318 70200 873374
rect 70000 873250 70200 873318
rect 70000 873194 70074 873250
rect 70130 873194 70200 873250
rect 70000 873126 70200 873194
rect 70000 873070 70074 873126
rect 70130 873070 70200 873126
rect 70000 873002 70200 873070
rect 70000 872946 70074 873002
rect 70130 872946 70200 873002
rect 70000 872878 70200 872946
rect 70000 872822 70074 872878
rect 70130 872822 70200 872878
rect 70000 872752 70200 872822
rect 707800 873732 708000 873802
rect 707800 873676 707870 873732
rect 707926 873676 708000 873732
rect 707800 873608 708000 873676
rect 707800 873552 707870 873608
rect 707926 873552 708000 873608
rect 707800 873484 708000 873552
rect 707800 873428 707870 873484
rect 707926 873428 708000 873484
rect 707800 873360 708000 873428
rect 707800 873304 707870 873360
rect 707926 873304 708000 873360
rect 707800 873236 708000 873304
rect 707800 873180 707870 873236
rect 707926 873180 708000 873236
rect 707800 873112 708000 873180
rect 707800 873056 707870 873112
rect 707926 873056 708000 873112
rect 707800 872988 708000 873056
rect 707800 872932 707870 872988
rect 707926 872932 708000 872988
rect 707800 872864 708000 872932
rect 707800 872808 707870 872864
rect 707926 872808 708000 872864
rect 707800 872740 708000 872808
rect 707800 872684 707870 872740
rect 707926 872684 708000 872740
rect 707800 872616 708000 872684
rect 707800 872560 707870 872616
rect 707926 872560 708000 872616
rect 707800 872492 708000 872560
rect 707800 872436 707870 872492
rect 707926 872436 708000 872492
rect 707800 872368 708000 872436
rect 707800 872312 707870 872368
rect 707926 872312 708000 872368
rect 707800 872244 708000 872312
rect 707800 872188 707870 872244
rect 707926 872188 708000 872244
rect 70000 872134 70200 872172
rect 70000 872078 70074 872134
rect 70130 872078 70200 872134
rect 70000 872010 70200 872078
rect 70000 871954 70074 872010
rect 70130 871954 70200 872010
rect 70000 871886 70200 871954
rect 70000 871830 70074 871886
rect 70130 871830 70200 871886
rect 70000 871762 70200 871830
rect 70000 871706 70074 871762
rect 70130 871706 70200 871762
rect 707800 872120 708000 872188
rect 707800 872064 707870 872120
rect 707926 872064 708000 872120
rect 707800 871996 708000 872064
rect 707800 871940 707870 871996
rect 707926 871940 708000 871996
rect 707800 871872 708000 871940
rect 707800 871816 707870 871872
rect 707926 871816 708000 871872
rect 707800 871752 708000 871816
rect 70000 871638 70200 871706
rect 70000 871582 70074 871638
rect 70130 871582 70200 871638
rect 70000 871514 70200 871582
rect 70000 871458 70074 871514
rect 70130 871458 70200 871514
rect 70000 871390 70200 871458
rect 70000 871334 70074 871390
rect 70130 871334 70200 871390
rect 70000 871266 70200 871334
rect 70000 871210 70074 871266
rect 70130 871210 70200 871266
rect 70000 871142 70200 871210
rect 70000 871086 70074 871142
rect 70130 871086 70200 871142
rect 70000 871018 70200 871086
rect 70000 870962 70074 871018
rect 70130 870962 70200 871018
rect 70000 870894 70200 870962
rect 70000 870838 70074 870894
rect 70130 870838 70200 870894
rect 70000 870770 70200 870838
rect 70000 870714 70074 870770
rect 70130 870714 70200 870770
rect 70000 870646 70200 870714
rect 70000 870590 70074 870646
rect 70130 870590 70200 870646
rect 70000 870522 70200 870590
rect 70000 870466 70074 870522
rect 70130 870466 70200 870522
rect 70000 870398 70200 870466
rect 70000 870342 70074 870398
rect 70130 870342 70200 870398
rect 70000 870272 70200 870342
rect 707800 871134 708000 871172
rect 707800 871078 707870 871134
rect 707926 871078 708000 871134
rect 707800 871010 708000 871078
rect 707800 870954 707870 871010
rect 707926 870954 708000 871010
rect 707800 870886 708000 870954
rect 707800 870830 707870 870886
rect 707926 870830 708000 870886
rect 707800 870762 708000 870830
rect 707800 870706 707870 870762
rect 707926 870706 708000 870762
rect 707800 870638 708000 870706
rect 707800 870582 707870 870638
rect 707926 870582 708000 870638
rect 707800 870514 708000 870582
rect 707800 870458 707870 870514
rect 707926 870458 708000 870514
rect 707800 870390 708000 870458
rect 707800 870334 707870 870390
rect 707926 870334 708000 870390
rect 707800 870266 708000 870334
rect 707800 870210 707870 870266
rect 707926 870210 708000 870266
rect 707800 870142 708000 870210
rect 707800 870086 707870 870142
rect 707926 870086 708000 870142
rect 707800 870018 708000 870086
rect 707800 869962 707870 870018
rect 707926 869962 708000 870018
rect 707800 869894 708000 869962
rect 707800 869838 707870 869894
rect 707926 869838 708000 869894
rect 707800 869770 708000 869838
rect 707800 869714 707870 869770
rect 707926 869714 708000 869770
rect 707800 869646 708000 869714
rect 707800 869590 707870 869646
rect 707926 869590 708000 869646
rect 707800 869522 708000 869590
rect 707800 869466 707870 869522
rect 707926 869466 708000 869522
rect 707800 869398 708000 869466
rect 707800 869342 707870 869398
rect 707926 869342 708000 869398
rect 707800 869272 708000 869342
rect 70000 843658 70200 843728
rect 70000 843602 70074 843658
rect 70130 843602 70200 843658
rect 70000 843534 70200 843602
rect 70000 843478 70074 843534
rect 70130 843478 70200 843534
rect 70000 843410 70200 843478
rect 70000 843354 70074 843410
rect 70130 843354 70200 843410
rect 70000 843286 70200 843354
rect 70000 843230 70074 843286
rect 70130 843230 70200 843286
rect 70000 843162 70200 843230
rect 70000 843106 70074 843162
rect 70130 843106 70200 843162
rect 70000 843038 70200 843106
rect 70000 842982 70074 843038
rect 70130 842982 70200 843038
rect 70000 842914 70200 842982
rect 70000 842858 70074 842914
rect 70130 842858 70200 842914
rect 70000 842790 70200 842858
rect 70000 842734 70074 842790
rect 70130 842734 70200 842790
rect 70000 842666 70200 842734
rect 70000 842610 70074 842666
rect 70130 842610 70200 842666
rect 70000 842542 70200 842610
rect 70000 842486 70074 842542
rect 70130 842486 70200 842542
rect 70000 842418 70200 842486
rect 70000 842362 70074 842418
rect 70130 842362 70200 842418
rect 70000 842294 70200 842362
rect 70000 842238 70074 842294
rect 70130 842238 70200 842294
rect 70000 842170 70200 842238
rect 70000 842114 70074 842170
rect 70130 842114 70200 842170
rect 70000 842046 70200 842114
rect 70000 841990 70074 842046
rect 70130 841990 70200 842046
rect 70000 841922 70200 841990
rect 70000 841866 70074 841922
rect 70130 841866 70200 841922
rect 70000 841828 70200 841866
rect 70000 841184 70200 841248
rect 70000 841128 70074 841184
rect 70130 841128 70200 841184
rect 70000 841060 70200 841128
rect 70000 841004 70074 841060
rect 70130 841004 70200 841060
rect 70000 840936 70200 841004
rect 70000 840880 70074 840936
rect 70130 840880 70200 840936
rect 70000 840812 70200 840880
rect 70000 840756 70074 840812
rect 70130 840756 70200 840812
rect 70000 840688 70200 840756
rect 70000 840632 70074 840688
rect 70130 840632 70200 840688
rect 70000 840564 70200 840632
rect 70000 840508 70074 840564
rect 70130 840508 70200 840564
rect 70000 840440 70200 840508
rect 70000 840384 70074 840440
rect 70130 840384 70200 840440
rect 70000 840316 70200 840384
rect 70000 840260 70074 840316
rect 70130 840260 70200 840316
rect 70000 840192 70200 840260
rect 70000 840136 70074 840192
rect 70130 840136 70200 840192
rect 70000 840068 70200 840136
rect 70000 840012 70074 840068
rect 70130 840012 70200 840068
rect 70000 839944 70200 840012
rect 70000 839888 70074 839944
rect 70130 839888 70200 839944
rect 70000 839820 70200 839888
rect 70000 839764 70074 839820
rect 70130 839764 70200 839820
rect 70000 839696 70200 839764
rect 70000 839640 70074 839696
rect 70130 839640 70200 839696
rect 70000 839572 70200 839640
rect 70000 839516 70074 839572
rect 70130 839516 70200 839572
rect 70000 839448 70200 839516
rect 70000 839392 70074 839448
rect 70130 839392 70200 839448
rect 70000 839324 70200 839392
rect 70000 839268 70074 839324
rect 70130 839268 70200 839324
rect 70000 839198 70200 839268
rect 70000 838814 70200 838878
rect 70000 838758 70074 838814
rect 70130 838758 70200 838814
rect 70000 838690 70200 838758
rect 70000 838634 70074 838690
rect 70130 838634 70200 838690
rect 70000 838566 70200 838634
rect 70000 838510 70074 838566
rect 70130 838510 70200 838566
rect 70000 838442 70200 838510
rect 70000 838386 70074 838442
rect 70130 838386 70200 838442
rect 70000 838318 70200 838386
rect 70000 838262 70074 838318
rect 70130 838262 70200 838318
rect 70000 838194 70200 838262
rect 70000 838138 70074 838194
rect 70130 838138 70200 838194
rect 70000 838070 70200 838138
rect 70000 838014 70074 838070
rect 70130 838014 70200 838070
rect 70000 837946 70200 838014
rect 70000 837890 70074 837946
rect 70130 837890 70200 837946
rect 70000 837822 70200 837890
rect 70000 837766 70074 837822
rect 70130 837766 70200 837822
rect 70000 837698 70200 837766
rect 70000 837642 70074 837698
rect 70130 837642 70200 837698
rect 70000 837574 70200 837642
rect 70000 837518 70074 837574
rect 70130 837518 70200 837574
rect 70000 837450 70200 837518
rect 70000 837394 70074 837450
rect 70130 837394 70200 837450
rect 70000 837326 70200 837394
rect 70000 837270 70074 837326
rect 70130 837270 70200 837326
rect 70000 837202 70200 837270
rect 70000 837146 70074 837202
rect 70130 837146 70200 837202
rect 70000 837078 70200 837146
rect 70000 837022 70074 837078
rect 70130 837022 70200 837078
rect 70000 836954 70200 837022
rect 70000 836898 70074 836954
rect 70130 836898 70200 836954
rect 70000 836828 70200 836898
rect 70000 836108 70200 836172
rect 70000 836052 70074 836108
rect 70130 836052 70200 836108
rect 70000 835984 70200 836052
rect 70000 835928 70074 835984
rect 70130 835928 70200 835984
rect 70000 835860 70200 835928
rect 70000 835804 70074 835860
rect 70130 835804 70200 835860
rect 70000 835736 70200 835804
rect 70000 835680 70074 835736
rect 70130 835680 70200 835736
rect 70000 835612 70200 835680
rect 70000 835556 70074 835612
rect 70130 835556 70200 835612
rect 70000 835488 70200 835556
rect 70000 835432 70074 835488
rect 70130 835432 70200 835488
rect 70000 835364 70200 835432
rect 70000 835308 70074 835364
rect 70130 835308 70200 835364
rect 70000 835240 70200 835308
rect 70000 835184 70074 835240
rect 70130 835184 70200 835240
rect 70000 835116 70200 835184
rect 70000 835060 70074 835116
rect 70130 835060 70200 835116
rect 70000 834992 70200 835060
rect 70000 834936 70074 834992
rect 70130 834936 70200 834992
rect 70000 834868 70200 834936
rect 70000 834812 70074 834868
rect 70130 834812 70200 834868
rect 70000 834744 70200 834812
rect 70000 834688 70074 834744
rect 70130 834688 70200 834744
rect 70000 834620 70200 834688
rect 70000 834564 70074 834620
rect 70130 834564 70200 834620
rect 70000 834496 70200 834564
rect 70000 834440 70074 834496
rect 70130 834440 70200 834496
rect 70000 834372 70200 834440
rect 70000 834316 70074 834372
rect 70130 834316 70200 834372
rect 70000 834248 70200 834316
rect 70000 834192 70074 834248
rect 70130 834192 70200 834248
rect 70000 834122 70200 834192
rect 70000 833738 70200 833802
rect 70000 833682 70074 833738
rect 70130 833682 70200 833738
rect 70000 833614 70200 833682
rect 70000 833558 70074 833614
rect 70130 833558 70200 833614
rect 70000 833490 70200 833558
rect 70000 833434 70074 833490
rect 70130 833434 70200 833490
rect 70000 833366 70200 833434
rect 70000 833310 70074 833366
rect 70130 833310 70200 833366
rect 70000 833242 70200 833310
rect 70000 833186 70074 833242
rect 70130 833186 70200 833242
rect 70000 833118 70200 833186
rect 70000 833062 70074 833118
rect 70130 833062 70200 833118
rect 70000 832994 70200 833062
rect 70000 832938 70074 832994
rect 70130 832938 70200 832994
rect 70000 832870 70200 832938
rect 70000 832814 70074 832870
rect 70130 832814 70200 832870
rect 70000 832746 70200 832814
rect 70000 832690 70074 832746
rect 70130 832690 70200 832746
rect 70000 832622 70200 832690
rect 70000 832566 70074 832622
rect 70130 832566 70200 832622
rect 70000 832498 70200 832566
rect 70000 832442 70074 832498
rect 70130 832442 70200 832498
rect 70000 832374 70200 832442
rect 70000 832318 70074 832374
rect 70130 832318 70200 832374
rect 70000 832250 70200 832318
rect 70000 832194 70074 832250
rect 70130 832194 70200 832250
rect 70000 832126 70200 832194
rect 70000 832070 70074 832126
rect 70130 832070 70200 832126
rect 70000 832002 70200 832070
rect 70000 831946 70074 832002
rect 70130 831946 70200 832002
rect 70000 831878 70200 831946
rect 70000 831822 70074 831878
rect 70130 831822 70200 831878
rect 70000 831752 70200 831822
rect 70000 831134 70200 831172
rect 70000 831078 70074 831134
rect 70130 831078 70200 831134
rect 70000 831010 70200 831078
rect 70000 830954 70074 831010
rect 70130 830954 70200 831010
rect 70000 830886 70200 830954
rect 70000 830830 70074 830886
rect 70130 830830 70200 830886
rect 70000 830762 70200 830830
rect 70000 830706 70074 830762
rect 70130 830706 70200 830762
rect 70000 830638 70200 830706
rect 70000 830582 70074 830638
rect 70130 830582 70200 830638
rect 70000 830514 70200 830582
rect 70000 830458 70074 830514
rect 70130 830458 70200 830514
rect 70000 830390 70200 830458
rect 70000 830334 70074 830390
rect 70130 830334 70200 830390
rect 70000 830266 70200 830334
rect 70000 830210 70074 830266
rect 70130 830210 70200 830266
rect 70000 830142 70200 830210
rect 70000 830086 70074 830142
rect 70130 830086 70200 830142
rect 70000 830018 70200 830086
rect 70000 829962 70074 830018
rect 70130 829962 70200 830018
rect 70000 829894 70200 829962
rect 70000 829838 70074 829894
rect 70130 829838 70200 829894
rect 70000 829770 70200 829838
rect 70000 829714 70074 829770
rect 70130 829714 70200 829770
rect 70000 829646 70200 829714
rect 70000 829590 70074 829646
rect 70130 829590 70200 829646
rect 70000 829522 70200 829590
rect 70000 829466 70074 829522
rect 70130 829466 70200 829522
rect 70000 829398 70200 829466
rect 70000 829342 70074 829398
rect 70130 829342 70200 829398
rect 70000 829272 70200 829342
rect 70000 802658 70200 802728
rect 70000 802602 70074 802658
rect 70130 802602 70200 802658
rect 70000 802534 70200 802602
rect 70000 802478 70074 802534
rect 70130 802478 70200 802534
rect 70000 802410 70200 802478
rect 70000 802354 70074 802410
rect 70130 802354 70200 802410
rect 70000 802286 70200 802354
rect 70000 802230 70074 802286
rect 70130 802230 70200 802286
rect 70000 802162 70200 802230
rect 70000 802106 70074 802162
rect 70130 802106 70200 802162
rect 70000 802038 70200 802106
rect 70000 801982 70074 802038
rect 70130 801982 70200 802038
rect 70000 801914 70200 801982
rect 70000 801858 70074 801914
rect 70130 801858 70200 801914
rect 70000 801790 70200 801858
rect 70000 801734 70074 801790
rect 70130 801734 70200 801790
rect 70000 801666 70200 801734
rect 70000 801610 70074 801666
rect 70130 801610 70200 801666
rect 70000 801542 70200 801610
rect 70000 801486 70074 801542
rect 70130 801486 70200 801542
rect 70000 801418 70200 801486
rect 70000 801362 70074 801418
rect 70130 801362 70200 801418
rect 70000 801294 70200 801362
rect 70000 801238 70074 801294
rect 70130 801238 70200 801294
rect 70000 801170 70200 801238
rect 70000 801114 70074 801170
rect 70130 801114 70200 801170
rect 70000 801046 70200 801114
rect 70000 800990 70074 801046
rect 70130 800990 70200 801046
rect 70000 800922 70200 800990
rect 70000 800866 70074 800922
rect 70130 800866 70200 800922
rect 70000 800828 70200 800866
rect 70000 800184 70200 800248
rect 70000 800128 70074 800184
rect 70130 800128 70200 800184
rect 70000 800060 70200 800128
rect 70000 800004 70074 800060
rect 70130 800004 70200 800060
rect 70000 799936 70200 800004
rect 70000 799880 70074 799936
rect 70130 799880 70200 799936
rect 70000 799812 70200 799880
rect 70000 799756 70074 799812
rect 70130 799756 70200 799812
rect 70000 799688 70200 799756
rect 70000 799632 70074 799688
rect 70130 799632 70200 799688
rect 70000 799564 70200 799632
rect 70000 799508 70074 799564
rect 70130 799508 70200 799564
rect 70000 799440 70200 799508
rect 70000 799384 70074 799440
rect 70130 799384 70200 799440
rect 70000 799316 70200 799384
rect 70000 799260 70074 799316
rect 70130 799260 70200 799316
rect 70000 799192 70200 799260
rect 70000 799136 70074 799192
rect 70130 799136 70200 799192
rect 70000 799068 70200 799136
rect 70000 799012 70074 799068
rect 70130 799012 70200 799068
rect 70000 798944 70200 799012
rect 70000 798888 70074 798944
rect 70130 798888 70200 798944
rect 70000 798820 70200 798888
rect 70000 798764 70074 798820
rect 70130 798764 70200 798820
rect 70000 798696 70200 798764
rect 70000 798640 70074 798696
rect 70130 798640 70200 798696
rect 70000 798572 70200 798640
rect 70000 798516 70074 798572
rect 70130 798516 70200 798572
rect 70000 798448 70200 798516
rect 70000 798392 70074 798448
rect 70130 798392 70200 798448
rect 70000 798324 70200 798392
rect 70000 798268 70074 798324
rect 70130 798268 70200 798324
rect 70000 798198 70200 798268
rect 70000 797814 70200 797878
rect 70000 797758 70074 797814
rect 70130 797758 70200 797814
rect 70000 797690 70200 797758
rect 70000 797634 70074 797690
rect 70130 797634 70200 797690
rect 70000 797566 70200 797634
rect 70000 797510 70074 797566
rect 70130 797510 70200 797566
rect 70000 797442 70200 797510
rect 70000 797386 70074 797442
rect 70130 797386 70200 797442
rect 70000 797318 70200 797386
rect 70000 797262 70074 797318
rect 70130 797262 70200 797318
rect 70000 797194 70200 797262
rect 70000 797138 70074 797194
rect 70130 797138 70200 797194
rect 70000 797070 70200 797138
rect 70000 797014 70074 797070
rect 70130 797014 70200 797070
rect 70000 796946 70200 797014
rect 70000 796890 70074 796946
rect 70130 796890 70200 796946
rect 70000 796822 70200 796890
rect 70000 796766 70074 796822
rect 70130 796766 70200 796822
rect 70000 796698 70200 796766
rect 70000 796642 70074 796698
rect 70130 796642 70200 796698
rect 70000 796574 70200 796642
rect 70000 796518 70074 796574
rect 70130 796518 70200 796574
rect 70000 796450 70200 796518
rect 70000 796394 70074 796450
rect 70130 796394 70200 796450
rect 70000 796326 70200 796394
rect 70000 796270 70074 796326
rect 70130 796270 70200 796326
rect 70000 796202 70200 796270
rect 70000 796146 70074 796202
rect 70130 796146 70200 796202
rect 70000 796078 70200 796146
rect 70000 796022 70074 796078
rect 70130 796022 70200 796078
rect 70000 795954 70200 796022
rect 70000 795898 70074 795954
rect 70130 795898 70200 795954
rect 70000 795828 70200 795898
rect 707800 797658 708000 797728
rect 707800 797602 707870 797658
rect 707926 797602 708000 797658
rect 707800 797534 708000 797602
rect 707800 797478 707870 797534
rect 707926 797478 708000 797534
rect 707800 797410 708000 797478
rect 707800 797354 707870 797410
rect 707926 797354 708000 797410
rect 707800 797286 708000 797354
rect 707800 797230 707870 797286
rect 707926 797230 708000 797286
rect 707800 797162 708000 797230
rect 707800 797106 707870 797162
rect 707926 797106 708000 797162
rect 707800 797038 708000 797106
rect 707800 796982 707870 797038
rect 707926 796982 708000 797038
rect 707800 796914 708000 796982
rect 707800 796858 707870 796914
rect 707926 796858 708000 796914
rect 707800 796790 708000 796858
rect 707800 796734 707870 796790
rect 707926 796734 708000 796790
rect 707800 796666 708000 796734
rect 707800 796610 707870 796666
rect 707926 796610 708000 796666
rect 707800 796542 708000 796610
rect 707800 796486 707870 796542
rect 707926 796486 708000 796542
rect 707800 796418 708000 796486
rect 707800 796362 707870 796418
rect 707926 796362 708000 796418
rect 707800 796294 708000 796362
rect 707800 796238 707870 796294
rect 707926 796238 708000 796294
rect 707800 796170 708000 796238
rect 707800 796114 707870 796170
rect 707926 796114 708000 796170
rect 707800 796046 708000 796114
rect 707800 795990 707870 796046
rect 707926 795990 708000 796046
rect 707800 795922 708000 795990
rect 707800 795866 707870 795922
rect 707926 795866 708000 795922
rect 707800 795828 708000 795866
rect 707800 795178 708000 795248
rect 70000 795108 70200 795172
rect 70000 795052 70074 795108
rect 70130 795052 70200 795108
rect 70000 794984 70200 795052
rect 70000 794928 70074 794984
rect 70130 794928 70200 794984
rect 70000 794860 70200 794928
rect 70000 794804 70074 794860
rect 70130 794804 70200 794860
rect 70000 794736 70200 794804
rect 70000 794680 70074 794736
rect 70130 794680 70200 794736
rect 70000 794612 70200 794680
rect 70000 794556 70074 794612
rect 70130 794556 70200 794612
rect 70000 794488 70200 794556
rect 70000 794432 70074 794488
rect 70130 794432 70200 794488
rect 70000 794364 70200 794432
rect 70000 794308 70074 794364
rect 70130 794308 70200 794364
rect 70000 794240 70200 794308
rect 70000 794184 70074 794240
rect 70130 794184 70200 794240
rect 70000 794116 70200 794184
rect 70000 794060 70074 794116
rect 70130 794060 70200 794116
rect 70000 793992 70200 794060
rect 70000 793936 70074 793992
rect 70130 793936 70200 793992
rect 70000 793868 70200 793936
rect 70000 793812 70074 793868
rect 70130 793812 70200 793868
rect 70000 793744 70200 793812
rect 70000 793688 70074 793744
rect 70130 793688 70200 793744
rect 70000 793620 70200 793688
rect 70000 793564 70074 793620
rect 70130 793564 70200 793620
rect 70000 793496 70200 793564
rect 70000 793440 70074 793496
rect 70130 793440 70200 793496
rect 70000 793372 70200 793440
rect 70000 793316 70074 793372
rect 70130 793316 70200 793372
rect 70000 793248 70200 793316
rect 70000 793192 70074 793248
rect 70130 793192 70200 793248
rect 707800 795122 707870 795178
rect 707926 795122 708000 795178
rect 707800 795054 708000 795122
rect 707800 794998 707870 795054
rect 707926 794998 708000 795054
rect 707800 794930 708000 794998
rect 707800 794874 707870 794930
rect 707926 794874 708000 794930
rect 707800 794806 708000 794874
rect 707800 794750 707870 794806
rect 707926 794750 708000 794806
rect 707800 794682 708000 794750
rect 707800 794626 707870 794682
rect 707926 794626 708000 794682
rect 707800 794558 708000 794626
rect 707800 794502 707870 794558
rect 707926 794502 708000 794558
rect 707800 794434 708000 794502
rect 707800 794378 707870 794434
rect 707926 794378 708000 794434
rect 707800 794310 708000 794378
rect 707800 794254 707870 794310
rect 707926 794254 708000 794310
rect 707800 794186 708000 794254
rect 707800 794130 707870 794186
rect 707926 794130 708000 794186
rect 707800 794062 708000 794130
rect 707800 794006 707870 794062
rect 707926 794006 708000 794062
rect 707800 793938 708000 794006
rect 707800 793882 707870 793938
rect 707926 793882 708000 793938
rect 707800 793814 708000 793882
rect 707800 793758 707870 793814
rect 707926 793758 708000 793814
rect 707800 793690 708000 793758
rect 707800 793634 707870 793690
rect 707926 793634 708000 793690
rect 707800 793566 708000 793634
rect 707800 793510 707870 793566
rect 707926 793510 708000 793566
rect 707800 793442 708000 793510
rect 707800 793386 707870 793442
rect 707926 793386 708000 793442
rect 707800 793318 708000 793386
rect 707800 793262 707870 793318
rect 707926 793262 708000 793318
rect 707800 793198 708000 793262
rect 70000 793122 70200 793192
rect 707800 792808 708000 792878
rect 70000 792738 70200 792802
rect 70000 792682 70074 792738
rect 70130 792682 70200 792738
rect 70000 792614 70200 792682
rect 70000 792558 70074 792614
rect 70130 792558 70200 792614
rect 70000 792490 70200 792558
rect 70000 792434 70074 792490
rect 70130 792434 70200 792490
rect 70000 792366 70200 792434
rect 70000 792310 70074 792366
rect 70130 792310 70200 792366
rect 70000 792242 70200 792310
rect 70000 792186 70074 792242
rect 70130 792186 70200 792242
rect 70000 792118 70200 792186
rect 70000 792062 70074 792118
rect 70130 792062 70200 792118
rect 70000 791994 70200 792062
rect 70000 791938 70074 791994
rect 70130 791938 70200 791994
rect 70000 791870 70200 791938
rect 70000 791814 70074 791870
rect 70130 791814 70200 791870
rect 70000 791746 70200 791814
rect 70000 791690 70074 791746
rect 70130 791690 70200 791746
rect 70000 791622 70200 791690
rect 70000 791566 70074 791622
rect 70130 791566 70200 791622
rect 70000 791498 70200 791566
rect 70000 791442 70074 791498
rect 70130 791442 70200 791498
rect 70000 791374 70200 791442
rect 70000 791318 70074 791374
rect 70130 791318 70200 791374
rect 70000 791250 70200 791318
rect 70000 791194 70074 791250
rect 70130 791194 70200 791250
rect 70000 791126 70200 791194
rect 70000 791070 70074 791126
rect 70130 791070 70200 791126
rect 70000 791002 70200 791070
rect 70000 790946 70074 791002
rect 70130 790946 70200 791002
rect 70000 790878 70200 790946
rect 70000 790822 70074 790878
rect 70130 790822 70200 790878
rect 707800 792752 707870 792808
rect 707926 792752 708000 792808
rect 707800 792684 708000 792752
rect 707800 792628 707870 792684
rect 707926 792628 708000 792684
rect 707800 792560 708000 792628
rect 707800 792504 707870 792560
rect 707926 792504 708000 792560
rect 707800 792436 708000 792504
rect 707800 792380 707870 792436
rect 707926 792380 708000 792436
rect 707800 792312 708000 792380
rect 707800 792256 707870 792312
rect 707926 792256 708000 792312
rect 707800 792188 708000 792256
rect 707800 792132 707870 792188
rect 707926 792132 708000 792188
rect 707800 792064 708000 792132
rect 707800 792008 707870 792064
rect 707926 792008 708000 792064
rect 707800 791940 708000 792008
rect 707800 791884 707870 791940
rect 707926 791884 708000 791940
rect 707800 791816 708000 791884
rect 707800 791760 707870 791816
rect 707926 791760 708000 791816
rect 707800 791692 708000 791760
rect 707800 791636 707870 791692
rect 707926 791636 708000 791692
rect 707800 791568 708000 791636
rect 707800 791512 707870 791568
rect 707926 791512 708000 791568
rect 707800 791444 708000 791512
rect 707800 791388 707870 791444
rect 707926 791388 708000 791444
rect 707800 791320 708000 791388
rect 707800 791264 707870 791320
rect 707926 791264 708000 791320
rect 707800 791196 708000 791264
rect 707800 791140 707870 791196
rect 707926 791140 708000 791196
rect 707800 791072 708000 791140
rect 707800 791016 707870 791072
rect 707926 791016 708000 791072
rect 707800 790948 708000 791016
rect 707800 790892 707870 790948
rect 707926 790892 708000 790948
rect 707800 790828 708000 790892
rect 70000 790752 70200 790822
rect 70000 790134 70200 790172
rect 70000 790078 70074 790134
rect 70130 790078 70200 790134
rect 70000 790010 70200 790078
rect 70000 789954 70074 790010
rect 70130 789954 70200 790010
rect 70000 789886 70200 789954
rect 70000 789830 70074 789886
rect 70130 789830 70200 789886
rect 70000 789762 70200 789830
rect 70000 789706 70074 789762
rect 70130 789706 70200 789762
rect 70000 789638 70200 789706
rect 70000 789582 70074 789638
rect 70130 789582 70200 789638
rect 70000 789514 70200 789582
rect 70000 789458 70074 789514
rect 70130 789458 70200 789514
rect 70000 789390 70200 789458
rect 70000 789334 70074 789390
rect 70130 789334 70200 789390
rect 70000 789266 70200 789334
rect 70000 789210 70074 789266
rect 70130 789210 70200 789266
rect 70000 789142 70200 789210
rect 70000 789086 70074 789142
rect 70130 789086 70200 789142
rect 70000 789018 70200 789086
rect 70000 788962 70074 789018
rect 70130 788962 70200 789018
rect 70000 788894 70200 788962
rect 70000 788838 70074 788894
rect 70130 788838 70200 788894
rect 70000 788770 70200 788838
rect 70000 788714 70074 788770
rect 70130 788714 70200 788770
rect 70000 788646 70200 788714
rect 70000 788590 70074 788646
rect 70130 788590 70200 788646
rect 70000 788522 70200 788590
rect 70000 788466 70074 788522
rect 70130 788466 70200 788522
rect 70000 788398 70200 788466
rect 70000 788342 70074 788398
rect 70130 788342 70200 788398
rect 70000 788272 70200 788342
rect 707800 790102 708000 790172
rect 707800 790046 707870 790102
rect 707926 790046 708000 790102
rect 707800 789978 708000 790046
rect 707800 789922 707870 789978
rect 707926 789922 708000 789978
rect 707800 789854 708000 789922
rect 707800 789798 707870 789854
rect 707926 789798 708000 789854
rect 707800 789730 708000 789798
rect 707800 789674 707870 789730
rect 707926 789674 708000 789730
rect 707800 789606 708000 789674
rect 707800 789550 707870 789606
rect 707926 789550 708000 789606
rect 707800 789482 708000 789550
rect 707800 789426 707870 789482
rect 707926 789426 708000 789482
rect 707800 789358 708000 789426
rect 707800 789302 707870 789358
rect 707926 789302 708000 789358
rect 707800 789234 708000 789302
rect 707800 789178 707870 789234
rect 707926 789178 708000 789234
rect 707800 789110 708000 789178
rect 707800 789054 707870 789110
rect 707926 789054 708000 789110
rect 707800 788986 708000 789054
rect 707800 788930 707870 788986
rect 707926 788930 708000 788986
rect 707800 788862 708000 788930
rect 707800 788806 707870 788862
rect 707926 788806 708000 788862
rect 707800 788738 708000 788806
rect 707800 788682 707870 788738
rect 707926 788682 708000 788738
rect 707800 788614 708000 788682
rect 707800 788558 707870 788614
rect 707926 788558 708000 788614
rect 707800 788490 708000 788558
rect 707800 788434 707870 788490
rect 707926 788434 708000 788490
rect 707800 788366 708000 788434
rect 707800 788310 707870 788366
rect 707926 788310 708000 788366
rect 707800 788242 708000 788310
rect 707800 788186 707870 788242
rect 707926 788186 708000 788242
rect 707800 788122 708000 788186
rect 707800 787732 708000 787802
rect 707800 787676 707870 787732
rect 707926 787676 708000 787732
rect 707800 787608 708000 787676
rect 707800 787552 707870 787608
rect 707926 787552 708000 787608
rect 707800 787484 708000 787552
rect 707800 787428 707870 787484
rect 707926 787428 708000 787484
rect 707800 787360 708000 787428
rect 707800 787304 707870 787360
rect 707926 787304 708000 787360
rect 707800 787236 708000 787304
rect 707800 787180 707870 787236
rect 707926 787180 708000 787236
rect 707800 787112 708000 787180
rect 707800 787056 707870 787112
rect 707926 787056 708000 787112
rect 707800 786988 708000 787056
rect 707800 786932 707870 786988
rect 707926 786932 708000 786988
rect 707800 786864 708000 786932
rect 707800 786808 707870 786864
rect 707926 786808 708000 786864
rect 707800 786740 708000 786808
rect 707800 786684 707870 786740
rect 707926 786684 708000 786740
rect 707800 786616 708000 786684
rect 707800 786560 707870 786616
rect 707926 786560 708000 786616
rect 707800 786492 708000 786560
rect 707800 786436 707870 786492
rect 707926 786436 708000 786492
rect 707800 786368 708000 786436
rect 707800 786312 707870 786368
rect 707926 786312 708000 786368
rect 707800 786244 708000 786312
rect 707800 786188 707870 786244
rect 707926 786188 708000 786244
rect 707800 786120 708000 786188
rect 707800 786064 707870 786120
rect 707926 786064 708000 786120
rect 707800 785996 708000 786064
rect 707800 785940 707870 785996
rect 707926 785940 708000 785996
rect 707800 785872 708000 785940
rect 707800 785816 707870 785872
rect 707926 785816 708000 785872
rect 707800 785752 708000 785816
rect 707800 785134 708000 785172
rect 707800 785078 707870 785134
rect 707926 785078 708000 785134
rect 707800 785010 708000 785078
rect 707800 784954 707870 785010
rect 707926 784954 708000 785010
rect 707800 784886 708000 784954
rect 707800 784830 707870 784886
rect 707926 784830 708000 784886
rect 707800 784762 708000 784830
rect 707800 784706 707870 784762
rect 707926 784706 708000 784762
rect 707800 784638 708000 784706
rect 707800 784582 707870 784638
rect 707926 784582 708000 784638
rect 707800 784514 708000 784582
rect 707800 784458 707870 784514
rect 707926 784458 708000 784514
rect 707800 784390 708000 784458
rect 707800 784334 707870 784390
rect 707926 784334 708000 784390
rect 707800 784266 708000 784334
rect 707800 784210 707870 784266
rect 707926 784210 708000 784266
rect 707800 784142 708000 784210
rect 707800 784086 707870 784142
rect 707926 784086 708000 784142
rect 707800 784018 708000 784086
rect 707800 783962 707870 784018
rect 707926 783962 708000 784018
rect 707800 783894 708000 783962
rect 707800 783838 707870 783894
rect 707926 783838 708000 783894
rect 707800 783770 708000 783838
rect 707800 783714 707870 783770
rect 707926 783714 708000 783770
rect 707800 783646 708000 783714
rect 707800 783590 707870 783646
rect 707926 783590 708000 783646
rect 707800 783522 708000 783590
rect 707800 783466 707870 783522
rect 707926 783466 708000 783522
rect 707800 783398 708000 783466
rect 707800 783342 707870 783398
rect 707926 783342 708000 783398
rect 707800 783272 708000 783342
rect 707800 496658 708000 496728
rect 707800 496602 707870 496658
rect 707926 496602 708000 496658
rect 707800 496534 708000 496602
rect 707800 496478 707870 496534
rect 707926 496478 708000 496534
rect 707800 496410 708000 496478
rect 707800 496354 707870 496410
rect 707926 496354 708000 496410
rect 707800 496286 708000 496354
rect 707800 496230 707870 496286
rect 707926 496230 708000 496286
rect 707800 496162 708000 496230
rect 707800 496106 707870 496162
rect 707926 496106 708000 496162
rect 707800 496038 708000 496106
rect 707800 495982 707870 496038
rect 707926 495982 708000 496038
rect 707800 495914 708000 495982
rect 707800 495858 707870 495914
rect 707926 495858 708000 495914
rect 707800 495790 708000 495858
rect 707800 495734 707870 495790
rect 707926 495734 708000 495790
rect 707800 495666 708000 495734
rect 707800 495610 707870 495666
rect 707926 495610 708000 495666
rect 707800 495542 708000 495610
rect 707800 495486 707870 495542
rect 707926 495486 708000 495542
rect 707800 495418 708000 495486
rect 707800 495362 707870 495418
rect 707926 495362 708000 495418
rect 707800 495294 708000 495362
rect 707800 495238 707870 495294
rect 707926 495238 708000 495294
rect 707800 495170 708000 495238
rect 707800 495114 707870 495170
rect 707926 495114 708000 495170
rect 707800 495046 708000 495114
rect 707800 494990 707870 495046
rect 707926 494990 708000 495046
rect 707800 494922 708000 494990
rect 707800 494866 707870 494922
rect 707926 494866 708000 494922
rect 707800 494828 708000 494866
rect 707800 494178 708000 494248
rect 707800 494122 707870 494178
rect 707926 494122 708000 494178
rect 707800 494054 708000 494122
rect 707800 493998 707870 494054
rect 707926 493998 708000 494054
rect 707800 493930 708000 493998
rect 707800 493874 707870 493930
rect 707926 493874 708000 493930
rect 707800 493806 708000 493874
rect 707800 493750 707870 493806
rect 707926 493750 708000 493806
rect 707800 493682 708000 493750
rect 707800 493626 707870 493682
rect 707926 493626 708000 493682
rect 707800 493558 708000 493626
rect 707800 493502 707870 493558
rect 707926 493502 708000 493558
rect 707800 493434 708000 493502
rect 707800 493378 707870 493434
rect 707926 493378 708000 493434
rect 707800 493310 708000 493378
rect 707800 493254 707870 493310
rect 707926 493254 708000 493310
rect 707800 493186 708000 493254
rect 707800 493130 707870 493186
rect 707926 493130 708000 493186
rect 707800 493062 708000 493130
rect 707800 493006 707870 493062
rect 707926 493006 708000 493062
rect 707800 492938 708000 493006
rect 707800 492882 707870 492938
rect 707926 492882 708000 492938
rect 707800 492814 708000 492882
rect 707800 492758 707870 492814
rect 707926 492758 708000 492814
rect 707800 492690 708000 492758
rect 707800 492634 707870 492690
rect 707926 492634 708000 492690
rect 707800 492566 708000 492634
rect 707800 492510 707870 492566
rect 707926 492510 708000 492566
rect 707800 492442 708000 492510
rect 707800 492386 707870 492442
rect 707926 492386 708000 492442
rect 707800 492318 708000 492386
rect 707800 492262 707870 492318
rect 707926 492262 708000 492318
rect 707800 492198 708000 492262
rect 707800 491808 708000 491878
rect 707800 491752 707870 491808
rect 707926 491752 708000 491808
rect 707800 491684 708000 491752
rect 707800 491628 707870 491684
rect 707926 491628 708000 491684
rect 707800 491560 708000 491628
rect 707800 491504 707870 491560
rect 707926 491504 708000 491560
rect 707800 491436 708000 491504
rect 707800 491380 707870 491436
rect 707926 491380 708000 491436
rect 707800 491312 708000 491380
rect 707800 491256 707870 491312
rect 707926 491256 708000 491312
rect 707800 491188 708000 491256
rect 707800 491132 707870 491188
rect 707926 491132 708000 491188
rect 707800 491064 708000 491132
rect 707800 491008 707870 491064
rect 707926 491008 708000 491064
rect 707800 490940 708000 491008
rect 707800 490884 707870 490940
rect 707926 490884 708000 490940
rect 707800 490816 708000 490884
rect 707800 490760 707870 490816
rect 707926 490760 708000 490816
rect 707800 490692 708000 490760
rect 707800 490636 707870 490692
rect 707926 490636 708000 490692
rect 707800 490568 708000 490636
rect 707800 490512 707870 490568
rect 707926 490512 708000 490568
rect 707800 490444 708000 490512
rect 707800 490388 707870 490444
rect 707926 490388 708000 490444
rect 707800 490320 708000 490388
rect 707800 490264 707870 490320
rect 707926 490264 708000 490320
rect 707800 490196 708000 490264
rect 707800 490140 707870 490196
rect 707926 490140 708000 490196
rect 707800 490072 708000 490140
rect 707800 490016 707870 490072
rect 707926 490016 708000 490072
rect 707800 489948 708000 490016
rect 707800 489892 707870 489948
rect 707926 489892 708000 489948
rect 707800 489828 708000 489892
rect 707800 489102 708000 489172
rect 707800 489046 707870 489102
rect 707926 489046 708000 489102
rect 707800 488978 708000 489046
rect 707800 488922 707870 488978
rect 707926 488922 708000 488978
rect 707800 488854 708000 488922
rect 707800 488798 707870 488854
rect 707926 488798 708000 488854
rect 707800 488730 708000 488798
rect 707800 488674 707870 488730
rect 707926 488674 708000 488730
rect 707800 488606 708000 488674
rect 707800 488550 707870 488606
rect 707926 488550 708000 488606
rect 707800 488482 708000 488550
rect 707800 488426 707870 488482
rect 707926 488426 708000 488482
rect 707800 488358 708000 488426
rect 707800 488302 707870 488358
rect 707926 488302 708000 488358
rect 707800 488234 708000 488302
rect 707800 488178 707870 488234
rect 707926 488178 708000 488234
rect 707800 488110 708000 488178
rect 707800 488054 707870 488110
rect 707926 488054 708000 488110
rect 707800 487986 708000 488054
rect 707800 487930 707870 487986
rect 707926 487930 708000 487986
rect 707800 487862 708000 487930
rect 707800 487806 707870 487862
rect 707926 487806 708000 487862
rect 707800 487738 708000 487806
rect 707800 487682 707870 487738
rect 707926 487682 708000 487738
rect 707800 487614 708000 487682
rect 707800 487558 707870 487614
rect 707926 487558 708000 487614
rect 707800 487490 708000 487558
rect 707800 487434 707870 487490
rect 707926 487434 708000 487490
rect 707800 487366 708000 487434
rect 707800 487310 707870 487366
rect 707926 487310 708000 487366
rect 707800 487242 708000 487310
rect 707800 487186 707870 487242
rect 707926 487186 708000 487242
rect 707800 487122 708000 487186
rect 707800 486732 708000 486802
rect 707800 486676 707870 486732
rect 707926 486676 708000 486732
rect 707800 486608 708000 486676
rect 707800 486552 707870 486608
rect 707926 486552 708000 486608
rect 707800 486484 708000 486552
rect 707800 486428 707870 486484
rect 707926 486428 708000 486484
rect 707800 486360 708000 486428
rect 707800 486304 707870 486360
rect 707926 486304 708000 486360
rect 707800 486236 708000 486304
rect 707800 486180 707870 486236
rect 707926 486180 708000 486236
rect 707800 486112 708000 486180
rect 707800 486056 707870 486112
rect 707926 486056 708000 486112
rect 707800 485988 708000 486056
rect 707800 485932 707870 485988
rect 707926 485932 708000 485988
rect 707800 485864 708000 485932
rect 707800 485808 707870 485864
rect 707926 485808 708000 485864
rect 707800 485740 708000 485808
rect 707800 485684 707870 485740
rect 707926 485684 708000 485740
rect 707800 485616 708000 485684
rect 707800 485560 707870 485616
rect 707926 485560 708000 485616
rect 707800 485492 708000 485560
rect 707800 485436 707870 485492
rect 707926 485436 708000 485492
rect 707800 485368 708000 485436
rect 707800 485312 707870 485368
rect 707926 485312 708000 485368
rect 707800 485244 708000 485312
rect 707800 485188 707870 485244
rect 707926 485188 708000 485244
rect 707800 485120 708000 485188
rect 707800 485064 707870 485120
rect 707926 485064 708000 485120
rect 707800 484996 708000 485064
rect 707800 484940 707870 484996
rect 707926 484940 708000 484996
rect 707800 484872 708000 484940
rect 707800 484816 707870 484872
rect 707926 484816 708000 484872
rect 707800 484752 708000 484816
rect 707800 484134 708000 484172
rect 707800 484078 707870 484134
rect 707926 484078 708000 484134
rect 707800 484010 708000 484078
rect 707800 483954 707870 484010
rect 707926 483954 708000 484010
rect 707800 483886 708000 483954
rect 707800 483830 707870 483886
rect 707926 483830 708000 483886
rect 707800 483762 708000 483830
rect 707800 483706 707870 483762
rect 707926 483706 708000 483762
rect 707800 483638 708000 483706
rect 707800 483582 707870 483638
rect 707926 483582 708000 483638
rect 707800 483514 708000 483582
rect 707800 483458 707870 483514
rect 707926 483458 708000 483514
rect 707800 483390 708000 483458
rect 707800 483334 707870 483390
rect 707926 483334 708000 483390
rect 707800 483266 708000 483334
rect 707800 483210 707870 483266
rect 707926 483210 708000 483266
rect 707800 483142 708000 483210
rect 707800 483086 707870 483142
rect 707926 483086 708000 483142
rect 707800 483018 708000 483086
rect 707800 482962 707870 483018
rect 707926 482962 708000 483018
rect 707800 482894 708000 482962
rect 707800 482838 707870 482894
rect 707926 482838 708000 482894
rect 707800 482770 708000 482838
rect 707800 482714 707870 482770
rect 707926 482714 708000 482770
rect 707800 482646 708000 482714
rect 707800 482590 707870 482646
rect 707926 482590 708000 482646
rect 707800 482522 708000 482590
rect 707800 482466 707870 482522
rect 707926 482466 708000 482522
rect 707800 482398 708000 482466
rect 707800 482342 707870 482398
rect 707926 482342 708000 482398
rect 707800 482272 708000 482342
rect 70000 474658 70200 474728
rect 70000 474602 70074 474658
rect 70130 474602 70200 474658
rect 70000 474534 70200 474602
rect 70000 474478 70074 474534
rect 70130 474478 70200 474534
rect 70000 474410 70200 474478
rect 70000 474354 70074 474410
rect 70130 474354 70200 474410
rect 70000 474286 70200 474354
rect 70000 474230 70074 474286
rect 70130 474230 70200 474286
rect 70000 474162 70200 474230
rect 70000 474106 70074 474162
rect 70130 474106 70200 474162
rect 70000 474038 70200 474106
rect 70000 473982 70074 474038
rect 70130 473982 70200 474038
rect 70000 473914 70200 473982
rect 70000 473858 70074 473914
rect 70130 473858 70200 473914
rect 70000 473790 70200 473858
rect 70000 473734 70074 473790
rect 70130 473734 70200 473790
rect 70000 473666 70200 473734
rect 70000 473610 70074 473666
rect 70130 473610 70200 473666
rect 70000 473542 70200 473610
rect 70000 473486 70074 473542
rect 70130 473486 70200 473542
rect 70000 473418 70200 473486
rect 70000 473362 70074 473418
rect 70130 473362 70200 473418
rect 70000 473294 70200 473362
rect 70000 473238 70074 473294
rect 70130 473238 70200 473294
rect 70000 473170 70200 473238
rect 70000 473114 70074 473170
rect 70130 473114 70200 473170
rect 70000 473046 70200 473114
rect 70000 472990 70074 473046
rect 70130 472990 70200 473046
rect 70000 472922 70200 472990
rect 70000 472866 70074 472922
rect 70130 472866 70200 472922
rect 70000 472828 70200 472866
rect 70000 472184 70200 472248
rect 70000 472128 70074 472184
rect 70130 472128 70200 472184
rect 70000 472060 70200 472128
rect 70000 472004 70074 472060
rect 70130 472004 70200 472060
rect 70000 471936 70200 472004
rect 70000 471880 70074 471936
rect 70130 471880 70200 471936
rect 70000 471812 70200 471880
rect 70000 471756 70074 471812
rect 70130 471756 70200 471812
rect 70000 471688 70200 471756
rect 70000 471632 70074 471688
rect 70130 471632 70200 471688
rect 70000 471564 70200 471632
rect 70000 471508 70074 471564
rect 70130 471508 70200 471564
rect 70000 471440 70200 471508
rect 70000 471384 70074 471440
rect 70130 471384 70200 471440
rect 70000 471316 70200 471384
rect 70000 471260 70074 471316
rect 70130 471260 70200 471316
rect 70000 471192 70200 471260
rect 70000 471136 70074 471192
rect 70130 471136 70200 471192
rect 70000 471068 70200 471136
rect 70000 471012 70074 471068
rect 70130 471012 70200 471068
rect 70000 470944 70200 471012
rect 70000 470888 70074 470944
rect 70130 470888 70200 470944
rect 70000 470820 70200 470888
rect 70000 470764 70074 470820
rect 70130 470764 70200 470820
rect 70000 470696 70200 470764
rect 70000 470640 70074 470696
rect 70130 470640 70200 470696
rect 70000 470572 70200 470640
rect 70000 470516 70074 470572
rect 70130 470516 70200 470572
rect 70000 470448 70200 470516
rect 70000 470392 70074 470448
rect 70130 470392 70200 470448
rect 70000 470324 70200 470392
rect 70000 470268 70074 470324
rect 70130 470268 70200 470324
rect 70000 470198 70200 470268
rect 70000 469814 70200 469878
rect 70000 469758 70074 469814
rect 70130 469758 70200 469814
rect 70000 469690 70200 469758
rect 70000 469634 70074 469690
rect 70130 469634 70200 469690
rect 70000 469566 70200 469634
rect 70000 469510 70074 469566
rect 70130 469510 70200 469566
rect 70000 469442 70200 469510
rect 70000 469386 70074 469442
rect 70130 469386 70200 469442
rect 70000 469318 70200 469386
rect 70000 469262 70074 469318
rect 70130 469262 70200 469318
rect 70000 469194 70200 469262
rect 70000 469138 70074 469194
rect 70130 469138 70200 469194
rect 70000 469070 70200 469138
rect 70000 469014 70074 469070
rect 70130 469014 70200 469070
rect 70000 468946 70200 469014
rect 70000 468890 70074 468946
rect 70130 468890 70200 468946
rect 70000 468822 70200 468890
rect 70000 468766 70074 468822
rect 70130 468766 70200 468822
rect 70000 468698 70200 468766
rect 70000 468642 70074 468698
rect 70130 468642 70200 468698
rect 70000 468574 70200 468642
rect 70000 468518 70074 468574
rect 70130 468518 70200 468574
rect 70000 468450 70200 468518
rect 70000 468394 70074 468450
rect 70130 468394 70200 468450
rect 70000 468326 70200 468394
rect 70000 468270 70074 468326
rect 70130 468270 70200 468326
rect 70000 468202 70200 468270
rect 70000 468146 70074 468202
rect 70130 468146 70200 468202
rect 70000 468078 70200 468146
rect 70000 468022 70074 468078
rect 70130 468022 70200 468078
rect 70000 467954 70200 468022
rect 70000 467898 70074 467954
rect 70130 467898 70200 467954
rect 70000 467828 70200 467898
rect 70000 467108 70200 467172
rect 70000 467052 70074 467108
rect 70130 467052 70200 467108
rect 70000 466984 70200 467052
rect 70000 466928 70074 466984
rect 70130 466928 70200 466984
rect 70000 466860 70200 466928
rect 70000 466804 70074 466860
rect 70130 466804 70200 466860
rect 70000 466736 70200 466804
rect 70000 466680 70074 466736
rect 70130 466680 70200 466736
rect 70000 466612 70200 466680
rect 70000 466556 70074 466612
rect 70130 466556 70200 466612
rect 70000 466488 70200 466556
rect 70000 466432 70074 466488
rect 70130 466432 70200 466488
rect 70000 466364 70200 466432
rect 70000 466308 70074 466364
rect 70130 466308 70200 466364
rect 70000 466240 70200 466308
rect 70000 466184 70074 466240
rect 70130 466184 70200 466240
rect 70000 466116 70200 466184
rect 70000 466060 70074 466116
rect 70130 466060 70200 466116
rect 70000 465992 70200 466060
rect 70000 465936 70074 465992
rect 70130 465936 70200 465992
rect 70000 465868 70200 465936
rect 70000 465812 70074 465868
rect 70130 465812 70200 465868
rect 70000 465744 70200 465812
rect 70000 465688 70074 465744
rect 70130 465688 70200 465744
rect 70000 465620 70200 465688
rect 70000 465564 70074 465620
rect 70130 465564 70200 465620
rect 70000 465496 70200 465564
rect 70000 465440 70074 465496
rect 70130 465440 70200 465496
rect 70000 465372 70200 465440
rect 70000 465316 70074 465372
rect 70130 465316 70200 465372
rect 70000 465248 70200 465316
rect 70000 465192 70074 465248
rect 70130 465192 70200 465248
rect 70000 465122 70200 465192
rect 70000 464738 70200 464802
rect 70000 464682 70074 464738
rect 70130 464682 70200 464738
rect 70000 464614 70200 464682
rect 70000 464558 70074 464614
rect 70130 464558 70200 464614
rect 70000 464490 70200 464558
rect 70000 464434 70074 464490
rect 70130 464434 70200 464490
rect 70000 464366 70200 464434
rect 70000 464310 70074 464366
rect 70130 464310 70200 464366
rect 70000 464242 70200 464310
rect 70000 464186 70074 464242
rect 70130 464186 70200 464242
rect 70000 464118 70200 464186
rect 70000 464062 70074 464118
rect 70130 464062 70200 464118
rect 70000 463994 70200 464062
rect 70000 463938 70074 463994
rect 70130 463938 70200 463994
rect 70000 463870 70200 463938
rect 70000 463814 70074 463870
rect 70130 463814 70200 463870
rect 70000 463746 70200 463814
rect 70000 463690 70074 463746
rect 70130 463690 70200 463746
rect 70000 463622 70200 463690
rect 70000 463566 70074 463622
rect 70130 463566 70200 463622
rect 70000 463498 70200 463566
rect 70000 463442 70074 463498
rect 70130 463442 70200 463498
rect 70000 463374 70200 463442
rect 70000 463318 70074 463374
rect 70130 463318 70200 463374
rect 70000 463250 70200 463318
rect 70000 463194 70074 463250
rect 70130 463194 70200 463250
rect 70000 463126 70200 463194
rect 70000 463070 70074 463126
rect 70130 463070 70200 463126
rect 70000 463002 70200 463070
rect 70000 462946 70074 463002
rect 70130 462946 70200 463002
rect 70000 462878 70200 462946
rect 70000 462822 70074 462878
rect 70130 462822 70200 462878
rect 70000 462752 70200 462822
rect 70000 462134 70200 462172
rect 70000 462078 70074 462134
rect 70130 462078 70200 462134
rect 70000 462010 70200 462078
rect 70000 461954 70074 462010
rect 70130 461954 70200 462010
rect 70000 461886 70200 461954
rect 70000 461830 70074 461886
rect 70130 461830 70200 461886
rect 70000 461762 70200 461830
rect 70000 461706 70074 461762
rect 70130 461706 70200 461762
rect 70000 461638 70200 461706
rect 70000 461582 70074 461638
rect 70130 461582 70200 461638
rect 70000 461514 70200 461582
rect 70000 461458 70074 461514
rect 70130 461458 70200 461514
rect 70000 461390 70200 461458
rect 70000 461334 70074 461390
rect 70130 461334 70200 461390
rect 70000 461266 70200 461334
rect 70000 461210 70074 461266
rect 70130 461210 70200 461266
rect 70000 461142 70200 461210
rect 70000 461086 70074 461142
rect 70130 461086 70200 461142
rect 70000 461018 70200 461086
rect 70000 460962 70074 461018
rect 70130 460962 70200 461018
rect 70000 460894 70200 460962
rect 70000 460838 70074 460894
rect 70130 460838 70200 460894
rect 70000 460770 70200 460838
rect 70000 460714 70074 460770
rect 70130 460714 70200 460770
rect 70000 460646 70200 460714
rect 70000 460590 70074 460646
rect 70130 460590 70200 460646
rect 70000 460522 70200 460590
rect 70000 460466 70074 460522
rect 70130 460466 70200 460522
rect 70000 460398 70200 460466
rect 70000 460342 70074 460398
rect 70130 460342 70200 460398
rect 70000 460272 70200 460342
rect 707801 453658 708001 453728
rect 707801 453602 707870 453658
rect 707926 453602 708001 453658
rect 707801 453534 708001 453602
rect 707801 453478 707870 453534
rect 707926 453478 708001 453534
rect 707801 453410 708001 453478
rect 707801 453354 707870 453410
rect 707926 453354 708001 453410
rect 707801 453286 708001 453354
rect 707801 453230 707870 453286
rect 707926 453230 708001 453286
rect 707801 453162 708001 453230
rect 707801 453106 707870 453162
rect 707926 453106 708001 453162
rect 707801 453038 708001 453106
rect 707801 452982 707870 453038
rect 707926 452982 708001 453038
rect 707801 452914 708001 452982
rect 707801 452858 707870 452914
rect 707926 452858 708001 452914
rect 707801 452790 708001 452858
rect 707801 452734 707870 452790
rect 707926 452734 708001 452790
rect 707801 452666 708001 452734
rect 707801 452610 707870 452666
rect 707926 452610 708001 452666
rect 707801 452542 708001 452610
rect 707801 452486 707870 452542
rect 707926 452486 708001 452542
rect 707801 452418 708001 452486
rect 707801 452362 707870 452418
rect 707926 452362 708001 452418
rect 707801 452294 708001 452362
rect 707801 452238 707870 452294
rect 707926 452238 708001 452294
rect 707801 452170 708001 452238
rect 707801 452114 707870 452170
rect 707926 452114 708001 452170
rect 707801 452046 708001 452114
rect 707801 451990 707870 452046
rect 707926 451990 708001 452046
rect 707801 451922 708001 451990
rect 707801 451866 707870 451922
rect 707926 451866 708001 451922
rect 707801 451828 708001 451866
rect 707801 451178 708001 451248
rect 707801 451122 707870 451178
rect 707926 451122 708001 451178
rect 707801 451054 708001 451122
rect 707801 450998 707870 451054
rect 707926 450998 708001 451054
rect 707801 450930 708001 450998
rect 707801 450874 707870 450930
rect 707926 450874 708001 450930
rect 707801 450806 708001 450874
rect 707801 450750 707870 450806
rect 707926 450750 708001 450806
rect 707801 450682 708001 450750
rect 707801 450626 707870 450682
rect 707926 450626 708001 450682
rect 707801 450558 708001 450626
rect 707801 450502 707870 450558
rect 707926 450502 708001 450558
rect 707801 450434 708001 450502
rect 707801 450378 707870 450434
rect 707926 450378 708001 450434
rect 707801 450310 708001 450378
rect 707801 450254 707870 450310
rect 707926 450254 708001 450310
rect 707801 450186 708001 450254
rect 707801 450130 707870 450186
rect 707926 450130 708001 450186
rect 707801 450062 708001 450130
rect 707801 450006 707870 450062
rect 707926 450006 708001 450062
rect 707801 449938 708001 450006
rect 707801 449882 707870 449938
rect 707926 449882 708001 449938
rect 707801 449814 708001 449882
rect 707801 449758 707870 449814
rect 707926 449758 708001 449814
rect 707801 449690 708001 449758
rect 707801 449634 707870 449690
rect 707926 449634 708001 449690
rect 707801 449566 708001 449634
rect 707801 449510 707870 449566
rect 707926 449510 708001 449566
rect 707801 449442 708001 449510
rect 707801 449386 707870 449442
rect 707926 449386 708001 449442
rect 707801 449318 708001 449386
rect 707801 449262 707870 449318
rect 707926 449262 708001 449318
rect 707801 449198 708001 449262
rect 707801 448808 708001 448878
rect 707801 448752 707870 448808
rect 707926 448752 708001 448808
rect 707801 448684 708001 448752
rect 707801 448628 707870 448684
rect 707926 448628 708001 448684
rect 707801 448560 708001 448628
rect 707801 448504 707870 448560
rect 707926 448504 708001 448560
rect 707801 448436 708001 448504
rect 707801 448380 707870 448436
rect 707926 448380 708001 448436
rect 707801 448312 708001 448380
rect 707801 448256 707870 448312
rect 707926 448256 708001 448312
rect 707801 448188 708001 448256
rect 707801 448132 707870 448188
rect 707926 448132 708001 448188
rect 707801 448064 708001 448132
rect 707801 448008 707870 448064
rect 707926 448008 708001 448064
rect 707801 447940 708001 448008
rect 707801 447884 707870 447940
rect 707926 447884 708001 447940
rect 707801 447816 708001 447884
rect 707801 447760 707870 447816
rect 707926 447760 708001 447816
rect 707801 447692 708001 447760
rect 707801 447636 707870 447692
rect 707926 447636 708001 447692
rect 707801 447568 708001 447636
rect 707801 447512 707870 447568
rect 707926 447512 708001 447568
rect 707801 447444 708001 447512
rect 707801 447388 707870 447444
rect 707926 447388 708001 447444
rect 707801 447320 708001 447388
rect 707801 447264 707870 447320
rect 707926 447264 708001 447320
rect 707801 447196 708001 447264
rect 707801 447140 707870 447196
rect 707926 447140 708001 447196
rect 707801 447072 708001 447140
rect 707801 447016 707870 447072
rect 707926 447016 708001 447072
rect 707801 446948 708001 447016
rect 707801 446892 707870 446948
rect 707926 446892 708001 446948
rect 707801 446828 708001 446892
rect 707801 446102 708001 446172
rect 707801 446046 707870 446102
rect 707926 446046 708001 446102
rect 707801 445978 708001 446046
rect 707801 445922 707870 445978
rect 707926 445922 708001 445978
rect 707801 445854 708001 445922
rect 707801 445798 707870 445854
rect 707926 445798 708001 445854
rect 707801 445730 708001 445798
rect 707801 445674 707870 445730
rect 707926 445674 708001 445730
rect 707801 445606 708001 445674
rect 707801 445550 707870 445606
rect 707926 445550 708001 445606
rect 707801 445482 708001 445550
rect 707801 445426 707870 445482
rect 707926 445426 708001 445482
rect 707801 445358 708001 445426
rect 707801 445302 707870 445358
rect 707926 445302 708001 445358
rect 707801 445234 708001 445302
rect 707801 445178 707870 445234
rect 707926 445178 708001 445234
rect 707801 445110 708001 445178
rect 707801 445054 707870 445110
rect 707926 445054 708001 445110
rect 707801 444986 708001 445054
rect 707801 444930 707870 444986
rect 707926 444930 708001 444986
rect 707801 444862 708001 444930
rect 707801 444806 707870 444862
rect 707926 444806 708001 444862
rect 707801 444738 708001 444806
rect 707801 444682 707870 444738
rect 707926 444682 708001 444738
rect 707801 444614 708001 444682
rect 707801 444558 707870 444614
rect 707926 444558 708001 444614
rect 707801 444490 708001 444558
rect 707801 444434 707870 444490
rect 707926 444434 708001 444490
rect 707801 444366 708001 444434
rect 707801 444310 707870 444366
rect 707926 444310 708001 444366
rect 707801 444242 708001 444310
rect 707801 444186 707870 444242
rect 707926 444186 708001 444242
rect 707801 444122 708001 444186
rect 707801 443732 708001 443802
rect 707801 443676 707870 443732
rect 707926 443676 708001 443732
rect 707801 443608 708001 443676
rect 707801 443552 707870 443608
rect 707926 443552 708001 443608
rect 707801 443484 708001 443552
rect 707801 443428 707870 443484
rect 707926 443428 708001 443484
rect 707801 443360 708001 443428
rect 707801 443304 707870 443360
rect 707926 443304 708001 443360
rect 707801 443236 708001 443304
rect 707801 443180 707870 443236
rect 707926 443180 708001 443236
rect 707801 443112 708001 443180
rect 707801 443056 707870 443112
rect 707926 443056 708001 443112
rect 707801 442988 708001 443056
rect 707801 442932 707870 442988
rect 707926 442932 708001 442988
rect 707801 442864 708001 442932
rect 707801 442808 707870 442864
rect 707926 442808 708001 442864
rect 707801 442740 708001 442808
rect 707801 442684 707870 442740
rect 707926 442684 708001 442740
rect 707801 442616 708001 442684
rect 707801 442560 707870 442616
rect 707926 442560 708001 442616
rect 707801 442492 708001 442560
rect 707801 442436 707870 442492
rect 707926 442436 708001 442492
rect 707801 442368 708001 442436
rect 707801 442312 707870 442368
rect 707926 442312 708001 442368
rect 707801 442244 708001 442312
rect 707801 442188 707870 442244
rect 707926 442188 708001 442244
rect 707801 442120 708001 442188
rect 707801 442064 707870 442120
rect 707926 442064 708001 442120
rect 707801 441996 708001 442064
rect 707801 441940 707870 441996
rect 707926 441940 708001 441996
rect 707801 441872 708001 441940
rect 707801 441816 707870 441872
rect 707926 441816 708001 441872
rect 707801 441752 708001 441816
rect 707801 441134 708001 441172
rect 707801 441078 707870 441134
rect 707926 441078 708001 441134
rect 707801 441010 708001 441078
rect 707801 440954 707870 441010
rect 707926 440954 708001 441010
rect 707801 440886 708001 440954
rect 707801 440830 707870 440886
rect 707926 440830 708001 440886
rect 707801 440762 708001 440830
rect 707801 440706 707870 440762
rect 707926 440706 708001 440762
rect 707801 440638 708001 440706
rect 707801 440582 707870 440638
rect 707926 440582 708001 440638
rect 707801 440514 708001 440582
rect 707801 440458 707870 440514
rect 707926 440458 708001 440514
rect 707801 440390 708001 440458
rect 707801 440334 707870 440390
rect 707926 440334 708001 440390
rect 707801 440266 708001 440334
rect 707801 440210 707870 440266
rect 707926 440210 708001 440266
rect 707801 440142 708001 440210
rect 707801 440086 707870 440142
rect 707926 440086 708001 440142
rect 707801 440018 708001 440086
rect 707801 439962 707870 440018
rect 707926 439962 708001 440018
rect 707801 439894 708001 439962
rect 707801 439838 707870 439894
rect 707926 439838 708001 439894
rect 707801 439770 708001 439838
rect 707801 439714 707870 439770
rect 707926 439714 708001 439770
rect 707801 439646 708001 439714
rect 707801 439590 707870 439646
rect 707926 439590 708001 439646
rect 707801 439522 708001 439590
rect 707801 439466 707870 439522
rect 707926 439466 708001 439522
rect 707801 439398 708001 439466
rect 707801 439342 707870 439398
rect 707926 439342 708001 439398
rect 707801 439272 708001 439342
rect 70000 433658 70200 433729
rect 70000 433602 70074 433658
rect 70130 433602 70200 433658
rect 70000 433534 70200 433602
rect 70000 433478 70074 433534
rect 70130 433478 70200 433534
rect 70000 433410 70200 433478
rect 70000 433354 70074 433410
rect 70130 433354 70200 433410
rect 70000 433286 70200 433354
rect 70000 433230 70074 433286
rect 70130 433230 70200 433286
rect 70000 433162 70200 433230
rect 70000 433106 70074 433162
rect 70130 433106 70200 433162
rect 70000 433038 70200 433106
rect 70000 432982 70074 433038
rect 70130 432982 70200 433038
rect 70000 432914 70200 432982
rect 70000 432858 70074 432914
rect 70130 432858 70200 432914
rect 70000 432790 70200 432858
rect 70000 432734 70074 432790
rect 70130 432734 70200 432790
rect 70000 432666 70200 432734
rect 70000 432610 70074 432666
rect 70130 432610 70200 432666
rect 70000 432542 70200 432610
rect 70000 432486 70074 432542
rect 70130 432486 70200 432542
rect 70000 432418 70200 432486
rect 70000 432362 70074 432418
rect 70130 432362 70200 432418
rect 70000 432294 70200 432362
rect 70000 432238 70074 432294
rect 70130 432238 70200 432294
rect 70000 432170 70200 432238
rect 70000 432114 70074 432170
rect 70130 432114 70200 432170
rect 70000 432046 70200 432114
rect 70000 431990 70074 432046
rect 70130 431990 70200 432046
rect 70000 431922 70200 431990
rect 70000 431866 70074 431922
rect 70130 431866 70200 431922
rect 70000 431829 70200 431866
rect 70000 431184 70200 431249
rect 70000 431128 70074 431184
rect 70130 431128 70200 431184
rect 70000 431060 70200 431128
rect 70000 431004 70074 431060
rect 70130 431004 70200 431060
rect 70000 430936 70200 431004
rect 70000 430880 70074 430936
rect 70130 430880 70200 430936
rect 70000 430812 70200 430880
rect 70000 430756 70074 430812
rect 70130 430756 70200 430812
rect 70000 430688 70200 430756
rect 70000 430632 70074 430688
rect 70130 430632 70200 430688
rect 70000 430564 70200 430632
rect 70000 430508 70074 430564
rect 70130 430508 70200 430564
rect 70000 430440 70200 430508
rect 70000 430384 70074 430440
rect 70130 430384 70200 430440
rect 70000 430316 70200 430384
rect 70000 430260 70074 430316
rect 70130 430260 70200 430316
rect 70000 430192 70200 430260
rect 70000 430136 70074 430192
rect 70130 430136 70200 430192
rect 70000 430068 70200 430136
rect 70000 430012 70074 430068
rect 70130 430012 70200 430068
rect 70000 429944 70200 430012
rect 70000 429888 70074 429944
rect 70130 429888 70200 429944
rect 70000 429820 70200 429888
rect 70000 429764 70074 429820
rect 70130 429764 70200 429820
rect 70000 429696 70200 429764
rect 70000 429640 70074 429696
rect 70130 429640 70200 429696
rect 70000 429572 70200 429640
rect 70000 429516 70074 429572
rect 70130 429516 70200 429572
rect 70000 429448 70200 429516
rect 70000 429392 70074 429448
rect 70130 429392 70200 429448
rect 70000 429324 70200 429392
rect 70000 429268 70074 429324
rect 70130 429268 70200 429324
rect 70000 429199 70200 429268
rect 70000 428814 70200 428879
rect 70000 428758 70074 428814
rect 70130 428758 70200 428814
rect 70000 428690 70200 428758
rect 70000 428634 70074 428690
rect 70130 428634 70200 428690
rect 70000 428566 70200 428634
rect 70000 428510 70074 428566
rect 70130 428510 70200 428566
rect 70000 428442 70200 428510
rect 70000 428386 70074 428442
rect 70130 428386 70200 428442
rect 70000 428318 70200 428386
rect 70000 428262 70074 428318
rect 70130 428262 70200 428318
rect 70000 428194 70200 428262
rect 70000 428138 70074 428194
rect 70130 428138 70200 428194
rect 70000 428070 70200 428138
rect 70000 428014 70074 428070
rect 70130 428014 70200 428070
rect 70000 427946 70200 428014
rect 70000 427890 70074 427946
rect 70130 427890 70200 427946
rect 70000 427822 70200 427890
rect 70000 427766 70074 427822
rect 70130 427766 70200 427822
rect 70000 427698 70200 427766
rect 70000 427642 70074 427698
rect 70130 427642 70200 427698
rect 70000 427574 70200 427642
rect 70000 427518 70074 427574
rect 70130 427518 70200 427574
rect 70000 427450 70200 427518
rect 70000 427394 70074 427450
rect 70130 427394 70200 427450
rect 70000 427326 70200 427394
rect 70000 427270 70074 427326
rect 70130 427270 70200 427326
rect 70000 427202 70200 427270
rect 70000 427146 70074 427202
rect 70130 427146 70200 427202
rect 70000 427078 70200 427146
rect 70000 427022 70074 427078
rect 70130 427022 70200 427078
rect 70000 426954 70200 427022
rect 70000 426898 70074 426954
rect 70130 426898 70200 426954
rect 70000 426829 70200 426898
rect 70000 426108 70200 426173
rect 70000 426052 70074 426108
rect 70130 426052 70200 426108
rect 70000 425984 70200 426052
rect 70000 425928 70074 425984
rect 70130 425928 70200 425984
rect 70000 425860 70200 425928
rect 70000 425804 70074 425860
rect 70130 425804 70200 425860
rect 70000 425736 70200 425804
rect 70000 425680 70074 425736
rect 70130 425680 70200 425736
rect 70000 425612 70200 425680
rect 70000 425556 70074 425612
rect 70130 425556 70200 425612
rect 70000 425488 70200 425556
rect 70000 425432 70074 425488
rect 70130 425432 70200 425488
rect 70000 425364 70200 425432
rect 70000 425308 70074 425364
rect 70130 425308 70200 425364
rect 70000 425240 70200 425308
rect 70000 425184 70074 425240
rect 70130 425184 70200 425240
rect 70000 425116 70200 425184
rect 70000 425060 70074 425116
rect 70130 425060 70200 425116
rect 70000 424992 70200 425060
rect 70000 424936 70074 424992
rect 70130 424936 70200 424992
rect 70000 424868 70200 424936
rect 70000 424812 70074 424868
rect 70130 424812 70200 424868
rect 70000 424744 70200 424812
rect 70000 424688 70074 424744
rect 70130 424688 70200 424744
rect 70000 424620 70200 424688
rect 70000 424564 70074 424620
rect 70130 424564 70200 424620
rect 70000 424496 70200 424564
rect 70000 424440 70074 424496
rect 70130 424440 70200 424496
rect 70000 424372 70200 424440
rect 70000 424316 70074 424372
rect 70130 424316 70200 424372
rect 70000 424248 70200 424316
rect 70000 424192 70074 424248
rect 70130 424192 70200 424248
rect 70000 424123 70200 424192
rect 70000 423738 70200 423803
rect 70000 423682 70074 423738
rect 70130 423682 70200 423738
rect 70000 423614 70200 423682
rect 70000 423558 70074 423614
rect 70130 423558 70200 423614
rect 70000 423490 70200 423558
rect 70000 423434 70074 423490
rect 70130 423434 70200 423490
rect 70000 423366 70200 423434
rect 70000 423310 70074 423366
rect 70130 423310 70200 423366
rect 70000 423242 70200 423310
rect 70000 423186 70074 423242
rect 70130 423186 70200 423242
rect 70000 423118 70200 423186
rect 70000 423062 70074 423118
rect 70130 423062 70200 423118
rect 70000 422994 70200 423062
rect 70000 422938 70074 422994
rect 70130 422938 70200 422994
rect 70000 422870 70200 422938
rect 70000 422814 70074 422870
rect 70130 422814 70200 422870
rect 70000 422746 70200 422814
rect 70000 422690 70074 422746
rect 70130 422690 70200 422746
rect 70000 422622 70200 422690
rect 70000 422566 70074 422622
rect 70130 422566 70200 422622
rect 70000 422498 70200 422566
rect 70000 422442 70074 422498
rect 70130 422442 70200 422498
rect 70000 422374 70200 422442
rect 70000 422318 70074 422374
rect 70130 422318 70200 422374
rect 70000 422250 70200 422318
rect 70000 422194 70074 422250
rect 70130 422194 70200 422250
rect 70000 422126 70200 422194
rect 70000 422070 70074 422126
rect 70130 422070 70200 422126
rect 70000 422002 70200 422070
rect 70000 421946 70074 422002
rect 70130 421946 70200 422002
rect 70000 421878 70200 421946
rect 70000 421822 70074 421878
rect 70130 421822 70200 421878
rect 70000 421753 70200 421822
rect 70000 421134 70200 421173
rect 70000 421078 70074 421134
rect 70130 421078 70200 421134
rect 70000 421010 70200 421078
rect 70000 420954 70074 421010
rect 70130 420954 70200 421010
rect 70000 420886 70200 420954
rect 70000 420830 70074 420886
rect 70130 420830 70200 420886
rect 70000 420762 70200 420830
rect 70000 420706 70074 420762
rect 70130 420706 70200 420762
rect 70000 420638 70200 420706
rect 70000 420582 70074 420638
rect 70130 420582 70200 420638
rect 70000 420514 70200 420582
rect 70000 420458 70074 420514
rect 70130 420458 70200 420514
rect 70000 420390 70200 420458
rect 70000 420334 70074 420390
rect 70130 420334 70200 420390
rect 70000 420266 70200 420334
rect 70000 420210 70074 420266
rect 70130 420210 70200 420266
rect 70000 420142 70200 420210
rect 70000 420086 70074 420142
rect 70130 420086 70200 420142
rect 70000 420018 70200 420086
rect 70000 419962 70074 420018
rect 70130 419962 70200 420018
rect 70000 419894 70200 419962
rect 70000 419838 70074 419894
rect 70130 419838 70200 419894
rect 70000 419770 70200 419838
rect 70000 419714 70074 419770
rect 70130 419714 70200 419770
rect 70000 419646 70200 419714
rect 70000 419590 70074 419646
rect 70130 419590 70200 419646
rect 70000 419522 70200 419590
rect 70000 419466 70074 419522
rect 70130 419466 70200 419522
rect 70000 419398 70200 419466
rect 70000 419342 70074 419398
rect 70130 419342 70200 419398
rect 70000 419273 70200 419342
rect 707800 410658 708000 410728
rect 707800 410602 707870 410658
rect 707926 410602 708000 410658
rect 707800 410534 708000 410602
rect 707800 410478 707870 410534
rect 707926 410478 708000 410534
rect 707800 410410 708000 410478
rect 707800 410354 707870 410410
rect 707926 410354 708000 410410
rect 707800 410286 708000 410354
rect 707800 410230 707870 410286
rect 707926 410230 708000 410286
rect 707800 410162 708000 410230
rect 707800 410106 707870 410162
rect 707926 410106 708000 410162
rect 707800 410038 708000 410106
rect 707800 409982 707870 410038
rect 707926 409982 708000 410038
rect 707800 409914 708000 409982
rect 707800 409858 707870 409914
rect 707926 409858 708000 409914
rect 707800 409790 708000 409858
rect 707800 409734 707870 409790
rect 707926 409734 708000 409790
rect 707800 409666 708000 409734
rect 707800 409610 707870 409666
rect 707926 409610 708000 409666
rect 707800 409542 708000 409610
rect 707800 409486 707870 409542
rect 707926 409486 708000 409542
rect 707800 409418 708000 409486
rect 707800 409362 707870 409418
rect 707926 409362 708000 409418
rect 707800 409294 708000 409362
rect 707800 409238 707870 409294
rect 707926 409238 708000 409294
rect 707800 409170 708000 409238
rect 707800 409114 707870 409170
rect 707926 409114 708000 409170
rect 707800 409046 708000 409114
rect 707800 408990 707870 409046
rect 707926 408990 708000 409046
rect 707800 408922 708000 408990
rect 707800 408866 707870 408922
rect 707926 408866 708000 408922
rect 707800 408828 708000 408866
rect 707800 408178 708000 408248
rect 707800 408122 707870 408178
rect 707926 408122 708000 408178
rect 707800 408054 708000 408122
rect 707800 407998 707870 408054
rect 707926 407998 708000 408054
rect 707800 407930 708000 407998
rect 707800 407874 707870 407930
rect 707926 407874 708000 407930
rect 707800 407806 708000 407874
rect 707800 407750 707870 407806
rect 707926 407750 708000 407806
rect 707800 407682 708000 407750
rect 707800 407626 707870 407682
rect 707926 407626 708000 407682
rect 707800 407558 708000 407626
rect 707800 407502 707870 407558
rect 707926 407502 708000 407558
rect 707800 407434 708000 407502
rect 707800 407378 707870 407434
rect 707926 407378 708000 407434
rect 707800 407310 708000 407378
rect 707800 407254 707870 407310
rect 707926 407254 708000 407310
rect 707800 407186 708000 407254
rect 707800 407130 707870 407186
rect 707926 407130 708000 407186
rect 707800 407062 708000 407130
rect 707800 407006 707870 407062
rect 707926 407006 708000 407062
rect 707800 406938 708000 407006
rect 707800 406882 707870 406938
rect 707926 406882 708000 406938
rect 707800 406814 708000 406882
rect 707800 406758 707870 406814
rect 707926 406758 708000 406814
rect 707800 406690 708000 406758
rect 707800 406634 707870 406690
rect 707926 406634 708000 406690
rect 707800 406566 708000 406634
rect 707800 406510 707870 406566
rect 707926 406510 708000 406566
rect 707800 406442 708000 406510
rect 707800 406386 707870 406442
rect 707926 406386 708000 406442
rect 707800 406318 708000 406386
rect 707800 406262 707870 406318
rect 707926 406262 708000 406318
rect 707800 406198 708000 406262
rect 707800 405808 708000 405878
rect 707800 405752 707870 405808
rect 707926 405752 708000 405808
rect 707800 405684 708000 405752
rect 707800 405628 707870 405684
rect 707926 405628 708000 405684
rect 707800 405560 708000 405628
rect 707800 405504 707870 405560
rect 707926 405504 708000 405560
rect 707800 405436 708000 405504
rect 707800 405380 707870 405436
rect 707926 405380 708000 405436
rect 707800 405312 708000 405380
rect 707800 405256 707870 405312
rect 707926 405256 708000 405312
rect 707800 405188 708000 405256
rect 707800 405132 707870 405188
rect 707926 405132 708000 405188
rect 707800 405064 708000 405132
rect 707800 405008 707870 405064
rect 707926 405008 708000 405064
rect 707800 404940 708000 405008
rect 707800 404884 707870 404940
rect 707926 404884 708000 404940
rect 707800 404816 708000 404884
rect 707800 404760 707870 404816
rect 707926 404760 708000 404816
rect 707800 404692 708000 404760
rect 707800 404636 707870 404692
rect 707926 404636 708000 404692
rect 707800 404568 708000 404636
rect 707800 404512 707870 404568
rect 707926 404512 708000 404568
rect 707800 404444 708000 404512
rect 707800 404388 707870 404444
rect 707926 404388 708000 404444
rect 707800 404320 708000 404388
rect 707800 404264 707870 404320
rect 707926 404264 708000 404320
rect 707800 404196 708000 404264
rect 707800 404140 707870 404196
rect 707926 404140 708000 404196
rect 707800 404072 708000 404140
rect 707800 404016 707870 404072
rect 707926 404016 708000 404072
rect 707800 403948 708000 404016
rect 707800 403892 707870 403948
rect 707926 403892 708000 403948
rect 707800 403828 708000 403892
rect 707800 403102 708000 403172
rect 707800 403046 707870 403102
rect 707926 403046 708000 403102
rect 707800 402978 708000 403046
rect 707800 402922 707870 402978
rect 707926 402922 708000 402978
rect 707800 402854 708000 402922
rect 707800 402798 707870 402854
rect 707926 402798 708000 402854
rect 707800 402730 708000 402798
rect 707800 402674 707870 402730
rect 707926 402674 708000 402730
rect 707800 402606 708000 402674
rect 707800 402550 707870 402606
rect 707926 402550 708000 402606
rect 707800 402482 708000 402550
rect 707800 402426 707870 402482
rect 707926 402426 708000 402482
rect 707800 402358 708000 402426
rect 707800 402302 707870 402358
rect 707926 402302 708000 402358
rect 707800 402234 708000 402302
rect 707800 402178 707870 402234
rect 707926 402178 708000 402234
rect 707800 402110 708000 402178
rect 707800 402054 707870 402110
rect 707926 402054 708000 402110
rect 707800 401986 708000 402054
rect 707800 401930 707870 401986
rect 707926 401930 708000 401986
rect 707800 401862 708000 401930
rect 707800 401806 707870 401862
rect 707926 401806 708000 401862
rect 707800 401738 708000 401806
rect 707800 401682 707870 401738
rect 707926 401682 708000 401738
rect 707800 401614 708000 401682
rect 707800 401558 707870 401614
rect 707926 401558 708000 401614
rect 707800 401490 708000 401558
rect 707800 401434 707870 401490
rect 707926 401434 708000 401490
rect 707800 401366 708000 401434
rect 707800 401310 707870 401366
rect 707926 401310 708000 401366
rect 707800 401242 708000 401310
rect 707800 401186 707870 401242
rect 707926 401186 708000 401242
rect 707800 401122 708000 401186
rect 707800 400732 708000 400802
rect 707800 400676 707870 400732
rect 707926 400676 708000 400732
rect 707800 400608 708000 400676
rect 707800 400552 707870 400608
rect 707926 400552 708000 400608
rect 707800 400484 708000 400552
rect 707800 400428 707870 400484
rect 707926 400428 708000 400484
rect 707800 400360 708000 400428
rect 707800 400304 707870 400360
rect 707926 400304 708000 400360
rect 707800 400236 708000 400304
rect 707800 400180 707870 400236
rect 707926 400180 708000 400236
rect 707800 400112 708000 400180
rect 707800 400056 707870 400112
rect 707926 400056 708000 400112
rect 707800 399988 708000 400056
rect 707800 399932 707870 399988
rect 707926 399932 708000 399988
rect 707800 399864 708000 399932
rect 707800 399808 707870 399864
rect 707926 399808 708000 399864
rect 707800 399740 708000 399808
rect 707800 399684 707870 399740
rect 707926 399684 708000 399740
rect 707800 399616 708000 399684
rect 707800 399560 707870 399616
rect 707926 399560 708000 399616
rect 707800 399492 708000 399560
rect 707800 399436 707870 399492
rect 707926 399436 708000 399492
rect 707800 399368 708000 399436
rect 707800 399312 707870 399368
rect 707926 399312 708000 399368
rect 707800 399244 708000 399312
rect 707800 399188 707870 399244
rect 707926 399188 708000 399244
rect 707800 399120 708000 399188
rect 707800 399064 707870 399120
rect 707926 399064 708000 399120
rect 707800 398996 708000 399064
rect 707800 398940 707870 398996
rect 707926 398940 708000 398996
rect 707800 398872 708000 398940
rect 707800 398816 707870 398872
rect 707926 398816 708000 398872
rect 707800 398752 708000 398816
rect 707800 398134 708000 398172
rect 707800 398078 707870 398134
rect 707926 398078 708000 398134
rect 707800 398010 708000 398078
rect 707800 397954 707870 398010
rect 707926 397954 708000 398010
rect 707800 397886 708000 397954
rect 707800 397830 707870 397886
rect 707926 397830 708000 397886
rect 707800 397762 708000 397830
rect 707800 397706 707870 397762
rect 707926 397706 708000 397762
rect 707800 397638 708000 397706
rect 707800 397582 707870 397638
rect 707926 397582 708000 397638
rect 707800 397514 708000 397582
rect 707800 397458 707870 397514
rect 707926 397458 708000 397514
rect 707800 397390 708000 397458
rect 707800 397334 707870 397390
rect 707926 397334 708000 397390
rect 707800 397266 708000 397334
rect 707800 397210 707870 397266
rect 707926 397210 708000 397266
rect 707800 397142 708000 397210
rect 707800 397086 707870 397142
rect 707926 397086 708000 397142
rect 707800 397018 708000 397086
rect 707800 396962 707870 397018
rect 707926 396962 708000 397018
rect 707800 396894 708000 396962
rect 707800 396838 707870 396894
rect 707926 396838 708000 396894
rect 707800 396770 708000 396838
rect 707800 396714 707870 396770
rect 707926 396714 708000 396770
rect 707800 396646 708000 396714
rect 707800 396590 707870 396646
rect 707926 396590 708000 396646
rect 707800 396522 708000 396590
rect 707800 396466 707870 396522
rect 707926 396466 708000 396522
rect 707800 396398 708000 396466
rect 707800 396342 707870 396398
rect 707926 396342 708000 396398
rect 707800 396272 708000 396342
rect 70000 146658 70200 146728
rect 70000 146602 70074 146658
rect 70130 146602 70200 146658
rect 70000 146534 70200 146602
rect 70000 146478 70074 146534
rect 70130 146478 70200 146534
rect 70000 146410 70200 146478
rect 70000 146354 70074 146410
rect 70130 146354 70200 146410
rect 70000 146286 70200 146354
rect 70000 146230 70074 146286
rect 70130 146230 70200 146286
rect 70000 146162 70200 146230
rect 70000 146106 70074 146162
rect 70130 146106 70200 146162
rect 70000 146038 70200 146106
rect 70000 145982 70074 146038
rect 70130 145982 70200 146038
rect 70000 145914 70200 145982
rect 70000 145858 70074 145914
rect 70130 145858 70200 145914
rect 70000 145790 70200 145858
rect 70000 145734 70074 145790
rect 70130 145734 70200 145790
rect 70000 145666 70200 145734
rect 70000 145610 70074 145666
rect 70130 145610 70200 145666
rect 70000 145542 70200 145610
rect 70000 145486 70074 145542
rect 70130 145486 70200 145542
rect 70000 145418 70200 145486
rect 70000 145362 70074 145418
rect 70130 145362 70200 145418
rect 70000 145294 70200 145362
rect 70000 145238 70074 145294
rect 70130 145238 70200 145294
rect 70000 145170 70200 145238
rect 70000 145114 70074 145170
rect 70130 145114 70200 145170
rect 70000 145046 70200 145114
rect 70000 144990 70074 145046
rect 70130 144990 70200 145046
rect 70000 144922 70200 144990
rect 70000 144866 70074 144922
rect 70130 144866 70200 144922
rect 70000 144828 70200 144866
rect 70000 144184 70200 144248
rect 70000 144128 70074 144184
rect 70130 144128 70200 144184
rect 70000 144060 70200 144128
rect 70000 144004 70074 144060
rect 70130 144004 70200 144060
rect 70000 143936 70200 144004
rect 70000 143880 70074 143936
rect 70130 143880 70200 143936
rect 70000 143812 70200 143880
rect 70000 143756 70074 143812
rect 70130 143756 70200 143812
rect 70000 143688 70200 143756
rect 70000 143632 70074 143688
rect 70130 143632 70200 143688
rect 70000 143564 70200 143632
rect 70000 143508 70074 143564
rect 70130 143508 70200 143564
rect 70000 143440 70200 143508
rect 70000 143384 70074 143440
rect 70130 143384 70200 143440
rect 70000 143316 70200 143384
rect 70000 143260 70074 143316
rect 70130 143260 70200 143316
rect 70000 143192 70200 143260
rect 70000 143136 70074 143192
rect 70130 143136 70200 143192
rect 70000 143068 70200 143136
rect 70000 143012 70074 143068
rect 70130 143012 70200 143068
rect 70000 142944 70200 143012
rect 70000 142888 70074 142944
rect 70130 142888 70200 142944
rect 70000 142820 70200 142888
rect 70000 142764 70074 142820
rect 70130 142764 70200 142820
rect 70000 142696 70200 142764
rect 70000 142640 70074 142696
rect 70130 142640 70200 142696
rect 70000 142572 70200 142640
rect 70000 142516 70074 142572
rect 70130 142516 70200 142572
rect 70000 142448 70200 142516
rect 70000 142392 70074 142448
rect 70130 142392 70200 142448
rect 70000 142324 70200 142392
rect 70000 142268 70074 142324
rect 70130 142268 70200 142324
rect 70000 142198 70200 142268
rect 70000 141814 70200 141878
rect 70000 141758 70074 141814
rect 70130 141758 70200 141814
rect 70000 141690 70200 141758
rect 70000 141634 70074 141690
rect 70130 141634 70200 141690
rect 70000 141566 70200 141634
rect 70000 141510 70074 141566
rect 70130 141510 70200 141566
rect 70000 141442 70200 141510
rect 70000 141386 70074 141442
rect 70130 141386 70200 141442
rect 70000 141318 70200 141386
rect 70000 141262 70074 141318
rect 70130 141262 70200 141318
rect 70000 141194 70200 141262
rect 70000 141138 70074 141194
rect 70130 141138 70200 141194
rect 70000 141070 70200 141138
rect 70000 141014 70074 141070
rect 70130 141014 70200 141070
rect 70000 140946 70200 141014
rect 70000 140890 70074 140946
rect 70130 140890 70200 140946
rect 70000 140822 70200 140890
rect 70000 140766 70074 140822
rect 70130 140766 70200 140822
rect 70000 140698 70200 140766
rect 70000 140642 70074 140698
rect 70130 140642 70200 140698
rect 70000 140574 70200 140642
rect 70000 140518 70074 140574
rect 70130 140518 70200 140574
rect 70000 140450 70200 140518
rect 70000 140394 70074 140450
rect 70130 140394 70200 140450
rect 70000 140326 70200 140394
rect 70000 140270 70074 140326
rect 70130 140270 70200 140326
rect 70000 140202 70200 140270
rect 70000 140146 70074 140202
rect 70130 140146 70200 140202
rect 70000 140078 70200 140146
rect 70000 140022 70074 140078
rect 70130 140022 70200 140078
rect 70000 139954 70200 140022
rect 70000 139898 70074 139954
rect 70130 139898 70200 139954
rect 70000 139828 70200 139898
rect 70000 139108 70200 139172
rect 70000 139052 70074 139108
rect 70130 139052 70200 139108
rect 70000 138984 70200 139052
rect 70000 138928 70074 138984
rect 70130 138928 70200 138984
rect 70000 138860 70200 138928
rect 70000 138804 70074 138860
rect 70130 138804 70200 138860
rect 70000 138736 70200 138804
rect 70000 138680 70074 138736
rect 70130 138680 70200 138736
rect 70000 138612 70200 138680
rect 70000 138556 70074 138612
rect 70130 138556 70200 138612
rect 70000 138488 70200 138556
rect 70000 138432 70074 138488
rect 70130 138432 70200 138488
rect 70000 138364 70200 138432
rect 70000 138308 70074 138364
rect 70130 138308 70200 138364
rect 70000 138240 70200 138308
rect 70000 138184 70074 138240
rect 70130 138184 70200 138240
rect 70000 138116 70200 138184
rect 70000 138060 70074 138116
rect 70130 138060 70200 138116
rect 70000 137992 70200 138060
rect 70000 137936 70074 137992
rect 70130 137936 70200 137992
rect 70000 137868 70200 137936
rect 70000 137812 70074 137868
rect 70130 137812 70200 137868
rect 70000 137744 70200 137812
rect 70000 137688 70074 137744
rect 70130 137688 70200 137744
rect 70000 137620 70200 137688
rect 70000 137564 70074 137620
rect 70130 137564 70200 137620
rect 70000 137496 70200 137564
rect 70000 137440 70074 137496
rect 70130 137440 70200 137496
rect 70000 137372 70200 137440
rect 70000 137316 70074 137372
rect 70130 137316 70200 137372
rect 70000 137248 70200 137316
rect 70000 137192 70074 137248
rect 70130 137192 70200 137248
rect 70000 137122 70200 137192
rect 70000 136738 70200 136802
rect 70000 136682 70074 136738
rect 70130 136682 70200 136738
rect 70000 136614 70200 136682
rect 70000 136558 70074 136614
rect 70130 136558 70200 136614
rect 70000 136490 70200 136558
rect 70000 136434 70074 136490
rect 70130 136434 70200 136490
rect 70000 136366 70200 136434
rect 70000 136310 70074 136366
rect 70130 136310 70200 136366
rect 70000 136242 70200 136310
rect 70000 136186 70074 136242
rect 70130 136186 70200 136242
rect 70000 136118 70200 136186
rect 70000 136062 70074 136118
rect 70130 136062 70200 136118
rect 70000 135994 70200 136062
rect 70000 135938 70074 135994
rect 70130 135938 70200 135994
rect 70000 135870 70200 135938
rect 70000 135814 70074 135870
rect 70130 135814 70200 135870
rect 70000 135746 70200 135814
rect 70000 135690 70074 135746
rect 70130 135690 70200 135746
rect 70000 135622 70200 135690
rect 70000 135566 70074 135622
rect 70130 135566 70200 135622
rect 70000 135498 70200 135566
rect 70000 135442 70074 135498
rect 70130 135442 70200 135498
rect 70000 135374 70200 135442
rect 70000 135318 70074 135374
rect 70130 135318 70200 135374
rect 70000 135250 70200 135318
rect 70000 135194 70074 135250
rect 70130 135194 70200 135250
rect 70000 135126 70200 135194
rect 70000 135070 70074 135126
rect 70130 135070 70200 135126
rect 70000 135002 70200 135070
rect 70000 134946 70074 135002
rect 70130 134946 70200 135002
rect 70000 134878 70200 134946
rect 70000 134822 70074 134878
rect 70130 134822 70200 134878
rect 70000 134752 70200 134822
rect 70000 134134 70200 134172
rect 70000 134078 70074 134134
rect 70130 134078 70200 134134
rect 70000 134010 70200 134078
rect 70000 133954 70074 134010
rect 70130 133954 70200 134010
rect 70000 133886 70200 133954
rect 70000 133830 70074 133886
rect 70130 133830 70200 133886
rect 70000 133762 70200 133830
rect 70000 133706 70074 133762
rect 70130 133706 70200 133762
rect 70000 133638 70200 133706
rect 70000 133582 70074 133638
rect 70130 133582 70200 133638
rect 70000 133514 70200 133582
rect 70000 133458 70074 133514
rect 70130 133458 70200 133514
rect 70000 133390 70200 133458
rect 70000 133334 70074 133390
rect 70130 133334 70200 133390
rect 70000 133266 70200 133334
rect 70000 133210 70074 133266
rect 70130 133210 70200 133266
rect 70000 133142 70200 133210
rect 70000 133086 70074 133142
rect 70130 133086 70200 133142
rect 70000 133018 70200 133086
rect 70000 132962 70074 133018
rect 70130 132962 70200 133018
rect 70000 132894 70200 132962
rect 70000 132838 70074 132894
rect 70130 132838 70200 132894
rect 70000 132770 70200 132838
rect 70000 132714 70074 132770
rect 70130 132714 70200 132770
rect 70000 132646 70200 132714
rect 70000 132590 70074 132646
rect 70130 132590 70200 132646
rect 70000 132522 70200 132590
rect 70000 132466 70074 132522
rect 70130 132466 70200 132522
rect 70000 132398 70200 132466
rect 70000 132342 70074 132398
rect 70130 132342 70200 132398
rect 70000 132272 70200 132342
rect 70000 105658 70200 105728
rect 70000 105602 70074 105658
rect 70130 105602 70200 105658
rect 70000 105534 70200 105602
rect 70000 105478 70074 105534
rect 70130 105478 70200 105534
rect 70000 105410 70200 105478
rect 70000 105354 70074 105410
rect 70130 105354 70200 105410
rect 70000 105286 70200 105354
rect 70000 105230 70074 105286
rect 70130 105230 70200 105286
rect 70000 105162 70200 105230
rect 70000 105106 70074 105162
rect 70130 105106 70200 105162
rect 70000 105038 70200 105106
rect 70000 104982 70074 105038
rect 70130 104982 70200 105038
rect 70000 104914 70200 104982
rect 70000 104858 70074 104914
rect 70130 104858 70200 104914
rect 70000 104790 70200 104858
rect 70000 104734 70074 104790
rect 70130 104734 70200 104790
rect 70000 104666 70200 104734
rect 70000 104610 70074 104666
rect 70130 104610 70200 104666
rect 70000 104542 70200 104610
rect 70000 104486 70074 104542
rect 70130 104486 70200 104542
rect 70000 104418 70200 104486
rect 70000 104362 70074 104418
rect 70130 104362 70200 104418
rect 70000 104294 70200 104362
rect 70000 104238 70074 104294
rect 70130 104238 70200 104294
rect 70000 104170 70200 104238
rect 70000 104114 70074 104170
rect 70130 104114 70200 104170
rect 70000 104046 70200 104114
rect 70000 103990 70074 104046
rect 70130 103990 70200 104046
rect 70000 103922 70200 103990
rect 70000 103866 70074 103922
rect 70130 103866 70200 103922
rect 70000 103828 70200 103866
rect 70000 103184 70200 103248
rect 70000 103128 70074 103184
rect 70130 103128 70200 103184
rect 70000 103060 70200 103128
rect 70000 103004 70074 103060
rect 70130 103004 70200 103060
rect 70000 102936 70200 103004
rect 70000 102880 70074 102936
rect 70130 102880 70200 102936
rect 70000 102812 70200 102880
rect 70000 102756 70074 102812
rect 70130 102756 70200 102812
rect 70000 102688 70200 102756
rect 70000 102632 70074 102688
rect 70130 102632 70200 102688
rect 70000 102564 70200 102632
rect 70000 102508 70074 102564
rect 70130 102508 70200 102564
rect 70000 102440 70200 102508
rect 70000 102384 70074 102440
rect 70130 102384 70200 102440
rect 70000 102316 70200 102384
rect 70000 102260 70074 102316
rect 70130 102260 70200 102316
rect 70000 102192 70200 102260
rect 70000 102136 70074 102192
rect 70130 102136 70200 102192
rect 70000 102068 70200 102136
rect 70000 102012 70074 102068
rect 70130 102012 70200 102068
rect 70000 101944 70200 102012
rect 70000 101888 70074 101944
rect 70130 101888 70200 101944
rect 70000 101820 70200 101888
rect 70000 101764 70074 101820
rect 70130 101764 70200 101820
rect 70000 101696 70200 101764
rect 70000 101640 70074 101696
rect 70130 101640 70200 101696
rect 70000 101572 70200 101640
rect 70000 101516 70074 101572
rect 70130 101516 70200 101572
rect 70000 101448 70200 101516
rect 70000 101392 70074 101448
rect 70130 101392 70200 101448
rect 70000 101324 70200 101392
rect 70000 101268 70074 101324
rect 70130 101268 70200 101324
rect 70000 101198 70200 101268
rect 70000 100814 70200 100878
rect 70000 100758 70074 100814
rect 70130 100758 70200 100814
rect 70000 100690 70200 100758
rect 70000 100634 70074 100690
rect 70130 100634 70200 100690
rect 70000 100566 70200 100634
rect 70000 100510 70074 100566
rect 70130 100510 70200 100566
rect 70000 100442 70200 100510
rect 70000 100386 70074 100442
rect 70130 100386 70200 100442
rect 70000 100318 70200 100386
rect 70000 100262 70074 100318
rect 70130 100262 70200 100318
rect 70000 100194 70200 100262
rect 70000 100138 70074 100194
rect 70130 100138 70200 100194
rect 70000 100070 70200 100138
rect 70000 100014 70074 100070
rect 70130 100014 70200 100070
rect 70000 99946 70200 100014
rect 70000 99890 70074 99946
rect 70130 99890 70200 99946
rect 70000 99822 70200 99890
rect 70000 99766 70074 99822
rect 70130 99766 70200 99822
rect 70000 99698 70200 99766
rect 70000 99642 70074 99698
rect 70130 99642 70200 99698
rect 70000 99574 70200 99642
rect 70000 99518 70074 99574
rect 70130 99518 70200 99574
rect 70000 99450 70200 99518
rect 70000 99394 70074 99450
rect 70130 99394 70200 99450
rect 70000 99326 70200 99394
rect 70000 99270 70074 99326
rect 70130 99270 70200 99326
rect 70000 99202 70200 99270
rect 70000 99146 70074 99202
rect 70130 99146 70200 99202
rect 70000 99078 70200 99146
rect 70000 99022 70074 99078
rect 70130 99022 70200 99078
rect 70000 98954 70200 99022
rect 70000 98898 70074 98954
rect 70130 98898 70200 98954
rect 70000 98828 70200 98898
rect 70000 98108 70200 98172
rect 70000 98052 70074 98108
rect 70130 98052 70200 98108
rect 70000 97984 70200 98052
rect 70000 97928 70074 97984
rect 70130 97928 70200 97984
rect 70000 97860 70200 97928
rect 70000 97804 70074 97860
rect 70130 97804 70200 97860
rect 70000 97736 70200 97804
rect 70000 97680 70074 97736
rect 70130 97680 70200 97736
rect 70000 97612 70200 97680
rect 70000 97556 70074 97612
rect 70130 97556 70200 97612
rect 70000 97488 70200 97556
rect 70000 97432 70074 97488
rect 70130 97432 70200 97488
rect 70000 97364 70200 97432
rect 70000 97308 70074 97364
rect 70130 97308 70200 97364
rect 70000 97240 70200 97308
rect 70000 97184 70074 97240
rect 70130 97184 70200 97240
rect 70000 97116 70200 97184
rect 70000 97060 70074 97116
rect 70130 97060 70200 97116
rect 70000 96992 70200 97060
rect 70000 96936 70074 96992
rect 70130 96936 70200 96992
rect 70000 96868 70200 96936
rect 70000 96812 70074 96868
rect 70130 96812 70200 96868
rect 70000 96744 70200 96812
rect 70000 96688 70074 96744
rect 70130 96688 70200 96744
rect 70000 96620 70200 96688
rect 70000 96564 70074 96620
rect 70130 96564 70200 96620
rect 70000 96496 70200 96564
rect 70000 96440 70074 96496
rect 70130 96440 70200 96496
rect 70000 96372 70200 96440
rect 70000 96316 70074 96372
rect 70130 96316 70200 96372
rect 70000 96248 70200 96316
rect 70000 96192 70074 96248
rect 70130 96192 70200 96248
rect 70000 96122 70200 96192
rect 70000 95738 70200 95802
rect 70000 95682 70074 95738
rect 70130 95682 70200 95738
rect 70000 95614 70200 95682
rect 70000 95558 70074 95614
rect 70130 95558 70200 95614
rect 70000 95490 70200 95558
rect 70000 95434 70074 95490
rect 70130 95434 70200 95490
rect 70000 95366 70200 95434
rect 70000 95310 70074 95366
rect 70130 95310 70200 95366
rect 70000 95242 70200 95310
rect 70000 95186 70074 95242
rect 70130 95186 70200 95242
rect 70000 95118 70200 95186
rect 70000 95062 70074 95118
rect 70130 95062 70200 95118
rect 70000 94994 70200 95062
rect 70000 94938 70074 94994
rect 70130 94938 70200 94994
rect 70000 94870 70200 94938
rect 70000 94814 70074 94870
rect 70130 94814 70200 94870
rect 70000 94746 70200 94814
rect 70000 94690 70074 94746
rect 70130 94690 70200 94746
rect 70000 94622 70200 94690
rect 70000 94566 70074 94622
rect 70130 94566 70200 94622
rect 70000 94498 70200 94566
rect 70000 94442 70074 94498
rect 70130 94442 70200 94498
rect 70000 94374 70200 94442
rect 70000 94318 70074 94374
rect 70130 94318 70200 94374
rect 70000 94250 70200 94318
rect 70000 94194 70074 94250
rect 70130 94194 70200 94250
rect 70000 94126 70200 94194
rect 70000 94070 70074 94126
rect 70130 94070 70200 94126
rect 70000 94002 70200 94070
rect 70000 93946 70074 94002
rect 70130 93946 70200 94002
rect 70000 93878 70200 93946
rect 70000 93822 70074 93878
rect 70130 93822 70200 93878
rect 70000 93752 70200 93822
rect 70000 93134 70200 93172
rect 70000 93078 70074 93134
rect 70130 93078 70200 93134
rect 70000 93010 70200 93078
rect 70000 92954 70074 93010
rect 70130 92954 70200 93010
rect 70000 92886 70200 92954
rect 70000 92830 70074 92886
rect 70130 92830 70200 92886
rect 70000 92762 70200 92830
rect 70000 92706 70074 92762
rect 70130 92706 70200 92762
rect 70000 92638 70200 92706
rect 70000 92582 70074 92638
rect 70130 92582 70200 92638
rect 70000 92514 70200 92582
rect 70000 92458 70074 92514
rect 70130 92458 70200 92514
rect 70000 92390 70200 92458
rect 70000 92334 70074 92390
rect 70130 92334 70200 92390
rect 70000 92266 70200 92334
rect 70000 92210 70074 92266
rect 70130 92210 70200 92266
rect 70000 92142 70200 92210
rect 70000 92086 70074 92142
rect 70130 92086 70200 92142
rect 70000 92018 70200 92086
rect 70000 91962 70074 92018
rect 70130 91962 70200 92018
rect 70000 91894 70200 91962
rect 70000 91838 70074 91894
rect 70130 91838 70200 91894
rect 70000 91770 70200 91838
rect 70000 91714 70074 91770
rect 70130 91714 70200 91770
rect 70000 91646 70200 91714
rect 70000 91590 70074 91646
rect 70130 91590 70200 91646
rect 70000 91522 70200 91590
rect 70000 91466 70074 91522
rect 70130 91466 70200 91522
rect 70000 91398 70200 91466
rect 70000 91342 70074 91398
rect 70130 91342 70200 91398
rect 70000 91272 70200 91342
rect 107272 70130 109172 70200
rect 107272 70074 107342 70130
rect 107398 70074 107466 70130
rect 107522 70074 107590 70130
rect 107646 70074 107714 70130
rect 107770 70074 107838 70130
rect 107894 70074 107962 70130
rect 108018 70074 108086 70130
rect 108142 70074 108210 70130
rect 108266 70074 108334 70130
rect 108390 70074 108458 70130
rect 108514 70074 108582 70130
rect 108638 70074 108706 70130
rect 108762 70074 108830 70130
rect 108886 70074 108954 70130
rect 109010 70074 109078 70130
rect 109134 70074 109172 70130
rect 107272 70000 109172 70074
rect 109752 70130 111802 70200
rect 109752 70074 109822 70130
rect 109878 70074 109946 70130
rect 110002 70074 110070 70130
rect 110126 70074 110194 70130
rect 110250 70074 110318 70130
rect 110374 70074 110442 70130
rect 110498 70074 110566 70130
rect 110622 70074 110690 70130
rect 110746 70074 110814 70130
rect 110870 70074 110938 70130
rect 110994 70074 111062 70130
rect 111118 70074 111186 70130
rect 111242 70074 111310 70130
rect 111366 70074 111434 70130
rect 111490 70074 111558 70130
rect 111614 70074 111682 70130
rect 111738 70074 111802 70130
rect 109752 70000 111802 70074
rect 112122 70130 114172 70200
rect 112122 70074 112192 70130
rect 112248 70074 112316 70130
rect 112372 70074 112440 70130
rect 112496 70074 112564 70130
rect 112620 70074 112688 70130
rect 112744 70074 112812 70130
rect 112868 70074 112936 70130
rect 112992 70074 113060 70130
rect 113116 70074 113184 70130
rect 113240 70074 113308 70130
rect 113364 70074 113432 70130
rect 113488 70074 113556 70130
rect 113612 70074 113680 70130
rect 113736 70074 113804 70130
rect 113860 70074 113928 70130
rect 113984 70074 114052 70130
rect 114108 70074 114172 70130
rect 112122 70000 114172 70074
rect 114828 70130 116878 70200
rect 114828 70074 114892 70130
rect 114948 70074 115016 70130
rect 115072 70074 115140 70130
rect 115196 70074 115264 70130
rect 115320 70074 115388 70130
rect 115444 70074 115512 70130
rect 115568 70074 115636 70130
rect 115692 70074 115760 70130
rect 115816 70074 115884 70130
rect 115940 70074 116008 70130
rect 116064 70074 116132 70130
rect 116188 70074 116256 70130
rect 116312 70074 116380 70130
rect 116436 70074 116504 70130
rect 116560 70074 116628 70130
rect 116684 70074 116752 70130
rect 116808 70074 116878 70130
rect 114828 70000 116878 70074
rect 117198 70130 119248 70200
rect 117198 70074 117262 70130
rect 117318 70074 117386 70130
rect 117442 70074 117510 70130
rect 117566 70074 117634 70130
rect 117690 70074 117758 70130
rect 117814 70074 117882 70130
rect 117938 70074 118006 70130
rect 118062 70074 118130 70130
rect 118186 70074 118254 70130
rect 118310 70074 118378 70130
rect 118434 70074 118502 70130
rect 118558 70074 118626 70130
rect 118682 70074 118750 70130
rect 118806 70074 118874 70130
rect 118930 70074 118998 70130
rect 119054 70074 119122 70130
rect 119178 70074 119248 70130
rect 117198 70000 119248 70074
rect 119828 70130 121728 70200
rect 119828 70074 119866 70130
rect 119922 70074 119990 70130
rect 120046 70074 120114 70130
rect 120170 70074 120238 70130
rect 120294 70074 120362 70130
rect 120418 70074 120486 70130
rect 120542 70074 120610 70130
rect 120666 70074 120734 70130
rect 120790 70074 120858 70130
rect 120914 70074 120982 70130
rect 121038 70074 121106 70130
rect 121162 70074 121230 70130
rect 121286 70074 121354 70130
rect 121410 70074 121478 70130
rect 121534 70074 121602 70130
rect 121658 70074 121728 70130
rect 119828 70000 121728 70074
rect 272272 70130 274172 70200
rect 272272 70074 272342 70130
rect 272398 70074 272466 70130
rect 272522 70074 272590 70130
rect 272646 70074 272714 70130
rect 272770 70074 272838 70130
rect 272894 70074 272962 70130
rect 273018 70074 273086 70130
rect 273142 70074 273210 70130
rect 273266 70074 273334 70130
rect 273390 70074 273458 70130
rect 273514 70074 273582 70130
rect 273638 70074 273706 70130
rect 273762 70074 273830 70130
rect 273886 70074 273954 70130
rect 274010 70074 274078 70130
rect 274134 70074 274172 70130
rect 272272 70000 274172 70074
rect 274752 70130 276802 70200
rect 274752 70074 274822 70130
rect 274878 70074 274946 70130
rect 275002 70074 275070 70130
rect 275126 70074 275194 70130
rect 275250 70074 275318 70130
rect 275374 70074 275442 70130
rect 275498 70074 275566 70130
rect 275622 70074 275690 70130
rect 275746 70074 275814 70130
rect 275870 70074 275938 70130
rect 275994 70074 276062 70130
rect 276118 70074 276186 70130
rect 276242 70074 276310 70130
rect 276366 70074 276434 70130
rect 276490 70074 276558 70130
rect 276614 70074 276682 70130
rect 276738 70074 276802 70130
rect 274752 70000 276802 70074
rect 277122 70130 279172 70200
rect 277122 70074 277192 70130
rect 277248 70074 277316 70130
rect 277372 70074 277440 70130
rect 277496 70074 277564 70130
rect 277620 70074 277688 70130
rect 277744 70074 277812 70130
rect 277868 70074 277936 70130
rect 277992 70074 278060 70130
rect 278116 70074 278184 70130
rect 278240 70074 278308 70130
rect 278364 70074 278432 70130
rect 278488 70074 278556 70130
rect 278612 70074 278680 70130
rect 278736 70074 278804 70130
rect 278860 70074 278928 70130
rect 278984 70074 279052 70130
rect 279108 70074 279172 70130
rect 277122 70000 279172 70074
rect 279828 70130 281878 70200
rect 279828 70074 279892 70130
rect 279948 70074 280016 70130
rect 280072 70074 280140 70130
rect 280196 70074 280264 70130
rect 280320 70074 280388 70130
rect 280444 70074 280512 70130
rect 280568 70074 280636 70130
rect 280692 70074 280760 70130
rect 280816 70074 280884 70130
rect 280940 70074 281008 70130
rect 281064 70074 281132 70130
rect 281188 70074 281256 70130
rect 281312 70074 281380 70130
rect 281436 70074 281504 70130
rect 281560 70074 281628 70130
rect 281684 70074 281752 70130
rect 281808 70074 281878 70130
rect 279828 70000 281878 70074
rect 282198 70130 284248 70200
rect 282198 70074 282262 70130
rect 282318 70074 282386 70130
rect 282442 70074 282510 70130
rect 282566 70074 282634 70130
rect 282690 70074 282758 70130
rect 282814 70074 282882 70130
rect 282938 70074 283006 70130
rect 283062 70074 283130 70130
rect 283186 70074 283254 70130
rect 283310 70074 283378 70130
rect 283434 70074 283502 70130
rect 283558 70074 283626 70130
rect 283682 70074 283750 70130
rect 283806 70074 283874 70130
rect 283930 70074 283998 70130
rect 284054 70074 284122 70130
rect 284178 70074 284248 70130
rect 282198 70000 284248 70074
rect 284828 70130 286728 70200
rect 284828 70074 284866 70130
rect 284922 70074 284990 70130
rect 285046 70074 285114 70130
rect 285170 70074 285238 70130
rect 285294 70074 285362 70130
rect 285418 70074 285486 70130
rect 285542 70074 285610 70130
rect 285666 70074 285734 70130
rect 285790 70074 285858 70130
rect 285914 70074 285982 70130
rect 286038 70074 286106 70130
rect 286162 70074 286230 70130
rect 286286 70074 286354 70130
rect 286410 70074 286478 70130
rect 286534 70074 286602 70130
rect 286658 70074 286728 70130
rect 284828 70000 286728 70074
rect 602272 70130 604172 70200
rect 602272 70074 602342 70130
rect 602398 70074 602466 70130
rect 602522 70074 602590 70130
rect 602646 70074 602714 70130
rect 602770 70074 602838 70130
rect 602894 70074 602962 70130
rect 603018 70074 603086 70130
rect 603142 70074 603210 70130
rect 603266 70074 603334 70130
rect 603390 70074 603458 70130
rect 603514 70074 603582 70130
rect 603638 70074 603706 70130
rect 603762 70074 603830 70130
rect 603886 70074 603954 70130
rect 604010 70074 604078 70130
rect 604134 70074 604172 70130
rect 602272 70000 604172 70074
rect 604752 70130 606802 70200
rect 604752 70074 604822 70130
rect 604878 70074 604946 70130
rect 605002 70074 605070 70130
rect 605126 70074 605194 70130
rect 605250 70074 605318 70130
rect 605374 70074 605442 70130
rect 605498 70074 605566 70130
rect 605622 70074 605690 70130
rect 605746 70074 605814 70130
rect 605870 70074 605938 70130
rect 605994 70074 606062 70130
rect 606118 70074 606186 70130
rect 606242 70074 606310 70130
rect 606366 70074 606434 70130
rect 606490 70074 606558 70130
rect 606614 70074 606682 70130
rect 606738 70074 606802 70130
rect 604752 70000 606802 70074
rect 607122 70130 609172 70200
rect 607122 70074 607192 70130
rect 607248 70074 607316 70130
rect 607372 70074 607440 70130
rect 607496 70074 607564 70130
rect 607620 70074 607688 70130
rect 607744 70074 607812 70130
rect 607868 70074 607936 70130
rect 607992 70074 608060 70130
rect 608116 70074 608184 70130
rect 608240 70074 608308 70130
rect 608364 70074 608432 70130
rect 608488 70074 608556 70130
rect 608612 70074 608680 70130
rect 608736 70074 608804 70130
rect 608860 70074 608928 70130
rect 608984 70074 609052 70130
rect 609108 70074 609172 70130
rect 607122 70000 609172 70074
rect 609828 70130 611878 70200
rect 609828 70074 609892 70130
rect 609948 70074 610016 70130
rect 610072 70074 610140 70130
rect 610196 70074 610264 70130
rect 610320 70074 610388 70130
rect 610444 70074 610512 70130
rect 610568 70074 610636 70130
rect 610692 70074 610760 70130
rect 610816 70074 610884 70130
rect 610940 70074 611008 70130
rect 611064 70074 611132 70130
rect 611188 70074 611256 70130
rect 611312 70074 611380 70130
rect 611436 70074 611504 70130
rect 611560 70074 611628 70130
rect 611684 70074 611752 70130
rect 611808 70074 611878 70130
rect 609828 70000 611878 70074
rect 612198 70130 614248 70200
rect 612198 70074 612262 70130
rect 612318 70074 612386 70130
rect 612442 70074 612510 70130
rect 612566 70074 612634 70130
rect 612690 70074 612758 70130
rect 612814 70074 612882 70130
rect 612938 70074 613006 70130
rect 613062 70074 613130 70130
rect 613186 70074 613254 70130
rect 613310 70074 613378 70130
rect 613434 70074 613502 70130
rect 613558 70074 613626 70130
rect 613682 70074 613750 70130
rect 613806 70074 613874 70130
rect 613930 70074 613998 70130
rect 614054 70074 614122 70130
rect 614178 70074 614248 70130
rect 612198 70000 614248 70074
rect 614828 70130 616728 70200
rect 614828 70074 614866 70130
rect 614922 70074 614990 70130
rect 615046 70074 615114 70130
rect 615170 70074 615238 70130
rect 615294 70074 615362 70130
rect 615418 70074 615486 70130
rect 615542 70074 615610 70130
rect 615666 70074 615734 70130
rect 615790 70074 615858 70130
rect 615914 70074 615982 70130
rect 616038 70074 616106 70130
rect 616162 70074 616230 70130
rect 616286 70074 616354 70130
rect 616410 70074 616478 70130
rect 616534 70074 616602 70130
rect 616658 70074 616728 70130
rect 614828 70000 616728 70074
rect 657272 70130 659172 70200
rect 657272 70074 657342 70130
rect 657398 70074 657466 70130
rect 657522 70074 657590 70130
rect 657646 70074 657714 70130
rect 657770 70074 657838 70130
rect 657894 70074 657962 70130
rect 658018 70074 658086 70130
rect 658142 70074 658210 70130
rect 658266 70074 658334 70130
rect 658390 70074 658458 70130
rect 658514 70074 658582 70130
rect 658638 70074 658706 70130
rect 658762 70074 658830 70130
rect 658886 70074 658954 70130
rect 659010 70074 659078 70130
rect 659134 70074 659172 70130
rect 657272 70000 659172 70074
rect 659752 70130 661802 70200
rect 659752 70074 659822 70130
rect 659878 70074 659946 70130
rect 660002 70074 660070 70130
rect 660126 70074 660194 70130
rect 660250 70074 660318 70130
rect 660374 70074 660442 70130
rect 660498 70074 660566 70130
rect 660622 70074 660690 70130
rect 660746 70074 660814 70130
rect 660870 70074 660938 70130
rect 660994 70074 661062 70130
rect 661118 70074 661186 70130
rect 661242 70074 661310 70130
rect 661366 70074 661434 70130
rect 661490 70074 661558 70130
rect 661614 70074 661682 70130
rect 661738 70074 661802 70130
rect 659752 70000 661802 70074
rect 662122 70130 664172 70200
rect 662122 70074 662192 70130
rect 662248 70074 662316 70130
rect 662372 70074 662440 70130
rect 662496 70074 662564 70130
rect 662620 70074 662688 70130
rect 662744 70074 662812 70130
rect 662868 70074 662936 70130
rect 662992 70074 663060 70130
rect 663116 70074 663184 70130
rect 663240 70074 663308 70130
rect 663364 70074 663432 70130
rect 663488 70074 663556 70130
rect 663612 70074 663680 70130
rect 663736 70074 663804 70130
rect 663860 70074 663928 70130
rect 663984 70074 664052 70130
rect 664108 70074 664172 70130
rect 662122 70000 664172 70074
rect 664828 70130 666878 70200
rect 664828 70074 664892 70130
rect 664948 70074 665016 70130
rect 665072 70074 665140 70130
rect 665196 70074 665264 70130
rect 665320 70074 665388 70130
rect 665444 70074 665512 70130
rect 665568 70074 665636 70130
rect 665692 70074 665760 70130
rect 665816 70074 665884 70130
rect 665940 70074 666008 70130
rect 666064 70074 666132 70130
rect 666188 70074 666256 70130
rect 666312 70074 666380 70130
rect 666436 70074 666504 70130
rect 666560 70074 666628 70130
rect 666684 70074 666752 70130
rect 666808 70074 666878 70130
rect 664828 70000 666878 70074
rect 667198 70130 669248 70200
rect 667198 70074 667262 70130
rect 667318 70074 667386 70130
rect 667442 70074 667510 70130
rect 667566 70074 667634 70130
rect 667690 70074 667758 70130
rect 667814 70074 667882 70130
rect 667938 70074 668006 70130
rect 668062 70074 668130 70130
rect 668186 70074 668254 70130
rect 668310 70074 668378 70130
rect 668434 70074 668502 70130
rect 668558 70074 668626 70130
rect 668682 70074 668750 70130
rect 668806 70074 668874 70130
rect 668930 70074 668998 70130
rect 669054 70074 669122 70130
rect 669178 70074 669248 70130
rect 667198 70000 669248 70074
rect 669828 70130 671728 70200
rect 669828 70074 669866 70130
rect 669922 70074 669990 70130
rect 670046 70074 670114 70130
rect 670170 70074 670238 70130
rect 670294 70074 670362 70130
rect 670418 70074 670486 70130
rect 670542 70074 670610 70130
rect 670666 70074 670734 70130
rect 670790 70074 670858 70130
rect 670914 70074 670982 70130
rect 671038 70074 671106 70130
rect 671162 70074 671230 70130
rect 671286 70074 671354 70130
rect 671410 70074 671478 70130
rect 671534 70074 671602 70130
rect 671658 70074 671728 70130
rect 669828 70000 671728 70074
<< via3 >>
rect 381342 949870 381398 949926
rect 381466 949870 381522 949926
rect 381590 949870 381646 949926
rect 381714 949870 381770 949926
rect 381838 949870 381894 949926
rect 381962 949870 382018 949926
rect 382086 949870 382142 949926
rect 382210 949870 382266 949926
rect 382334 949870 382390 949926
rect 382458 949870 382514 949926
rect 382582 949870 382638 949926
rect 382706 949870 382762 949926
rect 382830 949870 382886 949926
rect 382954 949870 383010 949926
rect 383078 949870 383134 949926
rect 383822 949870 383878 949926
rect 383946 949870 384002 949926
rect 384070 949870 384126 949926
rect 384194 949870 384250 949926
rect 384318 949870 384374 949926
rect 384442 949870 384498 949926
rect 384566 949870 384622 949926
rect 384690 949870 384746 949926
rect 384814 949870 384870 949926
rect 384938 949870 384994 949926
rect 385062 949870 385118 949926
rect 385186 949870 385242 949926
rect 385310 949870 385366 949926
rect 385434 949870 385490 949926
rect 385558 949870 385614 949926
rect 385682 949870 385738 949926
rect 386192 949870 386248 949926
rect 386316 949870 386372 949926
rect 386440 949870 386496 949926
rect 386564 949870 386620 949926
rect 386688 949870 386744 949926
rect 386812 949870 386868 949926
rect 386936 949870 386992 949926
rect 387060 949870 387116 949926
rect 387184 949870 387240 949926
rect 387308 949870 387364 949926
rect 387432 949870 387488 949926
rect 387556 949870 387612 949926
rect 387680 949870 387736 949926
rect 387804 949870 387860 949926
rect 387928 949870 387984 949926
rect 388052 949870 388108 949926
rect 388892 949870 388948 949926
rect 389016 949870 389072 949926
rect 389140 949870 389196 949926
rect 389264 949870 389320 949926
rect 389388 949870 389444 949926
rect 389512 949870 389568 949926
rect 389636 949870 389692 949926
rect 389760 949870 389816 949926
rect 389884 949870 389940 949926
rect 390008 949870 390064 949926
rect 390132 949870 390188 949926
rect 390256 949870 390312 949926
rect 390380 949870 390436 949926
rect 390504 949870 390560 949926
rect 390628 949870 390684 949926
rect 390752 949870 390808 949926
rect 391262 949870 391318 949926
rect 391386 949870 391442 949926
rect 391510 949870 391566 949926
rect 391634 949870 391690 949926
rect 391758 949870 391814 949926
rect 391882 949870 391938 949926
rect 392006 949870 392062 949926
rect 392130 949870 392186 949926
rect 392254 949870 392310 949926
rect 392378 949870 392434 949926
rect 392502 949870 392558 949926
rect 392626 949870 392682 949926
rect 392750 949870 392806 949926
rect 392874 949870 392930 949926
rect 392998 949870 393054 949926
rect 393122 949870 393178 949926
rect 393866 949870 393922 949926
rect 393990 949870 394046 949926
rect 394114 949870 394170 949926
rect 394238 949870 394294 949926
rect 394362 949870 394418 949926
rect 394486 949870 394542 949926
rect 394610 949870 394666 949926
rect 394734 949870 394790 949926
rect 394858 949870 394914 949926
rect 394982 949870 395038 949926
rect 395106 949870 395162 949926
rect 395230 949870 395286 949926
rect 395354 949870 395410 949926
rect 395478 949870 395534 949926
rect 395602 949870 395658 949926
rect 601342 949870 601398 949926
rect 601466 949870 601522 949926
rect 601590 949870 601646 949926
rect 601714 949870 601770 949926
rect 601838 949870 601894 949926
rect 601962 949870 602018 949926
rect 602086 949870 602142 949926
rect 602210 949870 602266 949926
rect 602334 949870 602390 949926
rect 602458 949870 602514 949926
rect 602582 949870 602638 949926
rect 602706 949870 602762 949926
rect 602830 949870 602886 949926
rect 602954 949870 603010 949926
rect 603078 949870 603134 949926
rect 603822 949870 603878 949926
rect 603946 949870 604002 949926
rect 604070 949870 604126 949926
rect 604194 949870 604250 949926
rect 604318 949870 604374 949926
rect 604442 949870 604498 949926
rect 604566 949870 604622 949926
rect 604690 949870 604746 949926
rect 604814 949870 604870 949926
rect 604938 949870 604994 949926
rect 605062 949870 605118 949926
rect 605186 949870 605242 949926
rect 605310 949870 605366 949926
rect 605434 949870 605490 949926
rect 605558 949870 605614 949926
rect 605682 949870 605738 949926
rect 606192 949870 606248 949926
rect 606316 949870 606372 949926
rect 606440 949870 606496 949926
rect 606564 949870 606620 949926
rect 606688 949870 606744 949926
rect 606812 949870 606868 949926
rect 606936 949870 606992 949926
rect 607060 949870 607116 949926
rect 607184 949870 607240 949926
rect 607308 949870 607364 949926
rect 607432 949870 607488 949926
rect 607556 949870 607612 949926
rect 607680 949870 607736 949926
rect 607804 949870 607860 949926
rect 607928 949870 607984 949926
rect 608052 949870 608108 949926
rect 608892 949870 608948 949926
rect 609016 949870 609072 949926
rect 609140 949870 609196 949926
rect 609264 949870 609320 949926
rect 609388 949870 609444 949926
rect 609512 949870 609568 949926
rect 609636 949870 609692 949926
rect 609760 949870 609816 949926
rect 609884 949870 609940 949926
rect 610008 949870 610064 949926
rect 610132 949870 610188 949926
rect 610256 949870 610312 949926
rect 610380 949870 610436 949926
rect 610504 949870 610560 949926
rect 610628 949870 610684 949926
rect 610752 949870 610808 949926
rect 611262 949870 611318 949926
rect 611386 949870 611442 949926
rect 611510 949870 611566 949926
rect 611634 949870 611690 949926
rect 611758 949870 611814 949926
rect 611882 949870 611938 949926
rect 612006 949870 612062 949926
rect 612130 949870 612186 949926
rect 612254 949870 612310 949926
rect 612378 949870 612434 949926
rect 612502 949870 612558 949926
rect 612626 949870 612682 949926
rect 612750 949870 612806 949926
rect 612874 949870 612930 949926
rect 612998 949870 613054 949926
rect 613122 949870 613178 949926
rect 613866 949870 613922 949926
rect 613990 949870 614046 949926
rect 614114 949870 614170 949926
rect 614238 949870 614294 949926
rect 614362 949870 614418 949926
rect 614486 949870 614542 949926
rect 614610 949870 614666 949926
rect 614734 949870 614790 949926
rect 614858 949870 614914 949926
rect 614982 949870 615038 949926
rect 615106 949870 615162 949926
rect 615230 949870 615286 949926
rect 615354 949870 615410 949926
rect 615478 949870 615534 949926
rect 615602 949870 615658 949926
rect 70074 884602 70130 884658
rect 70074 884478 70130 884534
rect 70074 884354 70130 884410
rect 70074 884230 70130 884286
rect 70074 884106 70130 884162
rect 70074 883982 70130 884038
rect 70074 883858 70130 883914
rect 70074 883734 70130 883790
rect 70074 883610 70130 883666
rect 70074 883486 70130 883542
rect 70074 883362 70130 883418
rect 70074 883238 70130 883294
rect 70074 883114 70130 883170
rect 70074 882990 70130 883046
rect 70074 882866 70130 882922
rect 707870 883602 707926 883658
rect 707870 883478 707926 883534
rect 707870 883354 707926 883410
rect 707870 883230 707926 883286
rect 707870 883106 707926 883162
rect 707870 882982 707926 883038
rect 707870 882858 707926 882914
rect 707870 882734 707926 882790
rect 707870 882610 707926 882666
rect 707870 882486 707926 882542
rect 707870 882362 707926 882418
rect 70074 882128 70130 882184
rect 70074 882004 70130 882060
rect 70074 881880 70130 881936
rect 707870 882238 707926 882294
rect 707870 882114 707926 882170
rect 707870 881990 707926 882046
rect 707870 881866 707926 881922
rect 70074 881756 70130 881812
rect 70074 881632 70130 881688
rect 70074 881508 70130 881564
rect 70074 881384 70130 881440
rect 70074 881260 70130 881316
rect 70074 881136 70130 881192
rect 70074 881012 70130 881068
rect 70074 880888 70130 880944
rect 70074 880764 70130 880820
rect 70074 880640 70130 880696
rect 70074 880516 70130 880572
rect 70074 880392 70130 880448
rect 70074 880268 70130 880324
rect 707870 881122 707926 881178
rect 707870 880998 707926 881054
rect 707870 880874 707926 880930
rect 707870 880750 707926 880806
rect 707870 880626 707926 880682
rect 707870 880502 707926 880558
rect 707870 880378 707926 880434
rect 707870 880254 707926 880310
rect 707870 880130 707926 880186
rect 707870 880006 707926 880062
rect 707870 879882 707926 879938
rect 70074 879758 70130 879814
rect 70074 879634 70130 879690
rect 70074 879510 70130 879566
rect 70074 879386 70130 879442
rect 70074 879262 70130 879318
rect 707870 879758 707926 879814
rect 707870 879634 707926 879690
rect 707870 879510 707926 879566
rect 707870 879386 707926 879442
rect 707870 879262 707926 879318
rect 70074 879138 70130 879194
rect 70074 879014 70130 879070
rect 70074 878890 70130 878946
rect 70074 878766 70130 878822
rect 70074 878642 70130 878698
rect 70074 878518 70130 878574
rect 70074 878394 70130 878450
rect 70074 878270 70130 878326
rect 70074 878146 70130 878202
rect 70074 878022 70130 878078
rect 70074 877898 70130 877954
rect 707870 878752 707926 878808
rect 707870 878628 707926 878684
rect 707870 878504 707926 878560
rect 707870 878380 707926 878436
rect 707870 878256 707926 878312
rect 707870 878132 707926 878188
rect 707870 878008 707926 878064
rect 707870 877884 707926 877940
rect 707870 877760 707926 877816
rect 707870 877636 707926 877692
rect 707870 877512 707926 877568
rect 707870 877388 707926 877444
rect 707870 877264 707926 877320
rect 70074 877052 70130 877108
rect 70074 876928 70130 876984
rect 70074 876804 70130 876860
rect 707870 877140 707926 877196
rect 707870 877016 707926 877072
rect 707870 876892 707926 876948
rect 70074 876680 70130 876736
rect 70074 876556 70130 876612
rect 70074 876432 70130 876488
rect 70074 876308 70130 876364
rect 70074 876184 70130 876240
rect 70074 876060 70130 876116
rect 70074 875936 70130 875992
rect 70074 875812 70130 875868
rect 70074 875688 70130 875744
rect 70074 875564 70130 875620
rect 70074 875440 70130 875496
rect 70074 875316 70130 875372
rect 70074 875192 70130 875248
rect 707870 876046 707926 876102
rect 707870 875922 707926 875978
rect 707870 875798 707926 875854
rect 707870 875674 707926 875730
rect 707870 875550 707926 875606
rect 707870 875426 707926 875482
rect 707870 875302 707926 875358
rect 707870 875178 707926 875234
rect 707870 875054 707926 875110
rect 707870 874930 707926 874986
rect 707870 874806 707926 874862
rect 70074 874682 70130 874738
rect 70074 874558 70130 874614
rect 70074 874434 70130 874490
rect 70074 874310 70130 874366
rect 70074 874186 70130 874242
rect 707870 874682 707926 874738
rect 707870 874558 707926 874614
rect 707870 874434 707926 874490
rect 707870 874310 707926 874366
rect 707870 874186 707926 874242
rect 70074 874062 70130 874118
rect 70074 873938 70130 873994
rect 70074 873814 70130 873870
rect 70074 873690 70130 873746
rect 70074 873566 70130 873622
rect 70074 873442 70130 873498
rect 70074 873318 70130 873374
rect 70074 873194 70130 873250
rect 70074 873070 70130 873126
rect 70074 872946 70130 873002
rect 70074 872822 70130 872878
rect 707870 873676 707926 873732
rect 707870 873552 707926 873608
rect 707870 873428 707926 873484
rect 707870 873304 707926 873360
rect 707870 873180 707926 873236
rect 707870 873056 707926 873112
rect 707870 872932 707926 872988
rect 707870 872808 707926 872864
rect 707870 872684 707926 872740
rect 707870 872560 707926 872616
rect 707870 872436 707926 872492
rect 707870 872312 707926 872368
rect 707870 872188 707926 872244
rect 70074 872078 70130 872134
rect 70074 871954 70130 872010
rect 70074 871830 70130 871886
rect 70074 871706 70130 871762
rect 707870 872064 707926 872120
rect 707870 871940 707926 871996
rect 707870 871816 707926 871872
rect 70074 871582 70130 871638
rect 70074 871458 70130 871514
rect 70074 871334 70130 871390
rect 70074 871210 70130 871266
rect 70074 871086 70130 871142
rect 70074 870962 70130 871018
rect 70074 870838 70130 870894
rect 70074 870714 70130 870770
rect 70074 870590 70130 870646
rect 70074 870466 70130 870522
rect 70074 870342 70130 870398
rect 707870 871078 707926 871134
rect 707870 870954 707926 871010
rect 707870 870830 707926 870886
rect 707870 870706 707926 870762
rect 707870 870582 707926 870638
rect 707870 870458 707926 870514
rect 707870 870334 707926 870390
rect 707870 870210 707926 870266
rect 707870 870086 707926 870142
rect 707870 869962 707926 870018
rect 707870 869838 707926 869894
rect 707870 869714 707926 869770
rect 707870 869590 707926 869646
rect 707870 869466 707926 869522
rect 707870 869342 707926 869398
rect 70074 843602 70130 843658
rect 70074 843478 70130 843534
rect 70074 843354 70130 843410
rect 70074 843230 70130 843286
rect 70074 843106 70130 843162
rect 70074 842982 70130 843038
rect 70074 842858 70130 842914
rect 70074 842734 70130 842790
rect 70074 842610 70130 842666
rect 70074 842486 70130 842542
rect 70074 842362 70130 842418
rect 70074 842238 70130 842294
rect 70074 842114 70130 842170
rect 70074 841990 70130 842046
rect 70074 841866 70130 841922
rect 70074 841128 70130 841184
rect 70074 841004 70130 841060
rect 70074 840880 70130 840936
rect 70074 840756 70130 840812
rect 70074 840632 70130 840688
rect 70074 840508 70130 840564
rect 70074 840384 70130 840440
rect 70074 840260 70130 840316
rect 70074 840136 70130 840192
rect 70074 840012 70130 840068
rect 70074 839888 70130 839944
rect 70074 839764 70130 839820
rect 70074 839640 70130 839696
rect 70074 839516 70130 839572
rect 70074 839392 70130 839448
rect 70074 839268 70130 839324
rect 70074 838758 70130 838814
rect 70074 838634 70130 838690
rect 70074 838510 70130 838566
rect 70074 838386 70130 838442
rect 70074 838262 70130 838318
rect 70074 838138 70130 838194
rect 70074 838014 70130 838070
rect 70074 837890 70130 837946
rect 70074 837766 70130 837822
rect 70074 837642 70130 837698
rect 70074 837518 70130 837574
rect 70074 837394 70130 837450
rect 70074 837270 70130 837326
rect 70074 837146 70130 837202
rect 70074 837022 70130 837078
rect 70074 836898 70130 836954
rect 70074 836052 70130 836108
rect 70074 835928 70130 835984
rect 70074 835804 70130 835860
rect 70074 835680 70130 835736
rect 70074 835556 70130 835612
rect 70074 835432 70130 835488
rect 70074 835308 70130 835364
rect 70074 835184 70130 835240
rect 70074 835060 70130 835116
rect 70074 834936 70130 834992
rect 70074 834812 70130 834868
rect 70074 834688 70130 834744
rect 70074 834564 70130 834620
rect 70074 834440 70130 834496
rect 70074 834316 70130 834372
rect 70074 834192 70130 834248
rect 70074 833682 70130 833738
rect 70074 833558 70130 833614
rect 70074 833434 70130 833490
rect 70074 833310 70130 833366
rect 70074 833186 70130 833242
rect 70074 833062 70130 833118
rect 70074 832938 70130 832994
rect 70074 832814 70130 832870
rect 70074 832690 70130 832746
rect 70074 832566 70130 832622
rect 70074 832442 70130 832498
rect 70074 832318 70130 832374
rect 70074 832194 70130 832250
rect 70074 832070 70130 832126
rect 70074 831946 70130 832002
rect 70074 831822 70130 831878
rect 70074 831078 70130 831134
rect 70074 830954 70130 831010
rect 70074 830830 70130 830886
rect 70074 830706 70130 830762
rect 70074 830582 70130 830638
rect 70074 830458 70130 830514
rect 70074 830334 70130 830390
rect 70074 830210 70130 830266
rect 70074 830086 70130 830142
rect 70074 829962 70130 830018
rect 70074 829838 70130 829894
rect 70074 829714 70130 829770
rect 70074 829590 70130 829646
rect 70074 829466 70130 829522
rect 70074 829342 70130 829398
rect 70074 802602 70130 802658
rect 70074 802478 70130 802534
rect 70074 802354 70130 802410
rect 70074 802230 70130 802286
rect 70074 802106 70130 802162
rect 70074 801982 70130 802038
rect 70074 801858 70130 801914
rect 70074 801734 70130 801790
rect 70074 801610 70130 801666
rect 70074 801486 70130 801542
rect 70074 801362 70130 801418
rect 70074 801238 70130 801294
rect 70074 801114 70130 801170
rect 70074 800990 70130 801046
rect 70074 800866 70130 800922
rect 70074 800128 70130 800184
rect 70074 800004 70130 800060
rect 70074 799880 70130 799936
rect 70074 799756 70130 799812
rect 70074 799632 70130 799688
rect 70074 799508 70130 799564
rect 70074 799384 70130 799440
rect 70074 799260 70130 799316
rect 70074 799136 70130 799192
rect 70074 799012 70130 799068
rect 70074 798888 70130 798944
rect 70074 798764 70130 798820
rect 70074 798640 70130 798696
rect 70074 798516 70130 798572
rect 70074 798392 70130 798448
rect 70074 798268 70130 798324
rect 70074 797758 70130 797814
rect 70074 797634 70130 797690
rect 70074 797510 70130 797566
rect 70074 797386 70130 797442
rect 70074 797262 70130 797318
rect 70074 797138 70130 797194
rect 70074 797014 70130 797070
rect 70074 796890 70130 796946
rect 70074 796766 70130 796822
rect 70074 796642 70130 796698
rect 70074 796518 70130 796574
rect 70074 796394 70130 796450
rect 70074 796270 70130 796326
rect 70074 796146 70130 796202
rect 70074 796022 70130 796078
rect 70074 795898 70130 795954
rect 707870 797602 707926 797658
rect 707870 797478 707926 797534
rect 707870 797354 707926 797410
rect 707870 797230 707926 797286
rect 707870 797106 707926 797162
rect 707870 796982 707926 797038
rect 707870 796858 707926 796914
rect 707870 796734 707926 796790
rect 707870 796610 707926 796666
rect 707870 796486 707926 796542
rect 707870 796362 707926 796418
rect 707870 796238 707926 796294
rect 707870 796114 707926 796170
rect 707870 795990 707926 796046
rect 707870 795866 707926 795922
rect 70074 795052 70130 795108
rect 70074 794928 70130 794984
rect 70074 794804 70130 794860
rect 70074 794680 70130 794736
rect 70074 794556 70130 794612
rect 70074 794432 70130 794488
rect 70074 794308 70130 794364
rect 70074 794184 70130 794240
rect 70074 794060 70130 794116
rect 70074 793936 70130 793992
rect 70074 793812 70130 793868
rect 70074 793688 70130 793744
rect 70074 793564 70130 793620
rect 70074 793440 70130 793496
rect 70074 793316 70130 793372
rect 70074 793192 70130 793248
rect 707870 795122 707926 795178
rect 707870 794998 707926 795054
rect 707870 794874 707926 794930
rect 707870 794750 707926 794806
rect 707870 794626 707926 794682
rect 707870 794502 707926 794558
rect 707870 794378 707926 794434
rect 707870 794254 707926 794310
rect 707870 794130 707926 794186
rect 707870 794006 707926 794062
rect 707870 793882 707926 793938
rect 707870 793758 707926 793814
rect 707870 793634 707926 793690
rect 707870 793510 707926 793566
rect 707870 793386 707926 793442
rect 707870 793262 707926 793318
rect 70074 792682 70130 792738
rect 70074 792558 70130 792614
rect 70074 792434 70130 792490
rect 70074 792310 70130 792366
rect 70074 792186 70130 792242
rect 70074 792062 70130 792118
rect 70074 791938 70130 791994
rect 70074 791814 70130 791870
rect 70074 791690 70130 791746
rect 70074 791566 70130 791622
rect 70074 791442 70130 791498
rect 70074 791318 70130 791374
rect 70074 791194 70130 791250
rect 70074 791070 70130 791126
rect 70074 790946 70130 791002
rect 70074 790822 70130 790878
rect 707870 792752 707926 792808
rect 707870 792628 707926 792684
rect 707870 792504 707926 792560
rect 707870 792380 707926 792436
rect 707870 792256 707926 792312
rect 707870 792132 707926 792188
rect 707870 792008 707926 792064
rect 707870 791884 707926 791940
rect 707870 791760 707926 791816
rect 707870 791636 707926 791692
rect 707870 791512 707926 791568
rect 707870 791388 707926 791444
rect 707870 791264 707926 791320
rect 707870 791140 707926 791196
rect 707870 791016 707926 791072
rect 707870 790892 707926 790948
rect 70074 790078 70130 790134
rect 70074 789954 70130 790010
rect 70074 789830 70130 789886
rect 70074 789706 70130 789762
rect 70074 789582 70130 789638
rect 70074 789458 70130 789514
rect 70074 789334 70130 789390
rect 70074 789210 70130 789266
rect 70074 789086 70130 789142
rect 70074 788962 70130 789018
rect 70074 788838 70130 788894
rect 70074 788714 70130 788770
rect 70074 788590 70130 788646
rect 70074 788466 70130 788522
rect 70074 788342 70130 788398
rect 707870 790046 707926 790102
rect 707870 789922 707926 789978
rect 707870 789798 707926 789854
rect 707870 789674 707926 789730
rect 707870 789550 707926 789606
rect 707870 789426 707926 789482
rect 707870 789302 707926 789358
rect 707870 789178 707926 789234
rect 707870 789054 707926 789110
rect 707870 788930 707926 788986
rect 707870 788806 707926 788862
rect 707870 788682 707926 788738
rect 707870 788558 707926 788614
rect 707870 788434 707926 788490
rect 707870 788310 707926 788366
rect 707870 788186 707926 788242
rect 707870 787676 707926 787732
rect 707870 787552 707926 787608
rect 707870 787428 707926 787484
rect 707870 787304 707926 787360
rect 707870 787180 707926 787236
rect 707870 787056 707926 787112
rect 707870 786932 707926 786988
rect 707870 786808 707926 786864
rect 707870 786684 707926 786740
rect 707870 786560 707926 786616
rect 707870 786436 707926 786492
rect 707870 786312 707926 786368
rect 707870 786188 707926 786244
rect 707870 786064 707926 786120
rect 707870 785940 707926 785996
rect 707870 785816 707926 785872
rect 707870 785078 707926 785134
rect 707870 784954 707926 785010
rect 707870 784830 707926 784886
rect 707870 784706 707926 784762
rect 707870 784582 707926 784638
rect 707870 784458 707926 784514
rect 707870 784334 707926 784390
rect 707870 784210 707926 784266
rect 707870 784086 707926 784142
rect 707870 783962 707926 784018
rect 707870 783838 707926 783894
rect 707870 783714 707926 783770
rect 707870 783590 707926 783646
rect 707870 783466 707926 783522
rect 707870 783342 707926 783398
rect 707870 496602 707926 496658
rect 707870 496478 707926 496534
rect 707870 496354 707926 496410
rect 707870 496230 707926 496286
rect 707870 496106 707926 496162
rect 707870 495982 707926 496038
rect 707870 495858 707926 495914
rect 707870 495734 707926 495790
rect 707870 495610 707926 495666
rect 707870 495486 707926 495542
rect 707870 495362 707926 495418
rect 707870 495238 707926 495294
rect 707870 495114 707926 495170
rect 707870 494990 707926 495046
rect 707870 494866 707926 494922
rect 707870 494122 707926 494178
rect 707870 493998 707926 494054
rect 707870 493874 707926 493930
rect 707870 493750 707926 493806
rect 707870 493626 707926 493682
rect 707870 493502 707926 493558
rect 707870 493378 707926 493434
rect 707870 493254 707926 493310
rect 707870 493130 707926 493186
rect 707870 493006 707926 493062
rect 707870 492882 707926 492938
rect 707870 492758 707926 492814
rect 707870 492634 707926 492690
rect 707870 492510 707926 492566
rect 707870 492386 707926 492442
rect 707870 492262 707926 492318
rect 707870 491752 707926 491808
rect 707870 491628 707926 491684
rect 707870 491504 707926 491560
rect 707870 491380 707926 491436
rect 707870 491256 707926 491312
rect 707870 491132 707926 491188
rect 707870 491008 707926 491064
rect 707870 490884 707926 490940
rect 707870 490760 707926 490816
rect 707870 490636 707926 490692
rect 707870 490512 707926 490568
rect 707870 490388 707926 490444
rect 707870 490264 707926 490320
rect 707870 490140 707926 490196
rect 707870 490016 707926 490072
rect 707870 489892 707926 489948
rect 707870 489046 707926 489102
rect 707870 488922 707926 488978
rect 707870 488798 707926 488854
rect 707870 488674 707926 488730
rect 707870 488550 707926 488606
rect 707870 488426 707926 488482
rect 707870 488302 707926 488358
rect 707870 488178 707926 488234
rect 707870 488054 707926 488110
rect 707870 487930 707926 487986
rect 707870 487806 707926 487862
rect 707870 487682 707926 487738
rect 707870 487558 707926 487614
rect 707870 487434 707926 487490
rect 707870 487310 707926 487366
rect 707870 487186 707926 487242
rect 707870 486676 707926 486732
rect 707870 486552 707926 486608
rect 707870 486428 707926 486484
rect 707870 486304 707926 486360
rect 707870 486180 707926 486236
rect 707870 486056 707926 486112
rect 707870 485932 707926 485988
rect 707870 485808 707926 485864
rect 707870 485684 707926 485740
rect 707870 485560 707926 485616
rect 707870 485436 707926 485492
rect 707870 485312 707926 485368
rect 707870 485188 707926 485244
rect 707870 485064 707926 485120
rect 707870 484940 707926 484996
rect 707870 484816 707926 484872
rect 707870 484078 707926 484134
rect 707870 483954 707926 484010
rect 707870 483830 707926 483886
rect 707870 483706 707926 483762
rect 707870 483582 707926 483638
rect 707870 483458 707926 483514
rect 707870 483334 707926 483390
rect 707870 483210 707926 483266
rect 707870 483086 707926 483142
rect 707870 482962 707926 483018
rect 707870 482838 707926 482894
rect 707870 482714 707926 482770
rect 707870 482590 707926 482646
rect 707870 482466 707926 482522
rect 707870 482342 707926 482398
rect 70074 474602 70130 474658
rect 70074 474478 70130 474534
rect 70074 474354 70130 474410
rect 70074 474230 70130 474286
rect 70074 474106 70130 474162
rect 70074 473982 70130 474038
rect 70074 473858 70130 473914
rect 70074 473734 70130 473790
rect 70074 473610 70130 473666
rect 70074 473486 70130 473542
rect 70074 473362 70130 473418
rect 70074 473238 70130 473294
rect 70074 473114 70130 473170
rect 70074 472990 70130 473046
rect 70074 472866 70130 472922
rect 70074 472128 70130 472184
rect 70074 472004 70130 472060
rect 70074 471880 70130 471936
rect 70074 471756 70130 471812
rect 70074 471632 70130 471688
rect 70074 471508 70130 471564
rect 70074 471384 70130 471440
rect 70074 471260 70130 471316
rect 70074 471136 70130 471192
rect 70074 471012 70130 471068
rect 70074 470888 70130 470944
rect 70074 470764 70130 470820
rect 70074 470640 70130 470696
rect 70074 470516 70130 470572
rect 70074 470392 70130 470448
rect 70074 470268 70130 470324
rect 70074 469758 70130 469814
rect 70074 469634 70130 469690
rect 70074 469510 70130 469566
rect 70074 469386 70130 469442
rect 70074 469262 70130 469318
rect 70074 469138 70130 469194
rect 70074 469014 70130 469070
rect 70074 468890 70130 468946
rect 70074 468766 70130 468822
rect 70074 468642 70130 468698
rect 70074 468518 70130 468574
rect 70074 468394 70130 468450
rect 70074 468270 70130 468326
rect 70074 468146 70130 468202
rect 70074 468022 70130 468078
rect 70074 467898 70130 467954
rect 70074 467052 70130 467108
rect 70074 466928 70130 466984
rect 70074 466804 70130 466860
rect 70074 466680 70130 466736
rect 70074 466556 70130 466612
rect 70074 466432 70130 466488
rect 70074 466308 70130 466364
rect 70074 466184 70130 466240
rect 70074 466060 70130 466116
rect 70074 465936 70130 465992
rect 70074 465812 70130 465868
rect 70074 465688 70130 465744
rect 70074 465564 70130 465620
rect 70074 465440 70130 465496
rect 70074 465316 70130 465372
rect 70074 465192 70130 465248
rect 70074 464682 70130 464738
rect 70074 464558 70130 464614
rect 70074 464434 70130 464490
rect 70074 464310 70130 464366
rect 70074 464186 70130 464242
rect 70074 464062 70130 464118
rect 70074 463938 70130 463994
rect 70074 463814 70130 463870
rect 70074 463690 70130 463746
rect 70074 463566 70130 463622
rect 70074 463442 70130 463498
rect 70074 463318 70130 463374
rect 70074 463194 70130 463250
rect 70074 463070 70130 463126
rect 70074 462946 70130 463002
rect 70074 462822 70130 462878
rect 70074 462078 70130 462134
rect 70074 461954 70130 462010
rect 70074 461830 70130 461886
rect 70074 461706 70130 461762
rect 70074 461582 70130 461638
rect 70074 461458 70130 461514
rect 70074 461334 70130 461390
rect 70074 461210 70130 461266
rect 70074 461086 70130 461142
rect 70074 460962 70130 461018
rect 70074 460838 70130 460894
rect 70074 460714 70130 460770
rect 70074 460590 70130 460646
rect 70074 460466 70130 460522
rect 70074 460342 70130 460398
rect 707870 453602 707926 453658
rect 707870 453478 707926 453534
rect 707870 453354 707926 453410
rect 707870 453230 707926 453286
rect 707870 453106 707926 453162
rect 707870 452982 707926 453038
rect 707870 452858 707926 452914
rect 707870 452734 707926 452790
rect 707870 452610 707926 452666
rect 707870 452486 707926 452542
rect 707870 452362 707926 452418
rect 707870 452238 707926 452294
rect 707870 452114 707926 452170
rect 707870 451990 707926 452046
rect 707870 451866 707926 451922
rect 707870 451122 707926 451178
rect 707870 450998 707926 451054
rect 707870 450874 707926 450930
rect 707870 450750 707926 450806
rect 707870 450626 707926 450682
rect 707870 450502 707926 450558
rect 707870 450378 707926 450434
rect 707870 450254 707926 450310
rect 707870 450130 707926 450186
rect 707870 450006 707926 450062
rect 707870 449882 707926 449938
rect 707870 449758 707926 449814
rect 707870 449634 707926 449690
rect 707870 449510 707926 449566
rect 707870 449386 707926 449442
rect 707870 449262 707926 449318
rect 707870 448752 707926 448808
rect 707870 448628 707926 448684
rect 707870 448504 707926 448560
rect 707870 448380 707926 448436
rect 707870 448256 707926 448312
rect 707870 448132 707926 448188
rect 707870 448008 707926 448064
rect 707870 447884 707926 447940
rect 707870 447760 707926 447816
rect 707870 447636 707926 447692
rect 707870 447512 707926 447568
rect 707870 447388 707926 447444
rect 707870 447264 707926 447320
rect 707870 447140 707926 447196
rect 707870 447016 707926 447072
rect 707870 446892 707926 446948
rect 707870 446046 707926 446102
rect 707870 445922 707926 445978
rect 707870 445798 707926 445854
rect 707870 445674 707926 445730
rect 707870 445550 707926 445606
rect 707870 445426 707926 445482
rect 707870 445302 707926 445358
rect 707870 445178 707926 445234
rect 707870 445054 707926 445110
rect 707870 444930 707926 444986
rect 707870 444806 707926 444862
rect 707870 444682 707926 444738
rect 707870 444558 707926 444614
rect 707870 444434 707926 444490
rect 707870 444310 707926 444366
rect 707870 444186 707926 444242
rect 707870 443676 707926 443732
rect 707870 443552 707926 443608
rect 707870 443428 707926 443484
rect 707870 443304 707926 443360
rect 707870 443180 707926 443236
rect 707870 443056 707926 443112
rect 707870 442932 707926 442988
rect 707870 442808 707926 442864
rect 707870 442684 707926 442740
rect 707870 442560 707926 442616
rect 707870 442436 707926 442492
rect 707870 442312 707926 442368
rect 707870 442188 707926 442244
rect 707870 442064 707926 442120
rect 707870 441940 707926 441996
rect 707870 441816 707926 441872
rect 707870 441078 707926 441134
rect 707870 440954 707926 441010
rect 707870 440830 707926 440886
rect 707870 440706 707926 440762
rect 707870 440582 707926 440638
rect 707870 440458 707926 440514
rect 707870 440334 707926 440390
rect 707870 440210 707926 440266
rect 707870 440086 707926 440142
rect 707870 439962 707926 440018
rect 707870 439838 707926 439894
rect 707870 439714 707926 439770
rect 707870 439590 707926 439646
rect 707870 439466 707926 439522
rect 707870 439342 707926 439398
rect 70074 433602 70130 433658
rect 70074 433478 70130 433534
rect 70074 433354 70130 433410
rect 70074 433230 70130 433286
rect 70074 433106 70130 433162
rect 70074 432982 70130 433038
rect 70074 432858 70130 432914
rect 70074 432734 70130 432790
rect 70074 432610 70130 432666
rect 70074 432486 70130 432542
rect 70074 432362 70130 432418
rect 70074 432238 70130 432294
rect 70074 432114 70130 432170
rect 70074 431990 70130 432046
rect 70074 431866 70130 431922
rect 70074 431128 70130 431184
rect 70074 431004 70130 431060
rect 70074 430880 70130 430936
rect 70074 430756 70130 430812
rect 70074 430632 70130 430688
rect 70074 430508 70130 430564
rect 70074 430384 70130 430440
rect 70074 430260 70130 430316
rect 70074 430136 70130 430192
rect 70074 430012 70130 430068
rect 70074 429888 70130 429944
rect 70074 429764 70130 429820
rect 70074 429640 70130 429696
rect 70074 429516 70130 429572
rect 70074 429392 70130 429448
rect 70074 429268 70130 429324
rect 70074 428758 70130 428814
rect 70074 428634 70130 428690
rect 70074 428510 70130 428566
rect 70074 428386 70130 428442
rect 70074 428262 70130 428318
rect 70074 428138 70130 428194
rect 70074 428014 70130 428070
rect 70074 427890 70130 427946
rect 70074 427766 70130 427822
rect 70074 427642 70130 427698
rect 70074 427518 70130 427574
rect 70074 427394 70130 427450
rect 70074 427270 70130 427326
rect 70074 427146 70130 427202
rect 70074 427022 70130 427078
rect 70074 426898 70130 426954
rect 70074 426052 70130 426108
rect 70074 425928 70130 425984
rect 70074 425804 70130 425860
rect 70074 425680 70130 425736
rect 70074 425556 70130 425612
rect 70074 425432 70130 425488
rect 70074 425308 70130 425364
rect 70074 425184 70130 425240
rect 70074 425060 70130 425116
rect 70074 424936 70130 424992
rect 70074 424812 70130 424868
rect 70074 424688 70130 424744
rect 70074 424564 70130 424620
rect 70074 424440 70130 424496
rect 70074 424316 70130 424372
rect 70074 424192 70130 424248
rect 70074 423682 70130 423738
rect 70074 423558 70130 423614
rect 70074 423434 70130 423490
rect 70074 423310 70130 423366
rect 70074 423186 70130 423242
rect 70074 423062 70130 423118
rect 70074 422938 70130 422994
rect 70074 422814 70130 422870
rect 70074 422690 70130 422746
rect 70074 422566 70130 422622
rect 70074 422442 70130 422498
rect 70074 422318 70130 422374
rect 70074 422194 70130 422250
rect 70074 422070 70130 422126
rect 70074 421946 70130 422002
rect 70074 421822 70130 421878
rect 70074 421078 70130 421134
rect 70074 420954 70130 421010
rect 70074 420830 70130 420886
rect 70074 420706 70130 420762
rect 70074 420582 70130 420638
rect 70074 420458 70130 420514
rect 70074 420334 70130 420390
rect 70074 420210 70130 420266
rect 70074 420086 70130 420142
rect 70074 419962 70130 420018
rect 70074 419838 70130 419894
rect 70074 419714 70130 419770
rect 70074 419590 70130 419646
rect 70074 419466 70130 419522
rect 70074 419342 70130 419398
rect 707870 410602 707926 410658
rect 707870 410478 707926 410534
rect 707870 410354 707926 410410
rect 707870 410230 707926 410286
rect 707870 410106 707926 410162
rect 707870 409982 707926 410038
rect 707870 409858 707926 409914
rect 707870 409734 707926 409790
rect 707870 409610 707926 409666
rect 707870 409486 707926 409542
rect 707870 409362 707926 409418
rect 707870 409238 707926 409294
rect 707870 409114 707926 409170
rect 707870 408990 707926 409046
rect 707870 408866 707926 408922
rect 707870 408122 707926 408178
rect 707870 407998 707926 408054
rect 707870 407874 707926 407930
rect 707870 407750 707926 407806
rect 707870 407626 707926 407682
rect 707870 407502 707926 407558
rect 707870 407378 707926 407434
rect 707870 407254 707926 407310
rect 707870 407130 707926 407186
rect 707870 407006 707926 407062
rect 707870 406882 707926 406938
rect 707870 406758 707926 406814
rect 707870 406634 707926 406690
rect 707870 406510 707926 406566
rect 707870 406386 707926 406442
rect 707870 406262 707926 406318
rect 707870 405752 707926 405808
rect 707870 405628 707926 405684
rect 707870 405504 707926 405560
rect 707870 405380 707926 405436
rect 707870 405256 707926 405312
rect 707870 405132 707926 405188
rect 707870 405008 707926 405064
rect 707870 404884 707926 404940
rect 707870 404760 707926 404816
rect 707870 404636 707926 404692
rect 707870 404512 707926 404568
rect 707870 404388 707926 404444
rect 707870 404264 707926 404320
rect 707870 404140 707926 404196
rect 707870 404016 707926 404072
rect 707870 403892 707926 403948
rect 707870 403046 707926 403102
rect 707870 402922 707926 402978
rect 707870 402798 707926 402854
rect 707870 402674 707926 402730
rect 707870 402550 707926 402606
rect 707870 402426 707926 402482
rect 707870 402302 707926 402358
rect 707870 402178 707926 402234
rect 707870 402054 707926 402110
rect 707870 401930 707926 401986
rect 707870 401806 707926 401862
rect 707870 401682 707926 401738
rect 707870 401558 707926 401614
rect 707870 401434 707926 401490
rect 707870 401310 707926 401366
rect 707870 401186 707926 401242
rect 707870 400676 707926 400732
rect 707870 400552 707926 400608
rect 707870 400428 707926 400484
rect 707870 400304 707926 400360
rect 707870 400180 707926 400236
rect 707870 400056 707926 400112
rect 707870 399932 707926 399988
rect 707870 399808 707926 399864
rect 707870 399684 707926 399740
rect 707870 399560 707926 399616
rect 707870 399436 707926 399492
rect 707870 399312 707926 399368
rect 707870 399188 707926 399244
rect 707870 399064 707926 399120
rect 707870 398940 707926 398996
rect 707870 398816 707926 398872
rect 707870 398078 707926 398134
rect 707870 397954 707926 398010
rect 707870 397830 707926 397886
rect 707870 397706 707926 397762
rect 707870 397582 707926 397638
rect 707870 397458 707926 397514
rect 707870 397334 707926 397390
rect 707870 397210 707926 397266
rect 707870 397086 707926 397142
rect 707870 396962 707926 397018
rect 707870 396838 707926 396894
rect 707870 396714 707926 396770
rect 707870 396590 707926 396646
rect 707870 396466 707926 396522
rect 707870 396342 707926 396398
rect 70074 146602 70130 146658
rect 70074 146478 70130 146534
rect 70074 146354 70130 146410
rect 70074 146230 70130 146286
rect 70074 146106 70130 146162
rect 70074 145982 70130 146038
rect 70074 145858 70130 145914
rect 70074 145734 70130 145790
rect 70074 145610 70130 145666
rect 70074 145486 70130 145542
rect 70074 145362 70130 145418
rect 70074 145238 70130 145294
rect 70074 145114 70130 145170
rect 70074 144990 70130 145046
rect 70074 144866 70130 144922
rect 70074 144128 70130 144184
rect 70074 144004 70130 144060
rect 70074 143880 70130 143936
rect 70074 143756 70130 143812
rect 70074 143632 70130 143688
rect 70074 143508 70130 143564
rect 70074 143384 70130 143440
rect 70074 143260 70130 143316
rect 70074 143136 70130 143192
rect 70074 143012 70130 143068
rect 70074 142888 70130 142944
rect 70074 142764 70130 142820
rect 70074 142640 70130 142696
rect 70074 142516 70130 142572
rect 70074 142392 70130 142448
rect 70074 142268 70130 142324
rect 70074 141758 70130 141814
rect 70074 141634 70130 141690
rect 70074 141510 70130 141566
rect 70074 141386 70130 141442
rect 70074 141262 70130 141318
rect 70074 141138 70130 141194
rect 70074 141014 70130 141070
rect 70074 140890 70130 140946
rect 70074 140766 70130 140822
rect 70074 140642 70130 140698
rect 70074 140518 70130 140574
rect 70074 140394 70130 140450
rect 70074 140270 70130 140326
rect 70074 140146 70130 140202
rect 70074 140022 70130 140078
rect 70074 139898 70130 139954
rect 70074 139052 70130 139108
rect 70074 138928 70130 138984
rect 70074 138804 70130 138860
rect 70074 138680 70130 138736
rect 70074 138556 70130 138612
rect 70074 138432 70130 138488
rect 70074 138308 70130 138364
rect 70074 138184 70130 138240
rect 70074 138060 70130 138116
rect 70074 137936 70130 137992
rect 70074 137812 70130 137868
rect 70074 137688 70130 137744
rect 70074 137564 70130 137620
rect 70074 137440 70130 137496
rect 70074 137316 70130 137372
rect 70074 137192 70130 137248
rect 70074 136682 70130 136738
rect 70074 136558 70130 136614
rect 70074 136434 70130 136490
rect 70074 136310 70130 136366
rect 70074 136186 70130 136242
rect 70074 136062 70130 136118
rect 70074 135938 70130 135994
rect 70074 135814 70130 135870
rect 70074 135690 70130 135746
rect 70074 135566 70130 135622
rect 70074 135442 70130 135498
rect 70074 135318 70130 135374
rect 70074 135194 70130 135250
rect 70074 135070 70130 135126
rect 70074 134946 70130 135002
rect 70074 134822 70130 134878
rect 70074 134078 70130 134134
rect 70074 133954 70130 134010
rect 70074 133830 70130 133886
rect 70074 133706 70130 133762
rect 70074 133582 70130 133638
rect 70074 133458 70130 133514
rect 70074 133334 70130 133390
rect 70074 133210 70130 133266
rect 70074 133086 70130 133142
rect 70074 132962 70130 133018
rect 70074 132838 70130 132894
rect 70074 132714 70130 132770
rect 70074 132590 70130 132646
rect 70074 132466 70130 132522
rect 70074 132342 70130 132398
rect 70074 105602 70130 105658
rect 70074 105478 70130 105534
rect 70074 105354 70130 105410
rect 70074 105230 70130 105286
rect 70074 105106 70130 105162
rect 70074 104982 70130 105038
rect 70074 104858 70130 104914
rect 70074 104734 70130 104790
rect 70074 104610 70130 104666
rect 70074 104486 70130 104542
rect 70074 104362 70130 104418
rect 70074 104238 70130 104294
rect 70074 104114 70130 104170
rect 70074 103990 70130 104046
rect 70074 103866 70130 103922
rect 70074 103128 70130 103184
rect 70074 103004 70130 103060
rect 70074 102880 70130 102936
rect 70074 102756 70130 102812
rect 70074 102632 70130 102688
rect 70074 102508 70130 102564
rect 70074 102384 70130 102440
rect 70074 102260 70130 102316
rect 70074 102136 70130 102192
rect 70074 102012 70130 102068
rect 70074 101888 70130 101944
rect 70074 101764 70130 101820
rect 70074 101640 70130 101696
rect 70074 101516 70130 101572
rect 70074 101392 70130 101448
rect 70074 101268 70130 101324
rect 70074 100758 70130 100814
rect 70074 100634 70130 100690
rect 70074 100510 70130 100566
rect 70074 100386 70130 100442
rect 70074 100262 70130 100318
rect 70074 100138 70130 100194
rect 70074 100014 70130 100070
rect 70074 99890 70130 99946
rect 70074 99766 70130 99822
rect 70074 99642 70130 99698
rect 70074 99518 70130 99574
rect 70074 99394 70130 99450
rect 70074 99270 70130 99326
rect 70074 99146 70130 99202
rect 70074 99022 70130 99078
rect 70074 98898 70130 98954
rect 70074 98052 70130 98108
rect 70074 97928 70130 97984
rect 70074 97804 70130 97860
rect 70074 97680 70130 97736
rect 70074 97556 70130 97612
rect 70074 97432 70130 97488
rect 70074 97308 70130 97364
rect 70074 97184 70130 97240
rect 70074 97060 70130 97116
rect 70074 96936 70130 96992
rect 70074 96812 70130 96868
rect 70074 96688 70130 96744
rect 70074 96564 70130 96620
rect 70074 96440 70130 96496
rect 70074 96316 70130 96372
rect 70074 96192 70130 96248
rect 70074 95682 70130 95738
rect 70074 95558 70130 95614
rect 70074 95434 70130 95490
rect 70074 95310 70130 95366
rect 70074 95186 70130 95242
rect 70074 95062 70130 95118
rect 70074 94938 70130 94994
rect 70074 94814 70130 94870
rect 70074 94690 70130 94746
rect 70074 94566 70130 94622
rect 70074 94442 70130 94498
rect 70074 94318 70130 94374
rect 70074 94194 70130 94250
rect 70074 94070 70130 94126
rect 70074 93946 70130 94002
rect 70074 93822 70130 93878
rect 70074 93078 70130 93134
rect 70074 92954 70130 93010
rect 70074 92830 70130 92886
rect 70074 92706 70130 92762
rect 70074 92582 70130 92638
rect 70074 92458 70130 92514
rect 70074 92334 70130 92390
rect 70074 92210 70130 92266
rect 70074 92086 70130 92142
rect 70074 91962 70130 92018
rect 70074 91838 70130 91894
rect 70074 91714 70130 91770
rect 70074 91590 70130 91646
rect 70074 91466 70130 91522
rect 70074 91342 70130 91398
rect 107342 70074 107398 70130
rect 107466 70074 107522 70130
rect 107590 70074 107646 70130
rect 107714 70074 107770 70130
rect 107838 70074 107894 70130
rect 107962 70074 108018 70130
rect 108086 70074 108142 70130
rect 108210 70074 108266 70130
rect 108334 70074 108390 70130
rect 108458 70074 108514 70130
rect 108582 70074 108638 70130
rect 108706 70074 108762 70130
rect 108830 70074 108886 70130
rect 108954 70074 109010 70130
rect 109078 70074 109134 70130
rect 109822 70074 109878 70130
rect 109946 70074 110002 70130
rect 110070 70074 110126 70130
rect 110194 70074 110250 70130
rect 110318 70074 110374 70130
rect 110442 70074 110498 70130
rect 110566 70074 110622 70130
rect 110690 70074 110746 70130
rect 110814 70074 110870 70130
rect 110938 70074 110994 70130
rect 111062 70074 111118 70130
rect 111186 70074 111242 70130
rect 111310 70074 111366 70130
rect 111434 70074 111490 70130
rect 111558 70074 111614 70130
rect 111682 70074 111738 70130
rect 112192 70074 112248 70130
rect 112316 70074 112372 70130
rect 112440 70074 112496 70130
rect 112564 70074 112620 70130
rect 112688 70074 112744 70130
rect 112812 70074 112868 70130
rect 112936 70074 112992 70130
rect 113060 70074 113116 70130
rect 113184 70074 113240 70130
rect 113308 70074 113364 70130
rect 113432 70074 113488 70130
rect 113556 70074 113612 70130
rect 113680 70074 113736 70130
rect 113804 70074 113860 70130
rect 113928 70074 113984 70130
rect 114052 70074 114108 70130
rect 114892 70074 114948 70130
rect 115016 70074 115072 70130
rect 115140 70074 115196 70130
rect 115264 70074 115320 70130
rect 115388 70074 115444 70130
rect 115512 70074 115568 70130
rect 115636 70074 115692 70130
rect 115760 70074 115816 70130
rect 115884 70074 115940 70130
rect 116008 70074 116064 70130
rect 116132 70074 116188 70130
rect 116256 70074 116312 70130
rect 116380 70074 116436 70130
rect 116504 70074 116560 70130
rect 116628 70074 116684 70130
rect 116752 70074 116808 70130
rect 117262 70074 117318 70130
rect 117386 70074 117442 70130
rect 117510 70074 117566 70130
rect 117634 70074 117690 70130
rect 117758 70074 117814 70130
rect 117882 70074 117938 70130
rect 118006 70074 118062 70130
rect 118130 70074 118186 70130
rect 118254 70074 118310 70130
rect 118378 70074 118434 70130
rect 118502 70074 118558 70130
rect 118626 70074 118682 70130
rect 118750 70074 118806 70130
rect 118874 70074 118930 70130
rect 118998 70074 119054 70130
rect 119122 70074 119178 70130
rect 119866 70074 119922 70130
rect 119990 70074 120046 70130
rect 120114 70074 120170 70130
rect 120238 70074 120294 70130
rect 120362 70074 120418 70130
rect 120486 70074 120542 70130
rect 120610 70074 120666 70130
rect 120734 70074 120790 70130
rect 120858 70074 120914 70130
rect 120982 70074 121038 70130
rect 121106 70074 121162 70130
rect 121230 70074 121286 70130
rect 121354 70074 121410 70130
rect 121478 70074 121534 70130
rect 121602 70074 121658 70130
rect 272342 70074 272398 70130
rect 272466 70074 272522 70130
rect 272590 70074 272646 70130
rect 272714 70074 272770 70130
rect 272838 70074 272894 70130
rect 272962 70074 273018 70130
rect 273086 70074 273142 70130
rect 273210 70074 273266 70130
rect 273334 70074 273390 70130
rect 273458 70074 273514 70130
rect 273582 70074 273638 70130
rect 273706 70074 273762 70130
rect 273830 70074 273886 70130
rect 273954 70074 274010 70130
rect 274078 70074 274134 70130
rect 274822 70074 274878 70130
rect 274946 70074 275002 70130
rect 275070 70074 275126 70130
rect 275194 70074 275250 70130
rect 275318 70074 275374 70130
rect 275442 70074 275498 70130
rect 275566 70074 275622 70130
rect 275690 70074 275746 70130
rect 275814 70074 275870 70130
rect 275938 70074 275994 70130
rect 276062 70074 276118 70130
rect 276186 70074 276242 70130
rect 276310 70074 276366 70130
rect 276434 70074 276490 70130
rect 276558 70074 276614 70130
rect 276682 70074 276738 70130
rect 277192 70074 277248 70130
rect 277316 70074 277372 70130
rect 277440 70074 277496 70130
rect 277564 70074 277620 70130
rect 277688 70074 277744 70130
rect 277812 70074 277868 70130
rect 277936 70074 277992 70130
rect 278060 70074 278116 70130
rect 278184 70074 278240 70130
rect 278308 70074 278364 70130
rect 278432 70074 278488 70130
rect 278556 70074 278612 70130
rect 278680 70074 278736 70130
rect 278804 70074 278860 70130
rect 278928 70074 278984 70130
rect 279052 70074 279108 70130
rect 279892 70074 279948 70130
rect 280016 70074 280072 70130
rect 280140 70074 280196 70130
rect 280264 70074 280320 70130
rect 280388 70074 280444 70130
rect 280512 70074 280568 70130
rect 280636 70074 280692 70130
rect 280760 70074 280816 70130
rect 280884 70074 280940 70130
rect 281008 70074 281064 70130
rect 281132 70074 281188 70130
rect 281256 70074 281312 70130
rect 281380 70074 281436 70130
rect 281504 70074 281560 70130
rect 281628 70074 281684 70130
rect 281752 70074 281808 70130
rect 282262 70074 282318 70130
rect 282386 70074 282442 70130
rect 282510 70074 282566 70130
rect 282634 70074 282690 70130
rect 282758 70074 282814 70130
rect 282882 70074 282938 70130
rect 283006 70074 283062 70130
rect 283130 70074 283186 70130
rect 283254 70074 283310 70130
rect 283378 70074 283434 70130
rect 283502 70074 283558 70130
rect 283626 70074 283682 70130
rect 283750 70074 283806 70130
rect 283874 70074 283930 70130
rect 283998 70074 284054 70130
rect 284122 70074 284178 70130
rect 284866 70074 284922 70130
rect 284990 70074 285046 70130
rect 285114 70074 285170 70130
rect 285238 70074 285294 70130
rect 285362 70074 285418 70130
rect 285486 70074 285542 70130
rect 285610 70074 285666 70130
rect 285734 70074 285790 70130
rect 285858 70074 285914 70130
rect 285982 70074 286038 70130
rect 286106 70074 286162 70130
rect 286230 70074 286286 70130
rect 286354 70074 286410 70130
rect 286478 70074 286534 70130
rect 286602 70074 286658 70130
rect 602342 70074 602398 70130
rect 602466 70074 602522 70130
rect 602590 70074 602646 70130
rect 602714 70074 602770 70130
rect 602838 70074 602894 70130
rect 602962 70074 603018 70130
rect 603086 70074 603142 70130
rect 603210 70074 603266 70130
rect 603334 70074 603390 70130
rect 603458 70074 603514 70130
rect 603582 70074 603638 70130
rect 603706 70074 603762 70130
rect 603830 70074 603886 70130
rect 603954 70074 604010 70130
rect 604078 70074 604134 70130
rect 604822 70074 604878 70130
rect 604946 70074 605002 70130
rect 605070 70074 605126 70130
rect 605194 70074 605250 70130
rect 605318 70074 605374 70130
rect 605442 70074 605498 70130
rect 605566 70074 605622 70130
rect 605690 70074 605746 70130
rect 605814 70074 605870 70130
rect 605938 70074 605994 70130
rect 606062 70074 606118 70130
rect 606186 70074 606242 70130
rect 606310 70074 606366 70130
rect 606434 70074 606490 70130
rect 606558 70074 606614 70130
rect 606682 70074 606738 70130
rect 607192 70074 607248 70130
rect 607316 70074 607372 70130
rect 607440 70074 607496 70130
rect 607564 70074 607620 70130
rect 607688 70074 607744 70130
rect 607812 70074 607868 70130
rect 607936 70074 607992 70130
rect 608060 70074 608116 70130
rect 608184 70074 608240 70130
rect 608308 70074 608364 70130
rect 608432 70074 608488 70130
rect 608556 70074 608612 70130
rect 608680 70074 608736 70130
rect 608804 70074 608860 70130
rect 608928 70074 608984 70130
rect 609052 70074 609108 70130
rect 609892 70074 609948 70130
rect 610016 70074 610072 70130
rect 610140 70074 610196 70130
rect 610264 70074 610320 70130
rect 610388 70074 610444 70130
rect 610512 70074 610568 70130
rect 610636 70074 610692 70130
rect 610760 70074 610816 70130
rect 610884 70074 610940 70130
rect 611008 70074 611064 70130
rect 611132 70074 611188 70130
rect 611256 70074 611312 70130
rect 611380 70074 611436 70130
rect 611504 70074 611560 70130
rect 611628 70074 611684 70130
rect 611752 70074 611808 70130
rect 612262 70074 612318 70130
rect 612386 70074 612442 70130
rect 612510 70074 612566 70130
rect 612634 70074 612690 70130
rect 612758 70074 612814 70130
rect 612882 70074 612938 70130
rect 613006 70074 613062 70130
rect 613130 70074 613186 70130
rect 613254 70074 613310 70130
rect 613378 70074 613434 70130
rect 613502 70074 613558 70130
rect 613626 70074 613682 70130
rect 613750 70074 613806 70130
rect 613874 70074 613930 70130
rect 613998 70074 614054 70130
rect 614122 70074 614178 70130
rect 614866 70074 614922 70130
rect 614990 70074 615046 70130
rect 615114 70074 615170 70130
rect 615238 70074 615294 70130
rect 615362 70074 615418 70130
rect 615486 70074 615542 70130
rect 615610 70074 615666 70130
rect 615734 70074 615790 70130
rect 615858 70074 615914 70130
rect 615982 70074 616038 70130
rect 616106 70074 616162 70130
rect 616230 70074 616286 70130
rect 616354 70074 616410 70130
rect 616478 70074 616534 70130
rect 616602 70074 616658 70130
rect 657342 70074 657398 70130
rect 657466 70074 657522 70130
rect 657590 70074 657646 70130
rect 657714 70074 657770 70130
rect 657838 70074 657894 70130
rect 657962 70074 658018 70130
rect 658086 70074 658142 70130
rect 658210 70074 658266 70130
rect 658334 70074 658390 70130
rect 658458 70074 658514 70130
rect 658582 70074 658638 70130
rect 658706 70074 658762 70130
rect 658830 70074 658886 70130
rect 658954 70074 659010 70130
rect 659078 70074 659134 70130
rect 659822 70074 659878 70130
rect 659946 70074 660002 70130
rect 660070 70074 660126 70130
rect 660194 70074 660250 70130
rect 660318 70074 660374 70130
rect 660442 70074 660498 70130
rect 660566 70074 660622 70130
rect 660690 70074 660746 70130
rect 660814 70074 660870 70130
rect 660938 70074 660994 70130
rect 661062 70074 661118 70130
rect 661186 70074 661242 70130
rect 661310 70074 661366 70130
rect 661434 70074 661490 70130
rect 661558 70074 661614 70130
rect 661682 70074 661738 70130
rect 662192 70074 662248 70130
rect 662316 70074 662372 70130
rect 662440 70074 662496 70130
rect 662564 70074 662620 70130
rect 662688 70074 662744 70130
rect 662812 70074 662868 70130
rect 662936 70074 662992 70130
rect 663060 70074 663116 70130
rect 663184 70074 663240 70130
rect 663308 70074 663364 70130
rect 663432 70074 663488 70130
rect 663556 70074 663612 70130
rect 663680 70074 663736 70130
rect 663804 70074 663860 70130
rect 663928 70074 663984 70130
rect 664052 70074 664108 70130
rect 664892 70074 664948 70130
rect 665016 70074 665072 70130
rect 665140 70074 665196 70130
rect 665264 70074 665320 70130
rect 665388 70074 665444 70130
rect 665512 70074 665568 70130
rect 665636 70074 665692 70130
rect 665760 70074 665816 70130
rect 665884 70074 665940 70130
rect 666008 70074 666064 70130
rect 666132 70074 666188 70130
rect 666256 70074 666312 70130
rect 666380 70074 666436 70130
rect 666504 70074 666560 70130
rect 666628 70074 666684 70130
rect 666752 70074 666808 70130
rect 667262 70074 667318 70130
rect 667386 70074 667442 70130
rect 667510 70074 667566 70130
rect 667634 70074 667690 70130
rect 667758 70074 667814 70130
rect 667882 70074 667938 70130
rect 668006 70074 668062 70130
rect 668130 70074 668186 70130
rect 668254 70074 668310 70130
rect 668378 70074 668434 70130
rect 668502 70074 668558 70130
rect 668626 70074 668682 70130
rect 668750 70074 668806 70130
rect 668874 70074 668930 70130
rect 668998 70074 669054 70130
rect 669122 70074 669178 70130
rect 669866 70074 669922 70130
rect 669990 70074 670046 70130
rect 670114 70074 670170 70130
rect 670238 70074 670294 70130
rect 670362 70074 670418 70130
rect 670486 70074 670542 70130
rect 670610 70074 670666 70130
rect 670734 70074 670790 70130
rect 670858 70074 670914 70130
rect 670982 70074 671038 70130
rect 671106 70074 671162 70130
rect 671230 70074 671286 70130
rect 671354 70074 671410 70130
rect 671478 70074 671534 70130
rect 671602 70074 671658 70130
<< metal4 >>
rect 381272 949926 383172 950000
rect 381272 949870 381342 949926
rect 381398 949870 381466 949926
rect 381522 949870 381590 949926
rect 381646 949870 381714 949926
rect 381770 949870 381838 949926
rect 381894 949870 381962 949926
rect 382018 949870 382086 949926
rect 382142 949870 382210 949926
rect 382266 949870 382334 949926
rect 382390 949870 382458 949926
rect 382514 949870 382582 949926
rect 382638 949870 382706 949926
rect 382762 949870 382830 949926
rect 382886 949870 382954 949926
rect 383010 949870 383078 949926
rect 383134 949870 383172 949926
rect 79078 946048 80078 946110
rect 79078 945992 79284 946048
rect 79340 945992 79584 946048
rect 79640 945992 79884 946048
rect 79940 945992 80078 946048
rect 77678 945633 78678 945710
rect 77678 945577 77847 945633
rect 77903 945577 78147 945633
rect 78203 945577 78447 945633
rect 78503 945577 78678 945633
rect 77678 942252 78678 945577
rect 77678 942196 77748 942252
rect 77804 942196 77872 942252
rect 77928 942196 77996 942252
rect 78052 942196 78120 942252
rect 78176 942196 78244 942252
rect 78300 942196 78368 942252
rect 78424 942196 78492 942252
rect 78548 942196 78678 942252
rect 77678 942128 78678 942196
rect 77678 942072 77748 942128
rect 77804 942072 77872 942128
rect 77928 942072 77996 942128
rect 78052 942072 78120 942128
rect 78176 942072 78244 942128
rect 78300 942072 78368 942128
rect 78424 942072 78492 942128
rect 78548 942072 78678 942128
rect 77678 942004 78678 942072
rect 77678 941948 77748 942004
rect 77804 941948 77872 942004
rect 77928 941948 77996 942004
rect 78052 941948 78120 942004
rect 78176 941948 78244 942004
rect 78300 941948 78368 942004
rect 78424 941948 78492 942004
rect 78548 941948 78678 942004
rect 77678 941880 78678 941948
rect 77678 941824 77748 941880
rect 77804 941824 77872 941880
rect 77928 941824 77996 941880
rect 78052 941824 78120 941880
rect 78176 941824 78244 941880
rect 78300 941824 78368 941880
rect 78424 941824 78492 941880
rect 78548 941824 78678 941880
rect 77678 941756 78678 941824
rect 77678 941700 77748 941756
rect 77804 941700 77872 941756
rect 77928 941700 77996 941756
rect 78052 941700 78120 941756
rect 78176 941700 78244 941756
rect 78300 941700 78368 941756
rect 78424 941700 78492 941756
rect 78548 941700 78678 941756
rect 77678 941632 78678 941700
rect 77678 941576 77748 941632
rect 77804 941576 77872 941632
rect 77928 941576 77996 941632
rect 78052 941576 78120 941632
rect 78176 941576 78244 941632
rect 78300 941576 78368 941632
rect 78424 941576 78492 941632
rect 78548 941576 78678 941632
rect 77678 941508 78678 941576
rect 77678 941452 77748 941508
rect 77804 941452 77872 941508
rect 77928 941452 77996 941508
rect 78052 941452 78120 941508
rect 78176 941452 78244 941508
rect 78300 941452 78368 941508
rect 78424 941452 78492 941508
rect 78548 941452 78678 941508
rect 77678 926102 78678 941452
rect 77678 926046 77900 926102
rect 77956 926046 78200 926102
rect 78256 926046 78500 926102
rect 78556 926046 78678 926102
rect 77678 919102 78678 926046
rect 77678 919046 77900 919102
rect 77956 919046 78200 919102
rect 78256 919046 78500 919102
rect 78556 919046 78678 919102
rect 77678 914429 78678 919046
rect 77678 914373 77800 914429
rect 77856 914373 78100 914429
rect 78156 914373 78400 914429
rect 78456 914373 78678 914429
rect 77678 914229 78678 914373
rect 77678 914173 77800 914229
rect 77856 914173 78100 914229
rect 78156 914173 78400 914229
rect 78456 914173 78678 914229
rect 77678 912102 78678 914173
rect 77678 912046 77900 912102
rect 77956 912046 78200 912102
rect 78256 912046 78500 912102
rect 78556 912046 78678 912102
rect 70000 884658 70200 884728
rect 70000 884602 70074 884658
rect 70130 884602 70200 884658
rect 70000 884534 70200 884602
rect 70000 884478 70074 884534
rect 70130 884478 70200 884534
rect 70000 884410 70200 884478
rect 70000 884354 70074 884410
rect 70130 884354 70200 884410
rect 70000 884286 70200 884354
rect 70000 884230 70074 884286
rect 70130 884230 70200 884286
rect 70000 884162 70200 884230
rect 70000 884106 70074 884162
rect 70130 884106 70200 884162
rect 70000 884038 70200 884106
rect 70000 883982 70074 884038
rect 70130 883982 70200 884038
rect 70000 883914 70200 883982
rect 70000 883858 70074 883914
rect 70130 883858 70200 883914
rect 70000 883790 70200 883858
rect 70000 883734 70074 883790
rect 70130 883734 70200 883790
rect 70000 883666 70200 883734
rect 70000 883610 70074 883666
rect 70130 883610 70200 883666
rect 70000 883542 70200 883610
rect 70000 883486 70074 883542
rect 70130 883486 70200 883542
rect 70000 883418 70200 883486
rect 70000 883362 70074 883418
rect 70130 883362 70200 883418
rect 70000 883294 70200 883362
rect 70000 883238 70074 883294
rect 70130 883238 70200 883294
rect 70000 883170 70200 883238
rect 70000 883114 70074 883170
rect 70130 883114 70200 883170
rect 70000 883046 70200 883114
rect 70000 882990 70074 883046
rect 70130 882990 70200 883046
rect 70000 882922 70200 882990
rect 70000 882866 70074 882922
rect 70130 882866 70200 882922
rect 70000 882828 70200 882866
rect 77678 884670 78678 912046
rect 77678 884614 77808 884670
rect 77864 884614 77932 884670
rect 77988 884614 78056 884670
rect 78112 884614 78180 884670
rect 78236 884614 78304 884670
rect 78360 884614 78428 884670
rect 78484 884614 78552 884670
rect 78608 884614 78678 884670
rect 77678 884546 78678 884614
rect 77678 884490 77808 884546
rect 77864 884490 77932 884546
rect 77988 884490 78056 884546
rect 78112 884490 78180 884546
rect 78236 884490 78304 884546
rect 78360 884490 78428 884546
rect 78484 884490 78552 884546
rect 78608 884490 78678 884546
rect 77678 884422 78678 884490
rect 77678 884366 77808 884422
rect 77864 884366 77932 884422
rect 77988 884366 78056 884422
rect 78112 884366 78180 884422
rect 78236 884366 78304 884422
rect 78360 884366 78428 884422
rect 78484 884366 78552 884422
rect 78608 884366 78678 884422
rect 77678 884298 78678 884366
rect 77678 884242 77808 884298
rect 77864 884242 77932 884298
rect 77988 884242 78056 884298
rect 78112 884242 78180 884298
rect 78236 884242 78304 884298
rect 78360 884242 78428 884298
rect 78484 884242 78552 884298
rect 78608 884242 78678 884298
rect 77678 884174 78678 884242
rect 77678 884118 77808 884174
rect 77864 884118 77932 884174
rect 77988 884118 78056 884174
rect 78112 884118 78180 884174
rect 78236 884118 78304 884174
rect 78360 884118 78428 884174
rect 78484 884118 78552 884174
rect 78608 884118 78678 884174
rect 77678 884050 78678 884118
rect 77678 883994 77808 884050
rect 77864 883994 77932 884050
rect 77988 883994 78056 884050
rect 78112 883994 78180 884050
rect 78236 883994 78304 884050
rect 78360 883994 78428 884050
rect 78484 883994 78552 884050
rect 78608 883994 78678 884050
rect 77678 883926 78678 883994
rect 77678 883870 77808 883926
rect 77864 883870 77932 883926
rect 77988 883870 78056 883926
rect 78112 883870 78180 883926
rect 78236 883870 78304 883926
rect 78360 883870 78428 883926
rect 78484 883870 78552 883926
rect 78608 883870 78678 883926
rect 77678 883802 78678 883870
rect 77678 883746 77808 883802
rect 77864 883746 77932 883802
rect 77988 883746 78056 883802
rect 78112 883746 78180 883802
rect 78236 883746 78304 883802
rect 78360 883746 78428 883802
rect 78484 883746 78552 883802
rect 78608 883746 78678 883802
rect 77678 883678 78678 883746
rect 77678 883622 77808 883678
rect 77864 883622 77932 883678
rect 77988 883622 78056 883678
rect 78112 883622 78180 883678
rect 78236 883622 78304 883678
rect 78360 883622 78428 883678
rect 78484 883622 78552 883678
rect 78608 883622 78678 883678
rect 77678 883554 78678 883622
rect 77678 883498 77808 883554
rect 77864 883498 77932 883554
rect 77988 883498 78056 883554
rect 78112 883498 78180 883554
rect 78236 883498 78304 883554
rect 78360 883498 78428 883554
rect 78484 883498 78552 883554
rect 78608 883498 78678 883554
rect 77678 883430 78678 883498
rect 77678 883374 77808 883430
rect 77864 883374 77932 883430
rect 77988 883374 78056 883430
rect 78112 883374 78180 883430
rect 78236 883374 78304 883430
rect 78360 883374 78428 883430
rect 78484 883374 78552 883430
rect 78608 883374 78678 883430
rect 77678 883306 78678 883374
rect 77678 883250 77808 883306
rect 77864 883250 77932 883306
rect 77988 883250 78056 883306
rect 78112 883250 78180 883306
rect 78236 883250 78304 883306
rect 78360 883250 78428 883306
rect 78484 883250 78552 883306
rect 78608 883250 78678 883306
rect 77678 883182 78678 883250
rect 77678 883126 77808 883182
rect 77864 883126 77932 883182
rect 77988 883126 78056 883182
rect 78112 883126 78180 883182
rect 78236 883126 78304 883182
rect 78360 883126 78428 883182
rect 78484 883126 78552 883182
rect 78608 883126 78678 883182
rect 77678 883058 78678 883126
rect 77678 883002 77808 883058
rect 77864 883002 77932 883058
rect 77988 883002 78056 883058
rect 78112 883002 78180 883058
rect 78236 883002 78304 883058
rect 78360 883002 78428 883058
rect 78484 883002 78552 883058
rect 78608 883002 78678 883058
rect 77678 882934 78678 883002
rect 77678 882878 77808 882934
rect 77864 882878 77932 882934
rect 77988 882878 78056 882934
rect 78112 882878 78180 882934
rect 78236 882878 78304 882934
rect 78360 882878 78428 882934
rect 78484 882878 78552 882934
rect 78608 882878 78678 882934
rect 70000 882184 70200 882248
rect 70000 882128 70074 882184
rect 70130 882128 70200 882184
rect 70000 882060 70200 882128
rect 70000 882004 70074 882060
rect 70130 882004 70200 882060
rect 70000 881936 70200 882004
rect 70000 881880 70074 881936
rect 70130 881880 70200 881936
rect 70000 881812 70200 881880
rect 70000 881756 70074 881812
rect 70130 881756 70200 881812
rect 70000 881688 70200 881756
rect 70000 881632 70074 881688
rect 70130 881632 70200 881688
rect 70000 881564 70200 881632
rect 70000 881508 70074 881564
rect 70130 881508 70200 881564
rect 70000 881440 70200 881508
rect 70000 881384 70074 881440
rect 70130 881384 70200 881440
rect 70000 881316 70200 881384
rect 70000 881260 70074 881316
rect 70130 881260 70200 881316
rect 70000 881192 70200 881260
rect 70000 881136 70074 881192
rect 70130 881136 70200 881192
rect 70000 881068 70200 881136
rect 70000 881012 70074 881068
rect 70130 881012 70200 881068
rect 70000 880944 70200 881012
rect 70000 880888 70074 880944
rect 70130 880888 70200 880944
rect 70000 880820 70200 880888
rect 70000 880764 70074 880820
rect 70130 880764 70200 880820
rect 70000 880696 70200 880764
rect 70000 880640 70074 880696
rect 70130 880640 70200 880696
rect 70000 880572 70200 880640
rect 70000 880516 70074 880572
rect 70130 880516 70200 880572
rect 70000 880448 70200 880516
rect 70000 880392 70074 880448
rect 70130 880392 70200 880448
rect 70000 880324 70200 880392
rect 70000 880268 70074 880324
rect 70130 880268 70200 880324
rect 70000 880198 70200 880268
rect 77678 882190 78678 882878
rect 77678 882134 77808 882190
rect 77864 882134 77932 882190
rect 77988 882134 78056 882190
rect 78112 882134 78180 882190
rect 78236 882134 78304 882190
rect 78360 882134 78428 882190
rect 78484 882134 78552 882190
rect 78608 882134 78678 882190
rect 77678 882066 78678 882134
rect 77678 882010 77808 882066
rect 77864 882010 77932 882066
rect 77988 882010 78056 882066
rect 78112 882010 78180 882066
rect 78236 882010 78304 882066
rect 78360 882010 78428 882066
rect 78484 882010 78552 882066
rect 78608 882010 78678 882066
rect 77678 881942 78678 882010
rect 77678 881886 77808 881942
rect 77864 881886 77932 881942
rect 77988 881886 78056 881942
rect 78112 881886 78180 881942
rect 78236 881886 78304 881942
rect 78360 881886 78428 881942
rect 78484 881886 78552 881942
rect 78608 881886 78678 881942
rect 77678 881818 78678 881886
rect 77678 881762 77808 881818
rect 77864 881762 77932 881818
rect 77988 881762 78056 881818
rect 78112 881762 78180 881818
rect 78236 881762 78304 881818
rect 78360 881762 78428 881818
rect 78484 881762 78552 881818
rect 78608 881762 78678 881818
rect 77678 881694 78678 881762
rect 77678 881638 77808 881694
rect 77864 881638 77932 881694
rect 77988 881638 78056 881694
rect 78112 881638 78180 881694
rect 78236 881638 78304 881694
rect 78360 881638 78428 881694
rect 78484 881638 78552 881694
rect 78608 881638 78678 881694
rect 77678 881570 78678 881638
rect 77678 881514 77808 881570
rect 77864 881514 77932 881570
rect 77988 881514 78056 881570
rect 78112 881514 78180 881570
rect 78236 881514 78304 881570
rect 78360 881514 78428 881570
rect 78484 881514 78552 881570
rect 78608 881514 78678 881570
rect 77678 881446 78678 881514
rect 77678 881390 77808 881446
rect 77864 881390 77932 881446
rect 77988 881390 78056 881446
rect 78112 881390 78180 881446
rect 78236 881390 78304 881446
rect 78360 881390 78428 881446
rect 78484 881390 78552 881446
rect 78608 881390 78678 881446
rect 77678 881322 78678 881390
rect 77678 881266 77808 881322
rect 77864 881266 77932 881322
rect 77988 881266 78056 881322
rect 78112 881266 78180 881322
rect 78236 881266 78304 881322
rect 78360 881266 78428 881322
rect 78484 881266 78552 881322
rect 78608 881266 78678 881322
rect 77678 881198 78678 881266
rect 77678 881142 77808 881198
rect 77864 881142 77932 881198
rect 77988 881142 78056 881198
rect 78112 881142 78180 881198
rect 78236 881142 78304 881198
rect 78360 881142 78428 881198
rect 78484 881142 78552 881198
rect 78608 881142 78678 881198
rect 77678 881074 78678 881142
rect 77678 881018 77808 881074
rect 77864 881018 77932 881074
rect 77988 881018 78056 881074
rect 78112 881018 78180 881074
rect 78236 881018 78304 881074
rect 78360 881018 78428 881074
rect 78484 881018 78552 881074
rect 78608 881018 78678 881074
rect 77678 880950 78678 881018
rect 77678 880894 77808 880950
rect 77864 880894 77932 880950
rect 77988 880894 78056 880950
rect 78112 880894 78180 880950
rect 78236 880894 78304 880950
rect 78360 880894 78428 880950
rect 78484 880894 78552 880950
rect 78608 880894 78678 880950
rect 77678 880826 78678 880894
rect 77678 880770 77808 880826
rect 77864 880770 77932 880826
rect 77988 880770 78056 880826
rect 78112 880770 78180 880826
rect 78236 880770 78304 880826
rect 78360 880770 78428 880826
rect 78484 880770 78552 880826
rect 78608 880770 78678 880826
rect 77678 880702 78678 880770
rect 77678 880646 77808 880702
rect 77864 880646 77932 880702
rect 77988 880646 78056 880702
rect 78112 880646 78180 880702
rect 78236 880646 78304 880702
rect 78360 880646 78428 880702
rect 78484 880646 78552 880702
rect 78608 880646 78678 880702
rect 77678 880578 78678 880646
rect 77678 880522 77808 880578
rect 77864 880522 77932 880578
rect 77988 880522 78056 880578
rect 78112 880522 78180 880578
rect 78236 880522 78304 880578
rect 78360 880522 78428 880578
rect 78484 880522 78552 880578
rect 78608 880522 78678 880578
rect 77678 880454 78678 880522
rect 77678 880398 77808 880454
rect 77864 880398 77932 880454
rect 77988 880398 78056 880454
rect 78112 880398 78180 880454
rect 78236 880398 78304 880454
rect 78360 880398 78428 880454
rect 78484 880398 78552 880454
rect 78608 880398 78678 880454
rect 77678 880330 78678 880398
rect 77678 880274 77808 880330
rect 77864 880274 77932 880330
rect 77988 880274 78056 880330
rect 78112 880274 78180 880330
rect 78236 880274 78304 880330
rect 78360 880274 78428 880330
rect 78484 880274 78552 880330
rect 78608 880274 78678 880330
rect 70000 879814 70200 879878
rect 70000 879758 70074 879814
rect 70130 879758 70200 879814
rect 70000 879690 70200 879758
rect 70000 879634 70074 879690
rect 70130 879634 70200 879690
rect 70000 879566 70200 879634
rect 70000 879510 70074 879566
rect 70130 879510 70200 879566
rect 70000 879442 70200 879510
rect 70000 879386 70074 879442
rect 70130 879386 70200 879442
rect 70000 879318 70200 879386
rect 70000 879262 70074 879318
rect 70130 879262 70200 879318
rect 70000 879194 70200 879262
rect 70000 879138 70074 879194
rect 70130 879138 70200 879194
rect 70000 879070 70200 879138
rect 70000 879014 70074 879070
rect 70130 879014 70200 879070
rect 70000 878946 70200 879014
rect 70000 878890 70074 878946
rect 70130 878890 70200 878946
rect 70000 878822 70200 878890
rect 70000 878766 70074 878822
rect 70130 878766 70200 878822
rect 70000 878698 70200 878766
rect 70000 878642 70074 878698
rect 70130 878642 70200 878698
rect 70000 878574 70200 878642
rect 70000 878518 70074 878574
rect 70130 878518 70200 878574
rect 70000 878450 70200 878518
rect 70000 878394 70074 878450
rect 70130 878394 70200 878450
rect 70000 878326 70200 878394
rect 70000 878270 70074 878326
rect 70130 878270 70200 878326
rect 70000 878202 70200 878270
rect 70000 878146 70074 878202
rect 70130 878146 70200 878202
rect 70000 878078 70200 878146
rect 70000 878022 70074 878078
rect 70130 878022 70200 878078
rect 70000 877954 70200 878022
rect 70000 877898 70074 877954
rect 70130 877898 70200 877954
rect 70000 877828 70200 877898
rect 77678 879820 78678 880274
rect 77678 879764 77808 879820
rect 77864 879764 77932 879820
rect 77988 879764 78056 879820
rect 78112 879764 78180 879820
rect 78236 879764 78304 879820
rect 78360 879764 78428 879820
rect 78484 879764 78552 879820
rect 78608 879764 78678 879820
rect 77678 879696 78678 879764
rect 77678 879640 77808 879696
rect 77864 879640 77932 879696
rect 77988 879640 78056 879696
rect 78112 879640 78180 879696
rect 78236 879640 78304 879696
rect 78360 879640 78428 879696
rect 78484 879640 78552 879696
rect 78608 879640 78678 879696
rect 77678 879572 78678 879640
rect 77678 879516 77808 879572
rect 77864 879516 77932 879572
rect 77988 879516 78056 879572
rect 78112 879516 78180 879572
rect 78236 879516 78304 879572
rect 78360 879516 78428 879572
rect 78484 879516 78552 879572
rect 78608 879516 78678 879572
rect 77678 879448 78678 879516
rect 77678 879392 77808 879448
rect 77864 879392 77932 879448
rect 77988 879392 78056 879448
rect 78112 879392 78180 879448
rect 78236 879392 78304 879448
rect 78360 879392 78428 879448
rect 78484 879392 78552 879448
rect 78608 879392 78678 879448
rect 77678 879324 78678 879392
rect 77678 879268 77808 879324
rect 77864 879268 77932 879324
rect 77988 879268 78056 879324
rect 78112 879268 78180 879324
rect 78236 879268 78304 879324
rect 78360 879268 78428 879324
rect 78484 879268 78552 879324
rect 78608 879268 78678 879324
rect 77678 879200 78678 879268
rect 77678 879144 77808 879200
rect 77864 879144 77932 879200
rect 77988 879144 78056 879200
rect 78112 879144 78180 879200
rect 78236 879144 78304 879200
rect 78360 879144 78428 879200
rect 78484 879144 78552 879200
rect 78608 879144 78678 879200
rect 77678 879076 78678 879144
rect 77678 879020 77808 879076
rect 77864 879020 77932 879076
rect 77988 879020 78056 879076
rect 78112 879020 78180 879076
rect 78236 879020 78304 879076
rect 78360 879020 78428 879076
rect 78484 879020 78552 879076
rect 78608 879020 78678 879076
rect 77678 878952 78678 879020
rect 77678 878896 77808 878952
rect 77864 878896 77932 878952
rect 77988 878896 78056 878952
rect 78112 878896 78180 878952
rect 78236 878896 78304 878952
rect 78360 878896 78428 878952
rect 78484 878896 78552 878952
rect 78608 878896 78678 878952
rect 77678 878828 78678 878896
rect 77678 878772 77808 878828
rect 77864 878772 77932 878828
rect 77988 878772 78056 878828
rect 78112 878772 78180 878828
rect 78236 878772 78304 878828
rect 78360 878772 78428 878828
rect 78484 878772 78552 878828
rect 78608 878772 78678 878828
rect 77678 878704 78678 878772
rect 77678 878648 77808 878704
rect 77864 878648 77932 878704
rect 77988 878648 78056 878704
rect 78112 878648 78180 878704
rect 78236 878648 78304 878704
rect 78360 878648 78428 878704
rect 78484 878648 78552 878704
rect 78608 878648 78678 878704
rect 77678 878580 78678 878648
rect 77678 878524 77808 878580
rect 77864 878524 77932 878580
rect 77988 878524 78056 878580
rect 78112 878524 78180 878580
rect 78236 878524 78304 878580
rect 78360 878524 78428 878580
rect 78484 878524 78552 878580
rect 78608 878524 78678 878580
rect 77678 878456 78678 878524
rect 77678 878400 77808 878456
rect 77864 878400 77932 878456
rect 77988 878400 78056 878456
rect 78112 878400 78180 878456
rect 78236 878400 78304 878456
rect 78360 878400 78428 878456
rect 78484 878400 78552 878456
rect 78608 878400 78678 878456
rect 77678 878332 78678 878400
rect 77678 878276 77808 878332
rect 77864 878276 77932 878332
rect 77988 878276 78056 878332
rect 78112 878276 78180 878332
rect 78236 878276 78304 878332
rect 78360 878276 78428 878332
rect 78484 878276 78552 878332
rect 78608 878276 78678 878332
rect 77678 878208 78678 878276
rect 77678 878152 77808 878208
rect 77864 878152 77932 878208
rect 77988 878152 78056 878208
rect 78112 878152 78180 878208
rect 78236 878152 78304 878208
rect 78360 878152 78428 878208
rect 78484 878152 78552 878208
rect 78608 878152 78678 878208
rect 77678 878084 78678 878152
rect 77678 878028 77808 878084
rect 77864 878028 77932 878084
rect 77988 878028 78056 878084
rect 78112 878028 78180 878084
rect 78236 878028 78304 878084
rect 78360 878028 78428 878084
rect 78484 878028 78552 878084
rect 78608 878028 78678 878084
rect 77678 877960 78678 878028
rect 77678 877904 77808 877960
rect 77864 877904 77932 877960
rect 77988 877904 78056 877960
rect 78112 877904 78180 877960
rect 78236 877904 78304 877960
rect 78360 877904 78428 877960
rect 78484 877904 78552 877960
rect 78608 877904 78678 877960
rect 70000 877108 70200 877172
rect 70000 877052 70074 877108
rect 70130 877052 70200 877108
rect 70000 876984 70200 877052
rect 70000 876928 70074 876984
rect 70130 876928 70200 876984
rect 70000 876860 70200 876928
rect 70000 876804 70074 876860
rect 70130 876804 70200 876860
rect 70000 876736 70200 876804
rect 70000 876680 70074 876736
rect 70130 876680 70200 876736
rect 70000 876612 70200 876680
rect 70000 876556 70074 876612
rect 70130 876556 70200 876612
rect 70000 876488 70200 876556
rect 70000 876432 70074 876488
rect 70130 876432 70200 876488
rect 70000 876364 70200 876432
rect 70000 876308 70074 876364
rect 70130 876308 70200 876364
rect 70000 876240 70200 876308
rect 70000 876184 70074 876240
rect 70130 876184 70200 876240
rect 70000 876116 70200 876184
rect 70000 876060 70074 876116
rect 70130 876060 70200 876116
rect 70000 875992 70200 876060
rect 70000 875936 70074 875992
rect 70130 875936 70200 875992
rect 70000 875868 70200 875936
rect 70000 875812 70074 875868
rect 70130 875812 70200 875868
rect 70000 875744 70200 875812
rect 70000 875688 70074 875744
rect 70130 875688 70200 875744
rect 70000 875620 70200 875688
rect 70000 875564 70074 875620
rect 70130 875564 70200 875620
rect 70000 875496 70200 875564
rect 70000 875440 70074 875496
rect 70130 875440 70200 875496
rect 70000 875372 70200 875440
rect 70000 875316 70074 875372
rect 70130 875316 70200 875372
rect 70000 875248 70200 875316
rect 70000 875192 70074 875248
rect 70130 875192 70200 875248
rect 70000 875122 70200 875192
rect 77678 877114 78678 877904
rect 77678 877058 77808 877114
rect 77864 877058 77932 877114
rect 77988 877058 78056 877114
rect 78112 877058 78180 877114
rect 78236 877058 78304 877114
rect 78360 877058 78428 877114
rect 78484 877058 78552 877114
rect 78608 877058 78678 877114
rect 77678 876990 78678 877058
rect 77678 876934 77808 876990
rect 77864 876934 77932 876990
rect 77988 876934 78056 876990
rect 78112 876934 78180 876990
rect 78236 876934 78304 876990
rect 78360 876934 78428 876990
rect 78484 876934 78552 876990
rect 78608 876934 78678 876990
rect 77678 876866 78678 876934
rect 77678 876810 77808 876866
rect 77864 876810 77932 876866
rect 77988 876810 78056 876866
rect 78112 876810 78180 876866
rect 78236 876810 78304 876866
rect 78360 876810 78428 876866
rect 78484 876810 78552 876866
rect 78608 876810 78678 876866
rect 77678 876742 78678 876810
rect 77678 876686 77808 876742
rect 77864 876686 77932 876742
rect 77988 876686 78056 876742
rect 78112 876686 78180 876742
rect 78236 876686 78304 876742
rect 78360 876686 78428 876742
rect 78484 876686 78552 876742
rect 78608 876686 78678 876742
rect 77678 876618 78678 876686
rect 77678 876562 77808 876618
rect 77864 876562 77932 876618
rect 77988 876562 78056 876618
rect 78112 876562 78180 876618
rect 78236 876562 78304 876618
rect 78360 876562 78428 876618
rect 78484 876562 78552 876618
rect 78608 876562 78678 876618
rect 77678 876494 78678 876562
rect 77678 876438 77808 876494
rect 77864 876438 77932 876494
rect 77988 876438 78056 876494
rect 78112 876438 78180 876494
rect 78236 876438 78304 876494
rect 78360 876438 78428 876494
rect 78484 876438 78552 876494
rect 78608 876438 78678 876494
rect 77678 876370 78678 876438
rect 77678 876314 77808 876370
rect 77864 876314 77932 876370
rect 77988 876314 78056 876370
rect 78112 876314 78180 876370
rect 78236 876314 78304 876370
rect 78360 876314 78428 876370
rect 78484 876314 78552 876370
rect 78608 876314 78678 876370
rect 77678 876246 78678 876314
rect 77678 876190 77808 876246
rect 77864 876190 77932 876246
rect 77988 876190 78056 876246
rect 78112 876190 78180 876246
rect 78236 876190 78304 876246
rect 78360 876190 78428 876246
rect 78484 876190 78552 876246
rect 78608 876190 78678 876246
rect 77678 876122 78678 876190
rect 77678 876066 77808 876122
rect 77864 876066 77932 876122
rect 77988 876066 78056 876122
rect 78112 876066 78180 876122
rect 78236 876066 78304 876122
rect 78360 876066 78428 876122
rect 78484 876066 78552 876122
rect 78608 876066 78678 876122
rect 77678 875998 78678 876066
rect 77678 875942 77808 875998
rect 77864 875942 77932 875998
rect 77988 875942 78056 875998
rect 78112 875942 78180 875998
rect 78236 875942 78304 875998
rect 78360 875942 78428 875998
rect 78484 875942 78552 875998
rect 78608 875942 78678 875998
rect 77678 875874 78678 875942
rect 77678 875818 77808 875874
rect 77864 875818 77932 875874
rect 77988 875818 78056 875874
rect 78112 875818 78180 875874
rect 78236 875818 78304 875874
rect 78360 875818 78428 875874
rect 78484 875818 78552 875874
rect 78608 875818 78678 875874
rect 77678 875750 78678 875818
rect 77678 875694 77808 875750
rect 77864 875694 77932 875750
rect 77988 875694 78056 875750
rect 78112 875694 78180 875750
rect 78236 875694 78304 875750
rect 78360 875694 78428 875750
rect 78484 875694 78552 875750
rect 78608 875694 78678 875750
rect 77678 875626 78678 875694
rect 77678 875570 77808 875626
rect 77864 875570 77932 875626
rect 77988 875570 78056 875626
rect 78112 875570 78180 875626
rect 78236 875570 78304 875626
rect 78360 875570 78428 875626
rect 78484 875570 78552 875626
rect 78608 875570 78678 875626
rect 77678 875502 78678 875570
rect 77678 875446 77808 875502
rect 77864 875446 77932 875502
rect 77988 875446 78056 875502
rect 78112 875446 78180 875502
rect 78236 875446 78304 875502
rect 78360 875446 78428 875502
rect 78484 875446 78552 875502
rect 78608 875446 78678 875502
rect 77678 875378 78678 875446
rect 77678 875322 77808 875378
rect 77864 875322 77932 875378
rect 77988 875322 78056 875378
rect 78112 875322 78180 875378
rect 78236 875322 78304 875378
rect 78360 875322 78428 875378
rect 78484 875322 78552 875378
rect 78608 875322 78678 875378
rect 77678 875254 78678 875322
rect 77678 875198 77808 875254
rect 77864 875198 77932 875254
rect 77988 875198 78056 875254
rect 78112 875198 78180 875254
rect 78236 875198 78304 875254
rect 78360 875198 78428 875254
rect 78484 875198 78552 875254
rect 78608 875198 78678 875254
rect 70000 874738 70200 874802
rect 70000 874682 70074 874738
rect 70130 874682 70200 874738
rect 70000 874614 70200 874682
rect 70000 874558 70074 874614
rect 70130 874558 70200 874614
rect 70000 874490 70200 874558
rect 70000 874434 70074 874490
rect 70130 874434 70200 874490
rect 70000 874366 70200 874434
rect 70000 874310 70074 874366
rect 70130 874310 70200 874366
rect 70000 874242 70200 874310
rect 70000 874186 70074 874242
rect 70130 874186 70200 874242
rect 70000 874118 70200 874186
rect 70000 874062 70074 874118
rect 70130 874062 70200 874118
rect 70000 873994 70200 874062
rect 70000 873938 70074 873994
rect 70130 873938 70200 873994
rect 70000 873870 70200 873938
rect 70000 873814 70074 873870
rect 70130 873814 70200 873870
rect 70000 873746 70200 873814
rect 70000 873690 70074 873746
rect 70130 873690 70200 873746
rect 70000 873622 70200 873690
rect 70000 873566 70074 873622
rect 70130 873566 70200 873622
rect 70000 873498 70200 873566
rect 70000 873442 70074 873498
rect 70130 873442 70200 873498
rect 70000 873374 70200 873442
rect 70000 873318 70074 873374
rect 70130 873318 70200 873374
rect 70000 873250 70200 873318
rect 70000 873194 70074 873250
rect 70130 873194 70200 873250
rect 70000 873126 70200 873194
rect 70000 873070 70074 873126
rect 70130 873070 70200 873126
rect 70000 873002 70200 873070
rect 70000 872946 70074 873002
rect 70130 872946 70200 873002
rect 70000 872878 70200 872946
rect 70000 872822 70074 872878
rect 70130 872822 70200 872878
rect 70000 872752 70200 872822
rect 77678 874744 78678 875198
rect 77678 874688 77808 874744
rect 77864 874688 77932 874744
rect 77988 874688 78056 874744
rect 78112 874688 78180 874744
rect 78236 874688 78304 874744
rect 78360 874688 78428 874744
rect 78484 874688 78552 874744
rect 78608 874688 78678 874744
rect 77678 874620 78678 874688
rect 77678 874564 77808 874620
rect 77864 874564 77932 874620
rect 77988 874564 78056 874620
rect 78112 874564 78180 874620
rect 78236 874564 78304 874620
rect 78360 874564 78428 874620
rect 78484 874564 78552 874620
rect 78608 874564 78678 874620
rect 77678 874496 78678 874564
rect 77678 874440 77808 874496
rect 77864 874440 77932 874496
rect 77988 874440 78056 874496
rect 78112 874440 78180 874496
rect 78236 874440 78304 874496
rect 78360 874440 78428 874496
rect 78484 874440 78552 874496
rect 78608 874440 78678 874496
rect 77678 874372 78678 874440
rect 77678 874316 77808 874372
rect 77864 874316 77932 874372
rect 77988 874316 78056 874372
rect 78112 874316 78180 874372
rect 78236 874316 78304 874372
rect 78360 874316 78428 874372
rect 78484 874316 78552 874372
rect 78608 874316 78678 874372
rect 77678 874248 78678 874316
rect 77678 874192 77808 874248
rect 77864 874192 77932 874248
rect 77988 874192 78056 874248
rect 78112 874192 78180 874248
rect 78236 874192 78304 874248
rect 78360 874192 78428 874248
rect 78484 874192 78552 874248
rect 78608 874192 78678 874248
rect 77678 874124 78678 874192
rect 77678 874068 77808 874124
rect 77864 874068 77932 874124
rect 77988 874068 78056 874124
rect 78112 874068 78180 874124
rect 78236 874068 78304 874124
rect 78360 874068 78428 874124
rect 78484 874068 78552 874124
rect 78608 874068 78678 874124
rect 77678 874000 78678 874068
rect 77678 873944 77808 874000
rect 77864 873944 77932 874000
rect 77988 873944 78056 874000
rect 78112 873944 78180 874000
rect 78236 873944 78304 874000
rect 78360 873944 78428 874000
rect 78484 873944 78552 874000
rect 78608 873944 78678 874000
rect 77678 873876 78678 873944
rect 77678 873820 77808 873876
rect 77864 873820 77932 873876
rect 77988 873820 78056 873876
rect 78112 873820 78180 873876
rect 78236 873820 78304 873876
rect 78360 873820 78428 873876
rect 78484 873820 78552 873876
rect 78608 873820 78678 873876
rect 77678 873752 78678 873820
rect 77678 873696 77808 873752
rect 77864 873696 77932 873752
rect 77988 873696 78056 873752
rect 78112 873696 78180 873752
rect 78236 873696 78304 873752
rect 78360 873696 78428 873752
rect 78484 873696 78552 873752
rect 78608 873696 78678 873752
rect 77678 873628 78678 873696
rect 77678 873572 77808 873628
rect 77864 873572 77932 873628
rect 77988 873572 78056 873628
rect 78112 873572 78180 873628
rect 78236 873572 78304 873628
rect 78360 873572 78428 873628
rect 78484 873572 78552 873628
rect 78608 873572 78678 873628
rect 77678 873504 78678 873572
rect 77678 873448 77808 873504
rect 77864 873448 77932 873504
rect 77988 873448 78056 873504
rect 78112 873448 78180 873504
rect 78236 873448 78304 873504
rect 78360 873448 78428 873504
rect 78484 873448 78552 873504
rect 78608 873448 78678 873504
rect 77678 873380 78678 873448
rect 77678 873324 77808 873380
rect 77864 873324 77932 873380
rect 77988 873324 78056 873380
rect 78112 873324 78180 873380
rect 78236 873324 78304 873380
rect 78360 873324 78428 873380
rect 78484 873324 78552 873380
rect 78608 873324 78678 873380
rect 77678 873256 78678 873324
rect 77678 873200 77808 873256
rect 77864 873200 77932 873256
rect 77988 873200 78056 873256
rect 78112 873200 78180 873256
rect 78236 873200 78304 873256
rect 78360 873200 78428 873256
rect 78484 873200 78552 873256
rect 78608 873200 78678 873256
rect 77678 873132 78678 873200
rect 77678 873076 77808 873132
rect 77864 873076 77932 873132
rect 77988 873076 78056 873132
rect 78112 873076 78180 873132
rect 78236 873076 78304 873132
rect 78360 873076 78428 873132
rect 78484 873076 78552 873132
rect 78608 873076 78678 873132
rect 77678 873008 78678 873076
rect 77678 872952 77808 873008
rect 77864 872952 77932 873008
rect 77988 872952 78056 873008
rect 78112 872952 78180 873008
rect 78236 872952 78304 873008
rect 78360 872952 78428 873008
rect 78484 872952 78552 873008
rect 78608 872952 78678 873008
rect 77678 872884 78678 872952
rect 77678 872828 77808 872884
rect 77864 872828 77932 872884
rect 77988 872828 78056 872884
rect 78112 872828 78180 872884
rect 78236 872828 78304 872884
rect 78360 872828 78428 872884
rect 78484 872828 78552 872884
rect 78608 872828 78678 872884
rect 70000 872134 70200 872172
rect 70000 872078 70074 872134
rect 70130 872078 70200 872134
rect 70000 872010 70200 872078
rect 70000 871954 70074 872010
rect 70130 871954 70200 872010
rect 70000 871886 70200 871954
rect 70000 871830 70074 871886
rect 70130 871830 70200 871886
rect 70000 871762 70200 871830
rect 70000 871706 70074 871762
rect 70130 871706 70200 871762
rect 70000 871638 70200 871706
rect 70000 871582 70074 871638
rect 70130 871582 70200 871638
rect 70000 871514 70200 871582
rect 70000 871458 70074 871514
rect 70130 871458 70200 871514
rect 70000 871390 70200 871458
rect 70000 871334 70074 871390
rect 70130 871334 70200 871390
rect 70000 871266 70200 871334
rect 70000 871210 70074 871266
rect 70130 871210 70200 871266
rect 70000 871142 70200 871210
rect 70000 871086 70074 871142
rect 70130 871086 70200 871142
rect 70000 871018 70200 871086
rect 70000 870962 70074 871018
rect 70130 870962 70200 871018
rect 70000 870894 70200 870962
rect 70000 870838 70074 870894
rect 70130 870838 70200 870894
rect 70000 870770 70200 870838
rect 70000 870714 70074 870770
rect 70130 870714 70200 870770
rect 70000 870646 70200 870714
rect 70000 870590 70074 870646
rect 70130 870590 70200 870646
rect 70000 870522 70200 870590
rect 70000 870466 70074 870522
rect 70130 870466 70200 870522
rect 70000 870398 70200 870466
rect 70000 870342 70074 870398
rect 70130 870342 70200 870398
rect 70000 870272 70200 870342
rect 77678 872140 78678 872828
rect 77678 872084 77808 872140
rect 77864 872084 77932 872140
rect 77988 872084 78056 872140
rect 78112 872084 78180 872140
rect 78236 872084 78304 872140
rect 78360 872084 78428 872140
rect 78484 872084 78552 872140
rect 78608 872084 78678 872140
rect 77678 872016 78678 872084
rect 77678 871960 77808 872016
rect 77864 871960 77932 872016
rect 77988 871960 78056 872016
rect 78112 871960 78180 872016
rect 78236 871960 78304 872016
rect 78360 871960 78428 872016
rect 78484 871960 78552 872016
rect 78608 871960 78678 872016
rect 77678 871892 78678 871960
rect 77678 871836 77808 871892
rect 77864 871836 77932 871892
rect 77988 871836 78056 871892
rect 78112 871836 78180 871892
rect 78236 871836 78304 871892
rect 78360 871836 78428 871892
rect 78484 871836 78552 871892
rect 78608 871836 78678 871892
rect 77678 871768 78678 871836
rect 77678 871712 77808 871768
rect 77864 871712 77932 871768
rect 77988 871712 78056 871768
rect 78112 871712 78180 871768
rect 78236 871712 78304 871768
rect 78360 871712 78428 871768
rect 78484 871712 78552 871768
rect 78608 871712 78678 871768
rect 77678 871644 78678 871712
rect 77678 871588 77808 871644
rect 77864 871588 77932 871644
rect 77988 871588 78056 871644
rect 78112 871588 78180 871644
rect 78236 871588 78304 871644
rect 78360 871588 78428 871644
rect 78484 871588 78552 871644
rect 78608 871588 78678 871644
rect 77678 871520 78678 871588
rect 77678 871464 77808 871520
rect 77864 871464 77932 871520
rect 77988 871464 78056 871520
rect 78112 871464 78180 871520
rect 78236 871464 78304 871520
rect 78360 871464 78428 871520
rect 78484 871464 78552 871520
rect 78608 871464 78678 871520
rect 77678 871396 78678 871464
rect 77678 871340 77808 871396
rect 77864 871340 77932 871396
rect 77988 871340 78056 871396
rect 78112 871340 78180 871396
rect 78236 871340 78304 871396
rect 78360 871340 78428 871396
rect 78484 871340 78552 871396
rect 78608 871340 78678 871396
rect 77678 871272 78678 871340
rect 77678 871216 77808 871272
rect 77864 871216 77932 871272
rect 77988 871216 78056 871272
rect 78112 871216 78180 871272
rect 78236 871216 78304 871272
rect 78360 871216 78428 871272
rect 78484 871216 78552 871272
rect 78608 871216 78678 871272
rect 77678 871148 78678 871216
rect 77678 871092 77808 871148
rect 77864 871092 77932 871148
rect 77988 871092 78056 871148
rect 78112 871092 78180 871148
rect 78236 871092 78304 871148
rect 78360 871092 78428 871148
rect 78484 871092 78552 871148
rect 78608 871092 78678 871148
rect 77678 871024 78678 871092
rect 77678 870968 77808 871024
rect 77864 870968 77932 871024
rect 77988 870968 78056 871024
rect 78112 870968 78180 871024
rect 78236 870968 78304 871024
rect 78360 870968 78428 871024
rect 78484 870968 78552 871024
rect 78608 870968 78678 871024
rect 77678 870900 78678 870968
rect 77678 870844 77808 870900
rect 77864 870844 77932 870900
rect 77988 870844 78056 870900
rect 78112 870844 78180 870900
rect 78236 870844 78304 870900
rect 78360 870844 78428 870900
rect 78484 870844 78552 870900
rect 78608 870844 78678 870900
rect 77678 870776 78678 870844
rect 77678 870720 77808 870776
rect 77864 870720 77932 870776
rect 77988 870720 78056 870776
rect 78112 870720 78180 870776
rect 78236 870720 78304 870776
rect 78360 870720 78428 870776
rect 78484 870720 78552 870776
rect 78608 870720 78678 870776
rect 77678 870652 78678 870720
rect 77678 870596 77808 870652
rect 77864 870596 77932 870652
rect 77988 870596 78056 870652
rect 78112 870596 78180 870652
rect 78236 870596 78304 870652
rect 78360 870596 78428 870652
rect 78484 870596 78552 870652
rect 78608 870596 78678 870652
rect 77678 870528 78678 870596
rect 77678 870472 77808 870528
rect 77864 870472 77932 870528
rect 77988 870472 78056 870528
rect 78112 870472 78180 870528
rect 78236 870472 78304 870528
rect 78360 870472 78428 870528
rect 78484 870472 78552 870528
rect 78608 870472 78678 870528
rect 77678 870404 78678 870472
rect 77678 870348 77808 870404
rect 77864 870348 77932 870404
rect 77988 870348 78056 870404
rect 78112 870348 78180 870404
rect 78236 870348 78304 870404
rect 78360 870348 78428 870404
rect 78484 870348 78552 870404
rect 78608 870348 78678 870404
rect 70000 843658 70200 843728
rect 70000 843602 70074 843658
rect 70130 843602 70200 843658
rect 70000 843534 70200 843602
rect 70000 843478 70074 843534
rect 70130 843478 70200 843534
rect 70000 843410 70200 843478
rect 70000 843354 70074 843410
rect 70130 843354 70200 843410
rect 70000 843286 70200 843354
rect 70000 843230 70074 843286
rect 70130 843230 70200 843286
rect 70000 843162 70200 843230
rect 70000 843106 70074 843162
rect 70130 843106 70200 843162
rect 70000 843038 70200 843106
rect 70000 842982 70074 843038
rect 70130 842982 70200 843038
rect 70000 842914 70200 842982
rect 70000 842858 70074 842914
rect 70130 842858 70200 842914
rect 70000 842790 70200 842858
rect 70000 842734 70074 842790
rect 70130 842734 70200 842790
rect 70000 842666 70200 842734
rect 70000 842610 70074 842666
rect 70130 842610 70200 842666
rect 70000 842542 70200 842610
rect 70000 842486 70074 842542
rect 70130 842486 70200 842542
rect 70000 842418 70200 842486
rect 70000 842362 70074 842418
rect 70130 842362 70200 842418
rect 70000 842294 70200 842362
rect 70000 842238 70074 842294
rect 70130 842238 70200 842294
rect 70000 842170 70200 842238
rect 70000 842114 70074 842170
rect 70130 842114 70200 842170
rect 70000 842046 70200 842114
rect 70000 841990 70074 842046
rect 70130 841990 70200 842046
rect 70000 841922 70200 841990
rect 70000 841866 70074 841922
rect 70130 841866 70200 841922
rect 70000 841828 70200 841866
rect 77678 843670 78678 870348
rect 77678 843614 77808 843670
rect 77864 843614 77932 843670
rect 77988 843614 78056 843670
rect 78112 843614 78180 843670
rect 78236 843614 78304 843670
rect 78360 843614 78428 843670
rect 78484 843614 78552 843670
rect 78608 843614 78678 843670
rect 77678 843546 78678 843614
rect 77678 843490 77808 843546
rect 77864 843490 77932 843546
rect 77988 843490 78056 843546
rect 78112 843490 78180 843546
rect 78236 843490 78304 843546
rect 78360 843490 78428 843546
rect 78484 843490 78552 843546
rect 78608 843490 78678 843546
rect 77678 843422 78678 843490
rect 77678 843366 77808 843422
rect 77864 843366 77932 843422
rect 77988 843366 78056 843422
rect 78112 843366 78180 843422
rect 78236 843366 78304 843422
rect 78360 843366 78428 843422
rect 78484 843366 78552 843422
rect 78608 843366 78678 843422
rect 77678 843298 78678 843366
rect 77678 843242 77808 843298
rect 77864 843242 77932 843298
rect 77988 843242 78056 843298
rect 78112 843242 78180 843298
rect 78236 843242 78304 843298
rect 78360 843242 78428 843298
rect 78484 843242 78552 843298
rect 78608 843242 78678 843298
rect 77678 843174 78678 843242
rect 77678 843118 77808 843174
rect 77864 843118 77932 843174
rect 77988 843118 78056 843174
rect 78112 843118 78180 843174
rect 78236 843118 78304 843174
rect 78360 843118 78428 843174
rect 78484 843118 78552 843174
rect 78608 843118 78678 843174
rect 77678 843050 78678 843118
rect 77678 842994 77808 843050
rect 77864 842994 77932 843050
rect 77988 842994 78056 843050
rect 78112 842994 78180 843050
rect 78236 842994 78304 843050
rect 78360 842994 78428 843050
rect 78484 842994 78552 843050
rect 78608 842994 78678 843050
rect 77678 842926 78678 842994
rect 77678 842870 77808 842926
rect 77864 842870 77932 842926
rect 77988 842870 78056 842926
rect 78112 842870 78180 842926
rect 78236 842870 78304 842926
rect 78360 842870 78428 842926
rect 78484 842870 78552 842926
rect 78608 842870 78678 842926
rect 77678 842802 78678 842870
rect 77678 842746 77808 842802
rect 77864 842746 77932 842802
rect 77988 842746 78056 842802
rect 78112 842746 78180 842802
rect 78236 842746 78304 842802
rect 78360 842746 78428 842802
rect 78484 842746 78552 842802
rect 78608 842746 78678 842802
rect 77678 842678 78678 842746
rect 77678 842622 77808 842678
rect 77864 842622 77932 842678
rect 77988 842622 78056 842678
rect 78112 842622 78180 842678
rect 78236 842622 78304 842678
rect 78360 842622 78428 842678
rect 78484 842622 78552 842678
rect 78608 842622 78678 842678
rect 77678 842554 78678 842622
rect 77678 842498 77808 842554
rect 77864 842498 77932 842554
rect 77988 842498 78056 842554
rect 78112 842498 78180 842554
rect 78236 842498 78304 842554
rect 78360 842498 78428 842554
rect 78484 842498 78552 842554
rect 78608 842498 78678 842554
rect 77678 842430 78678 842498
rect 77678 842374 77808 842430
rect 77864 842374 77932 842430
rect 77988 842374 78056 842430
rect 78112 842374 78180 842430
rect 78236 842374 78304 842430
rect 78360 842374 78428 842430
rect 78484 842374 78552 842430
rect 78608 842374 78678 842430
rect 77678 842306 78678 842374
rect 77678 842250 77808 842306
rect 77864 842250 77932 842306
rect 77988 842250 78056 842306
rect 78112 842250 78180 842306
rect 78236 842250 78304 842306
rect 78360 842250 78428 842306
rect 78484 842250 78552 842306
rect 78608 842250 78678 842306
rect 77678 842182 78678 842250
rect 77678 842126 77808 842182
rect 77864 842126 77932 842182
rect 77988 842126 78056 842182
rect 78112 842126 78180 842182
rect 78236 842126 78304 842182
rect 78360 842126 78428 842182
rect 78484 842126 78552 842182
rect 78608 842126 78678 842182
rect 77678 842058 78678 842126
rect 77678 842002 77808 842058
rect 77864 842002 77932 842058
rect 77988 842002 78056 842058
rect 78112 842002 78180 842058
rect 78236 842002 78304 842058
rect 78360 842002 78428 842058
rect 78484 842002 78552 842058
rect 78608 842002 78678 842058
rect 77678 841934 78678 842002
rect 77678 841878 77808 841934
rect 77864 841878 77932 841934
rect 77988 841878 78056 841934
rect 78112 841878 78180 841934
rect 78236 841878 78304 841934
rect 78360 841878 78428 841934
rect 78484 841878 78552 841934
rect 78608 841878 78678 841934
rect 70000 841184 70200 841248
rect 70000 841128 70074 841184
rect 70130 841128 70200 841184
rect 70000 841060 70200 841128
rect 70000 841004 70074 841060
rect 70130 841004 70200 841060
rect 70000 840936 70200 841004
rect 70000 840880 70074 840936
rect 70130 840880 70200 840936
rect 70000 840812 70200 840880
rect 70000 840756 70074 840812
rect 70130 840756 70200 840812
rect 70000 840688 70200 840756
rect 70000 840632 70074 840688
rect 70130 840632 70200 840688
rect 70000 840564 70200 840632
rect 70000 840508 70074 840564
rect 70130 840508 70200 840564
rect 70000 840440 70200 840508
rect 70000 840384 70074 840440
rect 70130 840384 70200 840440
rect 70000 840316 70200 840384
rect 70000 840260 70074 840316
rect 70130 840260 70200 840316
rect 70000 840192 70200 840260
rect 70000 840136 70074 840192
rect 70130 840136 70200 840192
rect 70000 840068 70200 840136
rect 70000 840012 70074 840068
rect 70130 840012 70200 840068
rect 70000 839944 70200 840012
rect 70000 839888 70074 839944
rect 70130 839888 70200 839944
rect 70000 839820 70200 839888
rect 70000 839764 70074 839820
rect 70130 839764 70200 839820
rect 70000 839696 70200 839764
rect 70000 839640 70074 839696
rect 70130 839640 70200 839696
rect 70000 839572 70200 839640
rect 70000 839516 70074 839572
rect 70130 839516 70200 839572
rect 70000 839448 70200 839516
rect 70000 839392 70074 839448
rect 70130 839392 70200 839448
rect 70000 839324 70200 839392
rect 70000 839268 70074 839324
rect 70130 839268 70200 839324
rect 70000 839198 70200 839268
rect 77678 841190 78678 841878
rect 77678 841134 77808 841190
rect 77864 841134 77932 841190
rect 77988 841134 78056 841190
rect 78112 841134 78180 841190
rect 78236 841134 78304 841190
rect 78360 841134 78428 841190
rect 78484 841134 78552 841190
rect 78608 841134 78678 841190
rect 77678 841066 78678 841134
rect 77678 841010 77808 841066
rect 77864 841010 77932 841066
rect 77988 841010 78056 841066
rect 78112 841010 78180 841066
rect 78236 841010 78304 841066
rect 78360 841010 78428 841066
rect 78484 841010 78552 841066
rect 78608 841010 78678 841066
rect 77678 840942 78678 841010
rect 77678 840886 77808 840942
rect 77864 840886 77932 840942
rect 77988 840886 78056 840942
rect 78112 840886 78180 840942
rect 78236 840886 78304 840942
rect 78360 840886 78428 840942
rect 78484 840886 78552 840942
rect 78608 840886 78678 840942
rect 77678 840818 78678 840886
rect 77678 840762 77808 840818
rect 77864 840762 77932 840818
rect 77988 840762 78056 840818
rect 78112 840762 78180 840818
rect 78236 840762 78304 840818
rect 78360 840762 78428 840818
rect 78484 840762 78552 840818
rect 78608 840762 78678 840818
rect 77678 840694 78678 840762
rect 77678 840638 77808 840694
rect 77864 840638 77932 840694
rect 77988 840638 78056 840694
rect 78112 840638 78180 840694
rect 78236 840638 78304 840694
rect 78360 840638 78428 840694
rect 78484 840638 78552 840694
rect 78608 840638 78678 840694
rect 77678 840570 78678 840638
rect 77678 840514 77808 840570
rect 77864 840514 77932 840570
rect 77988 840514 78056 840570
rect 78112 840514 78180 840570
rect 78236 840514 78304 840570
rect 78360 840514 78428 840570
rect 78484 840514 78552 840570
rect 78608 840514 78678 840570
rect 77678 840446 78678 840514
rect 77678 840390 77808 840446
rect 77864 840390 77932 840446
rect 77988 840390 78056 840446
rect 78112 840390 78180 840446
rect 78236 840390 78304 840446
rect 78360 840390 78428 840446
rect 78484 840390 78552 840446
rect 78608 840390 78678 840446
rect 77678 840322 78678 840390
rect 77678 840266 77808 840322
rect 77864 840266 77932 840322
rect 77988 840266 78056 840322
rect 78112 840266 78180 840322
rect 78236 840266 78304 840322
rect 78360 840266 78428 840322
rect 78484 840266 78552 840322
rect 78608 840266 78678 840322
rect 77678 840198 78678 840266
rect 77678 840142 77808 840198
rect 77864 840142 77932 840198
rect 77988 840142 78056 840198
rect 78112 840142 78180 840198
rect 78236 840142 78304 840198
rect 78360 840142 78428 840198
rect 78484 840142 78552 840198
rect 78608 840142 78678 840198
rect 77678 840074 78678 840142
rect 77678 840018 77808 840074
rect 77864 840018 77932 840074
rect 77988 840018 78056 840074
rect 78112 840018 78180 840074
rect 78236 840018 78304 840074
rect 78360 840018 78428 840074
rect 78484 840018 78552 840074
rect 78608 840018 78678 840074
rect 77678 839950 78678 840018
rect 77678 839894 77808 839950
rect 77864 839894 77932 839950
rect 77988 839894 78056 839950
rect 78112 839894 78180 839950
rect 78236 839894 78304 839950
rect 78360 839894 78428 839950
rect 78484 839894 78552 839950
rect 78608 839894 78678 839950
rect 77678 839826 78678 839894
rect 77678 839770 77808 839826
rect 77864 839770 77932 839826
rect 77988 839770 78056 839826
rect 78112 839770 78180 839826
rect 78236 839770 78304 839826
rect 78360 839770 78428 839826
rect 78484 839770 78552 839826
rect 78608 839770 78678 839826
rect 77678 839702 78678 839770
rect 77678 839646 77808 839702
rect 77864 839646 77932 839702
rect 77988 839646 78056 839702
rect 78112 839646 78180 839702
rect 78236 839646 78304 839702
rect 78360 839646 78428 839702
rect 78484 839646 78552 839702
rect 78608 839646 78678 839702
rect 77678 839578 78678 839646
rect 77678 839522 77808 839578
rect 77864 839522 77932 839578
rect 77988 839522 78056 839578
rect 78112 839522 78180 839578
rect 78236 839522 78304 839578
rect 78360 839522 78428 839578
rect 78484 839522 78552 839578
rect 78608 839522 78678 839578
rect 77678 839454 78678 839522
rect 77678 839398 77808 839454
rect 77864 839398 77932 839454
rect 77988 839398 78056 839454
rect 78112 839398 78180 839454
rect 78236 839398 78304 839454
rect 78360 839398 78428 839454
rect 78484 839398 78552 839454
rect 78608 839398 78678 839454
rect 77678 839330 78678 839398
rect 77678 839274 77808 839330
rect 77864 839274 77932 839330
rect 77988 839274 78056 839330
rect 78112 839274 78180 839330
rect 78236 839274 78304 839330
rect 78360 839274 78428 839330
rect 78484 839274 78552 839330
rect 78608 839274 78678 839330
rect 70000 838814 70200 838878
rect 70000 838758 70074 838814
rect 70130 838758 70200 838814
rect 70000 838690 70200 838758
rect 70000 838634 70074 838690
rect 70130 838634 70200 838690
rect 70000 838566 70200 838634
rect 70000 838510 70074 838566
rect 70130 838510 70200 838566
rect 70000 838442 70200 838510
rect 70000 838386 70074 838442
rect 70130 838386 70200 838442
rect 70000 838318 70200 838386
rect 70000 838262 70074 838318
rect 70130 838262 70200 838318
rect 70000 838194 70200 838262
rect 70000 838138 70074 838194
rect 70130 838138 70200 838194
rect 70000 838070 70200 838138
rect 70000 838014 70074 838070
rect 70130 838014 70200 838070
rect 70000 837946 70200 838014
rect 70000 837890 70074 837946
rect 70130 837890 70200 837946
rect 70000 837822 70200 837890
rect 70000 837766 70074 837822
rect 70130 837766 70200 837822
rect 70000 837698 70200 837766
rect 70000 837642 70074 837698
rect 70130 837642 70200 837698
rect 70000 837574 70200 837642
rect 70000 837518 70074 837574
rect 70130 837518 70200 837574
rect 70000 837450 70200 837518
rect 70000 837394 70074 837450
rect 70130 837394 70200 837450
rect 70000 837326 70200 837394
rect 70000 837270 70074 837326
rect 70130 837270 70200 837326
rect 70000 837202 70200 837270
rect 70000 837146 70074 837202
rect 70130 837146 70200 837202
rect 70000 837078 70200 837146
rect 70000 837022 70074 837078
rect 70130 837022 70200 837078
rect 70000 836954 70200 837022
rect 70000 836898 70074 836954
rect 70130 836898 70200 836954
rect 70000 836828 70200 836898
rect 77678 838820 78678 839274
rect 77678 838764 77808 838820
rect 77864 838764 77932 838820
rect 77988 838764 78056 838820
rect 78112 838764 78180 838820
rect 78236 838764 78304 838820
rect 78360 838764 78428 838820
rect 78484 838764 78552 838820
rect 78608 838764 78678 838820
rect 77678 838696 78678 838764
rect 77678 838640 77808 838696
rect 77864 838640 77932 838696
rect 77988 838640 78056 838696
rect 78112 838640 78180 838696
rect 78236 838640 78304 838696
rect 78360 838640 78428 838696
rect 78484 838640 78552 838696
rect 78608 838640 78678 838696
rect 77678 838572 78678 838640
rect 77678 838516 77808 838572
rect 77864 838516 77932 838572
rect 77988 838516 78056 838572
rect 78112 838516 78180 838572
rect 78236 838516 78304 838572
rect 78360 838516 78428 838572
rect 78484 838516 78552 838572
rect 78608 838516 78678 838572
rect 77678 838448 78678 838516
rect 77678 838392 77808 838448
rect 77864 838392 77932 838448
rect 77988 838392 78056 838448
rect 78112 838392 78180 838448
rect 78236 838392 78304 838448
rect 78360 838392 78428 838448
rect 78484 838392 78552 838448
rect 78608 838392 78678 838448
rect 77678 838324 78678 838392
rect 77678 838268 77808 838324
rect 77864 838268 77932 838324
rect 77988 838268 78056 838324
rect 78112 838268 78180 838324
rect 78236 838268 78304 838324
rect 78360 838268 78428 838324
rect 78484 838268 78552 838324
rect 78608 838268 78678 838324
rect 77678 838200 78678 838268
rect 77678 838144 77808 838200
rect 77864 838144 77932 838200
rect 77988 838144 78056 838200
rect 78112 838144 78180 838200
rect 78236 838144 78304 838200
rect 78360 838144 78428 838200
rect 78484 838144 78552 838200
rect 78608 838144 78678 838200
rect 77678 838076 78678 838144
rect 77678 838020 77808 838076
rect 77864 838020 77932 838076
rect 77988 838020 78056 838076
rect 78112 838020 78180 838076
rect 78236 838020 78304 838076
rect 78360 838020 78428 838076
rect 78484 838020 78552 838076
rect 78608 838020 78678 838076
rect 77678 837952 78678 838020
rect 77678 837896 77808 837952
rect 77864 837896 77932 837952
rect 77988 837896 78056 837952
rect 78112 837896 78180 837952
rect 78236 837896 78304 837952
rect 78360 837896 78428 837952
rect 78484 837896 78552 837952
rect 78608 837896 78678 837952
rect 77678 837828 78678 837896
rect 77678 837772 77808 837828
rect 77864 837772 77932 837828
rect 77988 837772 78056 837828
rect 78112 837772 78180 837828
rect 78236 837772 78304 837828
rect 78360 837772 78428 837828
rect 78484 837772 78552 837828
rect 78608 837772 78678 837828
rect 77678 837704 78678 837772
rect 77678 837648 77808 837704
rect 77864 837648 77932 837704
rect 77988 837648 78056 837704
rect 78112 837648 78180 837704
rect 78236 837648 78304 837704
rect 78360 837648 78428 837704
rect 78484 837648 78552 837704
rect 78608 837648 78678 837704
rect 77678 837580 78678 837648
rect 77678 837524 77808 837580
rect 77864 837524 77932 837580
rect 77988 837524 78056 837580
rect 78112 837524 78180 837580
rect 78236 837524 78304 837580
rect 78360 837524 78428 837580
rect 78484 837524 78552 837580
rect 78608 837524 78678 837580
rect 77678 837456 78678 837524
rect 77678 837400 77808 837456
rect 77864 837400 77932 837456
rect 77988 837400 78056 837456
rect 78112 837400 78180 837456
rect 78236 837400 78304 837456
rect 78360 837400 78428 837456
rect 78484 837400 78552 837456
rect 78608 837400 78678 837456
rect 77678 837332 78678 837400
rect 77678 837276 77808 837332
rect 77864 837276 77932 837332
rect 77988 837276 78056 837332
rect 78112 837276 78180 837332
rect 78236 837276 78304 837332
rect 78360 837276 78428 837332
rect 78484 837276 78552 837332
rect 78608 837276 78678 837332
rect 77678 837208 78678 837276
rect 77678 837152 77808 837208
rect 77864 837152 77932 837208
rect 77988 837152 78056 837208
rect 78112 837152 78180 837208
rect 78236 837152 78304 837208
rect 78360 837152 78428 837208
rect 78484 837152 78552 837208
rect 78608 837152 78678 837208
rect 77678 837084 78678 837152
rect 77678 837028 77808 837084
rect 77864 837028 77932 837084
rect 77988 837028 78056 837084
rect 78112 837028 78180 837084
rect 78236 837028 78304 837084
rect 78360 837028 78428 837084
rect 78484 837028 78552 837084
rect 78608 837028 78678 837084
rect 77678 836960 78678 837028
rect 77678 836904 77808 836960
rect 77864 836904 77932 836960
rect 77988 836904 78056 836960
rect 78112 836904 78180 836960
rect 78236 836904 78304 836960
rect 78360 836904 78428 836960
rect 78484 836904 78552 836960
rect 78608 836904 78678 836960
rect 70000 836108 70200 836172
rect 70000 836052 70074 836108
rect 70130 836052 70200 836108
rect 70000 835984 70200 836052
rect 70000 835928 70074 835984
rect 70130 835928 70200 835984
rect 70000 835860 70200 835928
rect 70000 835804 70074 835860
rect 70130 835804 70200 835860
rect 70000 835736 70200 835804
rect 70000 835680 70074 835736
rect 70130 835680 70200 835736
rect 70000 835612 70200 835680
rect 70000 835556 70074 835612
rect 70130 835556 70200 835612
rect 70000 835488 70200 835556
rect 70000 835432 70074 835488
rect 70130 835432 70200 835488
rect 70000 835364 70200 835432
rect 70000 835308 70074 835364
rect 70130 835308 70200 835364
rect 70000 835240 70200 835308
rect 70000 835184 70074 835240
rect 70130 835184 70200 835240
rect 70000 835116 70200 835184
rect 70000 835060 70074 835116
rect 70130 835060 70200 835116
rect 70000 834992 70200 835060
rect 70000 834936 70074 834992
rect 70130 834936 70200 834992
rect 70000 834868 70200 834936
rect 70000 834812 70074 834868
rect 70130 834812 70200 834868
rect 70000 834744 70200 834812
rect 70000 834688 70074 834744
rect 70130 834688 70200 834744
rect 70000 834620 70200 834688
rect 70000 834564 70074 834620
rect 70130 834564 70200 834620
rect 70000 834496 70200 834564
rect 70000 834440 70074 834496
rect 70130 834440 70200 834496
rect 70000 834372 70200 834440
rect 70000 834316 70074 834372
rect 70130 834316 70200 834372
rect 70000 834248 70200 834316
rect 70000 834192 70074 834248
rect 70130 834192 70200 834248
rect 70000 834122 70200 834192
rect 77678 836114 78678 836904
rect 77678 836058 77808 836114
rect 77864 836058 77932 836114
rect 77988 836058 78056 836114
rect 78112 836058 78180 836114
rect 78236 836058 78304 836114
rect 78360 836058 78428 836114
rect 78484 836058 78552 836114
rect 78608 836058 78678 836114
rect 77678 835990 78678 836058
rect 77678 835934 77808 835990
rect 77864 835934 77932 835990
rect 77988 835934 78056 835990
rect 78112 835934 78180 835990
rect 78236 835934 78304 835990
rect 78360 835934 78428 835990
rect 78484 835934 78552 835990
rect 78608 835934 78678 835990
rect 77678 835866 78678 835934
rect 77678 835810 77808 835866
rect 77864 835810 77932 835866
rect 77988 835810 78056 835866
rect 78112 835810 78180 835866
rect 78236 835810 78304 835866
rect 78360 835810 78428 835866
rect 78484 835810 78552 835866
rect 78608 835810 78678 835866
rect 77678 835742 78678 835810
rect 77678 835686 77808 835742
rect 77864 835686 77932 835742
rect 77988 835686 78056 835742
rect 78112 835686 78180 835742
rect 78236 835686 78304 835742
rect 78360 835686 78428 835742
rect 78484 835686 78552 835742
rect 78608 835686 78678 835742
rect 77678 835618 78678 835686
rect 77678 835562 77808 835618
rect 77864 835562 77932 835618
rect 77988 835562 78056 835618
rect 78112 835562 78180 835618
rect 78236 835562 78304 835618
rect 78360 835562 78428 835618
rect 78484 835562 78552 835618
rect 78608 835562 78678 835618
rect 77678 835494 78678 835562
rect 77678 835438 77808 835494
rect 77864 835438 77932 835494
rect 77988 835438 78056 835494
rect 78112 835438 78180 835494
rect 78236 835438 78304 835494
rect 78360 835438 78428 835494
rect 78484 835438 78552 835494
rect 78608 835438 78678 835494
rect 77678 835370 78678 835438
rect 77678 835314 77808 835370
rect 77864 835314 77932 835370
rect 77988 835314 78056 835370
rect 78112 835314 78180 835370
rect 78236 835314 78304 835370
rect 78360 835314 78428 835370
rect 78484 835314 78552 835370
rect 78608 835314 78678 835370
rect 77678 835246 78678 835314
rect 77678 835190 77808 835246
rect 77864 835190 77932 835246
rect 77988 835190 78056 835246
rect 78112 835190 78180 835246
rect 78236 835190 78304 835246
rect 78360 835190 78428 835246
rect 78484 835190 78552 835246
rect 78608 835190 78678 835246
rect 77678 835122 78678 835190
rect 77678 835066 77808 835122
rect 77864 835066 77932 835122
rect 77988 835066 78056 835122
rect 78112 835066 78180 835122
rect 78236 835066 78304 835122
rect 78360 835066 78428 835122
rect 78484 835066 78552 835122
rect 78608 835066 78678 835122
rect 77678 834998 78678 835066
rect 77678 834942 77808 834998
rect 77864 834942 77932 834998
rect 77988 834942 78056 834998
rect 78112 834942 78180 834998
rect 78236 834942 78304 834998
rect 78360 834942 78428 834998
rect 78484 834942 78552 834998
rect 78608 834942 78678 834998
rect 77678 834874 78678 834942
rect 77678 834818 77808 834874
rect 77864 834818 77932 834874
rect 77988 834818 78056 834874
rect 78112 834818 78180 834874
rect 78236 834818 78304 834874
rect 78360 834818 78428 834874
rect 78484 834818 78552 834874
rect 78608 834818 78678 834874
rect 77678 834750 78678 834818
rect 77678 834694 77808 834750
rect 77864 834694 77932 834750
rect 77988 834694 78056 834750
rect 78112 834694 78180 834750
rect 78236 834694 78304 834750
rect 78360 834694 78428 834750
rect 78484 834694 78552 834750
rect 78608 834694 78678 834750
rect 77678 834626 78678 834694
rect 77678 834570 77808 834626
rect 77864 834570 77932 834626
rect 77988 834570 78056 834626
rect 78112 834570 78180 834626
rect 78236 834570 78304 834626
rect 78360 834570 78428 834626
rect 78484 834570 78552 834626
rect 78608 834570 78678 834626
rect 77678 834502 78678 834570
rect 77678 834446 77808 834502
rect 77864 834446 77932 834502
rect 77988 834446 78056 834502
rect 78112 834446 78180 834502
rect 78236 834446 78304 834502
rect 78360 834446 78428 834502
rect 78484 834446 78552 834502
rect 78608 834446 78678 834502
rect 77678 834378 78678 834446
rect 77678 834322 77808 834378
rect 77864 834322 77932 834378
rect 77988 834322 78056 834378
rect 78112 834322 78180 834378
rect 78236 834322 78304 834378
rect 78360 834322 78428 834378
rect 78484 834322 78552 834378
rect 78608 834322 78678 834378
rect 77678 834254 78678 834322
rect 77678 834198 77808 834254
rect 77864 834198 77932 834254
rect 77988 834198 78056 834254
rect 78112 834198 78180 834254
rect 78236 834198 78304 834254
rect 78360 834198 78428 834254
rect 78484 834198 78552 834254
rect 78608 834198 78678 834254
rect 70000 833738 70200 833802
rect 70000 833682 70074 833738
rect 70130 833682 70200 833738
rect 70000 833614 70200 833682
rect 70000 833558 70074 833614
rect 70130 833558 70200 833614
rect 70000 833490 70200 833558
rect 70000 833434 70074 833490
rect 70130 833434 70200 833490
rect 70000 833366 70200 833434
rect 70000 833310 70074 833366
rect 70130 833310 70200 833366
rect 70000 833242 70200 833310
rect 70000 833186 70074 833242
rect 70130 833186 70200 833242
rect 70000 833118 70200 833186
rect 70000 833062 70074 833118
rect 70130 833062 70200 833118
rect 70000 832994 70200 833062
rect 70000 832938 70074 832994
rect 70130 832938 70200 832994
rect 70000 832870 70200 832938
rect 70000 832814 70074 832870
rect 70130 832814 70200 832870
rect 70000 832746 70200 832814
rect 70000 832690 70074 832746
rect 70130 832690 70200 832746
rect 70000 832622 70200 832690
rect 70000 832566 70074 832622
rect 70130 832566 70200 832622
rect 70000 832498 70200 832566
rect 70000 832442 70074 832498
rect 70130 832442 70200 832498
rect 70000 832374 70200 832442
rect 70000 832318 70074 832374
rect 70130 832318 70200 832374
rect 70000 832250 70200 832318
rect 70000 832194 70074 832250
rect 70130 832194 70200 832250
rect 70000 832126 70200 832194
rect 70000 832070 70074 832126
rect 70130 832070 70200 832126
rect 70000 832002 70200 832070
rect 70000 831946 70074 832002
rect 70130 831946 70200 832002
rect 70000 831878 70200 831946
rect 70000 831822 70074 831878
rect 70130 831822 70200 831878
rect 70000 831752 70200 831822
rect 77678 833744 78678 834198
rect 77678 833688 77808 833744
rect 77864 833688 77932 833744
rect 77988 833688 78056 833744
rect 78112 833688 78180 833744
rect 78236 833688 78304 833744
rect 78360 833688 78428 833744
rect 78484 833688 78552 833744
rect 78608 833688 78678 833744
rect 77678 833620 78678 833688
rect 77678 833564 77808 833620
rect 77864 833564 77932 833620
rect 77988 833564 78056 833620
rect 78112 833564 78180 833620
rect 78236 833564 78304 833620
rect 78360 833564 78428 833620
rect 78484 833564 78552 833620
rect 78608 833564 78678 833620
rect 77678 833496 78678 833564
rect 77678 833440 77808 833496
rect 77864 833440 77932 833496
rect 77988 833440 78056 833496
rect 78112 833440 78180 833496
rect 78236 833440 78304 833496
rect 78360 833440 78428 833496
rect 78484 833440 78552 833496
rect 78608 833440 78678 833496
rect 77678 833372 78678 833440
rect 77678 833316 77808 833372
rect 77864 833316 77932 833372
rect 77988 833316 78056 833372
rect 78112 833316 78180 833372
rect 78236 833316 78304 833372
rect 78360 833316 78428 833372
rect 78484 833316 78552 833372
rect 78608 833316 78678 833372
rect 77678 833248 78678 833316
rect 77678 833192 77808 833248
rect 77864 833192 77932 833248
rect 77988 833192 78056 833248
rect 78112 833192 78180 833248
rect 78236 833192 78304 833248
rect 78360 833192 78428 833248
rect 78484 833192 78552 833248
rect 78608 833192 78678 833248
rect 77678 833124 78678 833192
rect 77678 833068 77808 833124
rect 77864 833068 77932 833124
rect 77988 833068 78056 833124
rect 78112 833068 78180 833124
rect 78236 833068 78304 833124
rect 78360 833068 78428 833124
rect 78484 833068 78552 833124
rect 78608 833068 78678 833124
rect 77678 833000 78678 833068
rect 77678 832944 77808 833000
rect 77864 832944 77932 833000
rect 77988 832944 78056 833000
rect 78112 832944 78180 833000
rect 78236 832944 78304 833000
rect 78360 832944 78428 833000
rect 78484 832944 78552 833000
rect 78608 832944 78678 833000
rect 77678 832876 78678 832944
rect 77678 832820 77808 832876
rect 77864 832820 77932 832876
rect 77988 832820 78056 832876
rect 78112 832820 78180 832876
rect 78236 832820 78304 832876
rect 78360 832820 78428 832876
rect 78484 832820 78552 832876
rect 78608 832820 78678 832876
rect 77678 832752 78678 832820
rect 77678 832696 77808 832752
rect 77864 832696 77932 832752
rect 77988 832696 78056 832752
rect 78112 832696 78180 832752
rect 78236 832696 78304 832752
rect 78360 832696 78428 832752
rect 78484 832696 78552 832752
rect 78608 832696 78678 832752
rect 77678 832628 78678 832696
rect 77678 832572 77808 832628
rect 77864 832572 77932 832628
rect 77988 832572 78056 832628
rect 78112 832572 78180 832628
rect 78236 832572 78304 832628
rect 78360 832572 78428 832628
rect 78484 832572 78552 832628
rect 78608 832572 78678 832628
rect 77678 832504 78678 832572
rect 77678 832448 77808 832504
rect 77864 832448 77932 832504
rect 77988 832448 78056 832504
rect 78112 832448 78180 832504
rect 78236 832448 78304 832504
rect 78360 832448 78428 832504
rect 78484 832448 78552 832504
rect 78608 832448 78678 832504
rect 77678 832380 78678 832448
rect 77678 832324 77808 832380
rect 77864 832324 77932 832380
rect 77988 832324 78056 832380
rect 78112 832324 78180 832380
rect 78236 832324 78304 832380
rect 78360 832324 78428 832380
rect 78484 832324 78552 832380
rect 78608 832324 78678 832380
rect 77678 832256 78678 832324
rect 77678 832200 77808 832256
rect 77864 832200 77932 832256
rect 77988 832200 78056 832256
rect 78112 832200 78180 832256
rect 78236 832200 78304 832256
rect 78360 832200 78428 832256
rect 78484 832200 78552 832256
rect 78608 832200 78678 832256
rect 77678 832132 78678 832200
rect 77678 832076 77808 832132
rect 77864 832076 77932 832132
rect 77988 832076 78056 832132
rect 78112 832076 78180 832132
rect 78236 832076 78304 832132
rect 78360 832076 78428 832132
rect 78484 832076 78552 832132
rect 78608 832076 78678 832132
rect 77678 832008 78678 832076
rect 77678 831952 77808 832008
rect 77864 831952 77932 832008
rect 77988 831952 78056 832008
rect 78112 831952 78180 832008
rect 78236 831952 78304 832008
rect 78360 831952 78428 832008
rect 78484 831952 78552 832008
rect 78608 831952 78678 832008
rect 77678 831884 78678 831952
rect 77678 831828 77808 831884
rect 77864 831828 77932 831884
rect 77988 831828 78056 831884
rect 78112 831828 78180 831884
rect 78236 831828 78304 831884
rect 78360 831828 78428 831884
rect 78484 831828 78552 831884
rect 78608 831828 78678 831884
rect 70000 831134 70200 831172
rect 70000 831078 70074 831134
rect 70130 831078 70200 831134
rect 70000 831010 70200 831078
rect 70000 830954 70074 831010
rect 70130 830954 70200 831010
rect 70000 830886 70200 830954
rect 70000 830830 70074 830886
rect 70130 830830 70200 830886
rect 70000 830762 70200 830830
rect 70000 830706 70074 830762
rect 70130 830706 70200 830762
rect 70000 830638 70200 830706
rect 70000 830582 70074 830638
rect 70130 830582 70200 830638
rect 70000 830514 70200 830582
rect 70000 830458 70074 830514
rect 70130 830458 70200 830514
rect 70000 830390 70200 830458
rect 70000 830334 70074 830390
rect 70130 830334 70200 830390
rect 70000 830266 70200 830334
rect 70000 830210 70074 830266
rect 70130 830210 70200 830266
rect 70000 830142 70200 830210
rect 70000 830086 70074 830142
rect 70130 830086 70200 830142
rect 70000 830018 70200 830086
rect 70000 829962 70074 830018
rect 70130 829962 70200 830018
rect 70000 829894 70200 829962
rect 70000 829838 70074 829894
rect 70130 829838 70200 829894
rect 70000 829770 70200 829838
rect 70000 829714 70074 829770
rect 70130 829714 70200 829770
rect 70000 829646 70200 829714
rect 70000 829590 70074 829646
rect 70130 829590 70200 829646
rect 70000 829522 70200 829590
rect 70000 829466 70074 829522
rect 70130 829466 70200 829522
rect 70000 829398 70200 829466
rect 70000 829342 70074 829398
rect 70130 829342 70200 829398
rect 70000 829272 70200 829342
rect 77678 831140 78678 831828
rect 77678 831084 77808 831140
rect 77864 831084 77932 831140
rect 77988 831084 78056 831140
rect 78112 831084 78180 831140
rect 78236 831084 78304 831140
rect 78360 831084 78428 831140
rect 78484 831084 78552 831140
rect 78608 831084 78678 831140
rect 77678 831016 78678 831084
rect 77678 830960 77808 831016
rect 77864 830960 77932 831016
rect 77988 830960 78056 831016
rect 78112 830960 78180 831016
rect 78236 830960 78304 831016
rect 78360 830960 78428 831016
rect 78484 830960 78552 831016
rect 78608 830960 78678 831016
rect 77678 830892 78678 830960
rect 77678 830836 77808 830892
rect 77864 830836 77932 830892
rect 77988 830836 78056 830892
rect 78112 830836 78180 830892
rect 78236 830836 78304 830892
rect 78360 830836 78428 830892
rect 78484 830836 78552 830892
rect 78608 830836 78678 830892
rect 77678 830768 78678 830836
rect 77678 830712 77808 830768
rect 77864 830712 77932 830768
rect 77988 830712 78056 830768
rect 78112 830712 78180 830768
rect 78236 830712 78304 830768
rect 78360 830712 78428 830768
rect 78484 830712 78552 830768
rect 78608 830712 78678 830768
rect 77678 830644 78678 830712
rect 77678 830588 77808 830644
rect 77864 830588 77932 830644
rect 77988 830588 78056 830644
rect 78112 830588 78180 830644
rect 78236 830588 78304 830644
rect 78360 830588 78428 830644
rect 78484 830588 78552 830644
rect 78608 830588 78678 830644
rect 77678 830520 78678 830588
rect 77678 830464 77808 830520
rect 77864 830464 77932 830520
rect 77988 830464 78056 830520
rect 78112 830464 78180 830520
rect 78236 830464 78304 830520
rect 78360 830464 78428 830520
rect 78484 830464 78552 830520
rect 78608 830464 78678 830520
rect 77678 830396 78678 830464
rect 77678 830340 77808 830396
rect 77864 830340 77932 830396
rect 77988 830340 78056 830396
rect 78112 830340 78180 830396
rect 78236 830340 78304 830396
rect 78360 830340 78428 830396
rect 78484 830340 78552 830396
rect 78608 830340 78678 830396
rect 77678 830272 78678 830340
rect 77678 830216 77808 830272
rect 77864 830216 77932 830272
rect 77988 830216 78056 830272
rect 78112 830216 78180 830272
rect 78236 830216 78304 830272
rect 78360 830216 78428 830272
rect 78484 830216 78552 830272
rect 78608 830216 78678 830272
rect 77678 830148 78678 830216
rect 77678 830092 77808 830148
rect 77864 830092 77932 830148
rect 77988 830092 78056 830148
rect 78112 830092 78180 830148
rect 78236 830092 78304 830148
rect 78360 830092 78428 830148
rect 78484 830092 78552 830148
rect 78608 830092 78678 830148
rect 77678 830024 78678 830092
rect 77678 829968 77808 830024
rect 77864 829968 77932 830024
rect 77988 829968 78056 830024
rect 78112 829968 78180 830024
rect 78236 829968 78304 830024
rect 78360 829968 78428 830024
rect 78484 829968 78552 830024
rect 78608 829968 78678 830024
rect 77678 829900 78678 829968
rect 77678 829844 77808 829900
rect 77864 829844 77932 829900
rect 77988 829844 78056 829900
rect 78112 829844 78180 829900
rect 78236 829844 78304 829900
rect 78360 829844 78428 829900
rect 78484 829844 78552 829900
rect 78608 829844 78678 829900
rect 77678 829776 78678 829844
rect 77678 829720 77808 829776
rect 77864 829720 77932 829776
rect 77988 829720 78056 829776
rect 78112 829720 78180 829776
rect 78236 829720 78304 829776
rect 78360 829720 78428 829776
rect 78484 829720 78552 829776
rect 78608 829720 78678 829776
rect 77678 829652 78678 829720
rect 77678 829596 77808 829652
rect 77864 829596 77932 829652
rect 77988 829596 78056 829652
rect 78112 829596 78180 829652
rect 78236 829596 78304 829652
rect 78360 829596 78428 829652
rect 78484 829596 78552 829652
rect 78608 829596 78678 829652
rect 77678 829528 78678 829596
rect 77678 829472 77808 829528
rect 77864 829472 77932 829528
rect 77988 829472 78056 829528
rect 78112 829472 78180 829528
rect 78236 829472 78304 829528
rect 78360 829472 78428 829528
rect 78484 829472 78552 829528
rect 78608 829472 78678 829528
rect 77678 829404 78678 829472
rect 77678 829348 77808 829404
rect 77864 829348 77932 829404
rect 77988 829348 78056 829404
rect 78112 829348 78180 829404
rect 78236 829348 78304 829404
rect 78360 829348 78428 829404
rect 78484 829348 78552 829404
rect 78608 829348 78678 829404
rect 77678 806429 78678 829348
rect 77678 806373 77800 806429
rect 77856 806373 78100 806429
rect 78156 806373 78400 806429
rect 78456 806373 78678 806429
rect 77678 806229 78678 806373
rect 77678 806173 77800 806229
rect 77856 806173 78100 806229
rect 78156 806173 78400 806229
rect 78456 806173 78678 806229
rect 70000 802658 70200 802728
rect 70000 802602 70074 802658
rect 70130 802602 70200 802658
rect 70000 802534 70200 802602
rect 70000 802478 70074 802534
rect 70130 802478 70200 802534
rect 70000 802410 70200 802478
rect 70000 802354 70074 802410
rect 70130 802354 70200 802410
rect 70000 802286 70200 802354
rect 70000 802230 70074 802286
rect 70130 802230 70200 802286
rect 70000 802162 70200 802230
rect 70000 802106 70074 802162
rect 70130 802106 70200 802162
rect 70000 802038 70200 802106
rect 70000 801982 70074 802038
rect 70130 801982 70200 802038
rect 70000 801914 70200 801982
rect 70000 801858 70074 801914
rect 70130 801858 70200 801914
rect 70000 801790 70200 801858
rect 70000 801734 70074 801790
rect 70130 801734 70200 801790
rect 70000 801666 70200 801734
rect 70000 801610 70074 801666
rect 70130 801610 70200 801666
rect 70000 801542 70200 801610
rect 70000 801486 70074 801542
rect 70130 801486 70200 801542
rect 70000 801418 70200 801486
rect 70000 801362 70074 801418
rect 70130 801362 70200 801418
rect 70000 801294 70200 801362
rect 70000 801238 70074 801294
rect 70130 801238 70200 801294
rect 70000 801170 70200 801238
rect 70000 801114 70074 801170
rect 70130 801114 70200 801170
rect 70000 801046 70200 801114
rect 70000 800990 70074 801046
rect 70130 800990 70200 801046
rect 70000 800922 70200 800990
rect 70000 800866 70074 800922
rect 70130 800866 70200 800922
rect 70000 800828 70200 800866
rect 70000 800184 70200 800248
rect 70000 800128 70074 800184
rect 70130 800128 70200 800184
rect 70000 800060 70200 800128
rect 70000 800004 70074 800060
rect 70130 800004 70200 800060
rect 70000 799936 70200 800004
rect 70000 799880 70074 799936
rect 70130 799880 70200 799936
rect 70000 799812 70200 799880
rect 70000 799756 70074 799812
rect 70130 799756 70200 799812
rect 70000 799688 70200 799756
rect 70000 799632 70074 799688
rect 70130 799632 70200 799688
rect 70000 799564 70200 799632
rect 70000 799508 70074 799564
rect 70130 799508 70200 799564
rect 70000 799440 70200 799508
rect 70000 799384 70074 799440
rect 70130 799384 70200 799440
rect 70000 799316 70200 799384
rect 70000 799260 70074 799316
rect 70130 799260 70200 799316
rect 70000 799192 70200 799260
rect 70000 799136 70074 799192
rect 70130 799136 70200 799192
rect 70000 799068 70200 799136
rect 70000 799012 70074 799068
rect 70130 799012 70200 799068
rect 70000 798944 70200 799012
rect 70000 798888 70074 798944
rect 70130 798888 70200 798944
rect 70000 798820 70200 798888
rect 70000 798764 70074 798820
rect 70130 798764 70200 798820
rect 70000 798696 70200 798764
rect 70000 798640 70074 798696
rect 70130 798640 70200 798696
rect 70000 798572 70200 798640
rect 70000 798516 70074 798572
rect 70130 798516 70200 798572
rect 70000 798448 70200 798516
rect 70000 798392 70074 798448
rect 70130 798392 70200 798448
rect 70000 798324 70200 798392
rect 70000 798268 70074 798324
rect 70130 798268 70200 798324
rect 70000 798198 70200 798268
rect 70000 797814 70200 797878
rect 70000 797758 70074 797814
rect 70130 797758 70200 797814
rect 70000 797690 70200 797758
rect 70000 797634 70074 797690
rect 70130 797634 70200 797690
rect 70000 797566 70200 797634
rect 70000 797510 70074 797566
rect 70130 797510 70200 797566
rect 70000 797442 70200 797510
rect 70000 797386 70074 797442
rect 70130 797386 70200 797442
rect 70000 797318 70200 797386
rect 70000 797262 70074 797318
rect 70130 797262 70200 797318
rect 70000 797194 70200 797262
rect 70000 797138 70074 797194
rect 70130 797138 70200 797194
rect 70000 797070 70200 797138
rect 70000 797014 70074 797070
rect 70130 797014 70200 797070
rect 70000 796946 70200 797014
rect 70000 796890 70074 796946
rect 70130 796890 70200 796946
rect 70000 796822 70200 796890
rect 70000 796766 70074 796822
rect 70130 796766 70200 796822
rect 70000 796698 70200 796766
rect 70000 796642 70074 796698
rect 70130 796642 70200 796698
rect 70000 796574 70200 796642
rect 70000 796518 70074 796574
rect 70130 796518 70200 796574
rect 70000 796450 70200 796518
rect 70000 796394 70074 796450
rect 70130 796394 70200 796450
rect 70000 796326 70200 796394
rect 70000 796270 70074 796326
rect 70130 796270 70200 796326
rect 70000 796202 70200 796270
rect 70000 796146 70074 796202
rect 70130 796146 70200 796202
rect 70000 796078 70200 796146
rect 70000 796022 70074 796078
rect 70130 796022 70200 796078
rect 70000 795954 70200 796022
rect 70000 795898 70074 795954
rect 70130 795898 70200 795954
rect 70000 795828 70200 795898
rect 70000 795108 70200 795172
rect 70000 795052 70074 795108
rect 70130 795052 70200 795108
rect 70000 794984 70200 795052
rect 70000 794928 70074 794984
rect 70130 794928 70200 794984
rect 70000 794860 70200 794928
rect 70000 794804 70074 794860
rect 70130 794804 70200 794860
rect 70000 794736 70200 794804
rect 70000 794680 70074 794736
rect 70130 794680 70200 794736
rect 70000 794612 70200 794680
rect 70000 794556 70074 794612
rect 70130 794556 70200 794612
rect 70000 794488 70200 794556
rect 70000 794432 70074 794488
rect 70130 794432 70200 794488
rect 70000 794364 70200 794432
rect 70000 794308 70074 794364
rect 70130 794308 70200 794364
rect 70000 794240 70200 794308
rect 70000 794184 70074 794240
rect 70130 794184 70200 794240
rect 70000 794116 70200 794184
rect 70000 794060 70074 794116
rect 70130 794060 70200 794116
rect 70000 793992 70200 794060
rect 70000 793936 70074 793992
rect 70130 793936 70200 793992
rect 70000 793868 70200 793936
rect 70000 793812 70074 793868
rect 70130 793812 70200 793868
rect 70000 793744 70200 793812
rect 70000 793688 70074 793744
rect 70130 793688 70200 793744
rect 70000 793620 70200 793688
rect 70000 793564 70074 793620
rect 70130 793564 70200 793620
rect 70000 793496 70200 793564
rect 70000 793440 70074 793496
rect 70130 793440 70200 793496
rect 70000 793372 70200 793440
rect 70000 793316 70074 793372
rect 70130 793316 70200 793372
rect 70000 793248 70200 793316
rect 70000 793192 70074 793248
rect 70130 793192 70200 793248
rect 70000 793122 70200 793192
rect 70000 792738 70200 792802
rect 70000 792682 70074 792738
rect 70130 792682 70200 792738
rect 70000 792614 70200 792682
rect 70000 792558 70074 792614
rect 70130 792558 70200 792614
rect 70000 792490 70200 792558
rect 70000 792434 70074 792490
rect 70130 792434 70200 792490
rect 70000 792366 70200 792434
rect 70000 792310 70074 792366
rect 70130 792310 70200 792366
rect 70000 792242 70200 792310
rect 70000 792186 70074 792242
rect 70130 792186 70200 792242
rect 70000 792118 70200 792186
rect 70000 792062 70074 792118
rect 70130 792062 70200 792118
rect 70000 791994 70200 792062
rect 70000 791938 70074 791994
rect 70130 791938 70200 791994
rect 70000 791870 70200 791938
rect 70000 791814 70074 791870
rect 70130 791814 70200 791870
rect 70000 791746 70200 791814
rect 70000 791690 70074 791746
rect 70130 791690 70200 791746
rect 70000 791622 70200 791690
rect 70000 791566 70074 791622
rect 70130 791566 70200 791622
rect 70000 791498 70200 791566
rect 70000 791442 70074 791498
rect 70130 791442 70200 791498
rect 70000 791374 70200 791442
rect 70000 791318 70074 791374
rect 70130 791318 70200 791374
rect 70000 791250 70200 791318
rect 70000 791194 70074 791250
rect 70130 791194 70200 791250
rect 70000 791126 70200 791194
rect 70000 791070 70074 791126
rect 70130 791070 70200 791126
rect 70000 791002 70200 791070
rect 70000 790946 70074 791002
rect 70130 790946 70200 791002
rect 70000 790878 70200 790946
rect 70000 790822 70074 790878
rect 70130 790822 70200 790878
rect 70000 790752 70200 790822
rect 70000 790134 70200 790172
rect 70000 790078 70074 790134
rect 70130 790078 70200 790134
rect 70000 790010 70200 790078
rect 70000 789954 70074 790010
rect 70130 789954 70200 790010
rect 70000 789886 70200 789954
rect 70000 789830 70074 789886
rect 70130 789830 70200 789886
rect 70000 789762 70200 789830
rect 70000 789706 70074 789762
rect 70130 789706 70200 789762
rect 70000 789638 70200 789706
rect 70000 789582 70074 789638
rect 70130 789582 70200 789638
rect 70000 789514 70200 789582
rect 70000 789458 70074 789514
rect 70130 789458 70200 789514
rect 70000 789390 70200 789458
rect 70000 789334 70074 789390
rect 70130 789334 70200 789390
rect 70000 789266 70200 789334
rect 70000 789210 70074 789266
rect 70130 789210 70200 789266
rect 70000 789142 70200 789210
rect 70000 789086 70074 789142
rect 70130 789086 70200 789142
rect 70000 789018 70200 789086
rect 70000 788962 70074 789018
rect 70130 788962 70200 789018
rect 70000 788894 70200 788962
rect 70000 788838 70074 788894
rect 70130 788838 70200 788894
rect 70000 788770 70200 788838
rect 70000 788714 70074 788770
rect 70130 788714 70200 788770
rect 70000 788646 70200 788714
rect 70000 788590 70074 788646
rect 70130 788590 70200 788646
rect 70000 788522 70200 788590
rect 70000 788466 70074 788522
rect 70130 788466 70200 788522
rect 70000 788398 70200 788466
rect 70000 788342 70074 788398
rect 70130 788342 70200 788398
rect 70000 788272 70200 788342
rect 77678 781633 78678 806173
rect 77678 781577 77847 781633
rect 77903 781577 78147 781633
rect 78203 781577 78447 781633
rect 78503 781577 78678 781633
rect 77678 770429 78678 781577
rect 77678 770373 77800 770429
rect 77856 770373 78100 770429
rect 78156 770373 78400 770429
rect 78456 770373 78678 770429
rect 77678 770229 78678 770373
rect 77678 770173 77800 770229
rect 77856 770173 78100 770229
rect 78156 770173 78400 770229
rect 78456 770173 78678 770229
rect 77678 762102 78678 770173
rect 77678 762046 77900 762102
rect 77956 762046 78200 762102
rect 78256 762046 78500 762102
rect 78556 762046 78678 762102
rect 77678 755102 78678 762046
rect 77678 755046 77900 755102
rect 77956 755046 78200 755102
rect 78256 755046 78500 755102
rect 78556 755046 78678 755102
rect 77678 748102 78678 755046
rect 77678 748046 77900 748102
rect 77956 748046 78200 748102
rect 78256 748046 78500 748102
rect 78556 748046 78678 748102
rect 77678 740633 78678 748046
rect 77678 740577 77847 740633
rect 77903 740577 78147 740633
rect 78203 740577 78447 740633
rect 78503 740577 78678 740633
rect 77678 734429 78678 740577
rect 77678 734373 77800 734429
rect 77856 734373 78100 734429
rect 78156 734373 78400 734429
rect 78456 734373 78678 734429
rect 77678 734229 78678 734373
rect 77678 734173 77800 734229
rect 77856 734173 78100 734229
rect 78156 734173 78400 734229
rect 78456 734173 78678 734229
rect 77678 721102 78678 734173
rect 77678 721046 77900 721102
rect 77956 721046 78200 721102
rect 78256 721046 78500 721102
rect 78556 721046 78678 721102
rect 77678 714102 78678 721046
rect 77678 714046 77900 714102
rect 77956 714046 78200 714102
rect 78256 714046 78500 714102
rect 78556 714046 78678 714102
rect 77678 707102 78678 714046
rect 77678 707046 77900 707102
rect 77956 707046 78200 707102
rect 78256 707046 78500 707102
rect 78556 707046 78678 707102
rect 77678 699633 78678 707046
rect 77678 699577 77847 699633
rect 77903 699577 78147 699633
rect 78203 699577 78447 699633
rect 78503 699577 78678 699633
rect 77678 698429 78678 699577
rect 77678 698373 77800 698429
rect 77856 698373 78100 698429
rect 78156 698373 78400 698429
rect 78456 698373 78678 698429
rect 77678 698229 78678 698373
rect 77678 698173 77800 698229
rect 77856 698173 78100 698229
rect 78156 698173 78400 698229
rect 78456 698173 78678 698229
rect 77678 680102 78678 698173
rect 77678 680046 77900 680102
rect 77956 680046 78200 680102
rect 78256 680046 78500 680102
rect 78556 680046 78678 680102
rect 77678 673102 78678 680046
rect 77678 673046 77900 673102
rect 77956 673046 78200 673102
rect 78256 673046 78500 673102
rect 78556 673046 78678 673102
rect 77678 666102 78678 673046
rect 77678 666046 77900 666102
rect 77956 666046 78200 666102
rect 78256 666046 78500 666102
rect 78556 666046 78678 666102
rect 77678 662429 78678 666046
rect 77678 662373 77800 662429
rect 77856 662373 78100 662429
rect 78156 662373 78400 662429
rect 78456 662373 78678 662429
rect 77678 662229 78678 662373
rect 77678 662173 77800 662229
rect 77856 662173 78100 662229
rect 78156 662173 78400 662229
rect 78456 662173 78678 662229
rect 77678 658633 78678 662173
rect 77678 658577 77847 658633
rect 77903 658577 78147 658633
rect 78203 658577 78447 658633
rect 78503 658577 78678 658633
rect 77678 639102 78678 658577
rect 77678 639046 77900 639102
rect 77956 639046 78200 639102
rect 78256 639046 78500 639102
rect 78556 639046 78678 639102
rect 77678 632102 78678 639046
rect 77678 632046 77900 632102
rect 77956 632046 78200 632102
rect 78256 632046 78500 632102
rect 78556 632046 78678 632102
rect 77678 626429 78678 632046
rect 77678 626373 77800 626429
rect 77856 626373 78100 626429
rect 78156 626373 78400 626429
rect 78456 626373 78678 626429
rect 77678 626229 78678 626373
rect 77678 626173 77800 626229
rect 77856 626173 78100 626229
rect 78156 626173 78400 626229
rect 78456 626173 78678 626229
rect 77678 625102 78678 626173
rect 77678 625046 77900 625102
rect 77956 625046 78200 625102
rect 78256 625046 78500 625102
rect 78556 625046 78678 625102
rect 77678 617633 78678 625046
rect 77678 617577 77847 617633
rect 77903 617577 78147 617633
rect 78203 617577 78447 617633
rect 78503 617577 78678 617633
rect 77678 598102 78678 617577
rect 77678 598046 77900 598102
rect 77956 598046 78200 598102
rect 78256 598046 78500 598102
rect 78556 598046 78678 598102
rect 77678 591102 78678 598046
rect 77678 591046 77900 591102
rect 77956 591046 78200 591102
rect 78256 591046 78500 591102
rect 78556 591046 78678 591102
rect 77678 590429 78678 591046
rect 77678 590373 77800 590429
rect 77856 590373 78100 590429
rect 78156 590373 78400 590429
rect 78456 590373 78678 590429
rect 77678 590229 78678 590373
rect 77678 590173 77800 590229
rect 77856 590173 78100 590229
rect 78156 590173 78400 590229
rect 78456 590173 78678 590229
rect 77678 584102 78678 590173
rect 77678 584046 77900 584102
rect 77956 584046 78200 584102
rect 78256 584046 78500 584102
rect 78556 584046 78678 584102
rect 77678 576633 78678 584046
rect 77678 576577 77847 576633
rect 77903 576577 78147 576633
rect 78203 576577 78447 576633
rect 78503 576577 78678 576633
rect 77678 557102 78678 576577
rect 77678 557046 77900 557102
rect 77956 557046 78200 557102
rect 78256 557046 78500 557102
rect 78556 557046 78678 557102
rect 77678 554429 78678 557046
rect 77678 554373 77800 554429
rect 77856 554373 78100 554429
rect 78156 554373 78400 554429
rect 78456 554373 78678 554429
rect 77678 554229 78678 554373
rect 77678 554173 77800 554229
rect 77856 554173 78100 554229
rect 78156 554173 78400 554229
rect 78456 554173 78678 554229
rect 77678 550102 78678 554173
rect 77678 550046 77900 550102
rect 77956 550046 78200 550102
rect 78256 550046 78500 550102
rect 78556 550046 78678 550102
rect 77678 543102 78678 550046
rect 77678 543046 77900 543102
rect 77956 543046 78200 543102
rect 78256 543046 78500 543102
rect 78556 543046 78678 543102
rect 77678 535633 78678 543046
rect 77678 535577 77847 535633
rect 77903 535577 78147 535633
rect 78203 535577 78447 535633
rect 78503 535577 78678 535633
rect 77678 518429 78678 535577
rect 77678 518373 77800 518429
rect 77856 518373 78100 518429
rect 78156 518373 78400 518429
rect 78456 518373 78678 518429
rect 77678 518229 78678 518373
rect 77678 518173 77800 518229
rect 77856 518173 78100 518229
rect 78156 518173 78400 518229
rect 78456 518173 78678 518229
rect 77678 516102 78678 518173
rect 77678 516046 77900 516102
rect 77956 516046 78200 516102
rect 78256 516046 78500 516102
rect 78556 516046 78678 516102
rect 77678 509102 78678 516046
rect 77678 509046 77900 509102
rect 77956 509046 78200 509102
rect 78256 509046 78500 509102
rect 78556 509046 78678 509102
rect 77678 502102 78678 509046
rect 77678 502046 77900 502102
rect 77956 502046 78200 502102
rect 78256 502046 78500 502102
rect 78556 502046 78678 502102
rect 77678 482429 78678 502046
rect 77678 482373 77800 482429
rect 77856 482373 78100 482429
rect 78156 482373 78400 482429
rect 78456 482373 78678 482429
rect 77678 482229 78678 482373
rect 77678 482173 77800 482229
rect 77856 482173 78100 482229
rect 78156 482173 78400 482229
rect 78456 482173 78678 482229
rect 70000 474658 70200 474728
rect 70000 474602 70074 474658
rect 70130 474602 70200 474658
rect 70000 474534 70200 474602
rect 70000 474478 70074 474534
rect 70130 474478 70200 474534
rect 70000 474410 70200 474478
rect 70000 474354 70074 474410
rect 70130 474354 70200 474410
rect 70000 474286 70200 474354
rect 70000 474230 70074 474286
rect 70130 474230 70200 474286
rect 70000 474162 70200 474230
rect 70000 474106 70074 474162
rect 70130 474106 70200 474162
rect 70000 474038 70200 474106
rect 70000 473982 70074 474038
rect 70130 473982 70200 474038
rect 70000 473914 70200 473982
rect 70000 473858 70074 473914
rect 70130 473858 70200 473914
rect 70000 473790 70200 473858
rect 70000 473734 70074 473790
rect 70130 473734 70200 473790
rect 70000 473666 70200 473734
rect 70000 473610 70074 473666
rect 70130 473610 70200 473666
rect 70000 473542 70200 473610
rect 70000 473486 70074 473542
rect 70130 473486 70200 473542
rect 70000 473418 70200 473486
rect 70000 473362 70074 473418
rect 70130 473362 70200 473418
rect 70000 473294 70200 473362
rect 70000 473238 70074 473294
rect 70130 473238 70200 473294
rect 70000 473170 70200 473238
rect 70000 473114 70074 473170
rect 70130 473114 70200 473170
rect 70000 473046 70200 473114
rect 70000 472990 70074 473046
rect 70130 472990 70200 473046
rect 70000 472922 70200 472990
rect 70000 472866 70074 472922
rect 70130 472866 70200 472922
rect 70000 472828 70200 472866
rect 77678 474670 78678 482173
rect 77678 474614 77808 474670
rect 77864 474614 77932 474670
rect 77988 474614 78056 474670
rect 78112 474614 78180 474670
rect 78236 474614 78304 474670
rect 78360 474614 78428 474670
rect 78484 474614 78552 474670
rect 78608 474614 78678 474670
rect 77678 474546 78678 474614
rect 77678 474490 77808 474546
rect 77864 474490 77932 474546
rect 77988 474490 78056 474546
rect 78112 474490 78180 474546
rect 78236 474490 78304 474546
rect 78360 474490 78428 474546
rect 78484 474490 78552 474546
rect 78608 474490 78678 474546
rect 77678 474422 78678 474490
rect 77678 474366 77808 474422
rect 77864 474366 77932 474422
rect 77988 474366 78056 474422
rect 78112 474366 78180 474422
rect 78236 474366 78304 474422
rect 78360 474366 78428 474422
rect 78484 474366 78552 474422
rect 78608 474366 78678 474422
rect 77678 474298 78678 474366
rect 77678 474242 77808 474298
rect 77864 474242 77932 474298
rect 77988 474242 78056 474298
rect 78112 474242 78180 474298
rect 78236 474242 78304 474298
rect 78360 474242 78428 474298
rect 78484 474242 78552 474298
rect 78608 474242 78678 474298
rect 77678 474174 78678 474242
rect 77678 474118 77808 474174
rect 77864 474118 77932 474174
rect 77988 474118 78056 474174
rect 78112 474118 78180 474174
rect 78236 474118 78304 474174
rect 78360 474118 78428 474174
rect 78484 474118 78552 474174
rect 78608 474118 78678 474174
rect 77678 474050 78678 474118
rect 77678 473994 77808 474050
rect 77864 473994 77932 474050
rect 77988 473994 78056 474050
rect 78112 473994 78180 474050
rect 78236 473994 78304 474050
rect 78360 473994 78428 474050
rect 78484 473994 78552 474050
rect 78608 473994 78678 474050
rect 77678 473926 78678 473994
rect 77678 473870 77808 473926
rect 77864 473870 77932 473926
rect 77988 473870 78056 473926
rect 78112 473870 78180 473926
rect 78236 473870 78304 473926
rect 78360 473870 78428 473926
rect 78484 473870 78552 473926
rect 78608 473870 78678 473926
rect 77678 473802 78678 473870
rect 77678 473746 77808 473802
rect 77864 473746 77932 473802
rect 77988 473746 78056 473802
rect 78112 473746 78180 473802
rect 78236 473746 78304 473802
rect 78360 473746 78428 473802
rect 78484 473746 78552 473802
rect 78608 473746 78678 473802
rect 77678 473678 78678 473746
rect 77678 473622 77808 473678
rect 77864 473622 77932 473678
rect 77988 473622 78056 473678
rect 78112 473622 78180 473678
rect 78236 473622 78304 473678
rect 78360 473622 78428 473678
rect 78484 473622 78552 473678
rect 78608 473622 78678 473678
rect 77678 473554 78678 473622
rect 77678 473498 77808 473554
rect 77864 473498 77932 473554
rect 77988 473498 78056 473554
rect 78112 473498 78180 473554
rect 78236 473498 78304 473554
rect 78360 473498 78428 473554
rect 78484 473498 78552 473554
rect 78608 473498 78678 473554
rect 77678 473430 78678 473498
rect 77678 473374 77808 473430
rect 77864 473374 77932 473430
rect 77988 473374 78056 473430
rect 78112 473374 78180 473430
rect 78236 473374 78304 473430
rect 78360 473374 78428 473430
rect 78484 473374 78552 473430
rect 78608 473374 78678 473430
rect 77678 473306 78678 473374
rect 77678 473250 77808 473306
rect 77864 473250 77932 473306
rect 77988 473250 78056 473306
rect 78112 473250 78180 473306
rect 78236 473250 78304 473306
rect 78360 473250 78428 473306
rect 78484 473250 78552 473306
rect 78608 473250 78678 473306
rect 77678 473182 78678 473250
rect 77678 473126 77808 473182
rect 77864 473126 77932 473182
rect 77988 473126 78056 473182
rect 78112 473126 78180 473182
rect 78236 473126 78304 473182
rect 78360 473126 78428 473182
rect 78484 473126 78552 473182
rect 78608 473126 78678 473182
rect 77678 473058 78678 473126
rect 77678 473002 77808 473058
rect 77864 473002 77932 473058
rect 77988 473002 78056 473058
rect 78112 473002 78180 473058
rect 78236 473002 78304 473058
rect 78360 473002 78428 473058
rect 78484 473002 78552 473058
rect 78608 473002 78678 473058
rect 77678 472934 78678 473002
rect 77678 472878 77808 472934
rect 77864 472878 77932 472934
rect 77988 472878 78056 472934
rect 78112 472878 78180 472934
rect 78236 472878 78304 472934
rect 78360 472878 78428 472934
rect 78484 472878 78552 472934
rect 78608 472878 78678 472934
rect 70000 472184 70200 472248
rect 70000 472128 70074 472184
rect 70130 472128 70200 472184
rect 70000 472060 70200 472128
rect 70000 472004 70074 472060
rect 70130 472004 70200 472060
rect 70000 471936 70200 472004
rect 70000 471880 70074 471936
rect 70130 471880 70200 471936
rect 70000 471812 70200 471880
rect 70000 471756 70074 471812
rect 70130 471756 70200 471812
rect 70000 471688 70200 471756
rect 70000 471632 70074 471688
rect 70130 471632 70200 471688
rect 70000 471564 70200 471632
rect 70000 471508 70074 471564
rect 70130 471508 70200 471564
rect 70000 471440 70200 471508
rect 70000 471384 70074 471440
rect 70130 471384 70200 471440
rect 70000 471316 70200 471384
rect 70000 471260 70074 471316
rect 70130 471260 70200 471316
rect 70000 471192 70200 471260
rect 70000 471136 70074 471192
rect 70130 471136 70200 471192
rect 70000 471068 70200 471136
rect 70000 471012 70074 471068
rect 70130 471012 70200 471068
rect 70000 470944 70200 471012
rect 70000 470888 70074 470944
rect 70130 470888 70200 470944
rect 70000 470820 70200 470888
rect 70000 470764 70074 470820
rect 70130 470764 70200 470820
rect 70000 470696 70200 470764
rect 70000 470640 70074 470696
rect 70130 470640 70200 470696
rect 70000 470572 70200 470640
rect 70000 470516 70074 470572
rect 70130 470516 70200 470572
rect 70000 470448 70200 470516
rect 70000 470392 70074 470448
rect 70130 470392 70200 470448
rect 70000 470324 70200 470392
rect 70000 470268 70074 470324
rect 70130 470268 70200 470324
rect 70000 470198 70200 470268
rect 77678 472190 78678 472878
rect 77678 472134 77808 472190
rect 77864 472134 77932 472190
rect 77988 472134 78056 472190
rect 78112 472134 78180 472190
rect 78236 472134 78304 472190
rect 78360 472134 78428 472190
rect 78484 472134 78552 472190
rect 78608 472134 78678 472190
rect 77678 472066 78678 472134
rect 77678 472010 77808 472066
rect 77864 472010 77932 472066
rect 77988 472010 78056 472066
rect 78112 472010 78180 472066
rect 78236 472010 78304 472066
rect 78360 472010 78428 472066
rect 78484 472010 78552 472066
rect 78608 472010 78678 472066
rect 77678 471942 78678 472010
rect 77678 471886 77808 471942
rect 77864 471886 77932 471942
rect 77988 471886 78056 471942
rect 78112 471886 78180 471942
rect 78236 471886 78304 471942
rect 78360 471886 78428 471942
rect 78484 471886 78552 471942
rect 78608 471886 78678 471942
rect 77678 471818 78678 471886
rect 77678 471762 77808 471818
rect 77864 471762 77932 471818
rect 77988 471762 78056 471818
rect 78112 471762 78180 471818
rect 78236 471762 78304 471818
rect 78360 471762 78428 471818
rect 78484 471762 78552 471818
rect 78608 471762 78678 471818
rect 77678 471694 78678 471762
rect 77678 471638 77808 471694
rect 77864 471638 77932 471694
rect 77988 471638 78056 471694
rect 78112 471638 78180 471694
rect 78236 471638 78304 471694
rect 78360 471638 78428 471694
rect 78484 471638 78552 471694
rect 78608 471638 78678 471694
rect 77678 471570 78678 471638
rect 77678 471514 77808 471570
rect 77864 471514 77932 471570
rect 77988 471514 78056 471570
rect 78112 471514 78180 471570
rect 78236 471514 78304 471570
rect 78360 471514 78428 471570
rect 78484 471514 78552 471570
rect 78608 471514 78678 471570
rect 77678 471446 78678 471514
rect 77678 471390 77808 471446
rect 77864 471390 77932 471446
rect 77988 471390 78056 471446
rect 78112 471390 78180 471446
rect 78236 471390 78304 471446
rect 78360 471390 78428 471446
rect 78484 471390 78552 471446
rect 78608 471390 78678 471446
rect 77678 471322 78678 471390
rect 77678 471266 77808 471322
rect 77864 471266 77932 471322
rect 77988 471266 78056 471322
rect 78112 471266 78180 471322
rect 78236 471266 78304 471322
rect 78360 471266 78428 471322
rect 78484 471266 78552 471322
rect 78608 471266 78678 471322
rect 77678 471198 78678 471266
rect 77678 471142 77808 471198
rect 77864 471142 77932 471198
rect 77988 471142 78056 471198
rect 78112 471142 78180 471198
rect 78236 471142 78304 471198
rect 78360 471142 78428 471198
rect 78484 471142 78552 471198
rect 78608 471142 78678 471198
rect 77678 471074 78678 471142
rect 77678 471018 77808 471074
rect 77864 471018 77932 471074
rect 77988 471018 78056 471074
rect 78112 471018 78180 471074
rect 78236 471018 78304 471074
rect 78360 471018 78428 471074
rect 78484 471018 78552 471074
rect 78608 471018 78678 471074
rect 77678 470950 78678 471018
rect 77678 470894 77808 470950
rect 77864 470894 77932 470950
rect 77988 470894 78056 470950
rect 78112 470894 78180 470950
rect 78236 470894 78304 470950
rect 78360 470894 78428 470950
rect 78484 470894 78552 470950
rect 78608 470894 78678 470950
rect 77678 470826 78678 470894
rect 77678 470770 77808 470826
rect 77864 470770 77932 470826
rect 77988 470770 78056 470826
rect 78112 470770 78180 470826
rect 78236 470770 78304 470826
rect 78360 470770 78428 470826
rect 78484 470770 78552 470826
rect 78608 470770 78678 470826
rect 77678 470702 78678 470770
rect 77678 470646 77808 470702
rect 77864 470646 77932 470702
rect 77988 470646 78056 470702
rect 78112 470646 78180 470702
rect 78236 470646 78304 470702
rect 78360 470646 78428 470702
rect 78484 470646 78552 470702
rect 78608 470646 78678 470702
rect 77678 470578 78678 470646
rect 77678 470522 77808 470578
rect 77864 470522 77932 470578
rect 77988 470522 78056 470578
rect 78112 470522 78180 470578
rect 78236 470522 78304 470578
rect 78360 470522 78428 470578
rect 78484 470522 78552 470578
rect 78608 470522 78678 470578
rect 77678 470454 78678 470522
rect 77678 470398 77808 470454
rect 77864 470398 77932 470454
rect 77988 470398 78056 470454
rect 78112 470398 78180 470454
rect 78236 470398 78304 470454
rect 78360 470398 78428 470454
rect 78484 470398 78552 470454
rect 78608 470398 78678 470454
rect 77678 470330 78678 470398
rect 77678 470274 77808 470330
rect 77864 470274 77932 470330
rect 77988 470274 78056 470330
rect 78112 470274 78180 470330
rect 78236 470274 78304 470330
rect 78360 470274 78428 470330
rect 78484 470274 78552 470330
rect 78608 470274 78678 470330
rect 70000 469814 70200 469878
rect 70000 469758 70074 469814
rect 70130 469758 70200 469814
rect 70000 469690 70200 469758
rect 70000 469634 70074 469690
rect 70130 469634 70200 469690
rect 70000 469566 70200 469634
rect 70000 469510 70074 469566
rect 70130 469510 70200 469566
rect 70000 469442 70200 469510
rect 70000 469386 70074 469442
rect 70130 469386 70200 469442
rect 70000 469318 70200 469386
rect 70000 469262 70074 469318
rect 70130 469262 70200 469318
rect 70000 469194 70200 469262
rect 70000 469138 70074 469194
rect 70130 469138 70200 469194
rect 70000 469070 70200 469138
rect 70000 469014 70074 469070
rect 70130 469014 70200 469070
rect 70000 468946 70200 469014
rect 70000 468890 70074 468946
rect 70130 468890 70200 468946
rect 70000 468822 70200 468890
rect 70000 468766 70074 468822
rect 70130 468766 70200 468822
rect 70000 468698 70200 468766
rect 70000 468642 70074 468698
rect 70130 468642 70200 468698
rect 70000 468574 70200 468642
rect 70000 468518 70074 468574
rect 70130 468518 70200 468574
rect 70000 468450 70200 468518
rect 70000 468394 70074 468450
rect 70130 468394 70200 468450
rect 70000 468326 70200 468394
rect 70000 468270 70074 468326
rect 70130 468270 70200 468326
rect 70000 468202 70200 468270
rect 70000 468146 70074 468202
rect 70130 468146 70200 468202
rect 70000 468078 70200 468146
rect 70000 468022 70074 468078
rect 70130 468022 70200 468078
rect 70000 467954 70200 468022
rect 70000 467898 70074 467954
rect 70130 467898 70200 467954
rect 70000 467828 70200 467898
rect 77678 469820 78678 470274
rect 77678 469764 77808 469820
rect 77864 469764 77932 469820
rect 77988 469764 78056 469820
rect 78112 469764 78180 469820
rect 78236 469764 78304 469820
rect 78360 469764 78428 469820
rect 78484 469764 78552 469820
rect 78608 469764 78678 469820
rect 77678 469696 78678 469764
rect 77678 469640 77808 469696
rect 77864 469640 77932 469696
rect 77988 469640 78056 469696
rect 78112 469640 78180 469696
rect 78236 469640 78304 469696
rect 78360 469640 78428 469696
rect 78484 469640 78552 469696
rect 78608 469640 78678 469696
rect 77678 469572 78678 469640
rect 77678 469516 77808 469572
rect 77864 469516 77932 469572
rect 77988 469516 78056 469572
rect 78112 469516 78180 469572
rect 78236 469516 78304 469572
rect 78360 469516 78428 469572
rect 78484 469516 78552 469572
rect 78608 469516 78678 469572
rect 77678 469448 78678 469516
rect 77678 469392 77808 469448
rect 77864 469392 77932 469448
rect 77988 469392 78056 469448
rect 78112 469392 78180 469448
rect 78236 469392 78304 469448
rect 78360 469392 78428 469448
rect 78484 469392 78552 469448
rect 78608 469392 78678 469448
rect 77678 469324 78678 469392
rect 77678 469268 77808 469324
rect 77864 469268 77932 469324
rect 77988 469268 78056 469324
rect 78112 469268 78180 469324
rect 78236 469268 78304 469324
rect 78360 469268 78428 469324
rect 78484 469268 78552 469324
rect 78608 469268 78678 469324
rect 77678 469200 78678 469268
rect 77678 469144 77808 469200
rect 77864 469144 77932 469200
rect 77988 469144 78056 469200
rect 78112 469144 78180 469200
rect 78236 469144 78304 469200
rect 78360 469144 78428 469200
rect 78484 469144 78552 469200
rect 78608 469144 78678 469200
rect 77678 469076 78678 469144
rect 77678 469020 77808 469076
rect 77864 469020 77932 469076
rect 77988 469020 78056 469076
rect 78112 469020 78180 469076
rect 78236 469020 78304 469076
rect 78360 469020 78428 469076
rect 78484 469020 78552 469076
rect 78608 469020 78678 469076
rect 77678 468952 78678 469020
rect 77678 468896 77808 468952
rect 77864 468896 77932 468952
rect 77988 468896 78056 468952
rect 78112 468896 78180 468952
rect 78236 468896 78304 468952
rect 78360 468896 78428 468952
rect 78484 468896 78552 468952
rect 78608 468896 78678 468952
rect 77678 468828 78678 468896
rect 77678 468772 77808 468828
rect 77864 468772 77932 468828
rect 77988 468772 78056 468828
rect 78112 468772 78180 468828
rect 78236 468772 78304 468828
rect 78360 468772 78428 468828
rect 78484 468772 78552 468828
rect 78608 468772 78678 468828
rect 77678 468704 78678 468772
rect 77678 468648 77808 468704
rect 77864 468648 77932 468704
rect 77988 468648 78056 468704
rect 78112 468648 78180 468704
rect 78236 468648 78304 468704
rect 78360 468648 78428 468704
rect 78484 468648 78552 468704
rect 78608 468648 78678 468704
rect 77678 468580 78678 468648
rect 77678 468524 77808 468580
rect 77864 468524 77932 468580
rect 77988 468524 78056 468580
rect 78112 468524 78180 468580
rect 78236 468524 78304 468580
rect 78360 468524 78428 468580
rect 78484 468524 78552 468580
rect 78608 468524 78678 468580
rect 77678 468456 78678 468524
rect 77678 468400 77808 468456
rect 77864 468400 77932 468456
rect 77988 468400 78056 468456
rect 78112 468400 78180 468456
rect 78236 468400 78304 468456
rect 78360 468400 78428 468456
rect 78484 468400 78552 468456
rect 78608 468400 78678 468456
rect 77678 468332 78678 468400
rect 77678 468276 77808 468332
rect 77864 468276 77932 468332
rect 77988 468276 78056 468332
rect 78112 468276 78180 468332
rect 78236 468276 78304 468332
rect 78360 468276 78428 468332
rect 78484 468276 78552 468332
rect 78608 468276 78678 468332
rect 77678 468208 78678 468276
rect 77678 468152 77808 468208
rect 77864 468152 77932 468208
rect 77988 468152 78056 468208
rect 78112 468152 78180 468208
rect 78236 468152 78304 468208
rect 78360 468152 78428 468208
rect 78484 468152 78552 468208
rect 78608 468152 78678 468208
rect 77678 468084 78678 468152
rect 77678 468028 77808 468084
rect 77864 468028 77932 468084
rect 77988 468028 78056 468084
rect 78112 468028 78180 468084
rect 78236 468028 78304 468084
rect 78360 468028 78428 468084
rect 78484 468028 78552 468084
rect 78608 468028 78678 468084
rect 77678 467960 78678 468028
rect 77678 467904 77808 467960
rect 77864 467904 77932 467960
rect 77988 467904 78056 467960
rect 78112 467904 78180 467960
rect 78236 467904 78304 467960
rect 78360 467904 78428 467960
rect 78484 467904 78552 467960
rect 78608 467904 78678 467960
rect 70000 467108 70200 467172
rect 70000 467052 70074 467108
rect 70130 467052 70200 467108
rect 70000 466984 70200 467052
rect 70000 466928 70074 466984
rect 70130 466928 70200 466984
rect 70000 466860 70200 466928
rect 70000 466804 70074 466860
rect 70130 466804 70200 466860
rect 70000 466736 70200 466804
rect 70000 466680 70074 466736
rect 70130 466680 70200 466736
rect 70000 466612 70200 466680
rect 70000 466556 70074 466612
rect 70130 466556 70200 466612
rect 70000 466488 70200 466556
rect 70000 466432 70074 466488
rect 70130 466432 70200 466488
rect 70000 466364 70200 466432
rect 70000 466308 70074 466364
rect 70130 466308 70200 466364
rect 70000 466240 70200 466308
rect 70000 466184 70074 466240
rect 70130 466184 70200 466240
rect 70000 466116 70200 466184
rect 70000 466060 70074 466116
rect 70130 466060 70200 466116
rect 70000 465992 70200 466060
rect 70000 465936 70074 465992
rect 70130 465936 70200 465992
rect 70000 465868 70200 465936
rect 70000 465812 70074 465868
rect 70130 465812 70200 465868
rect 70000 465744 70200 465812
rect 70000 465688 70074 465744
rect 70130 465688 70200 465744
rect 70000 465620 70200 465688
rect 70000 465564 70074 465620
rect 70130 465564 70200 465620
rect 70000 465496 70200 465564
rect 70000 465440 70074 465496
rect 70130 465440 70200 465496
rect 70000 465372 70200 465440
rect 70000 465316 70074 465372
rect 70130 465316 70200 465372
rect 70000 465248 70200 465316
rect 70000 465192 70074 465248
rect 70130 465192 70200 465248
rect 70000 465122 70200 465192
rect 77678 467114 78678 467904
rect 77678 467058 77808 467114
rect 77864 467058 77932 467114
rect 77988 467058 78056 467114
rect 78112 467058 78180 467114
rect 78236 467058 78304 467114
rect 78360 467058 78428 467114
rect 78484 467058 78552 467114
rect 78608 467058 78678 467114
rect 77678 466990 78678 467058
rect 77678 466934 77808 466990
rect 77864 466934 77932 466990
rect 77988 466934 78056 466990
rect 78112 466934 78180 466990
rect 78236 466934 78304 466990
rect 78360 466934 78428 466990
rect 78484 466934 78552 466990
rect 78608 466934 78678 466990
rect 77678 466866 78678 466934
rect 77678 466810 77808 466866
rect 77864 466810 77932 466866
rect 77988 466810 78056 466866
rect 78112 466810 78180 466866
rect 78236 466810 78304 466866
rect 78360 466810 78428 466866
rect 78484 466810 78552 466866
rect 78608 466810 78678 466866
rect 77678 466742 78678 466810
rect 77678 466686 77808 466742
rect 77864 466686 77932 466742
rect 77988 466686 78056 466742
rect 78112 466686 78180 466742
rect 78236 466686 78304 466742
rect 78360 466686 78428 466742
rect 78484 466686 78552 466742
rect 78608 466686 78678 466742
rect 77678 466618 78678 466686
rect 77678 466562 77808 466618
rect 77864 466562 77932 466618
rect 77988 466562 78056 466618
rect 78112 466562 78180 466618
rect 78236 466562 78304 466618
rect 78360 466562 78428 466618
rect 78484 466562 78552 466618
rect 78608 466562 78678 466618
rect 77678 466494 78678 466562
rect 77678 466438 77808 466494
rect 77864 466438 77932 466494
rect 77988 466438 78056 466494
rect 78112 466438 78180 466494
rect 78236 466438 78304 466494
rect 78360 466438 78428 466494
rect 78484 466438 78552 466494
rect 78608 466438 78678 466494
rect 77678 466370 78678 466438
rect 77678 466314 77808 466370
rect 77864 466314 77932 466370
rect 77988 466314 78056 466370
rect 78112 466314 78180 466370
rect 78236 466314 78304 466370
rect 78360 466314 78428 466370
rect 78484 466314 78552 466370
rect 78608 466314 78678 466370
rect 77678 466246 78678 466314
rect 77678 466190 77808 466246
rect 77864 466190 77932 466246
rect 77988 466190 78056 466246
rect 78112 466190 78180 466246
rect 78236 466190 78304 466246
rect 78360 466190 78428 466246
rect 78484 466190 78552 466246
rect 78608 466190 78678 466246
rect 77678 466122 78678 466190
rect 77678 466066 77808 466122
rect 77864 466066 77932 466122
rect 77988 466066 78056 466122
rect 78112 466066 78180 466122
rect 78236 466066 78304 466122
rect 78360 466066 78428 466122
rect 78484 466066 78552 466122
rect 78608 466066 78678 466122
rect 77678 465998 78678 466066
rect 77678 465942 77808 465998
rect 77864 465942 77932 465998
rect 77988 465942 78056 465998
rect 78112 465942 78180 465998
rect 78236 465942 78304 465998
rect 78360 465942 78428 465998
rect 78484 465942 78552 465998
rect 78608 465942 78678 465998
rect 77678 465874 78678 465942
rect 77678 465818 77808 465874
rect 77864 465818 77932 465874
rect 77988 465818 78056 465874
rect 78112 465818 78180 465874
rect 78236 465818 78304 465874
rect 78360 465818 78428 465874
rect 78484 465818 78552 465874
rect 78608 465818 78678 465874
rect 77678 465750 78678 465818
rect 77678 465694 77808 465750
rect 77864 465694 77932 465750
rect 77988 465694 78056 465750
rect 78112 465694 78180 465750
rect 78236 465694 78304 465750
rect 78360 465694 78428 465750
rect 78484 465694 78552 465750
rect 78608 465694 78678 465750
rect 77678 465626 78678 465694
rect 77678 465570 77808 465626
rect 77864 465570 77932 465626
rect 77988 465570 78056 465626
rect 78112 465570 78180 465626
rect 78236 465570 78304 465626
rect 78360 465570 78428 465626
rect 78484 465570 78552 465626
rect 78608 465570 78678 465626
rect 77678 465502 78678 465570
rect 77678 465446 77808 465502
rect 77864 465446 77932 465502
rect 77988 465446 78056 465502
rect 78112 465446 78180 465502
rect 78236 465446 78304 465502
rect 78360 465446 78428 465502
rect 78484 465446 78552 465502
rect 78608 465446 78678 465502
rect 77678 465378 78678 465446
rect 77678 465322 77808 465378
rect 77864 465322 77932 465378
rect 77988 465322 78056 465378
rect 78112 465322 78180 465378
rect 78236 465322 78304 465378
rect 78360 465322 78428 465378
rect 78484 465322 78552 465378
rect 78608 465322 78678 465378
rect 77678 465254 78678 465322
rect 77678 465198 77808 465254
rect 77864 465198 77932 465254
rect 77988 465198 78056 465254
rect 78112 465198 78180 465254
rect 78236 465198 78304 465254
rect 78360 465198 78428 465254
rect 78484 465198 78552 465254
rect 78608 465198 78678 465254
rect 70000 464738 70200 464802
rect 70000 464682 70074 464738
rect 70130 464682 70200 464738
rect 70000 464614 70200 464682
rect 70000 464558 70074 464614
rect 70130 464558 70200 464614
rect 70000 464490 70200 464558
rect 70000 464434 70074 464490
rect 70130 464434 70200 464490
rect 70000 464366 70200 464434
rect 70000 464310 70074 464366
rect 70130 464310 70200 464366
rect 70000 464242 70200 464310
rect 70000 464186 70074 464242
rect 70130 464186 70200 464242
rect 70000 464118 70200 464186
rect 70000 464062 70074 464118
rect 70130 464062 70200 464118
rect 70000 463994 70200 464062
rect 70000 463938 70074 463994
rect 70130 463938 70200 463994
rect 70000 463870 70200 463938
rect 70000 463814 70074 463870
rect 70130 463814 70200 463870
rect 70000 463746 70200 463814
rect 70000 463690 70074 463746
rect 70130 463690 70200 463746
rect 70000 463622 70200 463690
rect 70000 463566 70074 463622
rect 70130 463566 70200 463622
rect 70000 463498 70200 463566
rect 70000 463442 70074 463498
rect 70130 463442 70200 463498
rect 70000 463374 70200 463442
rect 70000 463318 70074 463374
rect 70130 463318 70200 463374
rect 70000 463250 70200 463318
rect 70000 463194 70074 463250
rect 70130 463194 70200 463250
rect 70000 463126 70200 463194
rect 70000 463070 70074 463126
rect 70130 463070 70200 463126
rect 70000 463002 70200 463070
rect 70000 462946 70074 463002
rect 70130 462946 70200 463002
rect 70000 462878 70200 462946
rect 70000 462822 70074 462878
rect 70130 462822 70200 462878
rect 70000 462752 70200 462822
rect 77678 464744 78678 465198
rect 77678 464688 77808 464744
rect 77864 464688 77932 464744
rect 77988 464688 78056 464744
rect 78112 464688 78180 464744
rect 78236 464688 78304 464744
rect 78360 464688 78428 464744
rect 78484 464688 78552 464744
rect 78608 464688 78678 464744
rect 77678 464620 78678 464688
rect 77678 464564 77808 464620
rect 77864 464564 77932 464620
rect 77988 464564 78056 464620
rect 78112 464564 78180 464620
rect 78236 464564 78304 464620
rect 78360 464564 78428 464620
rect 78484 464564 78552 464620
rect 78608 464564 78678 464620
rect 77678 464496 78678 464564
rect 77678 464440 77808 464496
rect 77864 464440 77932 464496
rect 77988 464440 78056 464496
rect 78112 464440 78180 464496
rect 78236 464440 78304 464496
rect 78360 464440 78428 464496
rect 78484 464440 78552 464496
rect 78608 464440 78678 464496
rect 77678 464372 78678 464440
rect 77678 464316 77808 464372
rect 77864 464316 77932 464372
rect 77988 464316 78056 464372
rect 78112 464316 78180 464372
rect 78236 464316 78304 464372
rect 78360 464316 78428 464372
rect 78484 464316 78552 464372
rect 78608 464316 78678 464372
rect 77678 464248 78678 464316
rect 77678 464192 77808 464248
rect 77864 464192 77932 464248
rect 77988 464192 78056 464248
rect 78112 464192 78180 464248
rect 78236 464192 78304 464248
rect 78360 464192 78428 464248
rect 78484 464192 78552 464248
rect 78608 464192 78678 464248
rect 77678 464124 78678 464192
rect 77678 464068 77808 464124
rect 77864 464068 77932 464124
rect 77988 464068 78056 464124
rect 78112 464068 78180 464124
rect 78236 464068 78304 464124
rect 78360 464068 78428 464124
rect 78484 464068 78552 464124
rect 78608 464068 78678 464124
rect 77678 464000 78678 464068
rect 77678 463944 77808 464000
rect 77864 463944 77932 464000
rect 77988 463944 78056 464000
rect 78112 463944 78180 464000
rect 78236 463944 78304 464000
rect 78360 463944 78428 464000
rect 78484 463944 78552 464000
rect 78608 463944 78678 464000
rect 77678 463876 78678 463944
rect 77678 463820 77808 463876
rect 77864 463820 77932 463876
rect 77988 463820 78056 463876
rect 78112 463820 78180 463876
rect 78236 463820 78304 463876
rect 78360 463820 78428 463876
rect 78484 463820 78552 463876
rect 78608 463820 78678 463876
rect 77678 463752 78678 463820
rect 77678 463696 77808 463752
rect 77864 463696 77932 463752
rect 77988 463696 78056 463752
rect 78112 463696 78180 463752
rect 78236 463696 78304 463752
rect 78360 463696 78428 463752
rect 78484 463696 78552 463752
rect 78608 463696 78678 463752
rect 77678 463628 78678 463696
rect 77678 463572 77808 463628
rect 77864 463572 77932 463628
rect 77988 463572 78056 463628
rect 78112 463572 78180 463628
rect 78236 463572 78304 463628
rect 78360 463572 78428 463628
rect 78484 463572 78552 463628
rect 78608 463572 78678 463628
rect 77678 463504 78678 463572
rect 77678 463448 77808 463504
rect 77864 463448 77932 463504
rect 77988 463448 78056 463504
rect 78112 463448 78180 463504
rect 78236 463448 78304 463504
rect 78360 463448 78428 463504
rect 78484 463448 78552 463504
rect 78608 463448 78678 463504
rect 77678 463380 78678 463448
rect 77678 463324 77808 463380
rect 77864 463324 77932 463380
rect 77988 463324 78056 463380
rect 78112 463324 78180 463380
rect 78236 463324 78304 463380
rect 78360 463324 78428 463380
rect 78484 463324 78552 463380
rect 78608 463324 78678 463380
rect 77678 463256 78678 463324
rect 77678 463200 77808 463256
rect 77864 463200 77932 463256
rect 77988 463200 78056 463256
rect 78112 463200 78180 463256
rect 78236 463200 78304 463256
rect 78360 463200 78428 463256
rect 78484 463200 78552 463256
rect 78608 463200 78678 463256
rect 77678 463132 78678 463200
rect 77678 463076 77808 463132
rect 77864 463076 77932 463132
rect 77988 463076 78056 463132
rect 78112 463076 78180 463132
rect 78236 463076 78304 463132
rect 78360 463076 78428 463132
rect 78484 463076 78552 463132
rect 78608 463076 78678 463132
rect 77678 463008 78678 463076
rect 77678 462952 77808 463008
rect 77864 462952 77932 463008
rect 77988 462952 78056 463008
rect 78112 462952 78180 463008
rect 78236 462952 78304 463008
rect 78360 462952 78428 463008
rect 78484 462952 78552 463008
rect 78608 462952 78678 463008
rect 77678 462884 78678 462952
rect 77678 462828 77808 462884
rect 77864 462828 77932 462884
rect 77988 462828 78056 462884
rect 78112 462828 78180 462884
rect 78236 462828 78304 462884
rect 78360 462828 78428 462884
rect 78484 462828 78552 462884
rect 78608 462828 78678 462884
rect 70000 462134 70200 462172
rect 70000 462078 70074 462134
rect 70130 462078 70200 462134
rect 70000 462010 70200 462078
rect 70000 461954 70074 462010
rect 70130 461954 70200 462010
rect 70000 461886 70200 461954
rect 70000 461830 70074 461886
rect 70130 461830 70200 461886
rect 70000 461762 70200 461830
rect 70000 461706 70074 461762
rect 70130 461706 70200 461762
rect 70000 461638 70200 461706
rect 70000 461582 70074 461638
rect 70130 461582 70200 461638
rect 70000 461514 70200 461582
rect 70000 461458 70074 461514
rect 70130 461458 70200 461514
rect 70000 461390 70200 461458
rect 70000 461334 70074 461390
rect 70130 461334 70200 461390
rect 70000 461266 70200 461334
rect 70000 461210 70074 461266
rect 70130 461210 70200 461266
rect 70000 461142 70200 461210
rect 70000 461086 70074 461142
rect 70130 461086 70200 461142
rect 70000 461018 70200 461086
rect 70000 460962 70074 461018
rect 70130 460962 70200 461018
rect 70000 460894 70200 460962
rect 70000 460838 70074 460894
rect 70130 460838 70200 460894
rect 70000 460770 70200 460838
rect 70000 460714 70074 460770
rect 70130 460714 70200 460770
rect 70000 460646 70200 460714
rect 70000 460590 70074 460646
rect 70130 460590 70200 460646
rect 70000 460522 70200 460590
rect 70000 460466 70074 460522
rect 70130 460466 70200 460522
rect 70000 460398 70200 460466
rect 70000 460342 70074 460398
rect 70130 460342 70200 460398
rect 70000 460272 70200 460342
rect 77678 462140 78678 462828
rect 77678 462084 77808 462140
rect 77864 462084 77932 462140
rect 77988 462084 78056 462140
rect 78112 462084 78180 462140
rect 78236 462084 78304 462140
rect 78360 462084 78428 462140
rect 78484 462084 78552 462140
rect 78608 462084 78678 462140
rect 77678 462016 78678 462084
rect 77678 461960 77808 462016
rect 77864 461960 77932 462016
rect 77988 461960 78056 462016
rect 78112 461960 78180 462016
rect 78236 461960 78304 462016
rect 78360 461960 78428 462016
rect 78484 461960 78552 462016
rect 78608 461960 78678 462016
rect 77678 461892 78678 461960
rect 77678 461836 77808 461892
rect 77864 461836 77932 461892
rect 77988 461836 78056 461892
rect 78112 461836 78180 461892
rect 78236 461836 78304 461892
rect 78360 461836 78428 461892
rect 78484 461836 78552 461892
rect 78608 461836 78678 461892
rect 77678 461768 78678 461836
rect 77678 461712 77808 461768
rect 77864 461712 77932 461768
rect 77988 461712 78056 461768
rect 78112 461712 78180 461768
rect 78236 461712 78304 461768
rect 78360 461712 78428 461768
rect 78484 461712 78552 461768
rect 78608 461712 78678 461768
rect 77678 461644 78678 461712
rect 77678 461588 77808 461644
rect 77864 461588 77932 461644
rect 77988 461588 78056 461644
rect 78112 461588 78180 461644
rect 78236 461588 78304 461644
rect 78360 461588 78428 461644
rect 78484 461588 78552 461644
rect 78608 461588 78678 461644
rect 77678 461520 78678 461588
rect 77678 461464 77808 461520
rect 77864 461464 77932 461520
rect 77988 461464 78056 461520
rect 78112 461464 78180 461520
rect 78236 461464 78304 461520
rect 78360 461464 78428 461520
rect 78484 461464 78552 461520
rect 78608 461464 78678 461520
rect 77678 461396 78678 461464
rect 77678 461340 77808 461396
rect 77864 461340 77932 461396
rect 77988 461340 78056 461396
rect 78112 461340 78180 461396
rect 78236 461340 78304 461396
rect 78360 461340 78428 461396
rect 78484 461340 78552 461396
rect 78608 461340 78678 461396
rect 77678 461272 78678 461340
rect 77678 461216 77808 461272
rect 77864 461216 77932 461272
rect 77988 461216 78056 461272
rect 78112 461216 78180 461272
rect 78236 461216 78304 461272
rect 78360 461216 78428 461272
rect 78484 461216 78552 461272
rect 78608 461216 78678 461272
rect 77678 461148 78678 461216
rect 77678 461092 77808 461148
rect 77864 461092 77932 461148
rect 77988 461092 78056 461148
rect 78112 461092 78180 461148
rect 78236 461092 78304 461148
rect 78360 461092 78428 461148
rect 78484 461092 78552 461148
rect 78608 461092 78678 461148
rect 77678 461024 78678 461092
rect 77678 460968 77808 461024
rect 77864 460968 77932 461024
rect 77988 460968 78056 461024
rect 78112 460968 78180 461024
rect 78236 460968 78304 461024
rect 78360 460968 78428 461024
rect 78484 460968 78552 461024
rect 78608 460968 78678 461024
rect 77678 460900 78678 460968
rect 77678 460844 77808 460900
rect 77864 460844 77932 460900
rect 77988 460844 78056 460900
rect 78112 460844 78180 460900
rect 78236 460844 78304 460900
rect 78360 460844 78428 460900
rect 78484 460844 78552 460900
rect 78608 460844 78678 460900
rect 77678 460776 78678 460844
rect 77678 460720 77808 460776
rect 77864 460720 77932 460776
rect 77988 460720 78056 460776
rect 78112 460720 78180 460776
rect 78236 460720 78304 460776
rect 78360 460720 78428 460776
rect 78484 460720 78552 460776
rect 78608 460720 78678 460776
rect 77678 460652 78678 460720
rect 77678 460596 77808 460652
rect 77864 460596 77932 460652
rect 77988 460596 78056 460652
rect 78112 460596 78180 460652
rect 78236 460596 78304 460652
rect 78360 460596 78428 460652
rect 78484 460596 78552 460652
rect 78608 460596 78678 460652
rect 77678 460528 78678 460596
rect 77678 460472 77808 460528
rect 77864 460472 77932 460528
rect 77988 460472 78056 460528
rect 78112 460472 78180 460528
rect 78236 460472 78304 460528
rect 78360 460472 78428 460528
rect 78484 460472 78552 460528
rect 78608 460472 78678 460528
rect 77678 460404 78678 460472
rect 77678 460348 77808 460404
rect 77864 460348 77932 460404
rect 77988 460348 78056 460404
rect 78112 460348 78180 460404
rect 78236 460348 78304 460404
rect 78360 460348 78428 460404
rect 78484 460348 78552 460404
rect 78608 460348 78678 460404
rect 77678 446429 78678 460348
rect 77678 446373 77800 446429
rect 77856 446373 78100 446429
rect 78156 446373 78400 446429
rect 78456 446373 78678 446429
rect 77678 446229 78678 446373
rect 77678 446173 77800 446229
rect 77856 446173 78100 446229
rect 78156 446173 78400 446229
rect 78456 446173 78678 446229
rect 70000 433658 70200 433729
rect 70000 433602 70074 433658
rect 70130 433602 70200 433658
rect 70000 433534 70200 433602
rect 70000 433478 70074 433534
rect 70130 433478 70200 433534
rect 70000 433410 70200 433478
rect 70000 433354 70074 433410
rect 70130 433354 70200 433410
rect 70000 433286 70200 433354
rect 70000 433230 70074 433286
rect 70130 433230 70200 433286
rect 70000 433162 70200 433230
rect 70000 433106 70074 433162
rect 70130 433106 70200 433162
rect 70000 433038 70200 433106
rect 70000 432982 70074 433038
rect 70130 432982 70200 433038
rect 70000 432914 70200 432982
rect 70000 432858 70074 432914
rect 70130 432858 70200 432914
rect 70000 432790 70200 432858
rect 70000 432734 70074 432790
rect 70130 432734 70200 432790
rect 70000 432666 70200 432734
rect 70000 432610 70074 432666
rect 70130 432610 70200 432666
rect 70000 432542 70200 432610
rect 70000 432486 70074 432542
rect 70130 432486 70200 432542
rect 70000 432418 70200 432486
rect 70000 432362 70074 432418
rect 70130 432362 70200 432418
rect 70000 432294 70200 432362
rect 70000 432238 70074 432294
rect 70130 432238 70200 432294
rect 70000 432170 70200 432238
rect 70000 432114 70074 432170
rect 70130 432114 70200 432170
rect 70000 432046 70200 432114
rect 70000 431990 70074 432046
rect 70130 431990 70200 432046
rect 70000 431922 70200 431990
rect 70000 431866 70074 431922
rect 70130 431866 70200 431922
rect 70000 431829 70200 431866
rect 70000 431184 70200 431249
rect 70000 431128 70074 431184
rect 70130 431128 70200 431184
rect 70000 431060 70200 431128
rect 70000 431004 70074 431060
rect 70130 431004 70200 431060
rect 70000 430936 70200 431004
rect 70000 430880 70074 430936
rect 70130 430880 70200 430936
rect 70000 430812 70200 430880
rect 70000 430756 70074 430812
rect 70130 430756 70200 430812
rect 70000 430688 70200 430756
rect 70000 430632 70074 430688
rect 70130 430632 70200 430688
rect 70000 430564 70200 430632
rect 70000 430508 70074 430564
rect 70130 430508 70200 430564
rect 70000 430440 70200 430508
rect 70000 430384 70074 430440
rect 70130 430384 70200 430440
rect 70000 430316 70200 430384
rect 70000 430260 70074 430316
rect 70130 430260 70200 430316
rect 70000 430192 70200 430260
rect 70000 430136 70074 430192
rect 70130 430136 70200 430192
rect 70000 430068 70200 430136
rect 70000 430012 70074 430068
rect 70130 430012 70200 430068
rect 70000 429944 70200 430012
rect 70000 429888 70074 429944
rect 70130 429888 70200 429944
rect 70000 429820 70200 429888
rect 70000 429764 70074 429820
rect 70130 429764 70200 429820
rect 70000 429696 70200 429764
rect 70000 429640 70074 429696
rect 70130 429640 70200 429696
rect 70000 429572 70200 429640
rect 70000 429516 70074 429572
rect 70130 429516 70200 429572
rect 70000 429448 70200 429516
rect 70000 429392 70074 429448
rect 70130 429392 70200 429448
rect 70000 429324 70200 429392
rect 70000 429268 70074 429324
rect 70130 429268 70200 429324
rect 70000 429199 70200 429268
rect 70000 428814 70200 428879
rect 70000 428758 70074 428814
rect 70130 428758 70200 428814
rect 70000 428690 70200 428758
rect 70000 428634 70074 428690
rect 70130 428634 70200 428690
rect 70000 428566 70200 428634
rect 70000 428510 70074 428566
rect 70130 428510 70200 428566
rect 70000 428442 70200 428510
rect 70000 428386 70074 428442
rect 70130 428386 70200 428442
rect 70000 428318 70200 428386
rect 70000 428262 70074 428318
rect 70130 428262 70200 428318
rect 70000 428194 70200 428262
rect 70000 428138 70074 428194
rect 70130 428138 70200 428194
rect 70000 428070 70200 428138
rect 70000 428014 70074 428070
rect 70130 428014 70200 428070
rect 70000 427946 70200 428014
rect 70000 427890 70074 427946
rect 70130 427890 70200 427946
rect 70000 427822 70200 427890
rect 70000 427766 70074 427822
rect 70130 427766 70200 427822
rect 70000 427698 70200 427766
rect 70000 427642 70074 427698
rect 70130 427642 70200 427698
rect 70000 427574 70200 427642
rect 70000 427518 70074 427574
rect 70130 427518 70200 427574
rect 70000 427450 70200 427518
rect 70000 427394 70074 427450
rect 70130 427394 70200 427450
rect 70000 427326 70200 427394
rect 70000 427270 70074 427326
rect 70130 427270 70200 427326
rect 70000 427202 70200 427270
rect 70000 427146 70074 427202
rect 70130 427146 70200 427202
rect 70000 427078 70200 427146
rect 70000 427022 70074 427078
rect 70130 427022 70200 427078
rect 70000 426954 70200 427022
rect 70000 426898 70074 426954
rect 70130 426898 70200 426954
rect 70000 426829 70200 426898
rect 70000 426108 70200 426173
rect 70000 426052 70074 426108
rect 70130 426052 70200 426108
rect 70000 425984 70200 426052
rect 70000 425928 70074 425984
rect 70130 425928 70200 425984
rect 70000 425860 70200 425928
rect 70000 425804 70074 425860
rect 70130 425804 70200 425860
rect 70000 425736 70200 425804
rect 70000 425680 70074 425736
rect 70130 425680 70200 425736
rect 70000 425612 70200 425680
rect 70000 425556 70074 425612
rect 70130 425556 70200 425612
rect 70000 425488 70200 425556
rect 70000 425432 70074 425488
rect 70130 425432 70200 425488
rect 70000 425364 70200 425432
rect 70000 425308 70074 425364
rect 70130 425308 70200 425364
rect 70000 425240 70200 425308
rect 70000 425184 70074 425240
rect 70130 425184 70200 425240
rect 70000 425116 70200 425184
rect 70000 425060 70074 425116
rect 70130 425060 70200 425116
rect 70000 424992 70200 425060
rect 70000 424936 70074 424992
rect 70130 424936 70200 424992
rect 70000 424868 70200 424936
rect 70000 424812 70074 424868
rect 70130 424812 70200 424868
rect 70000 424744 70200 424812
rect 70000 424688 70074 424744
rect 70130 424688 70200 424744
rect 70000 424620 70200 424688
rect 70000 424564 70074 424620
rect 70130 424564 70200 424620
rect 70000 424496 70200 424564
rect 70000 424440 70074 424496
rect 70130 424440 70200 424496
rect 70000 424372 70200 424440
rect 70000 424316 70074 424372
rect 70130 424316 70200 424372
rect 70000 424248 70200 424316
rect 70000 424192 70074 424248
rect 70130 424192 70200 424248
rect 70000 424123 70200 424192
rect 70000 423738 70200 423803
rect 70000 423682 70074 423738
rect 70130 423682 70200 423738
rect 70000 423614 70200 423682
rect 70000 423558 70074 423614
rect 70130 423558 70200 423614
rect 70000 423490 70200 423558
rect 70000 423434 70074 423490
rect 70130 423434 70200 423490
rect 70000 423366 70200 423434
rect 70000 423310 70074 423366
rect 70130 423310 70200 423366
rect 70000 423242 70200 423310
rect 70000 423186 70074 423242
rect 70130 423186 70200 423242
rect 70000 423118 70200 423186
rect 70000 423062 70074 423118
rect 70130 423062 70200 423118
rect 70000 422994 70200 423062
rect 70000 422938 70074 422994
rect 70130 422938 70200 422994
rect 70000 422870 70200 422938
rect 70000 422814 70074 422870
rect 70130 422814 70200 422870
rect 70000 422746 70200 422814
rect 70000 422690 70074 422746
rect 70130 422690 70200 422746
rect 70000 422622 70200 422690
rect 70000 422566 70074 422622
rect 70130 422566 70200 422622
rect 70000 422498 70200 422566
rect 70000 422442 70074 422498
rect 70130 422442 70200 422498
rect 70000 422374 70200 422442
rect 70000 422318 70074 422374
rect 70130 422318 70200 422374
rect 70000 422250 70200 422318
rect 70000 422194 70074 422250
rect 70130 422194 70200 422250
rect 70000 422126 70200 422194
rect 70000 422070 70074 422126
rect 70130 422070 70200 422126
rect 70000 422002 70200 422070
rect 70000 421946 70074 422002
rect 70130 421946 70200 422002
rect 70000 421878 70200 421946
rect 70000 421822 70074 421878
rect 70130 421822 70200 421878
rect 70000 421753 70200 421822
rect 70000 421134 70200 421173
rect 70000 421078 70074 421134
rect 70130 421078 70200 421134
rect 70000 421010 70200 421078
rect 70000 420954 70074 421010
rect 70130 420954 70200 421010
rect 70000 420886 70200 420954
rect 70000 420830 70074 420886
rect 70130 420830 70200 420886
rect 70000 420762 70200 420830
rect 70000 420706 70074 420762
rect 70130 420706 70200 420762
rect 70000 420638 70200 420706
rect 70000 420582 70074 420638
rect 70130 420582 70200 420638
rect 70000 420514 70200 420582
rect 70000 420458 70074 420514
rect 70130 420458 70200 420514
rect 70000 420390 70200 420458
rect 70000 420334 70074 420390
rect 70130 420334 70200 420390
rect 70000 420266 70200 420334
rect 70000 420210 70074 420266
rect 70130 420210 70200 420266
rect 70000 420142 70200 420210
rect 70000 420086 70074 420142
rect 70130 420086 70200 420142
rect 70000 420018 70200 420086
rect 70000 419962 70074 420018
rect 70130 419962 70200 420018
rect 70000 419894 70200 419962
rect 70000 419838 70074 419894
rect 70130 419838 70200 419894
rect 70000 419770 70200 419838
rect 70000 419714 70074 419770
rect 70130 419714 70200 419770
rect 70000 419646 70200 419714
rect 70000 419590 70074 419646
rect 70130 419590 70200 419646
rect 70000 419522 70200 419590
rect 70000 419466 70074 419522
rect 70130 419466 70200 419522
rect 70000 419398 70200 419466
rect 70000 419342 70074 419398
rect 70130 419342 70200 419398
rect 70000 419273 70200 419342
rect 77678 412633 78678 446173
rect 77678 412577 77847 412633
rect 77903 412577 78147 412633
rect 78203 412577 78447 412633
rect 78503 412577 78678 412633
rect 77678 410429 78678 412577
rect 77678 410373 77800 410429
rect 77856 410373 78100 410429
rect 78156 410373 78400 410429
rect 78456 410373 78678 410429
rect 77678 410229 78678 410373
rect 77678 410173 77800 410229
rect 77856 410173 78100 410229
rect 78156 410173 78400 410229
rect 78456 410173 78678 410229
rect 77678 393102 78678 410173
rect 77678 393046 77900 393102
rect 77956 393046 78200 393102
rect 78256 393046 78500 393102
rect 78556 393046 78678 393102
rect 77678 386102 78678 393046
rect 77678 386046 77900 386102
rect 77956 386046 78200 386102
rect 78256 386046 78500 386102
rect 78556 386046 78678 386102
rect 77678 379102 78678 386046
rect 77678 379046 77900 379102
rect 77956 379046 78200 379102
rect 78256 379046 78500 379102
rect 78556 379046 78678 379102
rect 77678 374429 78678 379046
rect 77678 374373 77800 374429
rect 77856 374373 78100 374429
rect 78156 374373 78400 374429
rect 78456 374373 78678 374429
rect 77678 374229 78678 374373
rect 77678 374173 77800 374229
rect 77856 374173 78100 374229
rect 78156 374173 78400 374229
rect 78456 374173 78678 374229
rect 77678 371633 78678 374173
rect 77678 371577 77847 371633
rect 77903 371577 78147 371633
rect 78203 371577 78447 371633
rect 78503 371577 78678 371633
rect 77678 352102 78678 371577
rect 77678 352046 77900 352102
rect 77956 352046 78200 352102
rect 78256 352046 78500 352102
rect 78556 352046 78678 352102
rect 77678 345102 78678 352046
rect 77678 345046 77900 345102
rect 77956 345046 78200 345102
rect 78256 345046 78500 345102
rect 78556 345046 78678 345102
rect 77678 338429 78678 345046
rect 77678 338373 77800 338429
rect 77856 338373 78100 338429
rect 78156 338373 78400 338429
rect 78456 338373 78678 338429
rect 77678 338229 78678 338373
rect 77678 338173 77800 338229
rect 77856 338173 78100 338229
rect 78156 338173 78400 338229
rect 78456 338173 78678 338229
rect 77678 338102 78678 338173
rect 77678 338046 77900 338102
rect 77956 338046 78200 338102
rect 78256 338046 78500 338102
rect 78556 338046 78678 338102
rect 77678 330633 78678 338046
rect 77678 330577 77847 330633
rect 77903 330577 78147 330633
rect 78203 330577 78447 330633
rect 78503 330577 78678 330633
rect 77678 329640 78678 330577
rect 77678 329584 77808 329640
rect 77864 329584 77932 329640
rect 77988 329584 78056 329640
rect 78112 329584 78180 329640
rect 78236 329584 78304 329640
rect 78360 329584 78428 329640
rect 78484 329584 78552 329640
rect 78608 329584 78678 329640
rect 77678 329516 78678 329584
rect 77678 329460 77808 329516
rect 77864 329460 77932 329516
rect 77988 329460 78056 329516
rect 78112 329460 78180 329516
rect 78236 329460 78304 329516
rect 78360 329460 78428 329516
rect 78484 329460 78552 329516
rect 78608 329460 78678 329516
rect 77678 329392 78678 329460
rect 77678 329336 77808 329392
rect 77864 329336 77932 329392
rect 77988 329336 78056 329392
rect 78112 329336 78180 329392
rect 78236 329336 78304 329392
rect 78360 329336 78428 329392
rect 78484 329336 78552 329392
rect 78608 329336 78678 329392
rect 77678 329268 78678 329336
rect 77678 329212 77808 329268
rect 77864 329212 77932 329268
rect 77988 329212 78056 329268
rect 78112 329212 78180 329268
rect 78236 329212 78304 329268
rect 78360 329212 78428 329268
rect 78484 329212 78552 329268
rect 78608 329212 78678 329268
rect 77678 329144 78678 329212
rect 77678 329088 77808 329144
rect 77864 329088 77932 329144
rect 77988 329088 78056 329144
rect 78112 329088 78180 329144
rect 78236 329088 78304 329144
rect 78360 329088 78428 329144
rect 78484 329088 78552 329144
rect 78608 329088 78678 329144
rect 77678 329020 78678 329088
rect 77678 328964 77808 329020
rect 77864 328964 77932 329020
rect 77988 328964 78056 329020
rect 78112 328964 78180 329020
rect 78236 328964 78304 329020
rect 78360 328964 78428 329020
rect 78484 328964 78552 329020
rect 78608 328964 78678 329020
rect 77678 328896 78678 328964
rect 77678 328840 77808 328896
rect 77864 328840 77932 328896
rect 77988 328840 78056 328896
rect 78112 328840 78180 328896
rect 78236 328840 78304 328896
rect 78360 328840 78428 328896
rect 78484 328840 78552 328896
rect 78608 328840 78678 328896
rect 77678 311102 78678 328840
rect 77678 311046 77900 311102
rect 77956 311046 78200 311102
rect 78256 311046 78500 311102
rect 78556 311046 78678 311102
rect 77678 305786 78678 311046
rect 77678 305730 77808 305786
rect 77864 305730 77932 305786
rect 77988 305730 78056 305786
rect 78112 305730 78180 305786
rect 78236 305730 78304 305786
rect 78360 305730 78428 305786
rect 78484 305730 78552 305786
rect 78608 305730 78678 305786
rect 77678 305662 78678 305730
rect 77678 305606 77808 305662
rect 77864 305606 77932 305662
rect 77988 305606 78056 305662
rect 78112 305606 78180 305662
rect 78236 305606 78304 305662
rect 78360 305606 78428 305662
rect 78484 305606 78552 305662
rect 78608 305606 78678 305662
rect 77678 305538 78678 305606
rect 77678 305482 77808 305538
rect 77864 305482 77932 305538
rect 77988 305482 78056 305538
rect 78112 305482 78180 305538
rect 78236 305482 78304 305538
rect 78360 305482 78428 305538
rect 78484 305482 78552 305538
rect 78608 305482 78678 305538
rect 77678 305414 78678 305482
rect 77678 305358 77808 305414
rect 77864 305358 77932 305414
rect 77988 305358 78056 305414
rect 78112 305358 78180 305414
rect 78236 305358 78304 305414
rect 78360 305358 78428 305414
rect 78484 305358 78552 305414
rect 78608 305358 78678 305414
rect 77678 305290 78678 305358
rect 77678 305234 77808 305290
rect 77864 305234 77932 305290
rect 77988 305234 78056 305290
rect 78112 305234 78180 305290
rect 78236 305234 78304 305290
rect 78360 305234 78428 305290
rect 78484 305234 78552 305290
rect 78608 305234 78678 305290
rect 77678 305166 78678 305234
rect 77678 305110 77808 305166
rect 77864 305110 77932 305166
rect 77988 305110 78056 305166
rect 78112 305110 78180 305166
rect 78236 305110 78304 305166
rect 78360 305110 78428 305166
rect 78484 305110 78552 305166
rect 78608 305110 78678 305166
rect 77678 305042 78678 305110
rect 77678 304986 77808 305042
rect 77864 304986 77932 305042
rect 77988 304986 78056 305042
rect 78112 304986 78180 305042
rect 78236 304986 78304 305042
rect 78360 304986 78428 305042
rect 78484 304986 78552 305042
rect 78608 304986 78678 305042
rect 77678 304122 78678 304986
rect 77678 304066 77800 304122
rect 77856 304066 78100 304122
rect 78156 304066 78400 304122
rect 78456 304066 78678 304122
rect 77678 297102 78678 304066
rect 77678 297046 77900 297102
rect 77956 297046 78200 297102
rect 78256 297046 78500 297102
rect 78556 297046 78678 297102
rect 77678 289633 78678 297046
rect 77678 289577 77847 289633
rect 77903 289577 78147 289633
rect 78203 289577 78447 289633
rect 78503 289577 78678 289633
rect 77678 281972 78678 289577
rect 77678 281916 77808 281972
rect 77864 281916 77932 281972
rect 77988 281916 78056 281972
rect 78112 281916 78180 281972
rect 78236 281916 78304 281972
rect 78360 281916 78428 281972
rect 78484 281916 78552 281972
rect 78608 281916 78678 281972
rect 77678 281848 78678 281916
rect 77678 281792 77808 281848
rect 77864 281792 77932 281848
rect 77988 281792 78056 281848
rect 78112 281792 78180 281848
rect 78236 281792 78304 281848
rect 78360 281792 78428 281848
rect 78484 281792 78552 281848
rect 78608 281792 78678 281848
rect 77678 281724 78678 281792
rect 77678 281668 77808 281724
rect 77864 281668 77932 281724
rect 77988 281668 78056 281724
rect 78112 281668 78180 281724
rect 78236 281668 78304 281724
rect 78360 281668 78428 281724
rect 78484 281668 78552 281724
rect 78608 281668 78678 281724
rect 77678 281600 78678 281668
rect 77678 281544 77808 281600
rect 77864 281544 77932 281600
rect 77988 281544 78056 281600
rect 78112 281544 78180 281600
rect 78236 281544 78304 281600
rect 78360 281544 78428 281600
rect 78484 281544 78552 281600
rect 78608 281544 78678 281600
rect 77678 281476 78678 281544
rect 77678 281420 77808 281476
rect 77864 281420 77932 281476
rect 77988 281420 78056 281476
rect 78112 281420 78180 281476
rect 78236 281420 78304 281476
rect 78360 281420 78428 281476
rect 78484 281420 78552 281476
rect 78608 281420 78678 281476
rect 77678 281352 78678 281420
rect 77678 281296 77808 281352
rect 77864 281296 77932 281352
rect 77988 281296 78056 281352
rect 78112 281296 78180 281352
rect 78236 281296 78304 281352
rect 78360 281296 78428 281352
rect 78484 281296 78552 281352
rect 78608 281296 78678 281352
rect 77678 281228 78678 281296
rect 77678 281172 77808 281228
rect 77864 281172 77932 281228
rect 77988 281172 78056 281228
rect 78112 281172 78180 281228
rect 78236 281172 78304 281228
rect 78360 281172 78428 281228
rect 78484 281172 78552 281228
rect 78608 281172 78678 281228
rect 77678 270102 78678 281172
rect 77678 270046 77900 270102
rect 77956 270046 78200 270102
rect 78256 270046 78500 270102
rect 78556 270046 78678 270102
rect 77678 268372 78678 270046
rect 77678 268316 77748 268372
rect 77804 268316 77872 268372
rect 77928 268316 77996 268372
rect 78052 268316 78120 268372
rect 78176 268316 78244 268372
rect 78300 268316 78368 268372
rect 78424 268316 78492 268372
rect 78548 268316 78678 268372
rect 77678 268248 78678 268316
rect 77678 268192 77748 268248
rect 77804 268192 77872 268248
rect 77928 268192 77996 268248
rect 78052 268192 78120 268248
rect 78176 268192 78244 268248
rect 78300 268192 78368 268248
rect 78424 268192 78492 268248
rect 78548 268192 78678 268248
rect 77678 263102 78678 268192
rect 77678 263046 77900 263102
rect 77956 263046 78200 263102
rect 78256 263046 78500 263102
rect 78556 263046 78678 263102
rect 77678 256102 78678 263046
rect 77678 256046 77900 256102
rect 77956 256046 78200 256102
rect 78256 256046 78500 256102
rect 78556 256046 78678 256102
rect 77678 248633 78678 256046
rect 77678 248577 77847 248633
rect 77903 248577 78147 248633
rect 78203 248577 78447 248633
rect 78503 248577 78678 248633
rect 77678 242372 78678 248577
rect 77678 242316 77748 242372
rect 77804 242316 77872 242372
rect 77928 242316 77996 242372
rect 78052 242316 78120 242372
rect 78176 242316 78244 242372
rect 78300 242316 78368 242372
rect 78424 242316 78492 242372
rect 78548 242316 78678 242372
rect 77678 242248 78678 242316
rect 77678 242192 77748 242248
rect 77804 242192 77872 242248
rect 77928 242192 77996 242248
rect 78052 242192 78120 242248
rect 78176 242192 78244 242248
rect 78300 242192 78368 242248
rect 78424 242192 78492 242248
rect 78548 242192 78678 242248
rect 77678 229102 78678 242192
rect 77678 229046 77900 229102
rect 77956 229046 78200 229102
rect 78256 229046 78500 229102
rect 78556 229046 78678 229102
rect 77678 222102 78678 229046
rect 77678 222046 77900 222102
rect 77956 222046 78200 222102
rect 78256 222046 78500 222102
rect 78556 222046 78678 222102
rect 77678 216372 78678 222046
rect 77678 216316 77748 216372
rect 77804 216316 77872 216372
rect 77928 216316 77996 216372
rect 78052 216316 78120 216372
rect 78176 216316 78244 216372
rect 78300 216316 78368 216372
rect 78424 216316 78492 216372
rect 78548 216316 78678 216372
rect 77678 216248 78678 216316
rect 77678 216192 77748 216248
rect 77804 216192 77872 216248
rect 77928 216192 77996 216248
rect 78052 216192 78120 216248
rect 78176 216192 78244 216248
rect 78300 216192 78368 216248
rect 78424 216192 78492 216248
rect 78548 216192 78678 216248
rect 77678 215102 78678 216192
rect 77678 215046 77900 215102
rect 77956 215046 78200 215102
rect 78256 215046 78500 215102
rect 78556 215046 78678 215102
rect 77678 207633 78678 215046
rect 77678 207577 77847 207633
rect 77903 207577 78147 207633
rect 78203 207577 78447 207633
rect 78503 207577 78678 207633
rect 77678 190372 78678 207577
rect 77678 190316 77748 190372
rect 77804 190316 77872 190372
rect 77928 190316 77996 190372
rect 78052 190316 78120 190372
rect 78176 190316 78244 190372
rect 78300 190316 78368 190372
rect 78424 190316 78492 190372
rect 78548 190316 78678 190372
rect 77678 190248 78678 190316
rect 77678 190192 77748 190248
rect 77804 190192 77872 190248
rect 77928 190192 77996 190248
rect 78052 190192 78120 190248
rect 78176 190192 78244 190248
rect 78300 190192 78368 190248
rect 78424 190192 78492 190248
rect 78548 190192 78678 190248
rect 77678 188102 78678 190192
rect 77678 188046 77900 188102
rect 77956 188046 78200 188102
rect 78256 188046 78500 188102
rect 78556 188046 78678 188102
rect 77678 181102 78678 188046
rect 77678 181046 77900 181102
rect 77956 181046 78200 181102
rect 78256 181046 78500 181102
rect 78556 181046 78678 181102
rect 77678 174102 78678 181046
rect 77678 174046 77900 174102
rect 77956 174046 78200 174102
rect 78256 174046 78500 174102
rect 78556 174046 78678 174102
rect 77678 164372 78678 174046
rect 77678 164316 77748 164372
rect 77804 164316 77872 164372
rect 77928 164316 77996 164372
rect 78052 164316 78120 164372
rect 78176 164316 78244 164372
rect 78300 164316 78368 164372
rect 78424 164316 78492 164372
rect 78548 164316 78678 164372
rect 77678 164248 78678 164316
rect 77678 164192 77748 164248
rect 77804 164192 77872 164248
rect 77928 164192 77996 164248
rect 78052 164192 78120 164248
rect 78176 164192 78244 164248
rect 78300 164192 78368 164248
rect 78424 164192 78492 164248
rect 78548 164192 78678 164248
rect 70000 146658 70200 146728
rect 70000 146602 70074 146658
rect 70130 146602 70200 146658
rect 70000 146534 70200 146602
rect 70000 146478 70074 146534
rect 70130 146478 70200 146534
rect 70000 146410 70200 146478
rect 70000 146354 70074 146410
rect 70130 146354 70200 146410
rect 70000 146286 70200 146354
rect 70000 146230 70074 146286
rect 70130 146230 70200 146286
rect 70000 146162 70200 146230
rect 70000 146106 70074 146162
rect 70130 146106 70200 146162
rect 70000 146038 70200 146106
rect 70000 145982 70074 146038
rect 70130 145982 70200 146038
rect 70000 145914 70200 145982
rect 70000 145858 70074 145914
rect 70130 145858 70200 145914
rect 70000 145790 70200 145858
rect 70000 145734 70074 145790
rect 70130 145734 70200 145790
rect 70000 145666 70200 145734
rect 70000 145610 70074 145666
rect 70130 145610 70200 145666
rect 70000 145542 70200 145610
rect 70000 145486 70074 145542
rect 70130 145486 70200 145542
rect 70000 145418 70200 145486
rect 70000 145362 70074 145418
rect 70130 145362 70200 145418
rect 70000 145294 70200 145362
rect 70000 145238 70074 145294
rect 70130 145238 70200 145294
rect 70000 145170 70200 145238
rect 70000 145114 70074 145170
rect 70130 145114 70200 145170
rect 70000 145046 70200 145114
rect 70000 144990 70074 145046
rect 70130 144990 70200 145046
rect 70000 144922 70200 144990
rect 70000 144866 70074 144922
rect 70130 144866 70200 144922
rect 70000 144828 70200 144866
rect 77678 146670 78678 164192
rect 77678 146614 77808 146670
rect 77864 146614 77932 146670
rect 77988 146614 78056 146670
rect 78112 146614 78180 146670
rect 78236 146614 78304 146670
rect 78360 146614 78428 146670
rect 78484 146614 78552 146670
rect 78608 146614 78678 146670
rect 77678 146546 78678 146614
rect 77678 146490 77808 146546
rect 77864 146490 77932 146546
rect 77988 146490 78056 146546
rect 78112 146490 78180 146546
rect 78236 146490 78304 146546
rect 78360 146490 78428 146546
rect 78484 146490 78552 146546
rect 78608 146490 78678 146546
rect 77678 146422 78678 146490
rect 77678 146366 77808 146422
rect 77864 146366 77932 146422
rect 77988 146366 78056 146422
rect 78112 146366 78180 146422
rect 78236 146366 78304 146422
rect 78360 146366 78428 146422
rect 78484 146366 78552 146422
rect 78608 146366 78678 146422
rect 77678 146298 78678 146366
rect 77678 146242 77808 146298
rect 77864 146242 77932 146298
rect 77988 146242 78056 146298
rect 78112 146242 78180 146298
rect 78236 146242 78304 146298
rect 78360 146242 78428 146298
rect 78484 146242 78552 146298
rect 78608 146242 78678 146298
rect 77678 146174 78678 146242
rect 77678 146118 77808 146174
rect 77864 146118 77932 146174
rect 77988 146118 78056 146174
rect 78112 146118 78180 146174
rect 78236 146118 78304 146174
rect 78360 146118 78428 146174
rect 78484 146118 78552 146174
rect 78608 146118 78678 146174
rect 77678 146050 78678 146118
rect 77678 145994 77808 146050
rect 77864 145994 77932 146050
rect 77988 145994 78056 146050
rect 78112 145994 78180 146050
rect 78236 145994 78304 146050
rect 78360 145994 78428 146050
rect 78484 145994 78552 146050
rect 78608 145994 78678 146050
rect 77678 145926 78678 145994
rect 77678 145870 77808 145926
rect 77864 145870 77932 145926
rect 77988 145870 78056 145926
rect 78112 145870 78180 145926
rect 78236 145870 78304 145926
rect 78360 145870 78428 145926
rect 78484 145870 78552 145926
rect 78608 145870 78678 145926
rect 77678 145802 78678 145870
rect 77678 145746 77808 145802
rect 77864 145746 77932 145802
rect 77988 145746 78056 145802
rect 78112 145746 78180 145802
rect 78236 145746 78304 145802
rect 78360 145746 78428 145802
rect 78484 145746 78552 145802
rect 78608 145746 78678 145802
rect 77678 145678 78678 145746
rect 77678 145622 77808 145678
rect 77864 145622 77932 145678
rect 77988 145622 78056 145678
rect 78112 145622 78180 145678
rect 78236 145622 78304 145678
rect 78360 145622 78428 145678
rect 78484 145622 78552 145678
rect 78608 145622 78678 145678
rect 77678 145554 78678 145622
rect 77678 145498 77808 145554
rect 77864 145498 77932 145554
rect 77988 145498 78056 145554
rect 78112 145498 78180 145554
rect 78236 145498 78304 145554
rect 78360 145498 78428 145554
rect 78484 145498 78552 145554
rect 78608 145498 78678 145554
rect 77678 145430 78678 145498
rect 77678 145374 77808 145430
rect 77864 145374 77932 145430
rect 77988 145374 78056 145430
rect 78112 145374 78180 145430
rect 78236 145374 78304 145430
rect 78360 145374 78428 145430
rect 78484 145374 78552 145430
rect 78608 145374 78678 145430
rect 77678 145306 78678 145374
rect 77678 145250 77808 145306
rect 77864 145250 77932 145306
rect 77988 145250 78056 145306
rect 78112 145250 78180 145306
rect 78236 145250 78304 145306
rect 78360 145250 78428 145306
rect 78484 145250 78552 145306
rect 78608 145250 78678 145306
rect 77678 145182 78678 145250
rect 77678 145126 77808 145182
rect 77864 145126 77932 145182
rect 77988 145126 78056 145182
rect 78112 145126 78180 145182
rect 78236 145126 78304 145182
rect 78360 145126 78428 145182
rect 78484 145126 78552 145182
rect 78608 145126 78678 145182
rect 77678 145058 78678 145126
rect 77678 145002 77808 145058
rect 77864 145002 77932 145058
rect 77988 145002 78056 145058
rect 78112 145002 78180 145058
rect 78236 145002 78304 145058
rect 78360 145002 78428 145058
rect 78484 145002 78552 145058
rect 78608 145002 78678 145058
rect 77678 144934 78678 145002
rect 77678 144878 77808 144934
rect 77864 144878 77932 144934
rect 77988 144878 78056 144934
rect 78112 144878 78180 144934
rect 78236 144878 78304 144934
rect 78360 144878 78428 144934
rect 78484 144878 78552 144934
rect 78608 144878 78678 144934
rect 70000 144184 70200 144248
rect 70000 144128 70074 144184
rect 70130 144128 70200 144184
rect 70000 144060 70200 144128
rect 70000 144004 70074 144060
rect 70130 144004 70200 144060
rect 70000 143936 70200 144004
rect 70000 143880 70074 143936
rect 70130 143880 70200 143936
rect 70000 143812 70200 143880
rect 70000 143756 70074 143812
rect 70130 143756 70200 143812
rect 70000 143688 70200 143756
rect 70000 143632 70074 143688
rect 70130 143632 70200 143688
rect 70000 143564 70200 143632
rect 70000 143508 70074 143564
rect 70130 143508 70200 143564
rect 70000 143440 70200 143508
rect 70000 143384 70074 143440
rect 70130 143384 70200 143440
rect 70000 143316 70200 143384
rect 70000 143260 70074 143316
rect 70130 143260 70200 143316
rect 70000 143192 70200 143260
rect 70000 143136 70074 143192
rect 70130 143136 70200 143192
rect 70000 143068 70200 143136
rect 70000 143012 70074 143068
rect 70130 143012 70200 143068
rect 70000 142944 70200 143012
rect 70000 142888 70074 142944
rect 70130 142888 70200 142944
rect 70000 142820 70200 142888
rect 70000 142764 70074 142820
rect 70130 142764 70200 142820
rect 70000 142696 70200 142764
rect 70000 142640 70074 142696
rect 70130 142640 70200 142696
rect 70000 142572 70200 142640
rect 70000 142516 70074 142572
rect 70130 142516 70200 142572
rect 70000 142448 70200 142516
rect 70000 142392 70074 142448
rect 70130 142392 70200 142448
rect 70000 142324 70200 142392
rect 70000 142268 70074 142324
rect 70130 142268 70200 142324
rect 70000 142198 70200 142268
rect 77678 144190 78678 144878
rect 77678 144134 77808 144190
rect 77864 144134 77932 144190
rect 77988 144134 78056 144190
rect 78112 144134 78180 144190
rect 78236 144134 78304 144190
rect 78360 144134 78428 144190
rect 78484 144134 78552 144190
rect 78608 144134 78678 144190
rect 77678 144066 78678 144134
rect 77678 144010 77808 144066
rect 77864 144010 77932 144066
rect 77988 144010 78056 144066
rect 78112 144010 78180 144066
rect 78236 144010 78304 144066
rect 78360 144010 78428 144066
rect 78484 144010 78552 144066
rect 78608 144010 78678 144066
rect 77678 143942 78678 144010
rect 77678 143886 77808 143942
rect 77864 143886 77932 143942
rect 77988 143886 78056 143942
rect 78112 143886 78180 143942
rect 78236 143886 78304 143942
rect 78360 143886 78428 143942
rect 78484 143886 78552 143942
rect 78608 143886 78678 143942
rect 77678 143818 78678 143886
rect 77678 143762 77808 143818
rect 77864 143762 77932 143818
rect 77988 143762 78056 143818
rect 78112 143762 78180 143818
rect 78236 143762 78304 143818
rect 78360 143762 78428 143818
rect 78484 143762 78552 143818
rect 78608 143762 78678 143818
rect 77678 143694 78678 143762
rect 77678 143638 77808 143694
rect 77864 143638 77932 143694
rect 77988 143638 78056 143694
rect 78112 143638 78180 143694
rect 78236 143638 78304 143694
rect 78360 143638 78428 143694
rect 78484 143638 78552 143694
rect 78608 143638 78678 143694
rect 77678 143570 78678 143638
rect 77678 143514 77808 143570
rect 77864 143514 77932 143570
rect 77988 143514 78056 143570
rect 78112 143514 78180 143570
rect 78236 143514 78304 143570
rect 78360 143514 78428 143570
rect 78484 143514 78552 143570
rect 78608 143514 78678 143570
rect 77678 143446 78678 143514
rect 77678 143390 77808 143446
rect 77864 143390 77932 143446
rect 77988 143390 78056 143446
rect 78112 143390 78180 143446
rect 78236 143390 78304 143446
rect 78360 143390 78428 143446
rect 78484 143390 78552 143446
rect 78608 143390 78678 143446
rect 77678 143322 78678 143390
rect 77678 143266 77808 143322
rect 77864 143266 77932 143322
rect 77988 143266 78056 143322
rect 78112 143266 78180 143322
rect 78236 143266 78304 143322
rect 78360 143266 78428 143322
rect 78484 143266 78552 143322
rect 78608 143266 78678 143322
rect 77678 143198 78678 143266
rect 77678 143142 77808 143198
rect 77864 143142 77932 143198
rect 77988 143142 78056 143198
rect 78112 143142 78180 143198
rect 78236 143142 78304 143198
rect 78360 143142 78428 143198
rect 78484 143142 78552 143198
rect 78608 143142 78678 143198
rect 77678 143074 78678 143142
rect 77678 143018 77808 143074
rect 77864 143018 77932 143074
rect 77988 143018 78056 143074
rect 78112 143018 78180 143074
rect 78236 143018 78304 143074
rect 78360 143018 78428 143074
rect 78484 143018 78552 143074
rect 78608 143018 78678 143074
rect 77678 142950 78678 143018
rect 77678 142894 77808 142950
rect 77864 142894 77932 142950
rect 77988 142894 78056 142950
rect 78112 142894 78180 142950
rect 78236 142894 78304 142950
rect 78360 142894 78428 142950
rect 78484 142894 78552 142950
rect 78608 142894 78678 142950
rect 77678 142826 78678 142894
rect 77678 142770 77808 142826
rect 77864 142770 77932 142826
rect 77988 142770 78056 142826
rect 78112 142770 78180 142826
rect 78236 142770 78304 142826
rect 78360 142770 78428 142826
rect 78484 142770 78552 142826
rect 78608 142770 78678 142826
rect 77678 142702 78678 142770
rect 77678 142646 77808 142702
rect 77864 142646 77932 142702
rect 77988 142646 78056 142702
rect 78112 142646 78180 142702
rect 78236 142646 78304 142702
rect 78360 142646 78428 142702
rect 78484 142646 78552 142702
rect 78608 142646 78678 142702
rect 77678 142578 78678 142646
rect 77678 142522 77808 142578
rect 77864 142522 77932 142578
rect 77988 142522 78056 142578
rect 78112 142522 78180 142578
rect 78236 142522 78304 142578
rect 78360 142522 78428 142578
rect 78484 142522 78552 142578
rect 78608 142522 78678 142578
rect 77678 142454 78678 142522
rect 77678 142398 77808 142454
rect 77864 142398 77932 142454
rect 77988 142398 78056 142454
rect 78112 142398 78180 142454
rect 78236 142398 78304 142454
rect 78360 142398 78428 142454
rect 78484 142398 78552 142454
rect 78608 142398 78678 142454
rect 77678 142330 78678 142398
rect 77678 142274 77808 142330
rect 77864 142274 77932 142330
rect 77988 142274 78056 142330
rect 78112 142274 78180 142330
rect 78236 142274 78304 142330
rect 78360 142274 78428 142330
rect 78484 142274 78552 142330
rect 78608 142274 78678 142330
rect 70000 141814 70200 141878
rect 70000 141758 70074 141814
rect 70130 141758 70200 141814
rect 70000 141690 70200 141758
rect 70000 141634 70074 141690
rect 70130 141634 70200 141690
rect 70000 141566 70200 141634
rect 70000 141510 70074 141566
rect 70130 141510 70200 141566
rect 70000 141442 70200 141510
rect 70000 141386 70074 141442
rect 70130 141386 70200 141442
rect 70000 141318 70200 141386
rect 70000 141262 70074 141318
rect 70130 141262 70200 141318
rect 70000 141194 70200 141262
rect 70000 141138 70074 141194
rect 70130 141138 70200 141194
rect 70000 141070 70200 141138
rect 70000 141014 70074 141070
rect 70130 141014 70200 141070
rect 70000 140946 70200 141014
rect 70000 140890 70074 140946
rect 70130 140890 70200 140946
rect 70000 140822 70200 140890
rect 70000 140766 70074 140822
rect 70130 140766 70200 140822
rect 70000 140698 70200 140766
rect 70000 140642 70074 140698
rect 70130 140642 70200 140698
rect 70000 140574 70200 140642
rect 70000 140518 70074 140574
rect 70130 140518 70200 140574
rect 70000 140450 70200 140518
rect 70000 140394 70074 140450
rect 70130 140394 70200 140450
rect 70000 140326 70200 140394
rect 70000 140270 70074 140326
rect 70130 140270 70200 140326
rect 70000 140202 70200 140270
rect 70000 140146 70074 140202
rect 70130 140146 70200 140202
rect 70000 140078 70200 140146
rect 70000 140022 70074 140078
rect 70130 140022 70200 140078
rect 70000 139954 70200 140022
rect 70000 139898 70074 139954
rect 70130 139898 70200 139954
rect 70000 139828 70200 139898
rect 77678 141820 78678 142274
rect 77678 141764 77808 141820
rect 77864 141764 77932 141820
rect 77988 141764 78056 141820
rect 78112 141764 78180 141820
rect 78236 141764 78304 141820
rect 78360 141764 78428 141820
rect 78484 141764 78552 141820
rect 78608 141764 78678 141820
rect 77678 141696 78678 141764
rect 77678 141640 77808 141696
rect 77864 141640 77932 141696
rect 77988 141640 78056 141696
rect 78112 141640 78180 141696
rect 78236 141640 78304 141696
rect 78360 141640 78428 141696
rect 78484 141640 78552 141696
rect 78608 141640 78678 141696
rect 77678 141572 78678 141640
rect 77678 141516 77808 141572
rect 77864 141516 77932 141572
rect 77988 141516 78056 141572
rect 78112 141516 78180 141572
rect 78236 141516 78304 141572
rect 78360 141516 78428 141572
rect 78484 141516 78552 141572
rect 78608 141516 78678 141572
rect 77678 141448 78678 141516
rect 77678 141392 77808 141448
rect 77864 141392 77932 141448
rect 77988 141392 78056 141448
rect 78112 141392 78180 141448
rect 78236 141392 78304 141448
rect 78360 141392 78428 141448
rect 78484 141392 78552 141448
rect 78608 141392 78678 141448
rect 77678 141324 78678 141392
rect 77678 141268 77808 141324
rect 77864 141268 77932 141324
rect 77988 141268 78056 141324
rect 78112 141268 78180 141324
rect 78236 141268 78304 141324
rect 78360 141268 78428 141324
rect 78484 141268 78552 141324
rect 78608 141268 78678 141324
rect 77678 141200 78678 141268
rect 77678 141144 77808 141200
rect 77864 141144 77932 141200
rect 77988 141144 78056 141200
rect 78112 141144 78180 141200
rect 78236 141144 78304 141200
rect 78360 141144 78428 141200
rect 78484 141144 78552 141200
rect 78608 141144 78678 141200
rect 77678 141076 78678 141144
rect 77678 141020 77808 141076
rect 77864 141020 77932 141076
rect 77988 141020 78056 141076
rect 78112 141020 78180 141076
rect 78236 141020 78304 141076
rect 78360 141020 78428 141076
rect 78484 141020 78552 141076
rect 78608 141020 78678 141076
rect 77678 140952 78678 141020
rect 77678 140896 77808 140952
rect 77864 140896 77932 140952
rect 77988 140896 78056 140952
rect 78112 140896 78180 140952
rect 78236 140896 78304 140952
rect 78360 140896 78428 140952
rect 78484 140896 78552 140952
rect 78608 140896 78678 140952
rect 77678 140828 78678 140896
rect 77678 140772 77808 140828
rect 77864 140772 77932 140828
rect 77988 140772 78056 140828
rect 78112 140772 78180 140828
rect 78236 140772 78304 140828
rect 78360 140772 78428 140828
rect 78484 140772 78552 140828
rect 78608 140772 78678 140828
rect 77678 140704 78678 140772
rect 77678 140648 77808 140704
rect 77864 140648 77932 140704
rect 77988 140648 78056 140704
rect 78112 140648 78180 140704
rect 78236 140648 78304 140704
rect 78360 140648 78428 140704
rect 78484 140648 78552 140704
rect 78608 140648 78678 140704
rect 77678 140580 78678 140648
rect 77678 140524 77808 140580
rect 77864 140524 77932 140580
rect 77988 140524 78056 140580
rect 78112 140524 78180 140580
rect 78236 140524 78304 140580
rect 78360 140524 78428 140580
rect 78484 140524 78552 140580
rect 78608 140524 78678 140580
rect 77678 140456 78678 140524
rect 77678 140400 77808 140456
rect 77864 140400 77932 140456
rect 77988 140400 78056 140456
rect 78112 140400 78180 140456
rect 78236 140400 78304 140456
rect 78360 140400 78428 140456
rect 78484 140400 78552 140456
rect 78608 140400 78678 140456
rect 77678 140332 78678 140400
rect 77678 140276 77808 140332
rect 77864 140276 77932 140332
rect 77988 140276 78056 140332
rect 78112 140276 78180 140332
rect 78236 140276 78304 140332
rect 78360 140276 78428 140332
rect 78484 140276 78552 140332
rect 78608 140276 78678 140332
rect 77678 140208 78678 140276
rect 77678 140152 77808 140208
rect 77864 140152 77932 140208
rect 77988 140152 78056 140208
rect 78112 140152 78180 140208
rect 78236 140152 78304 140208
rect 78360 140152 78428 140208
rect 78484 140152 78552 140208
rect 78608 140152 78678 140208
rect 77678 140084 78678 140152
rect 77678 140028 77808 140084
rect 77864 140028 77932 140084
rect 77988 140028 78056 140084
rect 78112 140028 78180 140084
rect 78236 140028 78304 140084
rect 78360 140028 78428 140084
rect 78484 140028 78552 140084
rect 78608 140028 78678 140084
rect 77678 139960 78678 140028
rect 77678 139904 77808 139960
rect 77864 139904 77932 139960
rect 77988 139904 78056 139960
rect 78112 139904 78180 139960
rect 78236 139904 78304 139960
rect 78360 139904 78428 139960
rect 78484 139904 78552 139960
rect 78608 139904 78678 139960
rect 70000 139108 70200 139172
rect 70000 139052 70074 139108
rect 70130 139052 70200 139108
rect 70000 138984 70200 139052
rect 70000 138928 70074 138984
rect 70130 138928 70200 138984
rect 70000 138860 70200 138928
rect 70000 138804 70074 138860
rect 70130 138804 70200 138860
rect 70000 138736 70200 138804
rect 70000 138680 70074 138736
rect 70130 138680 70200 138736
rect 70000 138612 70200 138680
rect 70000 138556 70074 138612
rect 70130 138556 70200 138612
rect 70000 138488 70200 138556
rect 70000 138432 70074 138488
rect 70130 138432 70200 138488
rect 70000 138364 70200 138432
rect 70000 138308 70074 138364
rect 70130 138308 70200 138364
rect 70000 138240 70200 138308
rect 70000 138184 70074 138240
rect 70130 138184 70200 138240
rect 70000 138116 70200 138184
rect 70000 138060 70074 138116
rect 70130 138060 70200 138116
rect 70000 137992 70200 138060
rect 70000 137936 70074 137992
rect 70130 137936 70200 137992
rect 70000 137868 70200 137936
rect 70000 137812 70074 137868
rect 70130 137812 70200 137868
rect 70000 137744 70200 137812
rect 70000 137688 70074 137744
rect 70130 137688 70200 137744
rect 70000 137620 70200 137688
rect 70000 137564 70074 137620
rect 70130 137564 70200 137620
rect 70000 137496 70200 137564
rect 70000 137440 70074 137496
rect 70130 137440 70200 137496
rect 70000 137372 70200 137440
rect 70000 137316 70074 137372
rect 70130 137316 70200 137372
rect 70000 137248 70200 137316
rect 70000 137192 70074 137248
rect 70130 137192 70200 137248
rect 70000 137122 70200 137192
rect 77678 139114 78678 139904
rect 77678 139058 77808 139114
rect 77864 139058 77932 139114
rect 77988 139058 78056 139114
rect 78112 139058 78180 139114
rect 78236 139058 78304 139114
rect 78360 139058 78428 139114
rect 78484 139058 78552 139114
rect 78608 139058 78678 139114
rect 77678 138990 78678 139058
rect 77678 138934 77808 138990
rect 77864 138934 77932 138990
rect 77988 138934 78056 138990
rect 78112 138934 78180 138990
rect 78236 138934 78304 138990
rect 78360 138934 78428 138990
rect 78484 138934 78552 138990
rect 78608 138934 78678 138990
rect 77678 138866 78678 138934
rect 77678 138810 77808 138866
rect 77864 138810 77932 138866
rect 77988 138810 78056 138866
rect 78112 138810 78180 138866
rect 78236 138810 78304 138866
rect 78360 138810 78428 138866
rect 78484 138810 78552 138866
rect 78608 138810 78678 138866
rect 77678 138742 78678 138810
rect 77678 138686 77808 138742
rect 77864 138686 77932 138742
rect 77988 138686 78056 138742
rect 78112 138686 78180 138742
rect 78236 138686 78304 138742
rect 78360 138686 78428 138742
rect 78484 138686 78552 138742
rect 78608 138686 78678 138742
rect 77678 138618 78678 138686
rect 77678 138562 77808 138618
rect 77864 138562 77932 138618
rect 77988 138562 78056 138618
rect 78112 138562 78180 138618
rect 78236 138562 78304 138618
rect 78360 138562 78428 138618
rect 78484 138562 78552 138618
rect 78608 138562 78678 138618
rect 77678 138494 78678 138562
rect 77678 138438 77808 138494
rect 77864 138438 77932 138494
rect 77988 138438 78056 138494
rect 78112 138438 78180 138494
rect 78236 138438 78304 138494
rect 78360 138438 78428 138494
rect 78484 138438 78552 138494
rect 78608 138438 78678 138494
rect 77678 138370 78678 138438
rect 77678 138314 77808 138370
rect 77864 138314 77932 138370
rect 77988 138314 78056 138370
rect 78112 138314 78180 138370
rect 78236 138314 78304 138370
rect 78360 138314 78428 138370
rect 78484 138314 78552 138370
rect 78608 138314 78678 138370
rect 77678 138246 78678 138314
rect 77678 138190 77808 138246
rect 77864 138190 77932 138246
rect 77988 138190 78056 138246
rect 78112 138190 78180 138246
rect 78236 138190 78304 138246
rect 78360 138190 78428 138246
rect 78484 138190 78552 138246
rect 78608 138190 78678 138246
rect 77678 138122 78678 138190
rect 77678 138066 77808 138122
rect 77864 138066 77932 138122
rect 77988 138066 78056 138122
rect 78112 138066 78180 138122
rect 78236 138066 78304 138122
rect 78360 138066 78428 138122
rect 78484 138066 78552 138122
rect 78608 138066 78678 138122
rect 77678 137998 78678 138066
rect 77678 137942 77808 137998
rect 77864 137942 77932 137998
rect 77988 137942 78056 137998
rect 78112 137942 78180 137998
rect 78236 137942 78304 137998
rect 78360 137942 78428 137998
rect 78484 137942 78552 137998
rect 78608 137942 78678 137998
rect 77678 137874 78678 137942
rect 77678 137818 77808 137874
rect 77864 137818 77932 137874
rect 77988 137818 78056 137874
rect 78112 137818 78180 137874
rect 78236 137818 78304 137874
rect 78360 137818 78428 137874
rect 78484 137818 78552 137874
rect 78608 137818 78678 137874
rect 77678 137750 78678 137818
rect 77678 137694 77808 137750
rect 77864 137694 77932 137750
rect 77988 137694 78056 137750
rect 78112 137694 78180 137750
rect 78236 137694 78304 137750
rect 78360 137694 78428 137750
rect 78484 137694 78552 137750
rect 78608 137694 78678 137750
rect 77678 137626 78678 137694
rect 77678 137570 77808 137626
rect 77864 137570 77932 137626
rect 77988 137570 78056 137626
rect 78112 137570 78180 137626
rect 78236 137570 78304 137626
rect 78360 137570 78428 137626
rect 78484 137570 78552 137626
rect 78608 137570 78678 137626
rect 77678 137502 78678 137570
rect 77678 137446 77808 137502
rect 77864 137446 77932 137502
rect 77988 137446 78056 137502
rect 78112 137446 78180 137502
rect 78236 137446 78304 137502
rect 78360 137446 78428 137502
rect 78484 137446 78552 137502
rect 78608 137446 78678 137502
rect 77678 137378 78678 137446
rect 77678 137322 77808 137378
rect 77864 137322 77932 137378
rect 77988 137322 78056 137378
rect 78112 137322 78180 137378
rect 78236 137322 78304 137378
rect 78360 137322 78428 137378
rect 78484 137322 78552 137378
rect 78608 137322 78678 137378
rect 77678 137254 78678 137322
rect 77678 137198 77808 137254
rect 77864 137198 77932 137254
rect 77988 137198 78056 137254
rect 78112 137198 78180 137254
rect 78236 137198 78304 137254
rect 78360 137198 78428 137254
rect 78484 137198 78552 137254
rect 78608 137198 78678 137254
rect 70000 136738 70200 136802
rect 70000 136682 70074 136738
rect 70130 136682 70200 136738
rect 70000 136614 70200 136682
rect 70000 136558 70074 136614
rect 70130 136558 70200 136614
rect 70000 136490 70200 136558
rect 70000 136434 70074 136490
rect 70130 136434 70200 136490
rect 70000 136366 70200 136434
rect 70000 136310 70074 136366
rect 70130 136310 70200 136366
rect 70000 136242 70200 136310
rect 70000 136186 70074 136242
rect 70130 136186 70200 136242
rect 70000 136118 70200 136186
rect 70000 136062 70074 136118
rect 70130 136062 70200 136118
rect 70000 135994 70200 136062
rect 70000 135938 70074 135994
rect 70130 135938 70200 135994
rect 70000 135870 70200 135938
rect 70000 135814 70074 135870
rect 70130 135814 70200 135870
rect 70000 135746 70200 135814
rect 70000 135690 70074 135746
rect 70130 135690 70200 135746
rect 70000 135622 70200 135690
rect 70000 135566 70074 135622
rect 70130 135566 70200 135622
rect 70000 135498 70200 135566
rect 70000 135442 70074 135498
rect 70130 135442 70200 135498
rect 70000 135374 70200 135442
rect 70000 135318 70074 135374
rect 70130 135318 70200 135374
rect 70000 135250 70200 135318
rect 70000 135194 70074 135250
rect 70130 135194 70200 135250
rect 70000 135126 70200 135194
rect 70000 135070 70074 135126
rect 70130 135070 70200 135126
rect 70000 135002 70200 135070
rect 70000 134946 70074 135002
rect 70130 134946 70200 135002
rect 70000 134878 70200 134946
rect 70000 134822 70074 134878
rect 70130 134822 70200 134878
rect 70000 134752 70200 134822
rect 77678 136744 78678 137198
rect 77678 136688 77808 136744
rect 77864 136688 77932 136744
rect 77988 136688 78056 136744
rect 78112 136688 78180 136744
rect 78236 136688 78304 136744
rect 78360 136688 78428 136744
rect 78484 136688 78552 136744
rect 78608 136688 78678 136744
rect 77678 136620 78678 136688
rect 77678 136564 77808 136620
rect 77864 136564 77932 136620
rect 77988 136564 78056 136620
rect 78112 136564 78180 136620
rect 78236 136564 78304 136620
rect 78360 136564 78428 136620
rect 78484 136564 78552 136620
rect 78608 136564 78678 136620
rect 77678 136496 78678 136564
rect 77678 136440 77808 136496
rect 77864 136440 77932 136496
rect 77988 136440 78056 136496
rect 78112 136440 78180 136496
rect 78236 136440 78304 136496
rect 78360 136440 78428 136496
rect 78484 136440 78552 136496
rect 78608 136440 78678 136496
rect 77678 136372 78678 136440
rect 77678 136316 77808 136372
rect 77864 136316 77932 136372
rect 77988 136316 78056 136372
rect 78112 136316 78180 136372
rect 78236 136316 78304 136372
rect 78360 136316 78428 136372
rect 78484 136316 78552 136372
rect 78608 136316 78678 136372
rect 77678 136248 78678 136316
rect 77678 136192 77808 136248
rect 77864 136192 77932 136248
rect 77988 136192 78056 136248
rect 78112 136192 78180 136248
rect 78236 136192 78304 136248
rect 78360 136192 78428 136248
rect 78484 136192 78552 136248
rect 78608 136192 78678 136248
rect 77678 136124 78678 136192
rect 77678 136068 77808 136124
rect 77864 136068 77932 136124
rect 77988 136068 78056 136124
rect 78112 136068 78180 136124
rect 78236 136068 78304 136124
rect 78360 136068 78428 136124
rect 78484 136068 78552 136124
rect 78608 136068 78678 136124
rect 77678 136000 78678 136068
rect 77678 135944 77808 136000
rect 77864 135944 77932 136000
rect 77988 135944 78056 136000
rect 78112 135944 78180 136000
rect 78236 135944 78304 136000
rect 78360 135944 78428 136000
rect 78484 135944 78552 136000
rect 78608 135944 78678 136000
rect 77678 135876 78678 135944
rect 77678 135820 77808 135876
rect 77864 135820 77932 135876
rect 77988 135820 78056 135876
rect 78112 135820 78180 135876
rect 78236 135820 78304 135876
rect 78360 135820 78428 135876
rect 78484 135820 78552 135876
rect 78608 135820 78678 135876
rect 77678 135752 78678 135820
rect 77678 135696 77808 135752
rect 77864 135696 77932 135752
rect 77988 135696 78056 135752
rect 78112 135696 78180 135752
rect 78236 135696 78304 135752
rect 78360 135696 78428 135752
rect 78484 135696 78552 135752
rect 78608 135696 78678 135752
rect 77678 135628 78678 135696
rect 77678 135572 77808 135628
rect 77864 135572 77932 135628
rect 77988 135572 78056 135628
rect 78112 135572 78180 135628
rect 78236 135572 78304 135628
rect 78360 135572 78428 135628
rect 78484 135572 78552 135628
rect 78608 135572 78678 135628
rect 77678 135504 78678 135572
rect 77678 135448 77808 135504
rect 77864 135448 77932 135504
rect 77988 135448 78056 135504
rect 78112 135448 78180 135504
rect 78236 135448 78304 135504
rect 78360 135448 78428 135504
rect 78484 135448 78552 135504
rect 78608 135448 78678 135504
rect 77678 135380 78678 135448
rect 77678 135324 77808 135380
rect 77864 135324 77932 135380
rect 77988 135324 78056 135380
rect 78112 135324 78180 135380
rect 78236 135324 78304 135380
rect 78360 135324 78428 135380
rect 78484 135324 78552 135380
rect 78608 135324 78678 135380
rect 77678 135256 78678 135324
rect 77678 135200 77808 135256
rect 77864 135200 77932 135256
rect 77988 135200 78056 135256
rect 78112 135200 78180 135256
rect 78236 135200 78304 135256
rect 78360 135200 78428 135256
rect 78484 135200 78552 135256
rect 78608 135200 78678 135256
rect 77678 135132 78678 135200
rect 77678 135076 77808 135132
rect 77864 135076 77932 135132
rect 77988 135076 78056 135132
rect 78112 135076 78180 135132
rect 78236 135076 78304 135132
rect 78360 135076 78428 135132
rect 78484 135076 78552 135132
rect 78608 135076 78678 135132
rect 77678 135008 78678 135076
rect 77678 134952 77808 135008
rect 77864 134952 77932 135008
rect 77988 134952 78056 135008
rect 78112 134952 78180 135008
rect 78236 134952 78304 135008
rect 78360 134952 78428 135008
rect 78484 134952 78552 135008
rect 78608 134952 78678 135008
rect 77678 134884 78678 134952
rect 77678 134828 77808 134884
rect 77864 134828 77932 134884
rect 77988 134828 78056 134884
rect 78112 134828 78180 134884
rect 78236 134828 78304 134884
rect 78360 134828 78428 134884
rect 78484 134828 78552 134884
rect 78608 134828 78678 134884
rect 70000 134134 70200 134172
rect 70000 134078 70074 134134
rect 70130 134078 70200 134134
rect 70000 134010 70200 134078
rect 70000 133954 70074 134010
rect 70130 133954 70200 134010
rect 70000 133886 70200 133954
rect 70000 133830 70074 133886
rect 70130 133830 70200 133886
rect 70000 133762 70200 133830
rect 70000 133706 70074 133762
rect 70130 133706 70200 133762
rect 70000 133638 70200 133706
rect 70000 133582 70074 133638
rect 70130 133582 70200 133638
rect 70000 133514 70200 133582
rect 70000 133458 70074 133514
rect 70130 133458 70200 133514
rect 70000 133390 70200 133458
rect 70000 133334 70074 133390
rect 70130 133334 70200 133390
rect 70000 133266 70200 133334
rect 70000 133210 70074 133266
rect 70130 133210 70200 133266
rect 70000 133142 70200 133210
rect 70000 133086 70074 133142
rect 70130 133086 70200 133142
rect 70000 133018 70200 133086
rect 70000 132962 70074 133018
rect 70130 132962 70200 133018
rect 70000 132894 70200 132962
rect 70000 132838 70074 132894
rect 70130 132838 70200 132894
rect 70000 132770 70200 132838
rect 70000 132714 70074 132770
rect 70130 132714 70200 132770
rect 70000 132646 70200 132714
rect 70000 132590 70074 132646
rect 70130 132590 70200 132646
rect 70000 132522 70200 132590
rect 70000 132466 70074 132522
rect 70130 132466 70200 132522
rect 70000 132398 70200 132466
rect 70000 132342 70074 132398
rect 70130 132342 70200 132398
rect 70000 132272 70200 132342
rect 77678 134140 78678 134828
rect 77678 134084 77808 134140
rect 77864 134084 77932 134140
rect 77988 134084 78056 134140
rect 78112 134084 78180 134140
rect 78236 134084 78304 134140
rect 78360 134084 78428 134140
rect 78484 134084 78552 134140
rect 78608 134084 78678 134140
rect 77678 134016 78678 134084
rect 77678 133960 77808 134016
rect 77864 133960 77932 134016
rect 77988 133960 78056 134016
rect 78112 133960 78180 134016
rect 78236 133960 78304 134016
rect 78360 133960 78428 134016
rect 78484 133960 78552 134016
rect 78608 133960 78678 134016
rect 77678 133892 78678 133960
rect 77678 133836 77808 133892
rect 77864 133836 77932 133892
rect 77988 133836 78056 133892
rect 78112 133836 78180 133892
rect 78236 133836 78304 133892
rect 78360 133836 78428 133892
rect 78484 133836 78552 133892
rect 78608 133836 78678 133892
rect 77678 133768 78678 133836
rect 77678 133712 77808 133768
rect 77864 133712 77932 133768
rect 77988 133712 78056 133768
rect 78112 133712 78180 133768
rect 78236 133712 78304 133768
rect 78360 133712 78428 133768
rect 78484 133712 78552 133768
rect 78608 133712 78678 133768
rect 77678 133644 78678 133712
rect 77678 133588 77808 133644
rect 77864 133588 77932 133644
rect 77988 133588 78056 133644
rect 78112 133588 78180 133644
rect 78236 133588 78304 133644
rect 78360 133588 78428 133644
rect 78484 133588 78552 133644
rect 78608 133588 78678 133644
rect 77678 133520 78678 133588
rect 77678 133464 77808 133520
rect 77864 133464 77932 133520
rect 77988 133464 78056 133520
rect 78112 133464 78180 133520
rect 78236 133464 78304 133520
rect 78360 133464 78428 133520
rect 78484 133464 78552 133520
rect 78608 133464 78678 133520
rect 77678 133396 78678 133464
rect 77678 133340 77808 133396
rect 77864 133340 77932 133396
rect 77988 133340 78056 133396
rect 78112 133340 78180 133396
rect 78236 133340 78304 133396
rect 78360 133340 78428 133396
rect 78484 133340 78552 133396
rect 78608 133340 78678 133396
rect 77678 133272 78678 133340
rect 77678 133216 77808 133272
rect 77864 133216 77932 133272
rect 77988 133216 78056 133272
rect 78112 133216 78180 133272
rect 78236 133216 78304 133272
rect 78360 133216 78428 133272
rect 78484 133216 78552 133272
rect 78608 133216 78678 133272
rect 77678 133148 78678 133216
rect 77678 133092 77808 133148
rect 77864 133092 77932 133148
rect 77988 133092 78056 133148
rect 78112 133092 78180 133148
rect 78236 133092 78304 133148
rect 78360 133092 78428 133148
rect 78484 133092 78552 133148
rect 78608 133092 78678 133148
rect 77678 133024 78678 133092
rect 77678 132968 77808 133024
rect 77864 132968 77932 133024
rect 77988 132968 78056 133024
rect 78112 132968 78180 133024
rect 78236 132968 78304 133024
rect 78360 132968 78428 133024
rect 78484 132968 78552 133024
rect 78608 132968 78678 133024
rect 77678 132900 78678 132968
rect 77678 132844 77808 132900
rect 77864 132844 77932 132900
rect 77988 132844 78056 132900
rect 78112 132844 78180 132900
rect 78236 132844 78304 132900
rect 78360 132844 78428 132900
rect 78484 132844 78552 132900
rect 78608 132844 78678 132900
rect 77678 132776 78678 132844
rect 77678 132720 77808 132776
rect 77864 132720 77932 132776
rect 77988 132720 78056 132776
rect 78112 132720 78180 132776
rect 78236 132720 78304 132776
rect 78360 132720 78428 132776
rect 78484 132720 78552 132776
rect 78608 132720 78678 132776
rect 77678 132652 78678 132720
rect 77678 132596 77808 132652
rect 77864 132596 77932 132652
rect 77988 132596 78056 132652
rect 78112 132596 78180 132652
rect 78236 132596 78304 132652
rect 78360 132596 78428 132652
rect 78484 132596 78552 132652
rect 78608 132596 78678 132652
rect 77678 132528 78678 132596
rect 77678 132472 77808 132528
rect 77864 132472 77932 132528
rect 77988 132472 78056 132528
rect 78112 132472 78180 132528
rect 78236 132472 78304 132528
rect 78360 132472 78428 132528
rect 78484 132472 78552 132528
rect 78608 132472 78678 132528
rect 77678 132404 78678 132472
rect 77678 132348 77808 132404
rect 77864 132348 77932 132404
rect 77988 132348 78056 132404
rect 78112 132348 78180 132404
rect 78236 132348 78304 132404
rect 78360 132348 78428 132404
rect 78484 132348 78552 132404
rect 78608 132348 78678 132404
rect 77678 112372 78678 132348
rect 77678 112316 77748 112372
rect 77804 112316 77872 112372
rect 77928 112316 77996 112372
rect 78052 112316 78120 112372
rect 78176 112316 78244 112372
rect 78300 112316 78368 112372
rect 78424 112316 78492 112372
rect 78548 112316 78678 112372
rect 77678 112248 78678 112316
rect 77678 112192 77748 112248
rect 77804 112192 77872 112248
rect 77928 112192 77996 112248
rect 78052 112192 78120 112248
rect 78176 112192 78244 112248
rect 78300 112192 78368 112248
rect 78424 112192 78492 112248
rect 78548 112192 78678 112248
rect 70000 105658 70200 105728
rect 70000 105602 70074 105658
rect 70130 105602 70200 105658
rect 70000 105534 70200 105602
rect 70000 105478 70074 105534
rect 70130 105478 70200 105534
rect 70000 105410 70200 105478
rect 70000 105354 70074 105410
rect 70130 105354 70200 105410
rect 70000 105286 70200 105354
rect 70000 105230 70074 105286
rect 70130 105230 70200 105286
rect 70000 105162 70200 105230
rect 70000 105106 70074 105162
rect 70130 105106 70200 105162
rect 70000 105038 70200 105106
rect 70000 104982 70074 105038
rect 70130 104982 70200 105038
rect 70000 104914 70200 104982
rect 70000 104858 70074 104914
rect 70130 104858 70200 104914
rect 70000 104790 70200 104858
rect 70000 104734 70074 104790
rect 70130 104734 70200 104790
rect 70000 104666 70200 104734
rect 70000 104610 70074 104666
rect 70130 104610 70200 104666
rect 70000 104542 70200 104610
rect 70000 104486 70074 104542
rect 70130 104486 70200 104542
rect 70000 104418 70200 104486
rect 70000 104362 70074 104418
rect 70130 104362 70200 104418
rect 70000 104294 70200 104362
rect 70000 104238 70074 104294
rect 70130 104238 70200 104294
rect 70000 104170 70200 104238
rect 70000 104114 70074 104170
rect 70130 104114 70200 104170
rect 70000 104046 70200 104114
rect 70000 103990 70074 104046
rect 70130 103990 70200 104046
rect 70000 103922 70200 103990
rect 70000 103866 70074 103922
rect 70130 103866 70200 103922
rect 70000 103828 70200 103866
rect 77678 105670 78678 112192
rect 77678 105614 77808 105670
rect 77864 105614 77932 105670
rect 77988 105614 78056 105670
rect 78112 105614 78180 105670
rect 78236 105614 78304 105670
rect 78360 105614 78428 105670
rect 78484 105614 78552 105670
rect 78608 105614 78678 105670
rect 77678 105546 78678 105614
rect 77678 105490 77808 105546
rect 77864 105490 77932 105546
rect 77988 105490 78056 105546
rect 78112 105490 78180 105546
rect 78236 105490 78304 105546
rect 78360 105490 78428 105546
rect 78484 105490 78552 105546
rect 78608 105490 78678 105546
rect 77678 105422 78678 105490
rect 77678 105366 77808 105422
rect 77864 105366 77932 105422
rect 77988 105366 78056 105422
rect 78112 105366 78180 105422
rect 78236 105366 78304 105422
rect 78360 105366 78428 105422
rect 78484 105366 78552 105422
rect 78608 105366 78678 105422
rect 77678 105298 78678 105366
rect 77678 105242 77808 105298
rect 77864 105242 77932 105298
rect 77988 105242 78056 105298
rect 78112 105242 78180 105298
rect 78236 105242 78304 105298
rect 78360 105242 78428 105298
rect 78484 105242 78552 105298
rect 78608 105242 78678 105298
rect 77678 105174 78678 105242
rect 77678 105118 77808 105174
rect 77864 105118 77932 105174
rect 77988 105118 78056 105174
rect 78112 105118 78180 105174
rect 78236 105118 78304 105174
rect 78360 105118 78428 105174
rect 78484 105118 78552 105174
rect 78608 105118 78678 105174
rect 77678 105050 78678 105118
rect 77678 104994 77808 105050
rect 77864 104994 77932 105050
rect 77988 104994 78056 105050
rect 78112 104994 78180 105050
rect 78236 104994 78304 105050
rect 78360 104994 78428 105050
rect 78484 104994 78552 105050
rect 78608 104994 78678 105050
rect 77678 104926 78678 104994
rect 77678 104870 77808 104926
rect 77864 104870 77932 104926
rect 77988 104870 78056 104926
rect 78112 104870 78180 104926
rect 78236 104870 78304 104926
rect 78360 104870 78428 104926
rect 78484 104870 78552 104926
rect 78608 104870 78678 104926
rect 77678 104802 78678 104870
rect 77678 104746 77808 104802
rect 77864 104746 77932 104802
rect 77988 104746 78056 104802
rect 78112 104746 78180 104802
rect 78236 104746 78304 104802
rect 78360 104746 78428 104802
rect 78484 104746 78552 104802
rect 78608 104746 78678 104802
rect 77678 104678 78678 104746
rect 77678 104622 77808 104678
rect 77864 104622 77932 104678
rect 77988 104622 78056 104678
rect 78112 104622 78180 104678
rect 78236 104622 78304 104678
rect 78360 104622 78428 104678
rect 78484 104622 78552 104678
rect 78608 104622 78678 104678
rect 77678 104554 78678 104622
rect 77678 104498 77808 104554
rect 77864 104498 77932 104554
rect 77988 104498 78056 104554
rect 78112 104498 78180 104554
rect 78236 104498 78304 104554
rect 78360 104498 78428 104554
rect 78484 104498 78552 104554
rect 78608 104498 78678 104554
rect 77678 104430 78678 104498
rect 77678 104374 77808 104430
rect 77864 104374 77932 104430
rect 77988 104374 78056 104430
rect 78112 104374 78180 104430
rect 78236 104374 78304 104430
rect 78360 104374 78428 104430
rect 78484 104374 78552 104430
rect 78608 104374 78678 104430
rect 77678 104306 78678 104374
rect 77678 104250 77808 104306
rect 77864 104250 77932 104306
rect 77988 104250 78056 104306
rect 78112 104250 78180 104306
rect 78236 104250 78304 104306
rect 78360 104250 78428 104306
rect 78484 104250 78552 104306
rect 78608 104250 78678 104306
rect 77678 104182 78678 104250
rect 77678 104126 77808 104182
rect 77864 104126 77932 104182
rect 77988 104126 78056 104182
rect 78112 104126 78180 104182
rect 78236 104126 78304 104182
rect 78360 104126 78428 104182
rect 78484 104126 78552 104182
rect 78608 104126 78678 104182
rect 77678 104058 78678 104126
rect 77678 104002 77808 104058
rect 77864 104002 77932 104058
rect 77988 104002 78056 104058
rect 78112 104002 78180 104058
rect 78236 104002 78304 104058
rect 78360 104002 78428 104058
rect 78484 104002 78552 104058
rect 78608 104002 78678 104058
rect 77678 103934 78678 104002
rect 77678 103878 77808 103934
rect 77864 103878 77932 103934
rect 77988 103878 78056 103934
rect 78112 103878 78180 103934
rect 78236 103878 78304 103934
rect 78360 103878 78428 103934
rect 78484 103878 78552 103934
rect 78608 103878 78678 103934
rect 70000 103184 70200 103248
rect 70000 103128 70074 103184
rect 70130 103128 70200 103184
rect 70000 103060 70200 103128
rect 70000 103004 70074 103060
rect 70130 103004 70200 103060
rect 70000 102936 70200 103004
rect 70000 102880 70074 102936
rect 70130 102880 70200 102936
rect 70000 102812 70200 102880
rect 70000 102756 70074 102812
rect 70130 102756 70200 102812
rect 70000 102688 70200 102756
rect 70000 102632 70074 102688
rect 70130 102632 70200 102688
rect 70000 102564 70200 102632
rect 70000 102508 70074 102564
rect 70130 102508 70200 102564
rect 70000 102440 70200 102508
rect 70000 102384 70074 102440
rect 70130 102384 70200 102440
rect 70000 102316 70200 102384
rect 70000 102260 70074 102316
rect 70130 102260 70200 102316
rect 70000 102192 70200 102260
rect 70000 102136 70074 102192
rect 70130 102136 70200 102192
rect 70000 102068 70200 102136
rect 70000 102012 70074 102068
rect 70130 102012 70200 102068
rect 70000 101944 70200 102012
rect 70000 101888 70074 101944
rect 70130 101888 70200 101944
rect 70000 101820 70200 101888
rect 70000 101764 70074 101820
rect 70130 101764 70200 101820
rect 70000 101696 70200 101764
rect 70000 101640 70074 101696
rect 70130 101640 70200 101696
rect 70000 101572 70200 101640
rect 70000 101516 70074 101572
rect 70130 101516 70200 101572
rect 70000 101448 70200 101516
rect 70000 101392 70074 101448
rect 70130 101392 70200 101448
rect 70000 101324 70200 101392
rect 70000 101268 70074 101324
rect 70130 101268 70200 101324
rect 70000 101198 70200 101268
rect 77678 103190 78678 103878
rect 77678 103134 77808 103190
rect 77864 103134 77932 103190
rect 77988 103134 78056 103190
rect 78112 103134 78180 103190
rect 78236 103134 78304 103190
rect 78360 103134 78428 103190
rect 78484 103134 78552 103190
rect 78608 103134 78678 103190
rect 77678 103066 78678 103134
rect 77678 103010 77808 103066
rect 77864 103010 77932 103066
rect 77988 103010 78056 103066
rect 78112 103010 78180 103066
rect 78236 103010 78304 103066
rect 78360 103010 78428 103066
rect 78484 103010 78552 103066
rect 78608 103010 78678 103066
rect 77678 102942 78678 103010
rect 77678 102886 77808 102942
rect 77864 102886 77932 102942
rect 77988 102886 78056 102942
rect 78112 102886 78180 102942
rect 78236 102886 78304 102942
rect 78360 102886 78428 102942
rect 78484 102886 78552 102942
rect 78608 102886 78678 102942
rect 77678 102818 78678 102886
rect 77678 102762 77808 102818
rect 77864 102762 77932 102818
rect 77988 102762 78056 102818
rect 78112 102762 78180 102818
rect 78236 102762 78304 102818
rect 78360 102762 78428 102818
rect 78484 102762 78552 102818
rect 78608 102762 78678 102818
rect 77678 102694 78678 102762
rect 77678 102638 77808 102694
rect 77864 102638 77932 102694
rect 77988 102638 78056 102694
rect 78112 102638 78180 102694
rect 78236 102638 78304 102694
rect 78360 102638 78428 102694
rect 78484 102638 78552 102694
rect 78608 102638 78678 102694
rect 77678 102570 78678 102638
rect 77678 102514 77808 102570
rect 77864 102514 77932 102570
rect 77988 102514 78056 102570
rect 78112 102514 78180 102570
rect 78236 102514 78304 102570
rect 78360 102514 78428 102570
rect 78484 102514 78552 102570
rect 78608 102514 78678 102570
rect 77678 102446 78678 102514
rect 77678 102390 77808 102446
rect 77864 102390 77932 102446
rect 77988 102390 78056 102446
rect 78112 102390 78180 102446
rect 78236 102390 78304 102446
rect 78360 102390 78428 102446
rect 78484 102390 78552 102446
rect 78608 102390 78678 102446
rect 77678 102322 78678 102390
rect 77678 102266 77808 102322
rect 77864 102266 77932 102322
rect 77988 102266 78056 102322
rect 78112 102266 78180 102322
rect 78236 102266 78304 102322
rect 78360 102266 78428 102322
rect 78484 102266 78552 102322
rect 78608 102266 78678 102322
rect 77678 102198 78678 102266
rect 77678 102142 77808 102198
rect 77864 102142 77932 102198
rect 77988 102142 78056 102198
rect 78112 102142 78180 102198
rect 78236 102142 78304 102198
rect 78360 102142 78428 102198
rect 78484 102142 78552 102198
rect 78608 102142 78678 102198
rect 77678 102074 78678 102142
rect 77678 102018 77808 102074
rect 77864 102018 77932 102074
rect 77988 102018 78056 102074
rect 78112 102018 78180 102074
rect 78236 102018 78304 102074
rect 78360 102018 78428 102074
rect 78484 102018 78552 102074
rect 78608 102018 78678 102074
rect 77678 101950 78678 102018
rect 77678 101894 77808 101950
rect 77864 101894 77932 101950
rect 77988 101894 78056 101950
rect 78112 101894 78180 101950
rect 78236 101894 78304 101950
rect 78360 101894 78428 101950
rect 78484 101894 78552 101950
rect 78608 101894 78678 101950
rect 77678 101826 78678 101894
rect 77678 101770 77808 101826
rect 77864 101770 77932 101826
rect 77988 101770 78056 101826
rect 78112 101770 78180 101826
rect 78236 101770 78304 101826
rect 78360 101770 78428 101826
rect 78484 101770 78552 101826
rect 78608 101770 78678 101826
rect 77678 101702 78678 101770
rect 77678 101646 77808 101702
rect 77864 101646 77932 101702
rect 77988 101646 78056 101702
rect 78112 101646 78180 101702
rect 78236 101646 78304 101702
rect 78360 101646 78428 101702
rect 78484 101646 78552 101702
rect 78608 101646 78678 101702
rect 77678 101578 78678 101646
rect 77678 101522 77808 101578
rect 77864 101522 77932 101578
rect 77988 101522 78056 101578
rect 78112 101522 78180 101578
rect 78236 101522 78304 101578
rect 78360 101522 78428 101578
rect 78484 101522 78552 101578
rect 78608 101522 78678 101578
rect 77678 101454 78678 101522
rect 77678 101398 77808 101454
rect 77864 101398 77932 101454
rect 77988 101398 78056 101454
rect 78112 101398 78180 101454
rect 78236 101398 78304 101454
rect 78360 101398 78428 101454
rect 78484 101398 78552 101454
rect 78608 101398 78678 101454
rect 77678 101330 78678 101398
rect 77678 101274 77808 101330
rect 77864 101274 77932 101330
rect 77988 101274 78056 101330
rect 78112 101274 78180 101330
rect 78236 101274 78304 101330
rect 78360 101274 78428 101330
rect 78484 101274 78552 101330
rect 78608 101274 78678 101330
rect 70000 100814 70200 100878
rect 70000 100758 70074 100814
rect 70130 100758 70200 100814
rect 70000 100690 70200 100758
rect 70000 100634 70074 100690
rect 70130 100634 70200 100690
rect 70000 100566 70200 100634
rect 70000 100510 70074 100566
rect 70130 100510 70200 100566
rect 70000 100442 70200 100510
rect 70000 100386 70074 100442
rect 70130 100386 70200 100442
rect 70000 100318 70200 100386
rect 70000 100262 70074 100318
rect 70130 100262 70200 100318
rect 70000 100194 70200 100262
rect 70000 100138 70074 100194
rect 70130 100138 70200 100194
rect 70000 100070 70200 100138
rect 70000 100014 70074 100070
rect 70130 100014 70200 100070
rect 70000 99946 70200 100014
rect 70000 99890 70074 99946
rect 70130 99890 70200 99946
rect 70000 99822 70200 99890
rect 70000 99766 70074 99822
rect 70130 99766 70200 99822
rect 70000 99698 70200 99766
rect 70000 99642 70074 99698
rect 70130 99642 70200 99698
rect 70000 99574 70200 99642
rect 70000 99518 70074 99574
rect 70130 99518 70200 99574
rect 70000 99450 70200 99518
rect 70000 99394 70074 99450
rect 70130 99394 70200 99450
rect 70000 99326 70200 99394
rect 70000 99270 70074 99326
rect 70130 99270 70200 99326
rect 70000 99202 70200 99270
rect 70000 99146 70074 99202
rect 70130 99146 70200 99202
rect 70000 99078 70200 99146
rect 70000 99022 70074 99078
rect 70130 99022 70200 99078
rect 70000 98954 70200 99022
rect 70000 98898 70074 98954
rect 70130 98898 70200 98954
rect 70000 98828 70200 98898
rect 77678 100820 78678 101274
rect 77678 100764 77808 100820
rect 77864 100764 77932 100820
rect 77988 100764 78056 100820
rect 78112 100764 78180 100820
rect 78236 100764 78304 100820
rect 78360 100764 78428 100820
rect 78484 100764 78552 100820
rect 78608 100764 78678 100820
rect 77678 100696 78678 100764
rect 77678 100640 77808 100696
rect 77864 100640 77932 100696
rect 77988 100640 78056 100696
rect 78112 100640 78180 100696
rect 78236 100640 78304 100696
rect 78360 100640 78428 100696
rect 78484 100640 78552 100696
rect 78608 100640 78678 100696
rect 77678 100572 78678 100640
rect 77678 100516 77808 100572
rect 77864 100516 77932 100572
rect 77988 100516 78056 100572
rect 78112 100516 78180 100572
rect 78236 100516 78304 100572
rect 78360 100516 78428 100572
rect 78484 100516 78552 100572
rect 78608 100516 78678 100572
rect 77678 100448 78678 100516
rect 77678 100392 77808 100448
rect 77864 100392 77932 100448
rect 77988 100392 78056 100448
rect 78112 100392 78180 100448
rect 78236 100392 78304 100448
rect 78360 100392 78428 100448
rect 78484 100392 78552 100448
rect 78608 100392 78678 100448
rect 77678 100324 78678 100392
rect 77678 100268 77808 100324
rect 77864 100268 77932 100324
rect 77988 100268 78056 100324
rect 78112 100268 78180 100324
rect 78236 100268 78304 100324
rect 78360 100268 78428 100324
rect 78484 100268 78552 100324
rect 78608 100268 78678 100324
rect 77678 100200 78678 100268
rect 77678 100144 77808 100200
rect 77864 100144 77932 100200
rect 77988 100144 78056 100200
rect 78112 100144 78180 100200
rect 78236 100144 78304 100200
rect 78360 100144 78428 100200
rect 78484 100144 78552 100200
rect 78608 100144 78678 100200
rect 77678 100076 78678 100144
rect 77678 100020 77808 100076
rect 77864 100020 77932 100076
rect 77988 100020 78056 100076
rect 78112 100020 78180 100076
rect 78236 100020 78304 100076
rect 78360 100020 78428 100076
rect 78484 100020 78552 100076
rect 78608 100020 78678 100076
rect 77678 99952 78678 100020
rect 77678 99896 77808 99952
rect 77864 99896 77932 99952
rect 77988 99896 78056 99952
rect 78112 99896 78180 99952
rect 78236 99896 78304 99952
rect 78360 99896 78428 99952
rect 78484 99896 78552 99952
rect 78608 99896 78678 99952
rect 77678 99828 78678 99896
rect 77678 99772 77808 99828
rect 77864 99772 77932 99828
rect 77988 99772 78056 99828
rect 78112 99772 78180 99828
rect 78236 99772 78304 99828
rect 78360 99772 78428 99828
rect 78484 99772 78552 99828
rect 78608 99772 78678 99828
rect 77678 99704 78678 99772
rect 77678 99648 77808 99704
rect 77864 99648 77932 99704
rect 77988 99648 78056 99704
rect 78112 99648 78180 99704
rect 78236 99648 78304 99704
rect 78360 99648 78428 99704
rect 78484 99648 78552 99704
rect 78608 99648 78678 99704
rect 77678 99580 78678 99648
rect 77678 99524 77808 99580
rect 77864 99524 77932 99580
rect 77988 99524 78056 99580
rect 78112 99524 78180 99580
rect 78236 99524 78304 99580
rect 78360 99524 78428 99580
rect 78484 99524 78552 99580
rect 78608 99524 78678 99580
rect 77678 99456 78678 99524
rect 77678 99400 77808 99456
rect 77864 99400 77932 99456
rect 77988 99400 78056 99456
rect 78112 99400 78180 99456
rect 78236 99400 78304 99456
rect 78360 99400 78428 99456
rect 78484 99400 78552 99456
rect 78608 99400 78678 99456
rect 77678 99332 78678 99400
rect 77678 99276 77808 99332
rect 77864 99276 77932 99332
rect 77988 99276 78056 99332
rect 78112 99276 78180 99332
rect 78236 99276 78304 99332
rect 78360 99276 78428 99332
rect 78484 99276 78552 99332
rect 78608 99276 78678 99332
rect 77678 99208 78678 99276
rect 77678 99152 77808 99208
rect 77864 99152 77932 99208
rect 77988 99152 78056 99208
rect 78112 99152 78180 99208
rect 78236 99152 78304 99208
rect 78360 99152 78428 99208
rect 78484 99152 78552 99208
rect 78608 99152 78678 99208
rect 77678 99084 78678 99152
rect 77678 99028 77808 99084
rect 77864 99028 77932 99084
rect 77988 99028 78056 99084
rect 78112 99028 78180 99084
rect 78236 99028 78304 99084
rect 78360 99028 78428 99084
rect 78484 99028 78552 99084
rect 78608 99028 78678 99084
rect 77678 98960 78678 99028
rect 77678 98904 77808 98960
rect 77864 98904 77932 98960
rect 77988 98904 78056 98960
rect 78112 98904 78180 98960
rect 78236 98904 78304 98960
rect 78360 98904 78428 98960
rect 78484 98904 78552 98960
rect 78608 98904 78678 98960
rect 70000 98108 70200 98172
rect 70000 98052 70074 98108
rect 70130 98052 70200 98108
rect 70000 97984 70200 98052
rect 70000 97928 70074 97984
rect 70130 97928 70200 97984
rect 70000 97860 70200 97928
rect 70000 97804 70074 97860
rect 70130 97804 70200 97860
rect 70000 97736 70200 97804
rect 70000 97680 70074 97736
rect 70130 97680 70200 97736
rect 70000 97612 70200 97680
rect 70000 97556 70074 97612
rect 70130 97556 70200 97612
rect 70000 97488 70200 97556
rect 70000 97432 70074 97488
rect 70130 97432 70200 97488
rect 70000 97364 70200 97432
rect 70000 97308 70074 97364
rect 70130 97308 70200 97364
rect 70000 97240 70200 97308
rect 70000 97184 70074 97240
rect 70130 97184 70200 97240
rect 70000 97116 70200 97184
rect 70000 97060 70074 97116
rect 70130 97060 70200 97116
rect 70000 96992 70200 97060
rect 70000 96936 70074 96992
rect 70130 96936 70200 96992
rect 70000 96868 70200 96936
rect 70000 96812 70074 96868
rect 70130 96812 70200 96868
rect 70000 96744 70200 96812
rect 70000 96688 70074 96744
rect 70130 96688 70200 96744
rect 70000 96620 70200 96688
rect 70000 96564 70074 96620
rect 70130 96564 70200 96620
rect 70000 96496 70200 96564
rect 70000 96440 70074 96496
rect 70130 96440 70200 96496
rect 70000 96372 70200 96440
rect 70000 96316 70074 96372
rect 70130 96316 70200 96372
rect 70000 96248 70200 96316
rect 70000 96192 70074 96248
rect 70130 96192 70200 96248
rect 70000 96122 70200 96192
rect 77678 98114 78678 98904
rect 77678 98058 77808 98114
rect 77864 98058 77932 98114
rect 77988 98058 78056 98114
rect 78112 98058 78180 98114
rect 78236 98058 78304 98114
rect 78360 98058 78428 98114
rect 78484 98058 78552 98114
rect 78608 98058 78678 98114
rect 77678 97990 78678 98058
rect 77678 97934 77808 97990
rect 77864 97934 77932 97990
rect 77988 97934 78056 97990
rect 78112 97934 78180 97990
rect 78236 97934 78304 97990
rect 78360 97934 78428 97990
rect 78484 97934 78552 97990
rect 78608 97934 78678 97990
rect 77678 97866 78678 97934
rect 77678 97810 77808 97866
rect 77864 97810 77932 97866
rect 77988 97810 78056 97866
rect 78112 97810 78180 97866
rect 78236 97810 78304 97866
rect 78360 97810 78428 97866
rect 78484 97810 78552 97866
rect 78608 97810 78678 97866
rect 77678 97742 78678 97810
rect 77678 97686 77808 97742
rect 77864 97686 77932 97742
rect 77988 97686 78056 97742
rect 78112 97686 78180 97742
rect 78236 97686 78304 97742
rect 78360 97686 78428 97742
rect 78484 97686 78552 97742
rect 78608 97686 78678 97742
rect 77678 97618 78678 97686
rect 77678 97562 77808 97618
rect 77864 97562 77932 97618
rect 77988 97562 78056 97618
rect 78112 97562 78180 97618
rect 78236 97562 78304 97618
rect 78360 97562 78428 97618
rect 78484 97562 78552 97618
rect 78608 97562 78678 97618
rect 77678 97494 78678 97562
rect 77678 97438 77808 97494
rect 77864 97438 77932 97494
rect 77988 97438 78056 97494
rect 78112 97438 78180 97494
rect 78236 97438 78304 97494
rect 78360 97438 78428 97494
rect 78484 97438 78552 97494
rect 78608 97438 78678 97494
rect 77678 97370 78678 97438
rect 77678 97314 77808 97370
rect 77864 97314 77932 97370
rect 77988 97314 78056 97370
rect 78112 97314 78180 97370
rect 78236 97314 78304 97370
rect 78360 97314 78428 97370
rect 78484 97314 78552 97370
rect 78608 97314 78678 97370
rect 77678 97246 78678 97314
rect 77678 97190 77808 97246
rect 77864 97190 77932 97246
rect 77988 97190 78056 97246
rect 78112 97190 78180 97246
rect 78236 97190 78304 97246
rect 78360 97190 78428 97246
rect 78484 97190 78552 97246
rect 78608 97190 78678 97246
rect 77678 97122 78678 97190
rect 77678 97066 77808 97122
rect 77864 97066 77932 97122
rect 77988 97066 78056 97122
rect 78112 97066 78180 97122
rect 78236 97066 78304 97122
rect 78360 97066 78428 97122
rect 78484 97066 78552 97122
rect 78608 97066 78678 97122
rect 77678 96998 78678 97066
rect 77678 96942 77808 96998
rect 77864 96942 77932 96998
rect 77988 96942 78056 96998
rect 78112 96942 78180 96998
rect 78236 96942 78304 96998
rect 78360 96942 78428 96998
rect 78484 96942 78552 96998
rect 78608 96942 78678 96998
rect 77678 96874 78678 96942
rect 77678 96818 77808 96874
rect 77864 96818 77932 96874
rect 77988 96818 78056 96874
rect 78112 96818 78180 96874
rect 78236 96818 78304 96874
rect 78360 96818 78428 96874
rect 78484 96818 78552 96874
rect 78608 96818 78678 96874
rect 77678 96750 78678 96818
rect 77678 96694 77808 96750
rect 77864 96694 77932 96750
rect 77988 96694 78056 96750
rect 78112 96694 78180 96750
rect 78236 96694 78304 96750
rect 78360 96694 78428 96750
rect 78484 96694 78552 96750
rect 78608 96694 78678 96750
rect 77678 96626 78678 96694
rect 77678 96570 77808 96626
rect 77864 96570 77932 96626
rect 77988 96570 78056 96626
rect 78112 96570 78180 96626
rect 78236 96570 78304 96626
rect 78360 96570 78428 96626
rect 78484 96570 78552 96626
rect 78608 96570 78678 96626
rect 77678 96502 78678 96570
rect 77678 96446 77808 96502
rect 77864 96446 77932 96502
rect 77988 96446 78056 96502
rect 78112 96446 78180 96502
rect 78236 96446 78304 96502
rect 78360 96446 78428 96502
rect 78484 96446 78552 96502
rect 78608 96446 78678 96502
rect 77678 96378 78678 96446
rect 77678 96322 77808 96378
rect 77864 96322 77932 96378
rect 77988 96322 78056 96378
rect 78112 96322 78180 96378
rect 78236 96322 78304 96378
rect 78360 96322 78428 96378
rect 78484 96322 78552 96378
rect 78608 96322 78678 96378
rect 77678 96254 78678 96322
rect 77678 96198 77808 96254
rect 77864 96198 77932 96254
rect 77988 96198 78056 96254
rect 78112 96198 78180 96254
rect 78236 96198 78304 96254
rect 78360 96198 78428 96254
rect 78484 96198 78552 96254
rect 78608 96198 78678 96254
rect 70000 95738 70200 95802
rect 70000 95682 70074 95738
rect 70130 95682 70200 95738
rect 70000 95614 70200 95682
rect 70000 95558 70074 95614
rect 70130 95558 70200 95614
rect 70000 95490 70200 95558
rect 70000 95434 70074 95490
rect 70130 95434 70200 95490
rect 70000 95366 70200 95434
rect 70000 95310 70074 95366
rect 70130 95310 70200 95366
rect 70000 95242 70200 95310
rect 70000 95186 70074 95242
rect 70130 95186 70200 95242
rect 70000 95118 70200 95186
rect 70000 95062 70074 95118
rect 70130 95062 70200 95118
rect 70000 94994 70200 95062
rect 70000 94938 70074 94994
rect 70130 94938 70200 94994
rect 70000 94870 70200 94938
rect 70000 94814 70074 94870
rect 70130 94814 70200 94870
rect 70000 94746 70200 94814
rect 70000 94690 70074 94746
rect 70130 94690 70200 94746
rect 70000 94622 70200 94690
rect 70000 94566 70074 94622
rect 70130 94566 70200 94622
rect 70000 94498 70200 94566
rect 70000 94442 70074 94498
rect 70130 94442 70200 94498
rect 70000 94374 70200 94442
rect 70000 94318 70074 94374
rect 70130 94318 70200 94374
rect 70000 94250 70200 94318
rect 70000 94194 70074 94250
rect 70130 94194 70200 94250
rect 70000 94126 70200 94194
rect 70000 94070 70074 94126
rect 70130 94070 70200 94126
rect 70000 94002 70200 94070
rect 70000 93946 70074 94002
rect 70130 93946 70200 94002
rect 70000 93878 70200 93946
rect 70000 93822 70074 93878
rect 70130 93822 70200 93878
rect 70000 93752 70200 93822
rect 77678 95744 78678 96198
rect 77678 95688 77808 95744
rect 77864 95688 77932 95744
rect 77988 95688 78056 95744
rect 78112 95688 78180 95744
rect 78236 95688 78304 95744
rect 78360 95688 78428 95744
rect 78484 95688 78552 95744
rect 78608 95688 78678 95744
rect 77678 95620 78678 95688
rect 77678 95564 77808 95620
rect 77864 95564 77932 95620
rect 77988 95564 78056 95620
rect 78112 95564 78180 95620
rect 78236 95564 78304 95620
rect 78360 95564 78428 95620
rect 78484 95564 78552 95620
rect 78608 95564 78678 95620
rect 77678 95496 78678 95564
rect 77678 95440 77808 95496
rect 77864 95440 77932 95496
rect 77988 95440 78056 95496
rect 78112 95440 78180 95496
rect 78236 95440 78304 95496
rect 78360 95440 78428 95496
rect 78484 95440 78552 95496
rect 78608 95440 78678 95496
rect 77678 95372 78678 95440
rect 77678 95316 77808 95372
rect 77864 95316 77932 95372
rect 77988 95316 78056 95372
rect 78112 95316 78180 95372
rect 78236 95316 78304 95372
rect 78360 95316 78428 95372
rect 78484 95316 78552 95372
rect 78608 95316 78678 95372
rect 77678 95248 78678 95316
rect 77678 95192 77808 95248
rect 77864 95192 77932 95248
rect 77988 95192 78056 95248
rect 78112 95192 78180 95248
rect 78236 95192 78304 95248
rect 78360 95192 78428 95248
rect 78484 95192 78552 95248
rect 78608 95192 78678 95248
rect 77678 95124 78678 95192
rect 77678 95068 77808 95124
rect 77864 95068 77932 95124
rect 77988 95068 78056 95124
rect 78112 95068 78180 95124
rect 78236 95068 78304 95124
rect 78360 95068 78428 95124
rect 78484 95068 78552 95124
rect 78608 95068 78678 95124
rect 77678 95000 78678 95068
rect 77678 94944 77808 95000
rect 77864 94944 77932 95000
rect 77988 94944 78056 95000
rect 78112 94944 78180 95000
rect 78236 94944 78304 95000
rect 78360 94944 78428 95000
rect 78484 94944 78552 95000
rect 78608 94944 78678 95000
rect 77678 94876 78678 94944
rect 77678 94820 77808 94876
rect 77864 94820 77932 94876
rect 77988 94820 78056 94876
rect 78112 94820 78180 94876
rect 78236 94820 78304 94876
rect 78360 94820 78428 94876
rect 78484 94820 78552 94876
rect 78608 94820 78678 94876
rect 77678 94752 78678 94820
rect 77678 94696 77808 94752
rect 77864 94696 77932 94752
rect 77988 94696 78056 94752
rect 78112 94696 78180 94752
rect 78236 94696 78304 94752
rect 78360 94696 78428 94752
rect 78484 94696 78552 94752
rect 78608 94696 78678 94752
rect 77678 94628 78678 94696
rect 77678 94572 77808 94628
rect 77864 94572 77932 94628
rect 77988 94572 78056 94628
rect 78112 94572 78180 94628
rect 78236 94572 78304 94628
rect 78360 94572 78428 94628
rect 78484 94572 78552 94628
rect 78608 94572 78678 94628
rect 77678 94504 78678 94572
rect 77678 94448 77808 94504
rect 77864 94448 77932 94504
rect 77988 94448 78056 94504
rect 78112 94448 78180 94504
rect 78236 94448 78304 94504
rect 78360 94448 78428 94504
rect 78484 94448 78552 94504
rect 78608 94448 78678 94504
rect 77678 94380 78678 94448
rect 77678 94324 77808 94380
rect 77864 94324 77932 94380
rect 77988 94324 78056 94380
rect 78112 94324 78180 94380
rect 78236 94324 78304 94380
rect 78360 94324 78428 94380
rect 78484 94324 78552 94380
rect 78608 94324 78678 94380
rect 77678 94256 78678 94324
rect 77678 94200 77808 94256
rect 77864 94200 77932 94256
rect 77988 94200 78056 94256
rect 78112 94200 78180 94256
rect 78236 94200 78304 94256
rect 78360 94200 78428 94256
rect 78484 94200 78552 94256
rect 78608 94200 78678 94256
rect 77678 94132 78678 94200
rect 77678 94076 77808 94132
rect 77864 94076 77932 94132
rect 77988 94076 78056 94132
rect 78112 94076 78180 94132
rect 78236 94076 78304 94132
rect 78360 94076 78428 94132
rect 78484 94076 78552 94132
rect 78608 94076 78678 94132
rect 77678 94008 78678 94076
rect 77678 93952 77808 94008
rect 77864 93952 77932 94008
rect 77988 93952 78056 94008
rect 78112 93952 78180 94008
rect 78236 93952 78304 94008
rect 78360 93952 78428 94008
rect 78484 93952 78552 94008
rect 78608 93952 78678 94008
rect 77678 93884 78678 93952
rect 77678 93828 77808 93884
rect 77864 93828 77932 93884
rect 77988 93828 78056 93884
rect 78112 93828 78180 93884
rect 78236 93828 78304 93884
rect 78360 93828 78428 93884
rect 78484 93828 78552 93884
rect 78608 93828 78678 93884
rect 70000 93134 70200 93172
rect 70000 93078 70074 93134
rect 70130 93078 70200 93134
rect 70000 93010 70200 93078
rect 70000 92954 70074 93010
rect 70130 92954 70200 93010
rect 70000 92886 70200 92954
rect 70000 92830 70074 92886
rect 70130 92830 70200 92886
rect 70000 92762 70200 92830
rect 70000 92706 70074 92762
rect 70130 92706 70200 92762
rect 70000 92638 70200 92706
rect 70000 92582 70074 92638
rect 70130 92582 70200 92638
rect 70000 92514 70200 92582
rect 70000 92458 70074 92514
rect 70130 92458 70200 92514
rect 70000 92390 70200 92458
rect 70000 92334 70074 92390
rect 70130 92334 70200 92390
rect 70000 92266 70200 92334
rect 70000 92210 70074 92266
rect 70130 92210 70200 92266
rect 70000 92142 70200 92210
rect 70000 92086 70074 92142
rect 70130 92086 70200 92142
rect 70000 92018 70200 92086
rect 70000 91962 70074 92018
rect 70130 91962 70200 92018
rect 70000 91894 70200 91962
rect 70000 91838 70074 91894
rect 70130 91838 70200 91894
rect 70000 91770 70200 91838
rect 70000 91714 70074 91770
rect 70130 91714 70200 91770
rect 70000 91646 70200 91714
rect 70000 91590 70074 91646
rect 70130 91590 70200 91646
rect 70000 91522 70200 91590
rect 70000 91466 70074 91522
rect 70130 91466 70200 91522
rect 70000 91398 70200 91466
rect 70000 91342 70074 91398
rect 70130 91342 70200 91398
rect 70000 91272 70200 91342
rect 77678 93140 78678 93828
rect 77678 93084 77808 93140
rect 77864 93084 77932 93140
rect 77988 93084 78056 93140
rect 78112 93084 78180 93140
rect 78236 93084 78304 93140
rect 78360 93084 78428 93140
rect 78484 93084 78552 93140
rect 78608 93084 78678 93140
rect 77678 93016 78678 93084
rect 77678 92960 77808 93016
rect 77864 92960 77932 93016
rect 77988 92960 78056 93016
rect 78112 92960 78180 93016
rect 78236 92960 78304 93016
rect 78360 92960 78428 93016
rect 78484 92960 78552 93016
rect 78608 92960 78678 93016
rect 77678 92892 78678 92960
rect 77678 92836 77808 92892
rect 77864 92836 77932 92892
rect 77988 92836 78056 92892
rect 78112 92836 78180 92892
rect 78236 92836 78304 92892
rect 78360 92836 78428 92892
rect 78484 92836 78552 92892
rect 78608 92836 78678 92892
rect 77678 92768 78678 92836
rect 77678 92712 77808 92768
rect 77864 92712 77932 92768
rect 77988 92712 78056 92768
rect 78112 92712 78180 92768
rect 78236 92712 78304 92768
rect 78360 92712 78428 92768
rect 78484 92712 78552 92768
rect 78608 92712 78678 92768
rect 77678 92644 78678 92712
rect 77678 92588 77808 92644
rect 77864 92588 77932 92644
rect 77988 92588 78056 92644
rect 78112 92588 78180 92644
rect 78236 92588 78304 92644
rect 78360 92588 78428 92644
rect 78484 92588 78552 92644
rect 78608 92588 78678 92644
rect 77678 92520 78678 92588
rect 77678 92464 77808 92520
rect 77864 92464 77932 92520
rect 77988 92464 78056 92520
rect 78112 92464 78180 92520
rect 78236 92464 78304 92520
rect 78360 92464 78428 92520
rect 78484 92464 78552 92520
rect 78608 92464 78678 92520
rect 77678 92396 78678 92464
rect 77678 92340 77808 92396
rect 77864 92340 77932 92396
rect 77988 92340 78056 92396
rect 78112 92340 78180 92396
rect 78236 92340 78304 92396
rect 78360 92340 78428 92396
rect 78484 92340 78552 92396
rect 78608 92340 78678 92396
rect 77678 92272 78678 92340
rect 77678 92216 77808 92272
rect 77864 92216 77932 92272
rect 77988 92216 78056 92272
rect 78112 92216 78180 92272
rect 78236 92216 78304 92272
rect 78360 92216 78428 92272
rect 78484 92216 78552 92272
rect 78608 92216 78678 92272
rect 77678 92148 78678 92216
rect 77678 92092 77808 92148
rect 77864 92092 77932 92148
rect 77988 92092 78056 92148
rect 78112 92092 78180 92148
rect 78236 92092 78304 92148
rect 78360 92092 78428 92148
rect 78484 92092 78552 92148
rect 78608 92092 78678 92148
rect 77678 92024 78678 92092
rect 77678 91968 77808 92024
rect 77864 91968 77932 92024
rect 77988 91968 78056 92024
rect 78112 91968 78180 92024
rect 78236 91968 78304 92024
rect 78360 91968 78428 92024
rect 78484 91968 78552 92024
rect 78608 91968 78678 92024
rect 77678 91900 78678 91968
rect 77678 91844 77808 91900
rect 77864 91844 77932 91900
rect 77988 91844 78056 91900
rect 78112 91844 78180 91900
rect 78236 91844 78304 91900
rect 78360 91844 78428 91900
rect 78484 91844 78552 91900
rect 78608 91844 78678 91900
rect 77678 91776 78678 91844
rect 77678 91720 77808 91776
rect 77864 91720 77932 91776
rect 77988 91720 78056 91776
rect 78112 91720 78180 91776
rect 78236 91720 78304 91776
rect 78360 91720 78428 91776
rect 78484 91720 78552 91776
rect 78608 91720 78678 91776
rect 77678 91652 78678 91720
rect 77678 91596 77808 91652
rect 77864 91596 77932 91652
rect 77988 91596 78056 91652
rect 78112 91596 78180 91652
rect 78236 91596 78304 91652
rect 78360 91596 78428 91652
rect 78484 91596 78552 91652
rect 78608 91596 78678 91652
rect 77678 91528 78678 91596
rect 77678 91472 77808 91528
rect 77864 91472 77932 91528
rect 77988 91472 78056 91528
rect 78112 91472 78180 91528
rect 78236 91472 78304 91528
rect 78360 91472 78428 91528
rect 78484 91472 78552 91528
rect 78608 91472 78678 91528
rect 77678 91404 78678 91472
rect 77678 91348 77808 91404
rect 77864 91348 77932 91404
rect 77988 91348 78056 91404
rect 78112 91348 78180 91404
rect 78236 91348 78304 91404
rect 78360 91348 78428 91404
rect 78484 91348 78552 91404
rect 78608 91348 78678 91404
rect 77678 86372 78678 91348
rect 77678 86316 77748 86372
rect 77804 86316 77872 86372
rect 77928 86316 77996 86372
rect 78052 86316 78120 86372
rect 78176 86316 78244 86372
rect 78300 86316 78368 86372
rect 78424 86316 78492 86372
rect 78548 86316 78678 86372
rect 77678 86248 78678 86316
rect 77678 86192 77748 86248
rect 77804 86192 77872 86248
rect 77928 86192 77996 86248
rect 78052 86192 78120 86248
rect 78176 86192 78244 86248
rect 78300 86192 78368 86248
rect 78424 86192 78492 86248
rect 78548 86192 78678 86248
rect 77678 78608 78678 86192
rect 79078 940852 80078 945992
rect 140339 943565 140939 943885
rect 195339 943565 195939 943885
rect 250339 943565 250939 943885
rect 305339 943565 305939 943885
rect 360339 943565 360939 943885
rect 110424 943435 110744 943504
rect 110424 943379 110548 943435
rect 110604 943379 110744 943435
rect 79078 940796 79148 940852
rect 79204 940796 79272 940852
rect 79328 940796 79396 940852
rect 79452 940796 79520 940852
rect 79576 940796 79644 940852
rect 79700 940796 79768 940852
rect 79824 940796 79892 940852
rect 79948 940796 80078 940852
rect 79078 940728 80078 940796
rect 79078 940672 79148 940728
rect 79204 940672 79272 940728
rect 79328 940672 79396 940728
rect 79452 940672 79520 940728
rect 79576 940672 79644 940728
rect 79700 940672 79768 940728
rect 79824 940672 79892 940728
rect 79948 940672 80078 940728
rect 79078 940604 80078 940672
rect 79078 940548 79148 940604
rect 79204 940548 79272 940604
rect 79328 940548 79396 940604
rect 79452 940548 79520 940604
rect 79576 940548 79644 940604
rect 79700 940548 79768 940604
rect 79824 940548 79892 940604
rect 79948 940548 80078 940604
rect 79078 940480 80078 940548
rect 79078 940424 79148 940480
rect 79204 940424 79272 940480
rect 79328 940424 79396 940480
rect 79452 940424 79520 940480
rect 79576 940424 79644 940480
rect 79700 940424 79768 940480
rect 79824 940424 79892 940480
rect 79948 940424 80078 940480
rect 79078 940356 80078 940424
rect 79078 940300 79148 940356
rect 79204 940300 79272 940356
rect 79328 940300 79396 940356
rect 79452 940300 79520 940356
rect 79576 940300 79644 940356
rect 79700 940300 79768 940356
rect 79824 940300 79892 940356
rect 79948 940300 80078 940356
rect 79078 940232 80078 940300
rect 79078 940176 79148 940232
rect 79204 940176 79272 940232
rect 79328 940176 79396 940232
rect 79452 940176 79520 940232
rect 79576 940176 79644 940232
rect 79700 940176 79768 940232
rect 79824 940176 79892 940232
rect 79948 940176 80078 940232
rect 79078 940108 80078 940176
rect 79078 940052 79148 940108
rect 79204 940052 79272 940108
rect 79328 940052 79396 940108
rect 79452 940052 79520 940108
rect 79576 940052 79644 940108
rect 79700 940052 79768 940108
rect 79824 940052 79892 940108
rect 79948 940052 80078 940108
rect 79078 929622 80078 940052
rect 88006 942200 88626 942322
rect 88006 942144 88207 942200
rect 88263 942144 88407 942200
rect 88463 942144 88626 942200
rect 88006 941900 88626 942144
rect 88006 941844 88207 941900
rect 88263 941844 88407 941900
rect 88463 941844 88626 941900
rect 88006 941600 88626 941844
rect 88006 941544 88207 941600
rect 88263 941544 88407 941600
rect 88463 941544 88626 941600
rect 88006 933608 88626 941544
rect 106006 940800 106626 940922
rect 106006 940744 106207 940800
rect 106263 940744 106407 940800
rect 106463 940744 106626 940800
rect 106006 940500 106626 940744
rect 106006 940444 106207 940500
rect 106263 940444 106407 940500
rect 106463 940444 106626 940500
rect 106006 940200 106626 940444
rect 106006 940144 106207 940200
rect 106263 940144 106407 940200
rect 106463 940144 106626 940200
rect 106006 934568 106626 940144
rect 110424 940710 110744 943379
rect 110424 940654 110546 940710
rect 110602 940654 110744 940710
rect 110424 940410 110744 940654
rect 110424 940354 110546 940410
rect 110602 940354 110744 940410
rect 110424 940110 110744 940354
rect 110424 940054 110546 940110
rect 110602 940054 110744 940110
rect 110424 939922 110744 940054
rect 117424 943435 117744 943504
rect 117424 943379 117548 943435
rect 117604 943379 117744 943435
rect 117424 940710 117744 943379
rect 117424 940654 117546 940710
rect 117602 940654 117744 940710
rect 117424 940410 117744 940654
rect 117424 940354 117546 940410
rect 117602 940354 117744 940410
rect 117424 940110 117744 940354
rect 117424 940054 117546 940110
rect 117602 940054 117744 940110
rect 117424 939922 117744 940054
rect 124424 943435 124744 943504
rect 124424 943379 124548 943435
rect 124604 943379 124744 943435
rect 124424 940710 124744 943379
rect 140339 942153 140539 943085
rect 140339 942097 140406 942153
rect 140462 942097 140539 942153
rect 140339 941853 140539 942097
rect 140339 941797 140406 941853
rect 140462 941797 140539 941853
rect 140339 941553 140539 941797
rect 140339 941497 140406 941553
rect 140462 941497 140539 941553
rect 140339 941322 140539 941497
rect 124424 940654 124546 940710
rect 124602 940654 124744 940710
rect 124424 940410 124744 940654
rect 124424 940354 124546 940410
rect 124602 940354 124744 940410
rect 124424 940110 124744 940354
rect 124424 940054 124546 940110
rect 124602 940054 124744 940110
rect 124424 939922 124744 940054
rect 140739 940716 140939 943565
rect 165424 943435 165744 943504
rect 165424 943379 165548 943435
rect 165604 943379 165744 943435
rect 160006 942200 160626 942322
rect 160006 942144 160207 942200
rect 160263 942144 160407 942200
rect 160463 942144 160626 942200
rect 160006 941900 160626 942144
rect 160006 941844 160207 941900
rect 160263 941844 160407 941900
rect 160463 941844 160626 941900
rect 160006 941600 160626 941844
rect 160006 941544 160207 941600
rect 160263 941544 160407 941600
rect 160463 941544 160626 941600
rect 140739 940660 140821 940716
rect 140877 940660 140939 940716
rect 140739 940416 140939 940660
rect 140739 940360 140821 940416
rect 140877 940360 140939 940416
rect 140739 940116 140939 940360
rect 140739 940060 140821 940116
rect 140877 940060 140939 940116
rect 140739 939922 140939 940060
rect 142006 940800 142626 940922
rect 142006 940744 142207 940800
rect 142263 940744 142407 940800
rect 142463 940744 142626 940800
rect 142006 940500 142626 940744
rect 142006 940444 142207 940500
rect 142263 940444 142407 940500
rect 142463 940444 142626 940500
rect 142006 940200 142626 940444
rect 142006 940144 142207 940200
rect 142263 940144 142407 940200
rect 142463 940144 142626 940200
rect 142006 934568 142626 940144
rect 160006 933608 160626 941544
rect 165424 940710 165744 943379
rect 165424 940654 165546 940710
rect 165602 940654 165744 940710
rect 165424 940410 165744 940654
rect 165424 940354 165546 940410
rect 165602 940354 165744 940410
rect 165424 940110 165744 940354
rect 165424 940054 165546 940110
rect 165602 940054 165744 940110
rect 165424 939922 165744 940054
rect 172424 943435 172744 943504
rect 172424 943379 172548 943435
rect 172604 943379 172744 943435
rect 172424 940710 172744 943379
rect 179424 943435 179744 943504
rect 179424 943379 179548 943435
rect 179604 943379 179744 943435
rect 172424 940654 172546 940710
rect 172602 940654 172744 940710
rect 172424 940410 172744 940654
rect 172424 940354 172546 940410
rect 172602 940354 172744 940410
rect 172424 940110 172744 940354
rect 172424 940054 172546 940110
rect 172602 940054 172744 940110
rect 172424 939922 172744 940054
rect 178006 940800 178626 940922
rect 178006 940744 178207 940800
rect 178263 940744 178407 940800
rect 178463 940744 178626 940800
rect 178006 940500 178626 940744
rect 178006 940444 178207 940500
rect 178263 940444 178407 940500
rect 178463 940444 178626 940500
rect 178006 940200 178626 940444
rect 178006 940144 178207 940200
rect 178263 940144 178407 940200
rect 178463 940144 178626 940200
rect 178006 934568 178626 940144
rect 179424 940710 179744 943379
rect 195339 942153 195539 943085
rect 195339 942097 195406 942153
rect 195462 942097 195539 942153
rect 195339 941853 195539 942097
rect 195339 941797 195406 941853
rect 195462 941797 195539 941853
rect 195339 941553 195539 941797
rect 195339 941497 195406 941553
rect 195462 941497 195539 941553
rect 195339 941322 195539 941497
rect 179424 940654 179546 940710
rect 179602 940654 179744 940710
rect 179424 940410 179744 940654
rect 179424 940354 179546 940410
rect 179602 940354 179744 940410
rect 179424 940110 179744 940354
rect 179424 940054 179546 940110
rect 179602 940054 179744 940110
rect 179424 939922 179744 940054
rect 195739 940716 195939 943565
rect 220424 943435 220744 943504
rect 220424 943379 220548 943435
rect 220604 943379 220744 943435
rect 195739 940660 195821 940716
rect 195877 940660 195939 940716
rect 195739 940416 195939 940660
rect 195739 940360 195821 940416
rect 195877 940360 195939 940416
rect 195739 940116 195939 940360
rect 195739 940060 195821 940116
rect 195877 940060 195939 940116
rect 195739 939922 195939 940060
rect 214006 940800 214626 940922
rect 214006 940744 214207 940800
rect 214263 940744 214407 940800
rect 214463 940744 214626 940800
rect 214006 940500 214626 940744
rect 214006 940444 214207 940500
rect 214263 940444 214407 940500
rect 214463 940444 214626 940500
rect 214006 940200 214626 940444
rect 214006 940144 214207 940200
rect 214263 940144 214407 940200
rect 214463 940144 214626 940200
rect 214006 934568 214626 940144
rect 220424 940710 220744 943379
rect 220424 940654 220546 940710
rect 220602 940654 220744 940710
rect 220424 940410 220744 940654
rect 220424 940354 220546 940410
rect 220602 940354 220744 940410
rect 220424 940110 220744 940354
rect 220424 940054 220546 940110
rect 220602 940054 220744 940110
rect 220424 939922 220744 940054
rect 227424 943435 227744 943504
rect 227424 943379 227548 943435
rect 227604 943379 227744 943435
rect 227424 940710 227744 943379
rect 234424 943435 234744 943504
rect 234424 943379 234548 943435
rect 234604 943379 234744 943435
rect 227424 940654 227546 940710
rect 227602 940654 227744 940710
rect 227424 940410 227744 940654
rect 227424 940354 227546 940410
rect 227602 940354 227744 940410
rect 227424 940110 227744 940354
rect 227424 940054 227546 940110
rect 227602 940054 227744 940110
rect 227424 939922 227744 940054
rect 232006 942200 232626 942322
rect 232006 942144 232207 942200
rect 232263 942144 232407 942200
rect 232463 942144 232626 942200
rect 232006 941900 232626 942144
rect 232006 941844 232207 941900
rect 232263 941844 232407 941900
rect 232463 941844 232626 941900
rect 232006 941600 232626 941844
rect 232006 941544 232207 941600
rect 232263 941544 232407 941600
rect 232463 941544 232626 941600
rect 232006 933608 232626 941544
rect 234424 940710 234744 943379
rect 250339 942153 250539 943085
rect 250339 942097 250406 942153
rect 250462 942097 250539 942153
rect 250339 941853 250539 942097
rect 250339 941797 250406 941853
rect 250462 941797 250539 941853
rect 250339 941553 250539 941797
rect 250339 941497 250406 941553
rect 250462 941497 250539 941553
rect 250339 941322 250539 941497
rect 234424 940654 234546 940710
rect 234602 940654 234744 940710
rect 234424 940410 234744 940654
rect 234424 940354 234546 940410
rect 234602 940354 234744 940410
rect 234424 940110 234744 940354
rect 234424 940054 234546 940110
rect 234602 940054 234744 940110
rect 234424 939922 234744 940054
rect 250006 940800 250626 940922
rect 250006 940744 250207 940800
rect 250263 940744 250407 940800
rect 250463 940744 250626 940800
rect 250006 940500 250626 940744
rect 250006 940444 250207 940500
rect 250263 940444 250407 940500
rect 250463 940444 250626 940500
rect 250006 940200 250626 940444
rect 250006 940144 250207 940200
rect 250263 940144 250407 940200
rect 250463 940144 250626 940200
rect 250006 934568 250626 940144
rect 250739 940716 250939 943565
rect 275424 943435 275744 943504
rect 275424 943379 275548 943435
rect 275604 943379 275744 943435
rect 250739 940660 250821 940716
rect 250877 940660 250939 940716
rect 250739 940416 250939 940660
rect 250739 940360 250821 940416
rect 250877 940360 250939 940416
rect 250739 940116 250939 940360
rect 250739 940060 250821 940116
rect 250877 940060 250939 940116
rect 250739 939922 250939 940060
rect 268006 942200 268626 942322
rect 268006 942144 268207 942200
rect 268263 942144 268407 942200
rect 268463 942144 268626 942200
rect 268006 941900 268626 942144
rect 268006 941844 268207 941900
rect 268263 941844 268407 941900
rect 268463 941844 268626 941900
rect 268006 941600 268626 941844
rect 268006 941544 268207 941600
rect 268263 941544 268407 941600
rect 268463 941544 268626 941600
rect 268006 933608 268626 941544
rect 275424 940710 275744 943379
rect 275424 940654 275546 940710
rect 275602 940654 275744 940710
rect 275424 940410 275744 940654
rect 275424 940354 275546 940410
rect 275602 940354 275744 940410
rect 275424 940110 275744 940354
rect 275424 940054 275546 940110
rect 275602 940054 275744 940110
rect 275424 939922 275744 940054
rect 282424 943435 282744 943504
rect 282424 943379 282548 943435
rect 282604 943379 282744 943435
rect 282424 940710 282744 943379
rect 289424 943435 289744 943504
rect 289424 943379 289548 943435
rect 289604 943379 289744 943435
rect 282424 940654 282546 940710
rect 282602 940654 282744 940710
rect 282424 940410 282744 940654
rect 282424 940354 282546 940410
rect 282602 940354 282744 940410
rect 282424 940110 282744 940354
rect 282424 940054 282546 940110
rect 282602 940054 282744 940110
rect 282424 939922 282744 940054
rect 286006 940800 286626 940922
rect 286006 940744 286207 940800
rect 286263 940744 286407 940800
rect 286463 940744 286626 940800
rect 286006 940500 286626 940744
rect 286006 940444 286207 940500
rect 286263 940444 286407 940500
rect 286463 940444 286626 940500
rect 286006 940200 286626 940444
rect 286006 940144 286207 940200
rect 286263 940144 286407 940200
rect 286463 940144 286626 940200
rect 286006 934568 286626 940144
rect 289424 940710 289744 943379
rect 289424 940654 289546 940710
rect 289602 940654 289744 940710
rect 289424 940410 289744 940654
rect 289424 940354 289546 940410
rect 289602 940354 289744 940410
rect 289424 940110 289744 940354
rect 289424 940054 289546 940110
rect 289602 940054 289744 940110
rect 289424 939922 289744 940054
rect 304006 942200 304626 942322
rect 304006 942144 304207 942200
rect 304263 942144 304407 942200
rect 304463 942144 304626 942200
rect 304006 941900 304626 942144
rect 304006 941844 304207 941900
rect 304263 941844 304407 941900
rect 304463 941844 304626 941900
rect 304006 941600 304626 941844
rect 304006 941544 304207 941600
rect 304263 941544 304407 941600
rect 304463 941544 304626 941600
rect 304006 933608 304626 941544
rect 305339 942153 305539 943085
rect 305339 942097 305406 942153
rect 305462 942097 305539 942153
rect 305339 941853 305539 942097
rect 305339 941797 305406 941853
rect 305462 941797 305539 941853
rect 305339 941553 305539 941797
rect 305339 941497 305406 941553
rect 305462 941497 305539 941553
rect 305339 941322 305539 941497
rect 305739 940716 305939 943565
rect 330424 943435 330744 943504
rect 330424 943379 330548 943435
rect 330604 943379 330744 943435
rect 305739 940660 305821 940716
rect 305877 940660 305939 940716
rect 305739 940416 305939 940660
rect 305739 940360 305821 940416
rect 305877 940360 305939 940416
rect 305739 940116 305939 940360
rect 305739 940060 305821 940116
rect 305877 940060 305939 940116
rect 305739 939922 305939 940060
rect 322006 940800 322626 940922
rect 322006 940744 322207 940800
rect 322263 940744 322407 940800
rect 322463 940744 322626 940800
rect 322006 940500 322626 940744
rect 322006 940444 322207 940500
rect 322263 940444 322407 940500
rect 322463 940444 322626 940500
rect 322006 940200 322626 940444
rect 322006 940144 322207 940200
rect 322263 940144 322407 940200
rect 322463 940144 322626 940200
rect 322006 934568 322626 940144
rect 330424 940710 330744 943379
rect 330424 940654 330546 940710
rect 330602 940654 330744 940710
rect 330424 940410 330744 940654
rect 330424 940354 330546 940410
rect 330602 940354 330744 940410
rect 330424 940110 330744 940354
rect 330424 940054 330546 940110
rect 330602 940054 330744 940110
rect 330424 939922 330744 940054
rect 337424 943435 337744 943504
rect 337424 943379 337548 943435
rect 337604 943379 337744 943435
rect 337424 940710 337744 943379
rect 344424 943435 344744 943504
rect 344424 943379 344548 943435
rect 344604 943379 344744 943435
rect 337424 940654 337546 940710
rect 337602 940654 337744 940710
rect 337424 940410 337744 940654
rect 337424 940354 337546 940410
rect 337602 940354 337744 940410
rect 337424 940110 337744 940354
rect 337424 940054 337546 940110
rect 337602 940054 337744 940110
rect 337424 939922 337744 940054
rect 340006 942200 340626 942322
rect 340006 942144 340207 942200
rect 340263 942144 340407 942200
rect 340463 942144 340626 942200
rect 340006 941900 340626 942144
rect 340006 941844 340207 941900
rect 340263 941844 340407 941900
rect 340463 941844 340626 941900
rect 340006 941600 340626 941844
rect 340006 941544 340207 941600
rect 340263 941544 340407 941600
rect 340463 941544 340626 941600
rect 340006 933608 340626 941544
rect 344424 940710 344744 943379
rect 360339 942153 360539 943085
rect 360339 942097 360406 942153
rect 360462 942097 360539 942153
rect 360339 941853 360539 942097
rect 360339 941797 360406 941853
rect 360462 941797 360539 941853
rect 360339 941553 360539 941797
rect 360339 941497 360406 941553
rect 360462 941497 360539 941553
rect 360339 941322 360539 941497
rect 344424 940654 344546 940710
rect 344602 940654 344744 940710
rect 344424 940410 344744 940654
rect 344424 940354 344546 940410
rect 344602 940354 344744 940410
rect 344424 940110 344744 940354
rect 344424 940054 344546 940110
rect 344602 940054 344744 940110
rect 344424 939922 344744 940054
rect 358006 940800 358626 940922
rect 358006 940744 358207 940800
rect 358263 940744 358407 940800
rect 358463 940744 358626 940800
rect 358006 940500 358626 940744
rect 358006 940444 358207 940500
rect 358263 940444 358407 940500
rect 358463 940444 358626 940500
rect 358006 940200 358626 940444
rect 358006 940144 358207 940200
rect 358263 940144 358407 940200
rect 358463 940144 358626 940200
rect 358006 934568 358626 940144
rect 360739 940716 360939 943565
rect 360739 940660 360821 940716
rect 360877 940660 360939 940716
rect 360739 940416 360939 940660
rect 360739 940360 360821 940416
rect 360877 940360 360939 940416
rect 360739 940116 360939 940360
rect 360739 940060 360821 940116
rect 360877 940060 360939 940116
rect 360739 939922 360939 940060
rect 376006 942200 376626 942322
rect 376006 942144 376207 942200
rect 376263 942144 376407 942200
rect 376463 942144 376626 942200
rect 376006 941900 376626 942144
rect 376006 941844 376207 941900
rect 376263 941844 376407 941900
rect 376463 941844 376626 941900
rect 376006 941600 376626 941844
rect 376006 941544 376207 941600
rect 376263 941544 376407 941600
rect 376463 941544 376626 941600
rect 376006 933608 376626 941544
rect 381272 940792 383172 949870
rect 381272 940736 381348 940792
rect 381404 940736 381472 940792
rect 381528 940736 381596 940792
rect 381652 940736 381720 940792
rect 381776 940736 381844 940792
rect 381900 940736 381968 940792
rect 382024 940736 382092 940792
rect 382148 940736 382216 940792
rect 382272 940736 382340 940792
rect 382396 940736 382464 940792
rect 382520 940736 382588 940792
rect 382644 940736 382712 940792
rect 382768 940736 382836 940792
rect 382892 940736 382960 940792
rect 383016 940736 383084 940792
rect 383140 940736 383172 940792
rect 381272 940668 383172 940736
rect 381272 940612 381348 940668
rect 381404 940612 381472 940668
rect 381528 940612 381596 940668
rect 381652 940612 381720 940668
rect 381776 940612 381844 940668
rect 381900 940612 381968 940668
rect 382024 940612 382092 940668
rect 382148 940612 382216 940668
rect 382272 940612 382340 940668
rect 382396 940612 382464 940668
rect 382520 940612 382588 940668
rect 382644 940612 382712 940668
rect 382768 940612 382836 940668
rect 382892 940612 382960 940668
rect 383016 940612 383084 940668
rect 383140 940612 383172 940668
rect 381272 940544 383172 940612
rect 381272 940488 381348 940544
rect 381404 940488 381472 940544
rect 381528 940488 381596 940544
rect 381652 940488 381720 940544
rect 381776 940488 381844 940544
rect 381900 940488 381968 940544
rect 382024 940488 382092 940544
rect 382148 940488 382216 940544
rect 382272 940488 382340 940544
rect 382396 940488 382464 940544
rect 382520 940488 382588 940544
rect 382644 940488 382712 940544
rect 382768 940488 382836 940544
rect 382892 940488 382960 940544
rect 383016 940488 383084 940544
rect 383140 940488 383172 940544
rect 381272 940420 383172 940488
rect 381272 940364 381348 940420
rect 381404 940364 381472 940420
rect 381528 940364 381596 940420
rect 381652 940364 381720 940420
rect 381776 940364 381844 940420
rect 381900 940364 381968 940420
rect 382024 940364 382092 940420
rect 382148 940364 382216 940420
rect 382272 940364 382340 940420
rect 382396 940364 382464 940420
rect 382520 940364 382588 940420
rect 382644 940364 382712 940420
rect 382768 940364 382836 940420
rect 382892 940364 382960 940420
rect 383016 940364 383084 940420
rect 383140 940364 383172 940420
rect 381272 940296 383172 940364
rect 381272 940240 381348 940296
rect 381404 940240 381472 940296
rect 381528 940240 381596 940296
rect 381652 940240 381720 940296
rect 381776 940240 381844 940296
rect 381900 940240 381968 940296
rect 382024 940240 382092 940296
rect 382148 940240 382216 940296
rect 382272 940240 382340 940296
rect 382396 940240 382464 940296
rect 382520 940240 382588 940296
rect 382644 940240 382712 940296
rect 382768 940240 382836 940296
rect 382892 940240 382960 940296
rect 383016 940240 383084 940296
rect 383140 940240 383172 940296
rect 381272 940172 383172 940240
rect 381272 940116 381348 940172
rect 381404 940116 381472 940172
rect 381528 940116 381596 940172
rect 381652 940116 381720 940172
rect 381776 940116 381844 940172
rect 381900 940116 381968 940172
rect 382024 940116 382092 940172
rect 382148 940116 382216 940172
rect 382272 940116 382340 940172
rect 382396 940116 382464 940172
rect 382520 940116 382588 940172
rect 382644 940116 382712 940172
rect 382768 940116 382836 940172
rect 382892 940116 382960 940172
rect 383016 940116 383084 940172
rect 383140 940116 383172 940172
rect 381272 940048 383172 940116
rect 381272 939992 381348 940048
rect 381404 939992 381472 940048
rect 381528 939992 381596 940048
rect 381652 939992 381720 940048
rect 381776 939992 381844 940048
rect 381900 939992 381968 940048
rect 382024 939992 382092 940048
rect 382148 939992 382216 940048
rect 382272 939992 382340 940048
rect 382396 939992 382464 940048
rect 382520 939992 382588 940048
rect 382644 939992 382712 940048
rect 382768 939992 382836 940048
rect 382892 939992 382960 940048
rect 383016 939992 383084 940048
rect 383140 939992 383172 940048
rect 381272 939922 383172 939992
rect 383752 949926 385802 950000
rect 383752 949870 383822 949926
rect 383878 949870 383946 949926
rect 384002 949870 384070 949926
rect 384126 949870 384194 949926
rect 384250 949870 384318 949926
rect 384374 949870 384442 949926
rect 384498 949870 384566 949926
rect 384622 949870 384690 949926
rect 384746 949870 384814 949926
rect 384870 949870 384938 949926
rect 384994 949870 385062 949926
rect 385118 949870 385186 949926
rect 385242 949870 385310 949926
rect 385366 949870 385434 949926
rect 385490 949870 385558 949926
rect 385614 949870 385682 949926
rect 385738 949870 385802 949926
rect 383752 940792 385802 949870
rect 383752 940736 383828 940792
rect 383884 940736 383952 940792
rect 384008 940736 384076 940792
rect 384132 940736 384200 940792
rect 384256 940736 384324 940792
rect 384380 940736 384448 940792
rect 384504 940736 384572 940792
rect 384628 940736 384696 940792
rect 384752 940736 384820 940792
rect 384876 940736 384944 940792
rect 385000 940736 385068 940792
rect 385124 940736 385192 940792
rect 385248 940736 385316 940792
rect 385372 940736 385440 940792
rect 385496 940736 385564 940792
rect 385620 940736 385688 940792
rect 385744 940736 385802 940792
rect 383752 940668 385802 940736
rect 383752 940612 383828 940668
rect 383884 940612 383952 940668
rect 384008 940612 384076 940668
rect 384132 940612 384200 940668
rect 384256 940612 384324 940668
rect 384380 940612 384448 940668
rect 384504 940612 384572 940668
rect 384628 940612 384696 940668
rect 384752 940612 384820 940668
rect 384876 940612 384944 940668
rect 385000 940612 385068 940668
rect 385124 940612 385192 940668
rect 385248 940612 385316 940668
rect 385372 940612 385440 940668
rect 385496 940612 385564 940668
rect 385620 940612 385688 940668
rect 385744 940612 385802 940668
rect 383752 940544 385802 940612
rect 383752 940488 383828 940544
rect 383884 940488 383952 940544
rect 384008 940488 384076 940544
rect 384132 940488 384200 940544
rect 384256 940488 384324 940544
rect 384380 940488 384448 940544
rect 384504 940488 384572 940544
rect 384628 940488 384696 940544
rect 384752 940488 384820 940544
rect 384876 940488 384944 940544
rect 385000 940488 385068 940544
rect 385124 940488 385192 940544
rect 385248 940488 385316 940544
rect 385372 940488 385440 940544
rect 385496 940488 385564 940544
rect 385620 940488 385688 940544
rect 385744 940488 385802 940544
rect 383752 940420 385802 940488
rect 383752 940364 383828 940420
rect 383884 940364 383952 940420
rect 384008 940364 384076 940420
rect 384132 940364 384200 940420
rect 384256 940364 384324 940420
rect 384380 940364 384448 940420
rect 384504 940364 384572 940420
rect 384628 940364 384696 940420
rect 384752 940364 384820 940420
rect 384876 940364 384944 940420
rect 385000 940364 385068 940420
rect 385124 940364 385192 940420
rect 385248 940364 385316 940420
rect 385372 940364 385440 940420
rect 385496 940364 385564 940420
rect 385620 940364 385688 940420
rect 385744 940364 385802 940420
rect 383752 940296 385802 940364
rect 383752 940240 383828 940296
rect 383884 940240 383952 940296
rect 384008 940240 384076 940296
rect 384132 940240 384200 940296
rect 384256 940240 384324 940296
rect 384380 940240 384448 940296
rect 384504 940240 384572 940296
rect 384628 940240 384696 940296
rect 384752 940240 384820 940296
rect 384876 940240 384944 940296
rect 385000 940240 385068 940296
rect 385124 940240 385192 940296
rect 385248 940240 385316 940296
rect 385372 940240 385440 940296
rect 385496 940240 385564 940296
rect 385620 940240 385688 940296
rect 385744 940240 385802 940296
rect 383752 940172 385802 940240
rect 383752 940116 383828 940172
rect 383884 940116 383952 940172
rect 384008 940116 384076 940172
rect 384132 940116 384200 940172
rect 384256 940116 384324 940172
rect 384380 940116 384448 940172
rect 384504 940116 384572 940172
rect 384628 940116 384696 940172
rect 384752 940116 384820 940172
rect 384876 940116 384944 940172
rect 385000 940116 385068 940172
rect 385124 940116 385192 940172
rect 385248 940116 385316 940172
rect 385372 940116 385440 940172
rect 385496 940116 385564 940172
rect 385620 940116 385688 940172
rect 385744 940116 385802 940172
rect 383752 940048 385802 940116
rect 383752 939992 383828 940048
rect 383884 939992 383952 940048
rect 384008 939992 384076 940048
rect 384132 939992 384200 940048
rect 384256 939992 384324 940048
rect 384380 939992 384448 940048
rect 384504 939992 384572 940048
rect 384628 939992 384696 940048
rect 384752 939992 384820 940048
rect 384876 939992 384944 940048
rect 385000 939992 385068 940048
rect 385124 939992 385192 940048
rect 385248 939992 385316 940048
rect 385372 939992 385440 940048
rect 385496 939992 385564 940048
rect 385620 939992 385688 940048
rect 385744 939992 385802 940048
rect 383752 939922 385802 939992
rect 386122 949926 388172 950000
rect 386122 949870 386192 949926
rect 386248 949870 386316 949926
rect 386372 949870 386440 949926
rect 386496 949870 386564 949926
rect 386620 949870 386688 949926
rect 386744 949870 386812 949926
rect 386868 949870 386936 949926
rect 386992 949870 387060 949926
rect 387116 949870 387184 949926
rect 387240 949870 387308 949926
rect 387364 949870 387432 949926
rect 387488 949870 387556 949926
rect 387612 949870 387680 949926
rect 387736 949870 387804 949926
rect 387860 949870 387928 949926
rect 387984 949870 388052 949926
rect 388108 949870 388172 949926
rect 386122 940792 388172 949870
rect 386122 940736 386198 940792
rect 386254 940736 386322 940792
rect 386378 940736 386446 940792
rect 386502 940736 386570 940792
rect 386626 940736 386694 940792
rect 386750 940736 386818 940792
rect 386874 940736 386942 940792
rect 386998 940736 387066 940792
rect 387122 940736 387190 940792
rect 387246 940736 387314 940792
rect 387370 940736 387438 940792
rect 387494 940736 387562 940792
rect 387618 940736 387686 940792
rect 387742 940736 387810 940792
rect 387866 940736 387934 940792
rect 387990 940736 388058 940792
rect 388114 940736 388172 940792
rect 386122 940668 388172 940736
rect 386122 940612 386198 940668
rect 386254 940612 386322 940668
rect 386378 940612 386446 940668
rect 386502 940612 386570 940668
rect 386626 940612 386694 940668
rect 386750 940612 386818 940668
rect 386874 940612 386942 940668
rect 386998 940612 387066 940668
rect 387122 940612 387190 940668
rect 387246 940612 387314 940668
rect 387370 940612 387438 940668
rect 387494 940612 387562 940668
rect 387618 940612 387686 940668
rect 387742 940612 387810 940668
rect 387866 940612 387934 940668
rect 387990 940612 388058 940668
rect 388114 940612 388172 940668
rect 386122 940544 388172 940612
rect 386122 940488 386198 940544
rect 386254 940488 386322 940544
rect 386378 940488 386446 940544
rect 386502 940488 386570 940544
rect 386626 940488 386694 940544
rect 386750 940488 386818 940544
rect 386874 940488 386942 940544
rect 386998 940488 387066 940544
rect 387122 940488 387190 940544
rect 387246 940488 387314 940544
rect 387370 940488 387438 940544
rect 387494 940488 387562 940544
rect 387618 940488 387686 940544
rect 387742 940488 387810 940544
rect 387866 940488 387934 940544
rect 387990 940488 388058 940544
rect 388114 940488 388172 940544
rect 386122 940420 388172 940488
rect 386122 940364 386198 940420
rect 386254 940364 386322 940420
rect 386378 940364 386446 940420
rect 386502 940364 386570 940420
rect 386626 940364 386694 940420
rect 386750 940364 386818 940420
rect 386874 940364 386942 940420
rect 386998 940364 387066 940420
rect 387122 940364 387190 940420
rect 387246 940364 387314 940420
rect 387370 940364 387438 940420
rect 387494 940364 387562 940420
rect 387618 940364 387686 940420
rect 387742 940364 387810 940420
rect 387866 940364 387934 940420
rect 387990 940364 388058 940420
rect 388114 940364 388172 940420
rect 386122 940296 388172 940364
rect 386122 940240 386198 940296
rect 386254 940240 386322 940296
rect 386378 940240 386446 940296
rect 386502 940240 386570 940296
rect 386626 940240 386694 940296
rect 386750 940240 386818 940296
rect 386874 940240 386942 940296
rect 386998 940240 387066 940296
rect 387122 940240 387190 940296
rect 387246 940240 387314 940296
rect 387370 940240 387438 940296
rect 387494 940240 387562 940296
rect 387618 940240 387686 940296
rect 387742 940240 387810 940296
rect 387866 940240 387934 940296
rect 387990 940240 388058 940296
rect 388114 940240 388172 940296
rect 386122 940172 388172 940240
rect 386122 940116 386198 940172
rect 386254 940116 386322 940172
rect 386378 940116 386446 940172
rect 386502 940116 386570 940172
rect 386626 940116 386694 940172
rect 386750 940116 386818 940172
rect 386874 940116 386942 940172
rect 386998 940116 387066 940172
rect 387122 940116 387190 940172
rect 387246 940116 387314 940172
rect 387370 940116 387438 940172
rect 387494 940116 387562 940172
rect 387618 940116 387686 940172
rect 387742 940116 387810 940172
rect 387866 940116 387934 940172
rect 387990 940116 388058 940172
rect 388114 940116 388172 940172
rect 386122 940048 388172 940116
rect 386122 939992 386198 940048
rect 386254 939992 386322 940048
rect 386378 939992 386446 940048
rect 386502 939992 386570 940048
rect 386626 939992 386694 940048
rect 386750 939992 386818 940048
rect 386874 939992 386942 940048
rect 386998 939992 387066 940048
rect 387122 939992 387190 940048
rect 387246 939992 387314 940048
rect 387370 939992 387438 940048
rect 387494 939992 387562 940048
rect 387618 939992 387686 940048
rect 387742 939992 387810 940048
rect 387866 939992 387934 940048
rect 387990 939992 388058 940048
rect 388114 939992 388172 940048
rect 386122 939922 388172 939992
rect 388828 949926 390878 950000
rect 388828 949870 388892 949926
rect 388948 949870 389016 949926
rect 389072 949870 389140 949926
rect 389196 949870 389264 949926
rect 389320 949870 389388 949926
rect 389444 949870 389512 949926
rect 389568 949870 389636 949926
rect 389692 949870 389760 949926
rect 389816 949870 389884 949926
rect 389940 949870 390008 949926
rect 390064 949870 390132 949926
rect 390188 949870 390256 949926
rect 390312 949870 390380 949926
rect 390436 949870 390504 949926
rect 390560 949870 390628 949926
rect 390684 949870 390752 949926
rect 390808 949870 390878 949926
rect 388828 940792 390878 949870
rect 388828 940736 388904 940792
rect 388960 940736 389028 940792
rect 389084 940736 389152 940792
rect 389208 940736 389276 940792
rect 389332 940736 389400 940792
rect 389456 940736 389524 940792
rect 389580 940736 389648 940792
rect 389704 940736 389772 940792
rect 389828 940736 389896 940792
rect 389952 940736 390020 940792
rect 390076 940736 390144 940792
rect 390200 940736 390268 940792
rect 390324 940736 390392 940792
rect 390448 940736 390516 940792
rect 390572 940736 390640 940792
rect 390696 940736 390764 940792
rect 390820 940736 390878 940792
rect 388828 940668 390878 940736
rect 388828 940612 388904 940668
rect 388960 940612 389028 940668
rect 389084 940612 389152 940668
rect 389208 940612 389276 940668
rect 389332 940612 389400 940668
rect 389456 940612 389524 940668
rect 389580 940612 389648 940668
rect 389704 940612 389772 940668
rect 389828 940612 389896 940668
rect 389952 940612 390020 940668
rect 390076 940612 390144 940668
rect 390200 940612 390268 940668
rect 390324 940612 390392 940668
rect 390448 940612 390516 940668
rect 390572 940612 390640 940668
rect 390696 940612 390764 940668
rect 390820 940612 390878 940668
rect 388828 940544 390878 940612
rect 388828 940488 388904 940544
rect 388960 940488 389028 940544
rect 389084 940488 389152 940544
rect 389208 940488 389276 940544
rect 389332 940488 389400 940544
rect 389456 940488 389524 940544
rect 389580 940488 389648 940544
rect 389704 940488 389772 940544
rect 389828 940488 389896 940544
rect 389952 940488 390020 940544
rect 390076 940488 390144 940544
rect 390200 940488 390268 940544
rect 390324 940488 390392 940544
rect 390448 940488 390516 940544
rect 390572 940488 390640 940544
rect 390696 940488 390764 940544
rect 390820 940488 390878 940544
rect 388828 940420 390878 940488
rect 388828 940364 388904 940420
rect 388960 940364 389028 940420
rect 389084 940364 389152 940420
rect 389208 940364 389276 940420
rect 389332 940364 389400 940420
rect 389456 940364 389524 940420
rect 389580 940364 389648 940420
rect 389704 940364 389772 940420
rect 389828 940364 389896 940420
rect 389952 940364 390020 940420
rect 390076 940364 390144 940420
rect 390200 940364 390268 940420
rect 390324 940364 390392 940420
rect 390448 940364 390516 940420
rect 390572 940364 390640 940420
rect 390696 940364 390764 940420
rect 390820 940364 390878 940420
rect 388828 940296 390878 940364
rect 388828 940240 388904 940296
rect 388960 940240 389028 940296
rect 389084 940240 389152 940296
rect 389208 940240 389276 940296
rect 389332 940240 389400 940296
rect 389456 940240 389524 940296
rect 389580 940240 389648 940296
rect 389704 940240 389772 940296
rect 389828 940240 389896 940296
rect 389952 940240 390020 940296
rect 390076 940240 390144 940296
rect 390200 940240 390268 940296
rect 390324 940240 390392 940296
rect 390448 940240 390516 940296
rect 390572 940240 390640 940296
rect 390696 940240 390764 940296
rect 390820 940240 390878 940296
rect 388828 940172 390878 940240
rect 388828 940116 388904 940172
rect 388960 940116 389028 940172
rect 389084 940116 389152 940172
rect 389208 940116 389276 940172
rect 389332 940116 389400 940172
rect 389456 940116 389524 940172
rect 389580 940116 389648 940172
rect 389704 940116 389772 940172
rect 389828 940116 389896 940172
rect 389952 940116 390020 940172
rect 390076 940116 390144 940172
rect 390200 940116 390268 940172
rect 390324 940116 390392 940172
rect 390448 940116 390516 940172
rect 390572 940116 390640 940172
rect 390696 940116 390764 940172
rect 390820 940116 390878 940172
rect 388828 940048 390878 940116
rect 388828 939992 388904 940048
rect 388960 939992 389028 940048
rect 389084 939992 389152 940048
rect 389208 939992 389276 940048
rect 389332 939992 389400 940048
rect 389456 939992 389524 940048
rect 389580 939992 389648 940048
rect 389704 939992 389772 940048
rect 389828 939992 389896 940048
rect 389952 939992 390020 940048
rect 390076 939992 390144 940048
rect 390200 939992 390268 940048
rect 390324 939992 390392 940048
rect 390448 939992 390516 940048
rect 390572 939992 390640 940048
rect 390696 939992 390764 940048
rect 390820 939992 390878 940048
rect 388828 939922 390878 939992
rect 391198 949926 393248 950000
rect 391198 949870 391262 949926
rect 391318 949870 391386 949926
rect 391442 949870 391510 949926
rect 391566 949870 391634 949926
rect 391690 949870 391758 949926
rect 391814 949870 391882 949926
rect 391938 949870 392006 949926
rect 392062 949870 392130 949926
rect 392186 949870 392254 949926
rect 392310 949870 392378 949926
rect 392434 949870 392502 949926
rect 392558 949870 392626 949926
rect 392682 949870 392750 949926
rect 392806 949870 392874 949926
rect 392930 949870 392998 949926
rect 393054 949870 393122 949926
rect 393178 949870 393248 949926
rect 391198 940792 393248 949870
rect 391198 940736 391274 940792
rect 391330 940736 391398 940792
rect 391454 940736 391522 940792
rect 391578 940736 391646 940792
rect 391702 940736 391770 940792
rect 391826 940736 391894 940792
rect 391950 940736 392018 940792
rect 392074 940736 392142 940792
rect 392198 940736 392266 940792
rect 392322 940736 392390 940792
rect 392446 940736 392514 940792
rect 392570 940736 392638 940792
rect 392694 940736 392762 940792
rect 392818 940736 392886 940792
rect 392942 940736 393010 940792
rect 393066 940736 393134 940792
rect 393190 940736 393248 940792
rect 391198 940668 393248 940736
rect 391198 940612 391274 940668
rect 391330 940612 391398 940668
rect 391454 940612 391522 940668
rect 391578 940612 391646 940668
rect 391702 940612 391770 940668
rect 391826 940612 391894 940668
rect 391950 940612 392018 940668
rect 392074 940612 392142 940668
rect 392198 940612 392266 940668
rect 392322 940612 392390 940668
rect 392446 940612 392514 940668
rect 392570 940612 392638 940668
rect 392694 940612 392762 940668
rect 392818 940612 392886 940668
rect 392942 940612 393010 940668
rect 393066 940612 393134 940668
rect 393190 940612 393248 940668
rect 391198 940544 393248 940612
rect 391198 940488 391274 940544
rect 391330 940488 391398 940544
rect 391454 940488 391522 940544
rect 391578 940488 391646 940544
rect 391702 940488 391770 940544
rect 391826 940488 391894 940544
rect 391950 940488 392018 940544
rect 392074 940488 392142 940544
rect 392198 940488 392266 940544
rect 392322 940488 392390 940544
rect 392446 940488 392514 940544
rect 392570 940488 392638 940544
rect 392694 940488 392762 940544
rect 392818 940488 392886 940544
rect 392942 940488 393010 940544
rect 393066 940488 393134 940544
rect 393190 940488 393248 940544
rect 391198 940420 393248 940488
rect 391198 940364 391274 940420
rect 391330 940364 391398 940420
rect 391454 940364 391522 940420
rect 391578 940364 391646 940420
rect 391702 940364 391770 940420
rect 391826 940364 391894 940420
rect 391950 940364 392018 940420
rect 392074 940364 392142 940420
rect 392198 940364 392266 940420
rect 392322 940364 392390 940420
rect 392446 940364 392514 940420
rect 392570 940364 392638 940420
rect 392694 940364 392762 940420
rect 392818 940364 392886 940420
rect 392942 940364 393010 940420
rect 393066 940364 393134 940420
rect 393190 940364 393248 940420
rect 391198 940296 393248 940364
rect 391198 940240 391274 940296
rect 391330 940240 391398 940296
rect 391454 940240 391522 940296
rect 391578 940240 391646 940296
rect 391702 940240 391770 940296
rect 391826 940240 391894 940296
rect 391950 940240 392018 940296
rect 392074 940240 392142 940296
rect 392198 940240 392266 940296
rect 392322 940240 392390 940296
rect 392446 940240 392514 940296
rect 392570 940240 392638 940296
rect 392694 940240 392762 940296
rect 392818 940240 392886 940296
rect 392942 940240 393010 940296
rect 393066 940240 393134 940296
rect 393190 940240 393248 940296
rect 391198 940172 393248 940240
rect 391198 940116 391274 940172
rect 391330 940116 391398 940172
rect 391454 940116 391522 940172
rect 391578 940116 391646 940172
rect 391702 940116 391770 940172
rect 391826 940116 391894 940172
rect 391950 940116 392018 940172
rect 392074 940116 392142 940172
rect 392198 940116 392266 940172
rect 392322 940116 392390 940172
rect 392446 940116 392514 940172
rect 392570 940116 392638 940172
rect 392694 940116 392762 940172
rect 392818 940116 392886 940172
rect 392942 940116 393010 940172
rect 393066 940116 393134 940172
rect 393190 940116 393248 940172
rect 391198 940048 393248 940116
rect 391198 939992 391274 940048
rect 391330 939992 391398 940048
rect 391454 939992 391522 940048
rect 391578 939992 391646 940048
rect 391702 939992 391770 940048
rect 391826 939992 391894 940048
rect 391950 939992 392018 940048
rect 392074 939992 392142 940048
rect 392198 939992 392266 940048
rect 392322 939992 392390 940048
rect 392446 939992 392514 940048
rect 392570 939992 392638 940048
rect 392694 939992 392762 940048
rect 392818 939992 392886 940048
rect 392942 939992 393010 940048
rect 393066 939992 393134 940048
rect 393190 939992 393248 940048
rect 391198 939922 393248 939992
rect 393828 949926 395728 950000
rect 393828 949870 393866 949926
rect 393922 949870 393990 949926
rect 394046 949870 394114 949926
rect 394170 949870 394238 949926
rect 394294 949870 394362 949926
rect 394418 949870 394486 949926
rect 394542 949870 394610 949926
rect 394666 949870 394734 949926
rect 394790 949870 394858 949926
rect 394914 949870 394982 949926
rect 395038 949870 395106 949926
rect 395162 949870 395230 949926
rect 395286 949870 395354 949926
rect 395410 949870 395478 949926
rect 395534 949870 395602 949926
rect 395658 949870 395728 949926
rect 393828 940792 395728 949870
rect 601272 949926 603172 950000
rect 601272 949870 601342 949926
rect 601398 949870 601466 949926
rect 601522 949870 601590 949926
rect 601646 949870 601714 949926
rect 601770 949870 601838 949926
rect 601894 949870 601962 949926
rect 602018 949870 602086 949926
rect 602142 949870 602210 949926
rect 602266 949870 602334 949926
rect 602390 949870 602458 949926
rect 602514 949870 602582 949926
rect 602638 949870 602706 949926
rect 602762 949870 602830 949926
rect 602886 949870 602954 949926
rect 603010 949870 603078 949926
rect 603134 949870 603172 949926
rect 470339 943565 470939 943885
rect 525339 943565 525939 943885
rect 580339 943565 580939 943885
rect 440424 943435 440744 943504
rect 440424 943379 440548 943435
rect 440604 943379 440744 943435
rect 393828 940736 393878 940792
rect 393934 940736 394002 940792
rect 394058 940736 394126 940792
rect 394182 940736 394250 940792
rect 394306 940736 394374 940792
rect 394430 940736 394498 940792
rect 394554 940736 394622 940792
rect 394678 940736 394746 940792
rect 394802 940736 394870 940792
rect 394926 940736 394994 940792
rect 395050 940736 395118 940792
rect 395174 940736 395242 940792
rect 395298 940736 395366 940792
rect 395422 940736 395490 940792
rect 395546 940736 395614 940792
rect 395670 940736 395728 940792
rect 393828 940668 395728 940736
rect 393828 940612 393878 940668
rect 393934 940612 394002 940668
rect 394058 940612 394126 940668
rect 394182 940612 394250 940668
rect 394306 940612 394374 940668
rect 394430 940612 394498 940668
rect 394554 940612 394622 940668
rect 394678 940612 394746 940668
rect 394802 940612 394870 940668
rect 394926 940612 394994 940668
rect 395050 940612 395118 940668
rect 395174 940612 395242 940668
rect 395298 940612 395366 940668
rect 395422 940612 395490 940668
rect 395546 940612 395614 940668
rect 395670 940612 395728 940668
rect 393828 940544 395728 940612
rect 393828 940488 393878 940544
rect 393934 940488 394002 940544
rect 394058 940488 394126 940544
rect 394182 940488 394250 940544
rect 394306 940488 394374 940544
rect 394430 940488 394498 940544
rect 394554 940488 394622 940544
rect 394678 940488 394746 940544
rect 394802 940488 394870 940544
rect 394926 940488 394994 940544
rect 395050 940488 395118 940544
rect 395174 940488 395242 940544
rect 395298 940488 395366 940544
rect 395422 940488 395490 940544
rect 395546 940488 395614 940544
rect 395670 940488 395728 940544
rect 393828 940420 395728 940488
rect 393828 940364 393878 940420
rect 393934 940364 394002 940420
rect 394058 940364 394126 940420
rect 394182 940364 394250 940420
rect 394306 940364 394374 940420
rect 394430 940364 394498 940420
rect 394554 940364 394622 940420
rect 394678 940364 394746 940420
rect 394802 940364 394870 940420
rect 394926 940364 394994 940420
rect 395050 940364 395118 940420
rect 395174 940364 395242 940420
rect 395298 940364 395366 940420
rect 395422 940364 395490 940420
rect 395546 940364 395614 940420
rect 395670 940364 395728 940420
rect 393828 940296 395728 940364
rect 393828 940240 393878 940296
rect 393934 940240 394002 940296
rect 394058 940240 394126 940296
rect 394182 940240 394250 940296
rect 394306 940240 394374 940296
rect 394430 940240 394498 940296
rect 394554 940240 394622 940296
rect 394678 940240 394746 940296
rect 394802 940240 394870 940296
rect 394926 940240 394994 940296
rect 395050 940240 395118 940296
rect 395174 940240 395242 940296
rect 395298 940240 395366 940296
rect 395422 940240 395490 940296
rect 395546 940240 395614 940296
rect 395670 940240 395728 940296
rect 393828 940172 395728 940240
rect 393828 940116 393878 940172
rect 393934 940116 394002 940172
rect 394058 940116 394126 940172
rect 394182 940116 394250 940172
rect 394306 940116 394374 940172
rect 394430 940116 394498 940172
rect 394554 940116 394622 940172
rect 394678 940116 394746 940172
rect 394802 940116 394870 940172
rect 394926 940116 394994 940172
rect 395050 940116 395118 940172
rect 395174 940116 395242 940172
rect 395298 940116 395366 940172
rect 395422 940116 395490 940172
rect 395546 940116 395614 940172
rect 395670 940116 395728 940172
rect 393828 940048 395728 940116
rect 393828 939992 393878 940048
rect 393934 939992 394002 940048
rect 394058 939992 394126 940048
rect 394182 939992 394250 940048
rect 394306 939992 394374 940048
rect 394430 939992 394498 940048
rect 394554 939992 394622 940048
rect 394678 939992 394746 940048
rect 394802 939992 394870 940048
rect 394926 939992 394994 940048
rect 395050 939992 395118 940048
rect 395174 939992 395242 940048
rect 395298 939992 395366 940048
rect 395422 939992 395490 940048
rect 395546 939992 395614 940048
rect 395670 939992 395728 940048
rect 393828 939922 395728 939992
rect 412006 942200 412626 942322
rect 412006 942144 412207 942200
rect 412263 942144 412407 942200
rect 412463 942144 412626 942200
rect 412006 941900 412626 942144
rect 412006 941844 412207 941900
rect 412263 941844 412407 941900
rect 412463 941844 412626 941900
rect 412006 941600 412626 941844
rect 412006 941544 412207 941600
rect 412263 941544 412407 941600
rect 412463 941544 412626 941600
rect 394006 934568 394626 939922
rect 412006 933608 412626 941544
rect 430006 940800 430626 940922
rect 430006 940744 430207 940800
rect 430263 940744 430407 940800
rect 430463 940744 430626 940800
rect 430006 940500 430626 940744
rect 430006 940444 430207 940500
rect 430263 940444 430407 940500
rect 430463 940444 430626 940500
rect 430006 940200 430626 940444
rect 430006 940144 430207 940200
rect 430263 940144 430407 940200
rect 430463 940144 430626 940200
rect 430006 934568 430626 940144
rect 440424 940710 440744 943379
rect 440424 940654 440546 940710
rect 440602 940654 440744 940710
rect 440424 940410 440744 940654
rect 440424 940354 440546 940410
rect 440602 940354 440744 940410
rect 440424 940110 440744 940354
rect 440424 940054 440546 940110
rect 440602 940054 440744 940110
rect 440424 939922 440744 940054
rect 447424 943435 447744 943504
rect 447424 943379 447548 943435
rect 447604 943379 447744 943435
rect 447424 940710 447744 943379
rect 454424 943435 454744 943504
rect 454424 943379 454548 943435
rect 454604 943379 454744 943435
rect 447424 940654 447546 940710
rect 447602 940654 447744 940710
rect 447424 940410 447744 940654
rect 447424 940354 447546 940410
rect 447602 940354 447744 940410
rect 447424 940110 447744 940354
rect 447424 940054 447546 940110
rect 447602 940054 447744 940110
rect 447424 939922 447744 940054
rect 448006 942200 448626 942322
rect 448006 942144 448207 942200
rect 448263 942144 448407 942200
rect 448463 942144 448626 942200
rect 448006 941900 448626 942144
rect 448006 941844 448207 941900
rect 448263 941844 448407 941900
rect 448463 941844 448626 941900
rect 448006 941600 448626 941844
rect 448006 941544 448207 941600
rect 448263 941544 448407 941600
rect 448463 941544 448626 941600
rect 448006 933608 448626 941544
rect 454424 940710 454744 943379
rect 470339 942153 470539 943085
rect 470339 942097 470406 942153
rect 470462 942097 470539 942153
rect 470339 941853 470539 942097
rect 470339 941797 470406 941853
rect 470462 941797 470539 941853
rect 470339 941553 470539 941797
rect 470339 941497 470406 941553
rect 470462 941497 470539 941553
rect 470339 941322 470539 941497
rect 454424 940654 454546 940710
rect 454602 940654 454744 940710
rect 454424 940410 454744 940654
rect 454424 940354 454546 940410
rect 454602 940354 454744 940410
rect 454424 940110 454744 940354
rect 454424 940054 454546 940110
rect 454602 940054 454744 940110
rect 454424 939922 454744 940054
rect 466006 940800 466626 940922
rect 466006 940744 466207 940800
rect 466263 940744 466407 940800
rect 466463 940744 466626 940800
rect 466006 940500 466626 940744
rect 466006 940444 466207 940500
rect 466263 940444 466407 940500
rect 466463 940444 466626 940500
rect 466006 940200 466626 940444
rect 466006 940144 466207 940200
rect 466263 940144 466407 940200
rect 466463 940144 466626 940200
rect 466006 934568 466626 940144
rect 470739 940716 470939 943565
rect 495424 943435 495744 943504
rect 495424 943379 495548 943435
rect 495604 943379 495744 943435
rect 470739 940660 470821 940716
rect 470877 940660 470939 940716
rect 470739 940416 470939 940660
rect 470739 940360 470821 940416
rect 470877 940360 470939 940416
rect 470739 940116 470939 940360
rect 470739 940060 470821 940116
rect 470877 940060 470939 940116
rect 470739 939922 470939 940060
rect 484006 942200 484626 942322
rect 484006 942144 484207 942200
rect 484263 942144 484407 942200
rect 484463 942144 484626 942200
rect 484006 941900 484626 942144
rect 484006 941844 484207 941900
rect 484263 941844 484407 941900
rect 484463 941844 484626 941900
rect 484006 941600 484626 941844
rect 484006 941544 484207 941600
rect 484263 941544 484407 941600
rect 484463 941544 484626 941600
rect 484006 933608 484626 941544
rect 495424 940710 495744 943379
rect 502424 943435 502744 943504
rect 502424 943379 502548 943435
rect 502604 943379 502744 943435
rect 502424 940922 502744 943379
rect 495424 940654 495546 940710
rect 495602 940654 495744 940710
rect 495424 940410 495744 940654
rect 495424 940354 495546 940410
rect 495602 940354 495744 940410
rect 495424 940110 495744 940354
rect 495424 940054 495546 940110
rect 495602 940054 495744 940110
rect 495424 939922 495744 940054
rect 502006 940800 502744 940922
rect 502006 940744 502207 940800
rect 502263 940744 502407 940800
rect 502463 940744 502744 940800
rect 502006 940710 502744 940744
rect 502006 940654 502546 940710
rect 502602 940654 502744 940710
rect 502006 940500 502744 940654
rect 502006 940444 502207 940500
rect 502263 940444 502407 940500
rect 502463 940444 502744 940500
rect 502006 940410 502744 940444
rect 502006 940354 502546 940410
rect 502602 940354 502744 940410
rect 502006 940200 502744 940354
rect 502006 940144 502207 940200
rect 502263 940144 502407 940200
rect 502463 940144 502744 940200
rect 502006 940110 502744 940144
rect 502006 940054 502546 940110
rect 502602 940054 502744 940110
rect 502006 939922 502744 940054
rect 509424 943435 509744 943504
rect 509424 943379 509548 943435
rect 509604 943379 509744 943435
rect 509424 940710 509744 943379
rect 509424 940654 509546 940710
rect 509602 940654 509744 940710
rect 509424 940410 509744 940654
rect 509424 940354 509546 940410
rect 509602 940354 509744 940410
rect 509424 940110 509744 940354
rect 509424 940054 509546 940110
rect 509602 940054 509744 940110
rect 509424 939922 509744 940054
rect 520006 942200 520626 942322
rect 520006 942144 520207 942200
rect 520263 942144 520407 942200
rect 520463 942144 520626 942200
rect 520006 941900 520626 942144
rect 520006 941844 520207 941900
rect 520263 941844 520407 941900
rect 520463 941844 520626 941900
rect 520006 941600 520626 941844
rect 520006 941544 520207 941600
rect 520263 941544 520407 941600
rect 520463 941544 520626 941600
rect 502006 934568 502626 939922
rect 520006 933608 520626 941544
rect 525339 942153 525539 943085
rect 525339 942097 525406 942153
rect 525462 942097 525539 942153
rect 525339 941853 525539 942097
rect 525339 941797 525406 941853
rect 525462 941797 525539 941853
rect 525339 941553 525539 941797
rect 525339 941497 525406 941553
rect 525462 941497 525539 941553
rect 525339 941322 525539 941497
rect 525739 940716 525939 943565
rect 550424 943435 550744 943504
rect 550424 943379 550548 943435
rect 550604 943379 550744 943435
rect 525739 940660 525821 940716
rect 525877 940660 525939 940716
rect 525739 940416 525939 940660
rect 525739 940360 525821 940416
rect 525877 940360 525939 940416
rect 525739 940116 525939 940360
rect 525739 940060 525821 940116
rect 525877 940060 525939 940116
rect 525739 939922 525939 940060
rect 538006 940800 538626 940922
rect 538006 940744 538207 940800
rect 538263 940744 538407 940800
rect 538463 940744 538626 940800
rect 538006 940500 538626 940744
rect 538006 940444 538207 940500
rect 538263 940444 538407 940500
rect 538463 940444 538626 940500
rect 538006 940200 538626 940444
rect 538006 940144 538207 940200
rect 538263 940144 538407 940200
rect 538463 940144 538626 940200
rect 538006 934568 538626 940144
rect 550424 940710 550744 943379
rect 557424 943435 557744 943504
rect 557424 943379 557548 943435
rect 557604 943379 557744 943435
rect 550424 940654 550546 940710
rect 550602 940654 550744 940710
rect 550424 940410 550744 940654
rect 550424 940354 550546 940410
rect 550602 940354 550744 940410
rect 550424 940110 550744 940354
rect 550424 940054 550546 940110
rect 550602 940054 550744 940110
rect 550424 939922 550744 940054
rect 556006 942200 556626 942322
rect 556006 942144 556207 942200
rect 556263 942144 556407 942200
rect 556463 942144 556626 942200
rect 556006 941900 556626 942144
rect 556006 941844 556207 941900
rect 556263 941844 556407 941900
rect 556463 941844 556626 941900
rect 556006 941600 556626 941844
rect 556006 941544 556207 941600
rect 556263 941544 556407 941600
rect 556463 941544 556626 941600
rect 556006 933608 556626 941544
rect 557424 940710 557744 943379
rect 557424 940654 557546 940710
rect 557602 940654 557744 940710
rect 557424 940410 557744 940654
rect 557424 940354 557546 940410
rect 557602 940354 557744 940410
rect 557424 940110 557744 940354
rect 557424 940054 557546 940110
rect 557602 940054 557744 940110
rect 557424 939922 557744 940054
rect 564424 943435 564744 943504
rect 564424 943379 564548 943435
rect 564604 943379 564744 943435
rect 564424 940710 564744 943379
rect 580339 942153 580539 943085
rect 580339 942097 580406 942153
rect 580462 942097 580539 942153
rect 580339 941853 580539 942097
rect 580339 941797 580406 941853
rect 580462 941797 580539 941853
rect 580339 941553 580539 941797
rect 580339 941497 580406 941553
rect 580462 941497 580539 941553
rect 580339 941322 580539 941497
rect 564424 940654 564546 940710
rect 564602 940654 564744 940710
rect 564424 940410 564744 940654
rect 564424 940354 564546 940410
rect 564602 940354 564744 940410
rect 564424 940110 564744 940354
rect 564424 940054 564546 940110
rect 564602 940054 564744 940110
rect 564424 939922 564744 940054
rect 574006 940800 574626 940922
rect 574006 940744 574207 940800
rect 574263 940744 574407 940800
rect 574463 940744 574626 940800
rect 574006 940500 574626 940744
rect 574006 940444 574207 940500
rect 574263 940444 574407 940500
rect 574463 940444 574626 940500
rect 574006 940200 574626 940444
rect 574006 940144 574207 940200
rect 574263 940144 574407 940200
rect 574463 940144 574626 940200
rect 574006 934568 574626 940144
rect 580739 940716 580939 943565
rect 580739 940660 580821 940716
rect 580877 940660 580939 940716
rect 580739 940416 580939 940660
rect 580739 940360 580821 940416
rect 580877 940360 580939 940416
rect 580739 940116 580939 940360
rect 580739 940060 580821 940116
rect 580877 940060 580939 940116
rect 580739 939922 580939 940060
rect 592006 942200 592626 942322
rect 592006 942144 592207 942200
rect 592263 942144 592407 942200
rect 592463 942144 592626 942200
rect 592006 941900 592626 942144
rect 592006 941844 592207 941900
rect 592263 941844 592407 941900
rect 592463 941844 592626 941900
rect 592006 941600 592626 941844
rect 592006 941544 592207 941600
rect 592263 941544 592407 941600
rect 592463 941544 592626 941600
rect 592006 933608 592626 941544
rect 601272 940792 603172 949870
rect 601272 940736 601348 940792
rect 601404 940736 601472 940792
rect 601528 940736 601596 940792
rect 601652 940736 601720 940792
rect 601776 940736 601844 940792
rect 601900 940736 601968 940792
rect 602024 940736 602092 940792
rect 602148 940736 602216 940792
rect 602272 940736 602340 940792
rect 602396 940736 602464 940792
rect 602520 940736 602588 940792
rect 602644 940736 602712 940792
rect 602768 940736 602836 940792
rect 602892 940736 602960 940792
rect 603016 940736 603084 940792
rect 603140 940736 603172 940792
rect 601272 940668 603172 940736
rect 601272 940612 601348 940668
rect 601404 940612 601472 940668
rect 601528 940612 601596 940668
rect 601652 940612 601720 940668
rect 601776 940612 601844 940668
rect 601900 940612 601968 940668
rect 602024 940612 602092 940668
rect 602148 940612 602216 940668
rect 602272 940612 602340 940668
rect 602396 940612 602464 940668
rect 602520 940612 602588 940668
rect 602644 940612 602712 940668
rect 602768 940612 602836 940668
rect 602892 940612 602960 940668
rect 603016 940612 603084 940668
rect 603140 940612 603172 940668
rect 601272 940544 603172 940612
rect 601272 940488 601348 940544
rect 601404 940488 601472 940544
rect 601528 940488 601596 940544
rect 601652 940488 601720 940544
rect 601776 940488 601844 940544
rect 601900 940488 601968 940544
rect 602024 940488 602092 940544
rect 602148 940488 602216 940544
rect 602272 940488 602340 940544
rect 602396 940488 602464 940544
rect 602520 940488 602588 940544
rect 602644 940488 602712 940544
rect 602768 940488 602836 940544
rect 602892 940488 602960 940544
rect 603016 940488 603084 940544
rect 603140 940488 603172 940544
rect 601272 940420 603172 940488
rect 601272 940364 601348 940420
rect 601404 940364 601472 940420
rect 601528 940364 601596 940420
rect 601652 940364 601720 940420
rect 601776 940364 601844 940420
rect 601900 940364 601968 940420
rect 602024 940364 602092 940420
rect 602148 940364 602216 940420
rect 602272 940364 602340 940420
rect 602396 940364 602464 940420
rect 602520 940364 602588 940420
rect 602644 940364 602712 940420
rect 602768 940364 602836 940420
rect 602892 940364 602960 940420
rect 603016 940364 603084 940420
rect 603140 940364 603172 940420
rect 601272 940296 603172 940364
rect 601272 940240 601348 940296
rect 601404 940240 601472 940296
rect 601528 940240 601596 940296
rect 601652 940240 601720 940296
rect 601776 940240 601844 940296
rect 601900 940240 601968 940296
rect 602024 940240 602092 940296
rect 602148 940240 602216 940296
rect 602272 940240 602340 940296
rect 602396 940240 602464 940296
rect 602520 940240 602588 940296
rect 602644 940240 602712 940296
rect 602768 940240 602836 940296
rect 602892 940240 602960 940296
rect 603016 940240 603084 940296
rect 603140 940240 603172 940296
rect 601272 940172 603172 940240
rect 601272 940116 601348 940172
rect 601404 940116 601472 940172
rect 601528 940116 601596 940172
rect 601652 940116 601720 940172
rect 601776 940116 601844 940172
rect 601900 940116 601968 940172
rect 602024 940116 602092 940172
rect 602148 940116 602216 940172
rect 602272 940116 602340 940172
rect 602396 940116 602464 940172
rect 602520 940116 602588 940172
rect 602644 940116 602712 940172
rect 602768 940116 602836 940172
rect 602892 940116 602960 940172
rect 603016 940116 603084 940172
rect 603140 940116 603172 940172
rect 601272 940048 603172 940116
rect 601272 939992 601348 940048
rect 601404 939992 601472 940048
rect 601528 939992 601596 940048
rect 601652 939992 601720 940048
rect 601776 939992 601844 940048
rect 601900 939992 601968 940048
rect 602024 939992 602092 940048
rect 602148 939992 602216 940048
rect 602272 939992 602340 940048
rect 602396 939992 602464 940048
rect 602520 939992 602588 940048
rect 602644 939992 602712 940048
rect 602768 939992 602836 940048
rect 602892 939992 602960 940048
rect 603016 939992 603084 940048
rect 603140 939992 603172 940048
rect 601272 939922 603172 939992
rect 603752 949926 605802 950000
rect 603752 949870 603822 949926
rect 603878 949870 603946 949926
rect 604002 949870 604070 949926
rect 604126 949870 604194 949926
rect 604250 949870 604318 949926
rect 604374 949870 604442 949926
rect 604498 949870 604566 949926
rect 604622 949870 604690 949926
rect 604746 949870 604814 949926
rect 604870 949870 604938 949926
rect 604994 949870 605062 949926
rect 605118 949870 605186 949926
rect 605242 949870 605310 949926
rect 605366 949870 605434 949926
rect 605490 949870 605558 949926
rect 605614 949870 605682 949926
rect 605738 949870 605802 949926
rect 603752 940792 605802 949870
rect 603752 940736 603828 940792
rect 603884 940736 603952 940792
rect 604008 940736 604076 940792
rect 604132 940736 604200 940792
rect 604256 940736 604324 940792
rect 604380 940736 604448 940792
rect 604504 940736 604572 940792
rect 604628 940736 604696 940792
rect 604752 940736 604820 940792
rect 604876 940736 604944 940792
rect 605000 940736 605068 940792
rect 605124 940736 605192 940792
rect 605248 940736 605316 940792
rect 605372 940736 605440 940792
rect 605496 940736 605564 940792
rect 605620 940736 605688 940792
rect 605744 940736 605802 940792
rect 603752 940668 605802 940736
rect 603752 940612 603828 940668
rect 603884 940612 603952 940668
rect 604008 940612 604076 940668
rect 604132 940612 604200 940668
rect 604256 940612 604324 940668
rect 604380 940612 604448 940668
rect 604504 940612 604572 940668
rect 604628 940612 604696 940668
rect 604752 940612 604820 940668
rect 604876 940612 604944 940668
rect 605000 940612 605068 940668
rect 605124 940612 605192 940668
rect 605248 940612 605316 940668
rect 605372 940612 605440 940668
rect 605496 940612 605564 940668
rect 605620 940612 605688 940668
rect 605744 940612 605802 940668
rect 603752 940544 605802 940612
rect 603752 940488 603828 940544
rect 603884 940488 603952 940544
rect 604008 940488 604076 940544
rect 604132 940488 604200 940544
rect 604256 940488 604324 940544
rect 604380 940488 604448 940544
rect 604504 940488 604572 940544
rect 604628 940488 604696 940544
rect 604752 940488 604820 940544
rect 604876 940488 604944 940544
rect 605000 940488 605068 940544
rect 605124 940488 605192 940544
rect 605248 940488 605316 940544
rect 605372 940488 605440 940544
rect 605496 940488 605564 940544
rect 605620 940488 605688 940544
rect 605744 940488 605802 940544
rect 603752 940420 605802 940488
rect 603752 940364 603828 940420
rect 603884 940364 603952 940420
rect 604008 940364 604076 940420
rect 604132 940364 604200 940420
rect 604256 940364 604324 940420
rect 604380 940364 604448 940420
rect 604504 940364 604572 940420
rect 604628 940364 604696 940420
rect 604752 940364 604820 940420
rect 604876 940364 604944 940420
rect 605000 940364 605068 940420
rect 605124 940364 605192 940420
rect 605248 940364 605316 940420
rect 605372 940364 605440 940420
rect 605496 940364 605564 940420
rect 605620 940364 605688 940420
rect 605744 940364 605802 940420
rect 603752 940296 605802 940364
rect 603752 940240 603828 940296
rect 603884 940240 603952 940296
rect 604008 940240 604076 940296
rect 604132 940240 604200 940296
rect 604256 940240 604324 940296
rect 604380 940240 604448 940296
rect 604504 940240 604572 940296
rect 604628 940240 604696 940296
rect 604752 940240 604820 940296
rect 604876 940240 604944 940296
rect 605000 940240 605068 940296
rect 605124 940240 605192 940296
rect 605248 940240 605316 940296
rect 605372 940240 605440 940296
rect 605496 940240 605564 940296
rect 605620 940240 605688 940296
rect 605744 940240 605802 940296
rect 603752 940172 605802 940240
rect 603752 940116 603828 940172
rect 603884 940116 603952 940172
rect 604008 940116 604076 940172
rect 604132 940116 604200 940172
rect 604256 940116 604324 940172
rect 604380 940116 604448 940172
rect 604504 940116 604572 940172
rect 604628 940116 604696 940172
rect 604752 940116 604820 940172
rect 604876 940116 604944 940172
rect 605000 940116 605068 940172
rect 605124 940116 605192 940172
rect 605248 940116 605316 940172
rect 605372 940116 605440 940172
rect 605496 940116 605564 940172
rect 605620 940116 605688 940172
rect 605744 940116 605802 940172
rect 603752 940048 605802 940116
rect 603752 939992 603828 940048
rect 603884 939992 603952 940048
rect 604008 939992 604076 940048
rect 604132 939992 604200 940048
rect 604256 939992 604324 940048
rect 604380 939992 604448 940048
rect 604504 939992 604572 940048
rect 604628 939992 604696 940048
rect 604752 939992 604820 940048
rect 604876 939992 604944 940048
rect 605000 939992 605068 940048
rect 605124 939992 605192 940048
rect 605248 939992 605316 940048
rect 605372 939992 605440 940048
rect 605496 939992 605564 940048
rect 605620 939992 605688 940048
rect 605744 939992 605802 940048
rect 603752 939922 605802 939992
rect 606122 949926 608172 950000
rect 606122 949870 606192 949926
rect 606248 949870 606316 949926
rect 606372 949870 606440 949926
rect 606496 949870 606564 949926
rect 606620 949870 606688 949926
rect 606744 949870 606812 949926
rect 606868 949870 606936 949926
rect 606992 949870 607060 949926
rect 607116 949870 607184 949926
rect 607240 949870 607308 949926
rect 607364 949870 607432 949926
rect 607488 949870 607556 949926
rect 607612 949870 607680 949926
rect 607736 949870 607804 949926
rect 607860 949870 607928 949926
rect 607984 949870 608052 949926
rect 608108 949870 608172 949926
rect 606122 940792 608172 949870
rect 606122 940736 606198 940792
rect 606254 940736 606322 940792
rect 606378 940736 606446 940792
rect 606502 940736 606570 940792
rect 606626 940736 606694 940792
rect 606750 940736 606818 940792
rect 606874 940736 606942 940792
rect 606998 940736 607066 940792
rect 607122 940736 607190 940792
rect 607246 940736 607314 940792
rect 607370 940736 607438 940792
rect 607494 940736 607562 940792
rect 607618 940736 607686 940792
rect 607742 940736 607810 940792
rect 607866 940736 607934 940792
rect 607990 940736 608058 940792
rect 608114 940736 608172 940792
rect 606122 940668 608172 940736
rect 606122 940612 606198 940668
rect 606254 940612 606322 940668
rect 606378 940612 606446 940668
rect 606502 940612 606570 940668
rect 606626 940612 606694 940668
rect 606750 940612 606818 940668
rect 606874 940612 606942 940668
rect 606998 940612 607066 940668
rect 607122 940612 607190 940668
rect 607246 940612 607314 940668
rect 607370 940612 607438 940668
rect 607494 940612 607562 940668
rect 607618 940612 607686 940668
rect 607742 940612 607810 940668
rect 607866 940612 607934 940668
rect 607990 940612 608058 940668
rect 608114 940612 608172 940668
rect 606122 940544 608172 940612
rect 606122 940488 606198 940544
rect 606254 940488 606322 940544
rect 606378 940488 606446 940544
rect 606502 940488 606570 940544
rect 606626 940488 606694 940544
rect 606750 940488 606818 940544
rect 606874 940488 606942 940544
rect 606998 940488 607066 940544
rect 607122 940488 607190 940544
rect 607246 940488 607314 940544
rect 607370 940488 607438 940544
rect 607494 940488 607562 940544
rect 607618 940488 607686 940544
rect 607742 940488 607810 940544
rect 607866 940488 607934 940544
rect 607990 940488 608058 940544
rect 608114 940488 608172 940544
rect 606122 940420 608172 940488
rect 606122 940364 606198 940420
rect 606254 940364 606322 940420
rect 606378 940364 606446 940420
rect 606502 940364 606570 940420
rect 606626 940364 606694 940420
rect 606750 940364 606818 940420
rect 606874 940364 606942 940420
rect 606998 940364 607066 940420
rect 607122 940364 607190 940420
rect 607246 940364 607314 940420
rect 607370 940364 607438 940420
rect 607494 940364 607562 940420
rect 607618 940364 607686 940420
rect 607742 940364 607810 940420
rect 607866 940364 607934 940420
rect 607990 940364 608058 940420
rect 608114 940364 608172 940420
rect 606122 940296 608172 940364
rect 606122 940240 606198 940296
rect 606254 940240 606322 940296
rect 606378 940240 606446 940296
rect 606502 940240 606570 940296
rect 606626 940240 606694 940296
rect 606750 940240 606818 940296
rect 606874 940240 606942 940296
rect 606998 940240 607066 940296
rect 607122 940240 607190 940296
rect 607246 940240 607314 940296
rect 607370 940240 607438 940296
rect 607494 940240 607562 940296
rect 607618 940240 607686 940296
rect 607742 940240 607810 940296
rect 607866 940240 607934 940296
rect 607990 940240 608058 940296
rect 608114 940240 608172 940296
rect 606122 940172 608172 940240
rect 606122 940116 606198 940172
rect 606254 940116 606322 940172
rect 606378 940116 606446 940172
rect 606502 940116 606570 940172
rect 606626 940116 606694 940172
rect 606750 940116 606818 940172
rect 606874 940116 606942 940172
rect 606998 940116 607066 940172
rect 607122 940116 607190 940172
rect 607246 940116 607314 940172
rect 607370 940116 607438 940172
rect 607494 940116 607562 940172
rect 607618 940116 607686 940172
rect 607742 940116 607810 940172
rect 607866 940116 607934 940172
rect 607990 940116 608058 940172
rect 608114 940116 608172 940172
rect 606122 940048 608172 940116
rect 606122 939992 606198 940048
rect 606254 939992 606322 940048
rect 606378 939992 606446 940048
rect 606502 939992 606570 940048
rect 606626 939992 606694 940048
rect 606750 939992 606818 940048
rect 606874 939992 606942 940048
rect 606998 939992 607066 940048
rect 607122 939992 607190 940048
rect 607246 939992 607314 940048
rect 607370 939992 607438 940048
rect 607494 939992 607562 940048
rect 607618 939992 607686 940048
rect 607742 939992 607810 940048
rect 607866 939992 607934 940048
rect 607990 939992 608058 940048
rect 608114 939992 608172 940048
rect 606122 939922 608172 939992
rect 608828 949926 610878 950000
rect 608828 949870 608892 949926
rect 608948 949870 609016 949926
rect 609072 949870 609140 949926
rect 609196 949870 609264 949926
rect 609320 949870 609388 949926
rect 609444 949870 609512 949926
rect 609568 949870 609636 949926
rect 609692 949870 609760 949926
rect 609816 949870 609884 949926
rect 609940 949870 610008 949926
rect 610064 949870 610132 949926
rect 610188 949870 610256 949926
rect 610312 949870 610380 949926
rect 610436 949870 610504 949926
rect 610560 949870 610628 949926
rect 610684 949870 610752 949926
rect 610808 949870 610878 949926
rect 608828 940792 610878 949870
rect 608828 940736 608904 940792
rect 608960 940736 609028 940792
rect 609084 940736 609152 940792
rect 609208 940736 609276 940792
rect 609332 940736 609400 940792
rect 609456 940736 609524 940792
rect 609580 940736 609648 940792
rect 609704 940736 609772 940792
rect 609828 940736 609896 940792
rect 609952 940736 610020 940792
rect 610076 940736 610144 940792
rect 610200 940736 610268 940792
rect 610324 940736 610392 940792
rect 610448 940736 610516 940792
rect 610572 940736 610640 940792
rect 610696 940736 610764 940792
rect 610820 940736 610878 940792
rect 608828 940668 610878 940736
rect 608828 940612 608904 940668
rect 608960 940612 609028 940668
rect 609084 940612 609152 940668
rect 609208 940612 609276 940668
rect 609332 940612 609400 940668
rect 609456 940612 609524 940668
rect 609580 940612 609648 940668
rect 609704 940612 609772 940668
rect 609828 940612 609896 940668
rect 609952 940612 610020 940668
rect 610076 940612 610144 940668
rect 610200 940612 610268 940668
rect 610324 940612 610392 940668
rect 610448 940612 610516 940668
rect 610572 940612 610640 940668
rect 610696 940612 610764 940668
rect 610820 940612 610878 940668
rect 608828 940544 610878 940612
rect 608828 940488 608904 940544
rect 608960 940488 609028 940544
rect 609084 940488 609152 940544
rect 609208 940488 609276 940544
rect 609332 940488 609400 940544
rect 609456 940488 609524 940544
rect 609580 940488 609648 940544
rect 609704 940488 609772 940544
rect 609828 940488 609896 940544
rect 609952 940488 610020 940544
rect 610076 940488 610144 940544
rect 610200 940488 610268 940544
rect 610324 940488 610392 940544
rect 610448 940488 610516 940544
rect 610572 940488 610640 940544
rect 610696 940488 610764 940544
rect 610820 940488 610878 940544
rect 608828 940420 610878 940488
rect 608828 940364 608904 940420
rect 608960 940364 609028 940420
rect 609084 940364 609152 940420
rect 609208 940364 609276 940420
rect 609332 940364 609400 940420
rect 609456 940364 609524 940420
rect 609580 940364 609648 940420
rect 609704 940364 609772 940420
rect 609828 940364 609896 940420
rect 609952 940364 610020 940420
rect 610076 940364 610144 940420
rect 610200 940364 610268 940420
rect 610324 940364 610392 940420
rect 610448 940364 610516 940420
rect 610572 940364 610640 940420
rect 610696 940364 610764 940420
rect 610820 940364 610878 940420
rect 608828 940296 610878 940364
rect 608828 940240 608904 940296
rect 608960 940240 609028 940296
rect 609084 940240 609152 940296
rect 609208 940240 609276 940296
rect 609332 940240 609400 940296
rect 609456 940240 609524 940296
rect 609580 940240 609648 940296
rect 609704 940240 609772 940296
rect 609828 940240 609896 940296
rect 609952 940240 610020 940296
rect 610076 940240 610144 940296
rect 610200 940240 610268 940296
rect 610324 940240 610392 940296
rect 610448 940240 610516 940296
rect 610572 940240 610640 940296
rect 610696 940240 610764 940296
rect 610820 940240 610878 940296
rect 608828 940172 610878 940240
rect 608828 940116 608904 940172
rect 608960 940116 609028 940172
rect 609084 940116 609152 940172
rect 609208 940116 609276 940172
rect 609332 940116 609400 940172
rect 609456 940116 609524 940172
rect 609580 940116 609648 940172
rect 609704 940116 609772 940172
rect 609828 940116 609896 940172
rect 609952 940116 610020 940172
rect 610076 940116 610144 940172
rect 610200 940116 610268 940172
rect 610324 940116 610392 940172
rect 610448 940116 610516 940172
rect 610572 940116 610640 940172
rect 610696 940116 610764 940172
rect 610820 940116 610878 940172
rect 608828 940048 610878 940116
rect 608828 939992 608904 940048
rect 608960 939992 609028 940048
rect 609084 939992 609152 940048
rect 609208 939992 609276 940048
rect 609332 939992 609400 940048
rect 609456 939992 609524 940048
rect 609580 939992 609648 940048
rect 609704 939992 609772 940048
rect 609828 939992 609896 940048
rect 609952 939992 610020 940048
rect 610076 939992 610144 940048
rect 610200 939992 610268 940048
rect 610324 939992 610392 940048
rect 610448 939992 610516 940048
rect 610572 939992 610640 940048
rect 610696 939992 610764 940048
rect 610820 939992 610878 940048
rect 608828 939922 610878 939992
rect 611198 949926 613248 950000
rect 611198 949870 611262 949926
rect 611318 949870 611386 949926
rect 611442 949870 611510 949926
rect 611566 949870 611634 949926
rect 611690 949870 611758 949926
rect 611814 949870 611882 949926
rect 611938 949870 612006 949926
rect 612062 949870 612130 949926
rect 612186 949870 612254 949926
rect 612310 949870 612378 949926
rect 612434 949870 612502 949926
rect 612558 949870 612626 949926
rect 612682 949870 612750 949926
rect 612806 949870 612874 949926
rect 612930 949870 612998 949926
rect 613054 949870 613122 949926
rect 613178 949870 613248 949926
rect 611198 940792 613248 949870
rect 611198 940736 611274 940792
rect 611330 940736 611398 940792
rect 611454 940736 611522 940792
rect 611578 940736 611646 940792
rect 611702 940736 611770 940792
rect 611826 940736 611894 940792
rect 611950 940736 612018 940792
rect 612074 940736 612142 940792
rect 612198 940736 612266 940792
rect 612322 940736 612390 940792
rect 612446 940736 612514 940792
rect 612570 940736 612638 940792
rect 612694 940736 612762 940792
rect 612818 940736 612886 940792
rect 612942 940736 613010 940792
rect 613066 940736 613134 940792
rect 613190 940736 613248 940792
rect 611198 940668 613248 940736
rect 611198 940612 611274 940668
rect 611330 940612 611398 940668
rect 611454 940612 611522 940668
rect 611578 940612 611646 940668
rect 611702 940612 611770 940668
rect 611826 940612 611894 940668
rect 611950 940612 612018 940668
rect 612074 940612 612142 940668
rect 612198 940612 612266 940668
rect 612322 940612 612390 940668
rect 612446 940612 612514 940668
rect 612570 940612 612638 940668
rect 612694 940612 612762 940668
rect 612818 940612 612886 940668
rect 612942 940612 613010 940668
rect 613066 940612 613134 940668
rect 613190 940612 613248 940668
rect 611198 940544 613248 940612
rect 611198 940488 611274 940544
rect 611330 940488 611398 940544
rect 611454 940488 611522 940544
rect 611578 940488 611646 940544
rect 611702 940488 611770 940544
rect 611826 940488 611894 940544
rect 611950 940488 612018 940544
rect 612074 940488 612142 940544
rect 612198 940488 612266 940544
rect 612322 940488 612390 940544
rect 612446 940488 612514 940544
rect 612570 940488 612638 940544
rect 612694 940488 612762 940544
rect 612818 940488 612886 940544
rect 612942 940488 613010 940544
rect 613066 940488 613134 940544
rect 613190 940488 613248 940544
rect 611198 940420 613248 940488
rect 611198 940364 611274 940420
rect 611330 940364 611398 940420
rect 611454 940364 611522 940420
rect 611578 940364 611646 940420
rect 611702 940364 611770 940420
rect 611826 940364 611894 940420
rect 611950 940364 612018 940420
rect 612074 940364 612142 940420
rect 612198 940364 612266 940420
rect 612322 940364 612390 940420
rect 612446 940364 612514 940420
rect 612570 940364 612638 940420
rect 612694 940364 612762 940420
rect 612818 940364 612886 940420
rect 612942 940364 613010 940420
rect 613066 940364 613134 940420
rect 613190 940364 613248 940420
rect 611198 940296 613248 940364
rect 611198 940240 611274 940296
rect 611330 940240 611398 940296
rect 611454 940240 611522 940296
rect 611578 940240 611646 940296
rect 611702 940240 611770 940296
rect 611826 940240 611894 940296
rect 611950 940240 612018 940296
rect 612074 940240 612142 940296
rect 612198 940240 612266 940296
rect 612322 940240 612390 940296
rect 612446 940240 612514 940296
rect 612570 940240 612638 940296
rect 612694 940240 612762 940296
rect 612818 940240 612886 940296
rect 612942 940240 613010 940296
rect 613066 940240 613134 940296
rect 613190 940240 613248 940296
rect 611198 940172 613248 940240
rect 611198 940116 611274 940172
rect 611330 940116 611398 940172
rect 611454 940116 611522 940172
rect 611578 940116 611646 940172
rect 611702 940116 611770 940172
rect 611826 940116 611894 940172
rect 611950 940116 612018 940172
rect 612074 940116 612142 940172
rect 612198 940116 612266 940172
rect 612322 940116 612390 940172
rect 612446 940116 612514 940172
rect 612570 940116 612638 940172
rect 612694 940116 612762 940172
rect 612818 940116 612886 940172
rect 612942 940116 613010 940172
rect 613066 940116 613134 940172
rect 613190 940116 613248 940172
rect 611198 940048 613248 940116
rect 611198 939992 611274 940048
rect 611330 939992 611398 940048
rect 611454 939992 611522 940048
rect 611578 939992 611646 940048
rect 611702 939992 611770 940048
rect 611826 939992 611894 940048
rect 611950 939992 612018 940048
rect 612074 939992 612142 940048
rect 612198 939992 612266 940048
rect 612322 939992 612390 940048
rect 612446 939992 612514 940048
rect 612570 939992 612638 940048
rect 612694 939992 612762 940048
rect 612818 939992 612886 940048
rect 612942 939992 613010 940048
rect 613066 939992 613134 940048
rect 613190 939992 613248 940048
rect 611198 939922 613248 939992
rect 613828 949926 615728 950000
rect 613828 949870 613866 949926
rect 613922 949870 613990 949926
rect 614046 949870 614114 949926
rect 614170 949870 614238 949926
rect 614294 949870 614362 949926
rect 614418 949870 614486 949926
rect 614542 949870 614610 949926
rect 614666 949870 614734 949926
rect 614790 949870 614858 949926
rect 614914 949870 614982 949926
rect 615038 949870 615106 949926
rect 615162 949870 615230 949926
rect 615286 949870 615354 949926
rect 615410 949870 615478 949926
rect 615534 949870 615602 949926
rect 615658 949870 615728 949926
rect 613828 940792 615728 949870
rect 690339 943565 690939 943885
rect 660424 943435 660744 943504
rect 660424 943379 660548 943435
rect 660604 943379 660744 943435
rect 613828 940736 613878 940792
rect 613934 940736 614002 940792
rect 614058 940736 614126 940792
rect 614182 940736 614250 940792
rect 614306 940736 614374 940792
rect 614430 940736 614498 940792
rect 614554 940736 614622 940792
rect 614678 940736 614746 940792
rect 614802 940736 614870 940792
rect 614926 940736 614994 940792
rect 615050 940736 615118 940792
rect 615174 940736 615242 940792
rect 615298 940736 615366 940792
rect 615422 940736 615490 940792
rect 615546 940736 615614 940792
rect 615670 940736 615728 940792
rect 613828 940668 615728 940736
rect 613828 940612 613878 940668
rect 613934 940612 614002 940668
rect 614058 940612 614126 940668
rect 614182 940612 614250 940668
rect 614306 940612 614374 940668
rect 614430 940612 614498 940668
rect 614554 940612 614622 940668
rect 614678 940612 614746 940668
rect 614802 940612 614870 940668
rect 614926 940612 614994 940668
rect 615050 940612 615118 940668
rect 615174 940612 615242 940668
rect 615298 940612 615366 940668
rect 615422 940612 615490 940668
rect 615546 940612 615614 940668
rect 615670 940612 615728 940668
rect 613828 940544 615728 940612
rect 613828 940488 613878 940544
rect 613934 940488 614002 940544
rect 614058 940488 614126 940544
rect 614182 940488 614250 940544
rect 614306 940488 614374 940544
rect 614430 940488 614498 940544
rect 614554 940488 614622 940544
rect 614678 940488 614746 940544
rect 614802 940488 614870 940544
rect 614926 940488 614994 940544
rect 615050 940488 615118 940544
rect 615174 940488 615242 940544
rect 615298 940488 615366 940544
rect 615422 940488 615490 940544
rect 615546 940488 615614 940544
rect 615670 940488 615728 940544
rect 613828 940420 615728 940488
rect 613828 940364 613878 940420
rect 613934 940364 614002 940420
rect 614058 940364 614126 940420
rect 614182 940364 614250 940420
rect 614306 940364 614374 940420
rect 614430 940364 614498 940420
rect 614554 940364 614622 940420
rect 614678 940364 614746 940420
rect 614802 940364 614870 940420
rect 614926 940364 614994 940420
rect 615050 940364 615118 940420
rect 615174 940364 615242 940420
rect 615298 940364 615366 940420
rect 615422 940364 615490 940420
rect 615546 940364 615614 940420
rect 615670 940364 615728 940420
rect 613828 940296 615728 940364
rect 613828 940240 613878 940296
rect 613934 940240 614002 940296
rect 614058 940240 614126 940296
rect 614182 940240 614250 940296
rect 614306 940240 614374 940296
rect 614430 940240 614498 940296
rect 614554 940240 614622 940296
rect 614678 940240 614746 940296
rect 614802 940240 614870 940296
rect 614926 940240 614994 940296
rect 615050 940240 615118 940296
rect 615174 940240 615242 940296
rect 615298 940240 615366 940296
rect 615422 940240 615490 940296
rect 615546 940240 615614 940296
rect 615670 940240 615728 940296
rect 613828 940172 615728 940240
rect 613828 940116 613878 940172
rect 613934 940116 614002 940172
rect 614058 940116 614126 940172
rect 614182 940116 614250 940172
rect 614306 940116 614374 940172
rect 614430 940116 614498 940172
rect 614554 940116 614622 940172
rect 614678 940116 614746 940172
rect 614802 940116 614870 940172
rect 614926 940116 614994 940172
rect 615050 940116 615118 940172
rect 615174 940116 615242 940172
rect 615298 940116 615366 940172
rect 615422 940116 615490 940172
rect 615546 940116 615614 940172
rect 615670 940116 615728 940172
rect 613828 940048 615728 940116
rect 613828 939992 613878 940048
rect 613934 939992 614002 940048
rect 614058 939992 614126 940048
rect 614182 939992 614250 940048
rect 614306 939992 614374 940048
rect 614430 939992 614498 940048
rect 614554 939992 614622 940048
rect 614678 939992 614746 940048
rect 614802 939992 614870 940048
rect 614926 939992 614994 940048
rect 615050 939992 615118 940048
rect 615174 939992 615242 940048
rect 615298 939992 615366 940048
rect 615422 939992 615490 940048
rect 615546 939992 615614 940048
rect 615670 939992 615728 940048
rect 613828 939922 615728 939992
rect 628006 942200 628626 942322
rect 628006 942144 628207 942200
rect 628263 942144 628407 942200
rect 628463 942144 628626 942200
rect 628006 941900 628626 942144
rect 628006 941844 628207 941900
rect 628263 941844 628407 941900
rect 628463 941844 628626 941900
rect 628006 941600 628626 941844
rect 628006 941544 628207 941600
rect 628263 941544 628407 941600
rect 628463 941544 628626 941600
rect 610006 934568 610626 939922
rect 628006 933608 628626 941544
rect 646006 940800 646626 940922
rect 646006 940744 646207 940800
rect 646263 940744 646407 940800
rect 646463 940744 646626 940800
rect 646006 940500 646626 940744
rect 646006 940444 646207 940500
rect 646263 940444 646407 940500
rect 646463 940444 646626 940500
rect 646006 940200 646626 940444
rect 646006 940144 646207 940200
rect 646263 940144 646407 940200
rect 646463 940144 646626 940200
rect 646006 934568 646626 940144
rect 660424 940710 660744 943379
rect 667424 943435 667744 943504
rect 667424 943379 667548 943435
rect 667604 943379 667744 943435
rect 660424 940654 660546 940710
rect 660602 940654 660744 940710
rect 660424 940410 660744 940654
rect 660424 940354 660546 940410
rect 660602 940354 660744 940410
rect 660424 940110 660744 940354
rect 660424 940054 660546 940110
rect 660602 940054 660744 940110
rect 660424 939922 660744 940054
rect 664006 942200 664626 942322
rect 664006 942144 664207 942200
rect 664263 942144 664407 942200
rect 664463 942144 664626 942200
rect 664006 941900 664626 942144
rect 664006 941844 664207 941900
rect 664263 941844 664407 941900
rect 664463 941844 664626 941900
rect 664006 941600 664626 941844
rect 664006 941544 664207 941600
rect 664263 941544 664407 941600
rect 664463 941544 664626 941600
rect 664006 933608 664626 941544
rect 667424 940710 667744 943379
rect 667424 940654 667546 940710
rect 667602 940654 667744 940710
rect 667424 940410 667744 940654
rect 667424 940354 667546 940410
rect 667602 940354 667744 940410
rect 667424 940110 667744 940354
rect 667424 940054 667546 940110
rect 667602 940054 667744 940110
rect 667424 939922 667744 940054
rect 674424 943435 674744 943504
rect 674424 943379 674548 943435
rect 674604 943379 674744 943435
rect 674424 940710 674744 943379
rect 690339 942153 690539 943085
rect 690339 942097 690406 942153
rect 690462 942097 690539 942153
rect 690339 941853 690539 942097
rect 690339 941797 690406 941853
rect 690462 941797 690539 941853
rect 690339 941553 690539 941797
rect 690339 941497 690406 941553
rect 690462 941497 690539 941553
rect 690339 941322 690539 941497
rect 674424 940654 674546 940710
rect 674602 940654 674744 940710
rect 674424 940410 674744 940654
rect 674424 940354 674546 940410
rect 674602 940354 674744 940410
rect 674424 940110 674744 940354
rect 674424 940054 674546 940110
rect 674602 940054 674744 940110
rect 674424 939922 674744 940054
rect 682006 940800 682626 940922
rect 682006 940744 682207 940800
rect 682263 940744 682407 940800
rect 682463 940744 682626 940800
rect 682006 940500 682626 940744
rect 682006 940444 682207 940500
rect 682263 940444 682407 940500
rect 682463 940444 682626 940500
rect 682006 940200 682626 940444
rect 682006 940144 682207 940200
rect 682263 940144 682407 940200
rect 682463 940144 682626 940200
rect 682006 934568 682626 940144
rect 690739 940716 690939 943565
rect 699322 942192 700322 942322
rect 699322 942136 699452 942192
rect 699508 942136 699576 942192
rect 699632 942136 699700 942192
rect 699756 942136 699824 942192
rect 699880 942136 699948 942192
rect 700004 942136 700072 942192
rect 700128 942136 700196 942192
rect 700252 942136 700322 942192
rect 699322 942068 700322 942136
rect 699322 942012 699452 942068
rect 699508 942012 699576 942068
rect 699632 942012 699700 942068
rect 699756 942012 699824 942068
rect 699880 942012 699948 942068
rect 700004 942012 700072 942068
rect 700128 942012 700196 942068
rect 700252 942012 700322 942068
rect 699322 941944 700322 942012
rect 699322 941888 699452 941944
rect 699508 941888 699576 941944
rect 699632 941888 699700 941944
rect 699756 941888 699824 941944
rect 699880 941888 699948 941944
rect 700004 941888 700072 941944
rect 700128 941888 700196 941944
rect 700252 941888 700322 941944
rect 699322 941820 700322 941888
rect 699322 941764 699452 941820
rect 699508 941764 699576 941820
rect 699632 941764 699700 941820
rect 699756 941764 699824 941820
rect 699880 941764 699948 941820
rect 700004 941764 700072 941820
rect 700128 941764 700196 941820
rect 700252 941764 700322 941820
rect 699322 941696 700322 941764
rect 699322 941640 699452 941696
rect 699508 941640 699576 941696
rect 699632 941640 699700 941696
rect 699756 941640 699824 941696
rect 699880 941640 699948 941696
rect 700004 941640 700072 941696
rect 700128 941640 700196 941696
rect 700252 941640 700322 941696
rect 699322 941572 700322 941640
rect 699322 941516 699452 941572
rect 699508 941516 699576 941572
rect 699632 941516 699700 941572
rect 699756 941516 699824 941572
rect 699880 941516 699948 941572
rect 700004 941516 700072 941572
rect 700128 941516 700196 941572
rect 700252 941516 700322 941572
rect 699322 941448 700322 941516
rect 699322 941392 699452 941448
rect 699508 941392 699576 941448
rect 699632 941392 699700 941448
rect 699756 941392 699824 941448
rect 699880 941392 699948 941448
rect 700004 941392 700072 941448
rect 700128 941392 700196 941448
rect 700252 941392 700322 941448
rect 690739 940660 690821 940716
rect 690877 940660 690939 940716
rect 690739 940416 690939 940660
rect 690739 940360 690821 940416
rect 690877 940360 690939 940416
rect 690739 940116 690939 940360
rect 690739 940060 690821 940116
rect 690877 940060 690939 940116
rect 690739 939922 690939 940060
rect 697922 940792 698922 940922
rect 697922 940736 698052 940792
rect 698108 940736 698176 940792
rect 698232 940736 698300 940792
rect 698356 940736 698424 940792
rect 698480 940736 698548 940792
rect 698604 940736 698672 940792
rect 698728 940736 698796 940792
rect 698852 940736 698922 940792
rect 697922 940668 698922 940736
rect 697922 940612 698052 940668
rect 698108 940612 698176 940668
rect 698232 940612 698300 940668
rect 698356 940612 698424 940668
rect 698480 940612 698548 940668
rect 698604 940612 698672 940668
rect 698728 940612 698796 940668
rect 698852 940612 698922 940668
rect 697922 940544 698922 940612
rect 697922 940488 698052 940544
rect 698108 940488 698176 940544
rect 698232 940488 698300 940544
rect 698356 940488 698424 940544
rect 698480 940488 698548 940544
rect 698604 940488 698672 940544
rect 698728 940488 698796 940544
rect 698852 940488 698922 940544
rect 697922 940420 698922 940488
rect 697922 940364 698052 940420
rect 698108 940364 698176 940420
rect 698232 940364 698300 940420
rect 698356 940364 698424 940420
rect 698480 940364 698548 940420
rect 698604 940364 698672 940420
rect 698728 940364 698796 940420
rect 698852 940364 698922 940420
rect 697922 940296 698922 940364
rect 697922 940240 698052 940296
rect 698108 940240 698176 940296
rect 698232 940240 698300 940296
rect 698356 940240 698424 940296
rect 698480 940240 698548 940296
rect 698604 940240 698672 940296
rect 698728 940240 698796 940296
rect 698852 940240 698922 940296
rect 697922 940172 698922 940240
rect 697922 940116 698052 940172
rect 698108 940116 698176 940172
rect 698232 940116 698300 940172
rect 698356 940116 698424 940172
rect 698480 940116 698548 940172
rect 698604 940116 698672 940172
rect 698728 940116 698796 940172
rect 698852 940116 698922 940172
rect 697922 940048 698922 940116
rect 697922 939992 698052 940048
rect 698108 939992 698176 940048
rect 698232 939992 698300 940048
rect 698356 939992 698424 940048
rect 698480 939992 698548 940048
rect 698604 939992 698672 940048
rect 698728 939992 698796 940048
rect 698852 939992 698922 940048
rect 79078 929566 79300 929622
rect 79356 929566 79600 929622
rect 79656 929566 79900 929622
rect 79956 929566 80078 929622
rect 79078 922622 80078 929566
rect 79078 922566 79300 922622
rect 79356 922566 79600 922622
rect 79656 922566 79900 922622
rect 79956 922566 80078 922622
rect 79078 915622 80078 922566
rect 79078 915566 79300 915622
rect 79356 915566 79600 915622
rect 79656 915566 79900 915622
rect 79956 915566 80078 915622
rect 79078 896429 80078 915566
rect 79078 896373 79200 896429
rect 79256 896373 79500 896429
rect 79556 896373 79800 896429
rect 79856 896373 80078 896429
rect 79078 896229 80078 896373
rect 79078 896173 79200 896229
rect 79256 896173 79500 896229
rect 79556 896173 79800 896229
rect 79856 896173 80078 896229
rect 79078 860429 80078 896173
rect 79078 860373 79200 860429
rect 79256 860373 79500 860429
rect 79556 860373 79800 860429
rect 79856 860373 80078 860429
rect 79078 860229 80078 860373
rect 79078 860173 79200 860229
rect 79256 860173 79500 860229
rect 79556 860173 79800 860229
rect 79856 860173 80078 860229
rect 79078 824429 80078 860173
rect 79078 824373 79200 824429
rect 79256 824373 79500 824429
rect 79556 824373 79800 824429
rect 79856 824373 80078 824429
rect 79078 824229 80078 824373
rect 79078 824173 79200 824229
rect 79256 824173 79500 824229
rect 79556 824173 79800 824229
rect 79856 824173 80078 824229
rect 79078 802670 80078 824173
rect 79078 802614 79208 802670
rect 79264 802614 79332 802670
rect 79388 802614 79456 802670
rect 79512 802614 79580 802670
rect 79636 802614 79704 802670
rect 79760 802614 79828 802670
rect 79884 802614 79952 802670
rect 80008 802614 80078 802670
rect 79078 802546 80078 802614
rect 79078 802490 79208 802546
rect 79264 802490 79332 802546
rect 79388 802490 79456 802546
rect 79512 802490 79580 802546
rect 79636 802490 79704 802546
rect 79760 802490 79828 802546
rect 79884 802490 79952 802546
rect 80008 802490 80078 802546
rect 79078 802422 80078 802490
rect 79078 802366 79208 802422
rect 79264 802366 79332 802422
rect 79388 802366 79456 802422
rect 79512 802366 79580 802422
rect 79636 802366 79704 802422
rect 79760 802366 79828 802422
rect 79884 802366 79952 802422
rect 80008 802366 80078 802422
rect 79078 802298 80078 802366
rect 79078 802242 79208 802298
rect 79264 802242 79332 802298
rect 79388 802242 79456 802298
rect 79512 802242 79580 802298
rect 79636 802242 79704 802298
rect 79760 802242 79828 802298
rect 79884 802242 79952 802298
rect 80008 802242 80078 802298
rect 79078 802174 80078 802242
rect 79078 802118 79208 802174
rect 79264 802118 79332 802174
rect 79388 802118 79456 802174
rect 79512 802118 79580 802174
rect 79636 802118 79704 802174
rect 79760 802118 79828 802174
rect 79884 802118 79952 802174
rect 80008 802118 80078 802174
rect 79078 802050 80078 802118
rect 79078 801994 79208 802050
rect 79264 801994 79332 802050
rect 79388 801994 79456 802050
rect 79512 801994 79580 802050
rect 79636 801994 79704 802050
rect 79760 801994 79828 802050
rect 79884 801994 79952 802050
rect 80008 801994 80078 802050
rect 79078 801926 80078 801994
rect 79078 801870 79208 801926
rect 79264 801870 79332 801926
rect 79388 801870 79456 801926
rect 79512 801870 79580 801926
rect 79636 801870 79704 801926
rect 79760 801870 79828 801926
rect 79884 801870 79952 801926
rect 80008 801870 80078 801926
rect 79078 801802 80078 801870
rect 79078 801746 79208 801802
rect 79264 801746 79332 801802
rect 79388 801746 79456 801802
rect 79512 801746 79580 801802
rect 79636 801746 79704 801802
rect 79760 801746 79828 801802
rect 79884 801746 79952 801802
rect 80008 801746 80078 801802
rect 79078 801678 80078 801746
rect 79078 801622 79208 801678
rect 79264 801622 79332 801678
rect 79388 801622 79456 801678
rect 79512 801622 79580 801678
rect 79636 801622 79704 801678
rect 79760 801622 79828 801678
rect 79884 801622 79952 801678
rect 80008 801622 80078 801678
rect 79078 801554 80078 801622
rect 79078 801498 79208 801554
rect 79264 801498 79332 801554
rect 79388 801498 79456 801554
rect 79512 801498 79580 801554
rect 79636 801498 79704 801554
rect 79760 801498 79828 801554
rect 79884 801498 79952 801554
rect 80008 801498 80078 801554
rect 79078 801430 80078 801498
rect 79078 801374 79208 801430
rect 79264 801374 79332 801430
rect 79388 801374 79456 801430
rect 79512 801374 79580 801430
rect 79636 801374 79704 801430
rect 79760 801374 79828 801430
rect 79884 801374 79952 801430
rect 80008 801374 80078 801430
rect 79078 801306 80078 801374
rect 79078 801250 79208 801306
rect 79264 801250 79332 801306
rect 79388 801250 79456 801306
rect 79512 801250 79580 801306
rect 79636 801250 79704 801306
rect 79760 801250 79828 801306
rect 79884 801250 79952 801306
rect 80008 801250 80078 801306
rect 79078 801182 80078 801250
rect 79078 801126 79208 801182
rect 79264 801126 79332 801182
rect 79388 801126 79456 801182
rect 79512 801126 79580 801182
rect 79636 801126 79704 801182
rect 79760 801126 79828 801182
rect 79884 801126 79952 801182
rect 80008 801126 80078 801182
rect 79078 801058 80078 801126
rect 79078 801002 79208 801058
rect 79264 801002 79332 801058
rect 79388 801002 79456 801058
rect 79512 801002 79580 801058
rect 79636 801002 79704 801058
rect 79760 801002 79828 801058
rect 79884 801002 79952 801058
rect 80008 801002 80078 801058
rect 79078 800934 80078 801002
rect 79078 800878 79208 800934
rect 79264 800878 79332 800934
rect 79388 800878 79456 800934
rect 79512 800878 79580 800934
rect 79636 800878 79704 800934
rect 79760 800878 79828 800934
rect 79884 800878 79952 800934
rect 80008 800878 80078 800934
rect 79078 800190 80078 800878
rect 79078 800134 79208 800190
rect 79264 800134 79332 800190
rect 79388 800134 79456 800190
rect 79512 800134 79580 800190
rect 79636 800134 79704 800190
rect 79760 800134 79828 800190
rect 79884 800134 79952 800190
rect 80008 800134 80078 800190
rect 79078 800066 80078 800134
rect 79078 800010 79208 800066
rect 79264 800010 79332 800066
rect 79388 800010 79456 800066
rect 79512 800010 79580 800066
rect 79636 800010 79704 800066
rect 79760 800010 79828 800066
rect 79884 800010 79952 800066
rect 80008 800010 80078 800066
rect 79078 799942 80078 800010
rect 79078 799886 79208 799942
rect 79264 799886 79332 799942
rect 79388 799886 79456 799942
rect 79512 799886 79580 799942
rect 79636 799886 79704 799942
rect 79760 799886 79828 799942
rect 79884 799886 79952 799942
rect 80008 799886 80078 799942
rect 79078 799818 80078 799886
rect 79078 799762 79208 799818
rect 79264 799762 79332 799818
rect 79388 799762 79456 799818
rect 79512 799762 79580 799818
rect 79636 799762 79704 799818
rect 79760 799762 79828 799818
rect 79884 799762 79952 799818
rect 80008 799762 80078 799818
rect 79078 799694 80078 799762
rect 79078 799638 79208 799694
rect 79264 799638 79332 799694
rect 79388 799638 79456 799694
rect 79512 799638 79580 799694
rect 79636 799638 79704 799694
rect 79760 799638 79828 799694
rect 79884 799638 79952 799694
rect 80008 799638 80078 799694
rect 79078 799570 80078 799638
rect 79078 799514 79208 799570
rect 79264 799514 79332 799570
rect 79388 799514 79456 799570
rect 79512 799514 79580 799570
rect 79636 799514 79704 799570
rect 79760 799514 79828 799570
rect 79884 799514 79952 799570
rect 80008 799514 80078 799570
rect 79078 799446 80078 799514
rect 79078 799390 79208 799446
rect 79264 799390 79332 799446
rect 79388 799390 79456 799446
rect 79512 799390 79580 799446
rect 79636 799390 79704 799446
rect 79760 799390 79828 799446
rect 79884 799390 79952 799446
rect 80008 799390 80078 799446
rect 79078 799322 80078 799390
rect 79078 799266 79208 799322
rect 79264 799266 79332 799322
rect 79388 799266 79456 799322
rect 79512 799266 79580 799322
rect 79636 799266 79704 799322
rect 79760 799266 79828 799322
rect 79884 799266 79952 799322
rect 80008 799266 80078 799322
rect 79078 799198 80078 799266
rect 79078 799142 79208 799198
rect 79264 799142 79332 799198
rect 79388 799142 79456 799198
rect 79512 799142 79580 799198
rect 79636 799142 79704 799198
rect 79760 799142 79828 799198
rect 79884 799142 79952 799198
rect 80008 799142 80078 799198
rect 79078 799074 80078 799142
rect 79078 799018 79208 799074
rect 79264 799018 79332 799074
rect 79388 799018 79456 799074
rect 79512 799018 79580 799074
rect 79636 799018 79704 799074
rect 79760 799018 79828 799074
rect 79884 799018 79952 799074
rect 80008 799018 80078 799074
rect 79078 798950 80078 799018
rect 79078 798894 79208 798950
rect 79264 798894 79332 798950
rect 79388 798894 79456 798950
rect 79512 798894 79580 798950
rect 79636 798894 79704 798950
rect 79760 798894 79828 798950
rect 79884 798894 79952 798950
rect 80008 798894 80078 798950
rect 79078 798826 80078 798894
rect 79078 798770 79208 798826
rect 79264 798770 79332 798826
rect 79388 798770 79456 798826
rect 79512 798770 79580 798826
rect 79636 798770 79704 798826
rect 79760 798770 79828 798826
rect 79884 798770 79952 798826
rect 80008 798770 80078 798826
rect 79078 798702 80078 798770
rect 79078 798646 79208 798702
rect 79264 798646 79332 798702
rect 79388 798646 79456 798702
rect 79512 798646 79580 798702
rect 79636 798646 79704 798702
rect 79760 798646 79828 798702
rect 79884 798646 79952 798702
rect 80008 798646 80078 798702
rect 79078 798578 80078 798646
rect 79078 798522 79208 798578
rect 79264 798522 79332 798578
rect 79388 798522 79456 798578
rect 79512 798522 79580 798578
rect 79636 798522 79704 798578
rect 79760 798522 79828 798578
rect 79884 798522 79952 798578
rect 80008 798522 80078 798578
rect 79078 798454 80078 798522
rect 79078 798398 79208 798454
rect 79264 798398 79332 798454
rect 79388 798398 79456 798454
rect 79512 798398 79580 798454
rect 79636 798398 79704 798454
rect 79760 798398 79828 798454
rect 79884 798398 79952 798454
rect 80008 798398 80078 798454
rect 79078 798330 80078 798398
rect 79078 798274 79208 798330
rect 79264 798274 79332 798330
rect 79388 798274 79456 798330
rect 79512 798274 79580 798330
rect 79636 798274 79704 798330
rect 79760 798274 79828 798330
rect 79884 798274 79952 798330
rect 80008 798274 80078 798330
rect 79078 797820 80078 798274
rect 79078 797764 79208 797820
rect 79264 797764 79332 797820
rect 79388 797764 79456 797820
rect 79512 797764 79580 797820
rect 79636 797764 79704 797820
rect 79760 797764 79828 797820
rect 79884 797764 79952 797820
rect 80008 797764 80078 797820
rect 79078 797696 80078 797764
rect 79078 797640 79208 797696
rect 79264 797640 79332 797696
rect 79388 797640 79456 797696
rect 79512 797640 79580 797696
rect 79636 797640 79704 797696
rect 79760 797640 79828 797696
rect 79884 797640 79952 797696
rect 80008 797640 80078 797696
rect 79078 797572 80078 797640
rect 79078 797516 79208 797572
rect 79264 797516 79332 797572
rect 79388 797516 79456 797572
rect 79512 797516 79580 797572
rect 79636 797516 79704 797572
rect 79760 797516 79828 797572
rect 79884 797516 79952 797572
rect 80008 797516 80078 797572
rect 79078 797448 80078 797516
rect 79078 797392 79208 797448
rect 79264 797392 79332 797448
rect 79388 797392 79456 797448
rect 79512 797392 79580 797448
rect 79636 797392 79704 797448
rect 79760 797392 79828 797448
rect 79884 797392 79952 797448
rect 80008 797392 80078 797448
rect 79078 797324 80078 797392
rect 79078 797268 79208 797324
rect 79264 797268 79332 797324
rect 79388 797268 79456 797324
rect 79512 797268 79580 797324
rect 79636 797268 79704 797324
rect 79760 797268 79828 797324
rect 79884 797268 79952 797324
rect 80008 797268 80078 797324
rect 79078 797200 80078 797268
rect 79078 797144 79208 797200
rect 79264 797144 79332 797200
rect 79388 797144 79456 797200
rect 79512 797144 79580 797200
rect 79636 797144 79704 797200
rect 79760 797144 79828 797200
rect 79884 797144 79952 797200
rect 80008 797144 80078 797200
rect 79078 797076 80078 797144
rect 79078 797020 79208 797076
rect 79264 797020 79332 797076
rect 79388 797020 79456 797076
rect 79512 797020 79580 797076
rect 79636 797020 79704 797076
rect 79760 797020 79828 797076
rect 79884 797020 79952 797076
rect 80008 797020 80078 797076
rect 79078 796952 80078 797020
rect 79078 796896 79208 796952
rect 79264 796896 79332 796952
rect 79388 796896 79456 796952
rect 79512 796896 79580 796952
rect 79636 796896 79704 796952
rect 79760 796896 79828 796952
rect 79884 796896 79952 796952
rect 80008 796896 80078 796952
rect 79078 796828 80078 796896
rect 79078 796772 79208 796828
rect 79264 796772 79332 796828
rect 79388 796772 79456 796828
rect 79512 796772 79580 796828
rect 79636 796772 79704 796828
rect 79760 796772 79828 796828
rect 79884 796772 79952 796828
rect 80008 796772 80078 796828
rect 79078 796704 80078 796772
rect 79078 796648 79208 796704
rect 79264 796648 79332 796704
rect 79388 796648 79456 796704
rect 79512 796648 79580 796704
rect 79636 796648 79704 796704
rect 79760 796648 79828 796704
rect 79884 796648 79952 796704
rect 80008 796648 80078 796704
rect 79078 796580 80078 796648
rect 79078 796524 79208 796580
rect 79264 796524 79332 796580
rect 79388 796524 79456 796580
rect 79512 796524 79580 796580
rect 79636 796524 79704 796580
rect 79760 796524 79828 796580
rect 79884 796524 79952 796580
rect 80008 796524 80078 796580
rect 79078 796456 80078 796524
rect 79078 796400 79208 796456
rect 79264 796400 79332 796456
rect 79388 796400 79456 796456
rect 79512 796400 79580 796456
rect 79636 796400 79704 796456
rect 79760 796400 79828 796456
rect 79884 796400 79952 796456
rect 80008 796400 80078 796456
rect 79078 796332 80078 796400
rect 79078 796276 79208 796332
rect 79264 796276 79332 796332
rect 79388 796276 79456 796332
rect 79512 796276 79580 796332
rect 79636 796276 79704 796332
rect 79760 796276 79828 796332
rect 79884 796276 79952 796332
rect 80008 796276 80078 796332
rect 79078 796208 80078 796276
rect 79078 796152 79208 796208
rect 79264 796152 79332 796208
rect 79388 796152 79456 796208
rect 79512 796152 79580 796208
rect 79636 796152 79704 796208
rect 79760 796152 79828 796208
rect 79884 796152 79952 796208
rect 80008 796152 80078 796208
rect 79078 796084 80078 796152
rect 79078 796028 79208 796084
rect 79264 796028 79332 796084
rect 79388 796028 79456 796084
rect 79512 796028 79580 796084
rect 79636 796028 79704 796084
rect 79760 796028 79828 796084
rect 79884 796028 79952 796084
rect 80008 796028 80078 796084
rect 79078 795960 80078 796028
rect 79078 795904 79208 795960
rect 79264 795904 79332 795960
rect 79388 795904 79456 795960
rect 79512 795904 79580 795960
rect 79636 795904 79704 795960
rect 79760 795904 79828 795960
rect 79884 795904 79952 795960
rect 80008 795904 80078 795960
rect 79078 795114 80078 795904
rect 79078 795058 79208 795114
rect 79264 795058 79332 795114
rect 79388 795058 79456 795114
rect 79512 795058 79580 795114
rect 79636 795058 79704 795114
rect 79760 795058 79828 795114
rect 79884 795058 79952 795114
rect 80008 795058 80078 795114
rect 79078 794990 80078 795058
rect 79078 794934 79208 794990
rect 79264 794934 79332 794990
rect 79388 794934 79456 794990
rect 79512 794934 79580 794990
rect 79636 794934 79704 794990
rect 79760 794934 79828 794990
rect 79884 794934 79952 794990
rect 80008 794934 80078 794990
rect 79078 794866 80078 794934
rect 79078 794810 79208 794866
rect 79264 794810 79332 794866
rect 79388 794810 79456 794866
rect 79512 794810 79580 794866
rect 79636 794810 79704 794866
rect 79760 794810 79828 794866
rect 79884 794810 79952 794866
rect 80008 794810 80078 794866
rect 79078 794742 80078 794810
rect 79078 794686 79208 794742
rect 79264 794686 79332 794742
rect 79388 794686 79456 794742
rect 79512 794686 79580 794742
rect 79636 794686 79704 794742
rect 79760 794686 79828 794742
rect 79884 794686 79952 794742
rect 80008 794686 80078 794742
rect 79078 794618 80078 794686
rect 79078 794562 79208 794618
rect 79264 794562 79332 794618
rect 79388 794562 79456 794618
rect 79512 794562 79580 794618
rect 79636 794562 79704 794618
rect 79760 794562 79828 794618
rect 79884 794562 79952 794618
rect 80008 794562 80078 794618
rect 79078 794494 80078 794562
rect 79078 794438 79208 794494
rect 79264 794438 79332 794494
rect 79388 794438 79456 794494
rect 79512 794438 79580 794494
rect 79636 794438 79704 794494
rect 79760 794438 79828 794494
rect 79884 794438 79952 794494
rect 80008 794438 80078 794494
rect 79078 794370 80078 794438
rect 79078 794314 79208 794370
rect 79264 794314 79332 794370
rect 79388 794314 79456 794370
rect 79512 794314 79580 794370
rect 79636 794314 79704 794370
rect 79760 794314 79828 794370
rect 79884 794314 79952 794370
rect 80008 794314 80078 794370
rect 79078 794246 80078 794314
rect 79078 794190 79208 794246
rect 79264 794190 79332 794246
rect 79388 794190 79456 794246
rect 79512 794190 79580 794246
rect 79636 794190 79704 794246
rect 79760 794190 79828 794246
rect 79884 794190 79952 794246
rect 80008 794190 80078 794246
rect 79078 794122 80078 794190
rect 79078 794066 79208 794122
rect 79264 794066 79332 794122
rect 79388 794066 79456 794122
rect 79512 794066 79580 794122
rect 79636 794066 79704 794122
rect 79760 794066 79828 794122
rect 79884 794066 79952 794122
rect 80008 794066 80078 794122
rect 79078 793998 80078 794066
rect 79078 793942 79208 793998
rect 79264 793942 79332 793998
rect 79388 793942 79456 793998
rect 79512 793942 79580 793998
rect 79636 793942 79704 793998
rect 79760 793942 79828 793998
rect 79884 793942 79952 793998
rect 80008 793942 80078 793998
rect 79078 793874 80078 793942
rect 79078 793818 79208 793874
rect 79264 793818 79332 793874
rect 79388 793818 79456 793874
rect 79512 793818 79580 793874
rect 79636 793818 79704 793874
rect 79760 793818 79828 793874
rect 79884 793818 79952 793874
rect 80008 793818 80078 793874
rect 79078 793750 80078 793818
rect 79078 793694 79208 793750
rect 79264 793694 79332 793750
rect 79388 793694 79456 793750
rect 79512 793694 79580 793750
rect 79636 793694 79704 793750
rect 79760 793694 79828 793750
rect 79884 793694 79952 793750
rect 80008 793694 80078 793750
rect 79078 793626 80078 793694
rect 79078 793570 79208 793626
rect 79264 793570 79332 793626
rect 79388 793570 79456 793626
rect 79512 793570 79580 793626
rect 79636 793570 79704 793626
rect 79760 793570 79828 793626
rect 79884 793570 79952 793626
rect 80008 793570 80078 793626
rect 79078 793502 80078 793570
rect 79078 793446 79208 793502
rect 79264 793446 79332 793502
rect 79388 793446 79456 793502
rect 79512 793446 79580 793502
rect 79636 793446 79704 793502
rect 79760 793446 79828 793502
rect 79884 793446 79952 793502
rect 80008 793446 80078 793502
rect 79078 793378 80078 793446
rect 79078 793322 79208 793378
rect 79264 793322 79332 793378
rect 79388 793322 79456 793378
rect 79512 793322 79580 793378
rect 79636 793322 79704 793378
rect 79760 793322 79828 793378
rect 79884 793322 79952 793378
rect 80008 793322 80078 793378
rect 79078 793254 80078 793322
rect 79078 793198 79208 793254
rect 79264 793198 79332 793254
rect 79388 793198 79456 793254
rect 79512 793198 79580 793254
rect 79636 793198 79704 793254
rect 79760 793198 79828 793254
rect 79884 793198 79952 793254
rect 80008 793198 80078 793254
rect 79078 792744 80078 793198
rect 79078 792688 79208 792744
rect 79264 792688 79332 792744
rect 79388 792688 79456 792744
rect 79512 792688 79580 792744
rect 79636 792688 79704 792744
rect 79760 792688 79828 792744
rect 79884 792688 79952 792744
rect 80008 792688 80078 792744
rect 79078 792620 80078 792688
rect 79078 792564 79208 792620
rect 79264 792564 79332 792620
rect 79388 792564 79456 792620
rect 79512 792564 79580 792620
rect 79636 792564 79704 792620
rect 79760 792564 79828 792620
rect 79884 792564 79952 792620
rect 80008 792564 80078 792620
rect 79078 792496 80078 792564
rect 79078 792440 79208 792496
rect 79264 792440 79332 792496
rect 79388 792440 79456 792496
rect 79512 792440 79580 792496
rect 79636 792440 79704 792496
rect 79760 792440 79828 792496
rect 79884 792440 79952 792496
rect 80008 792440 80078 792496
rect 79078 792372 80078 792440
rect 79078 792316 79208 792372
rect 79264 792316 79332 792372
rect 79388 792316 79456 792372
rect 79512 792316 79580 792372
rect 79636 792316 79704 792372
rect 79760 792316 79828 792372
rect 79884 792316 79952 792372
rect 80008 792316 80078 792372
rect 79078 792248 80078 792316
rect 79078 792192 79208 792248
rect 79264 792192 79332 792248
rect 79388 792192 79456 792248
rect 79512 792192 79580 792248
rect 79636 792192 79704 792248
rect 79760 792192 79828 792248
rect 79884 792192 79952 792248
rect 80008 792192 80078 792248
rect 79078 792124 80078 792192
rect 79078 792068 79208 792124
rect 79264 792068 79332 792124
rect 79388 792068 79456 792124
rect 79512 792068 79580 792124
rect 79636 792068 79704 792124
rect 79760 792068 79828 792124
rect 79884 792068 79952 792124
rect 80008 792068 80078 792124
rect 79078 792000 80078 792068
rect 79078 791944 79208 792000
rect 79264 791944 79332 792000
rect 79388 791944 79456 792000
rect 79512 791944 79580 792000
rect 79636 791944 79704 792000
rect 79760 791944 79828 792000
rect 79884 791944 79952 792000
rect 80008 791944 80078 792000
rect 79078 791876 80078 791944
rect 79078 791820 79208 791876
rect 79264 791820 79332 791876
rect 79388 791820 79456 791876
rect 79512 791820 79580 791876
rect 79636 791820 79704 791876
rect 79760 791820 79828 791876
rect 79884 791820 79952 791876
rect 80008 791820 80078 791876
rect 79078 791752 80078 791820
rect 79078 791696 79208 791752
rect 79264 791696 79332 791752
rect 79388 791696 79456 791752
rect 79512 791696 79580 791752
rect 79636 791696 79704 791752
rect 79760 791696 79828 791752
rect 79884 791696 79952 791752
rect 80008 791696 80078 791752
rect 79078 791628 80078 791696
rect 79078 791572 79208 791628
rect 79264 791572 79332 791628
rect 79388 791572 79456 791628
rect 79512 791572 79580 791628
rect 79636 791572 79704 791628
rect 79760 791572 79828 791628
rect 79884 791572 79952 791628
rect 80008 791572 80078 791628
rect 79078 791504 80078 791572
rect 79078 791448 79208 791504
rect 79264 791448 79332 791504
rect 79388 791448 79456 791504
rect 79512 791448 79580 791504
rect 79636 791448 79704 791504
rect 79760 791448 79828 791504
rect 79884 791448 79952 791504
rect 80008 791448 80078 791504
rect 79078 791380 80078 791448
rect 79078 791324 79208 791380
rect 79264 791324 79332 791380
rect 79388 791324 79456 791380
rect 79512 791324 79580 791380
rect 79636 791324 79704 791380
rect 79760 791324 79828 791380
rect 79884 791324 79952 791380
rect 80008 791324 80078 791380
rect 79078 791256 80078 791324
rect 79078 791200 79208 791256
rect 79264 791200 79332 791256
rect 79388 791200 79456 791256
rect 79512 791200 79580 791256
rect 79636 791200 79704 791256
rect 79760 791200 79828 791256
rect 79884 791200 79952 791256
rect 80008 791200 80078 791256
rect 79078 791132 80078 791200
rect 79078 791076 79208 791132
rect 79264 791076 79332 791132
rect 79388 791076 79456 791132
rect 79512 791076 79580 791132
rect 79636 791076 79704 791132
rect 79760 791076 79828 791132
rect 79884 791076 79952 791132
rect 80008 791076 80078 791132
rect 79078 791008 80078 791076
rect 79078 790952 79208 791008
rect 79264 790952 79332 791008
rect 79388 790952 79456 791008
rect 79512 790952 79580 791008
rect 79636 790952 79704 791008
rect 79760 790952 79828 791008
rect 79884 790952 79952 791008
rect 80008 790952 80078 791008
rect 79078 790884 80078 790952
rect 79078 790828 79208 790884
rect 79264 790828 79332 790884
rect 79388 790828 79456 790884
rect 79512 790828 79580 790884
rect 79636 790828 79704 790884
rect 79760 790828 79828 790884
rect 79884 790828 79952 790884
rect 80008 790828 80078 790884
rect 79078 790140 80078 790828
rect 79078 790084 79208 790140
rect 79264 790084 79332 790140
rect 79388 790084 79456 790140
rect 79512 790084 79580 790140
rect 79636 790084 79704 790140
rect 79760 790084 79828 790140
rect 79884 790084 79952 790140
rect 80008 790084 80078 790140
rect 79078 790016 80078 790084
rect 79078 789960 79208 790016
rect 79264 789960 79332 790016
rect 79388 789960 79456 790016
rect 79512 789960 79580 790016
rect 79636 789960 79704 790016
rect 79760 789960 79828 790016
rect 79884 789960 79952 790016
rect 80008 789960 80078 790016
rect 79078 789892 80078 789960
rect 79078 789836 79208 789892
rect 79264 789836 79332 789892
rect 79388 789836 79456 789892
rect 79512 789836 79580 789892
rect 79636 789836 79704 789892
rect 79760 789836 79828 789892
rect 79884 789836 79952 789892
rect 80008 789836 80078 789892
rect 79078 789768 80078 789836
rect 79078 789712 79208 789768
rect 79264 789712 79332 789768
rect 79388 789712 79456 789768
rect 79512 789712 79580 789768
rect 79636 789712 79704 789768
rect 79760 789712 79828 789768
rect 79884 789712 79952 789768
rect 80008 789712 80078 789768
rect 79078 789644 80078 789712
rect 79078 789588 79208 789644
rect 79264 789588 79332 789644
rect 79388 789588 79456 789644
rect 79512 789588 79580 789644
rect 79636 789588 79704 789644
rect 79760 789588 79828 789644
rect 79884 789588 79952 789644
rect 80008 789588 80078 789644
rect 79078 789520 80078 789588
rect 79078 789464 79208 789520
rect 79264 789464 79332 789520
rect 79388 789464 79456 789520
rect 79512 789464 79580 789520
rect 79636 789464 79704 789520
rect 79760 789464 79828 789520
rect 79884 789464 79952 789520
rect 80008 789464 80078 789520
rect 79078 789396 80078 789464
rect 79078 789340 79208 789396
rect 79264 789340 79332 789396
rect 79388 789340 79456 789396
rect 79512 789340 79580 789396
rect 79636 789340 79704 789396
rect 79760 789340 79828 789396
rect 79884 789340 79952 789396
rect 80008 789340 80078 789396
rect 79078 789272 80078 789340
rect 79078 789216 79208 789272
rect 79264 789216 79332 789272
rect 79388 789216 79456 789272
rect 79512 789216 79580 789272
rect 79636 789216 79704 789272
rect 79760 789216 79828 789272
rect 79884 789216 79952 789272
rect 80008 789216 80078 789272
rect 79078 789148 80078 789216
rect 79078 789092 79208 789148
rect 79264 789092 79332 789148
rect 79388 789092 79456 789148
rect 79512 789092 79580 789148
rect 79636 789092 79704 789148
rect 79760 789092 79828 789148
rect 79884 789092 79952 789148
rect 80008 789092 80078 789148
rect 79078 789024 80078 789092
rect 79078 788968 79208 789024
rect 79264 788968 79332 789024
rect 79388 788968 79456 789024
rect 79512 788968 79580 789024
rect 79636 788968 79704 789024
rect 79760 788968 79828 789024
rect 79884 788968 79952 789024
rect 80008 788968 80078 789024
rect 79078 788900 80078 788968
rect 79078 788844 79208 788900
rect 79264 788844 79332 788900
rect 79388 788844 79456 788900
rect 79512 788844 79580 788900
rect 79636 788844 79704 788900
rect 79760 788844 79828 788900
rect 79884 788844 79952 788900
rect 80008 788844 80078 788900
rect 79078 788776 80078 788844
rect 79078 788720 79208 788776
rect 79264 788720 79332 788776
rect 79388 788720 79456 788776
rect 79512 788720 79580 788776
rect 79636 788720 79704 788776
rect 79760 788720 79828 788776
rect 79884 788720 79952 788776
rect 80008 788720 80078 788776
rect 79078 788652 80078 788720
rect 79078 788596 79208 788652
rect 79264 788596 79332 788652
rect 79388 788596 79456 788652
rect 79512 788596 79580 788652
rect 79636 788596 79704 788652
rect 79760 788596 79828 788652
rect 79884 788596 79952 788652
rect 80008 788596 80078 788652
rect 79078 788528 80078 788596
rect 79078 788472 79208 788528
rect 79264 788472 79332 788528
rect 79388 788472 79456 788528
rect 79512 788472 79580 788528
rect 79636 788472 79704 788528
rect 79760 788472 79828 788528
rect 79884 788472 79952 788528
rect 80008 788472 80078 788528
rect 79078 788404 80078 788472
rect 79078 788348 79208 788404
rect 79264 788348 79332 788404
rect 79388 788348 79456 788404
rect 79512 788348 79580 788404
rect 79636 788348 79704 788404
rect 79760 788348 79828 788404
rect 79884 788348 79952 788404
rect 80008 788348 80078 788404
rect 79078 782048 80078 788348
rect 79078 781992 79284 782048
rect 79340 781992 79584 782048
rect 79640 781992 79884 782048
rect 79940 781992 80078 782048
rect 79078 765622 80078 781992
rect 79078 765566 79300 765622
rect 79356 765566 79600 765622
rect 79656 765566 79900 765622
rect 79956 765566 80078 765622
rect 79078 758622 80078 765566
rect 79078 758566 79300 758622
rect 79356 758566 79600 758622
rect 79656 758566 79900 758622
rect 79956 758566 80078 758622
rect 79078 752429 80078 758566
rect 79078 752373 79200 752429
rect 79256 752373 79500 752429
rect 79556 752373 79800 752429
rect 79856 752373 80078 752429
rect 79078 752229 80078 752373
rect 79078 752173 79200 752229
rect 79256 752173 79500 752229
rect 79556 752173 79800 752229
rect 79856 752173 80078 752229
rect 79078 751622 80078 752173
rect 79078 751566 79300 751622
rect 79356 751566 79600 751622
rect 79656 751566 79900 751622
rect 79956 751566 80078 751622
rect 79078 741048 80078 751566
rect 79078 740992 79284 741048
rect 79340 740992 79584 741048
rect 79640 740992 79884 741048
rect 79940 740992 80078 741048
rect 79078 724622 80078 740992
rect 79078 724566 79300 724622
rect 79356 724566 79600 724622
rect 79656 724566 79900 724622
rect 79956 724566 80078 724622
rect 79078 717622 80078 724566
rect 79078 717566 79300 717622
rect 79356 717566 79600 717622
rect 79656 717566 79900 717622
rect 79956 717566 80078 717622
rect 79078 716429 80078 717566
rect 79078 716373 79200 716429
rect 79256 716373 79500 716429
rect 79556 716373 79800 716429
rect 79856 716373 80078 716429
rect 79078 716229 80078 716373
rect 79078 716173 79200 716229
rect 79256 716173 79500 716229
rect 79556 716173 79800 716229
rect 79856 716173 80078 716229
rect 79078 710622 80078 716173
rect 79078 710566 79300 710622
rect 79356 710566 79600 710622
rect 79656 710566 79900 710622
rect 79956 710566 80078 710622
rect 79078 700048 80078 710566
rect 79078 699992 79284 700048
rect 79340 699992 79584 700048
rect 79640 699992 79884 700048
rect 79940 699992 80078 700048
rect 79078 683622 80078 699992
rect 79078 683566 79300 683622
rect 79356 683566 79600 683622
rect 79656 683566 79900 683622
rect 79956 683566 80078 683622
rect 79078 680429 80078 683566
rect 79078 680373 79200 680429
rect 79256 680373 79500 680429
rect 79556 680373 79800 680429
rect 79856 680373 80078 680429
rect 79078 680229 80078 680373
rect 79078 680173 79200 680229
rect 79256 680173 79500 680229
rect 79556 680173 79800 680229
rect 79856 680173 80078 680229
rect 79078 676622 80078 680173
rect 79078 676566 79300 676622
rect 79356 676566 79600 676622
rect 79656 676566 79900 676622
rect 79956 676566 80078 676622
rect 79078 669622 80078 676566
rect 79078 669566 79300 669622
rect 79356 669566 79600 669622
rect 79656 669566 79900 669622
rect 79956 669566 80078 669622
rect 79078 659048 80078 669566
rect 79078 658992 79284 659048
rect 79340 658992 79584 659048
rect 79640 658992 79884 659048
rect 79940 658992 80078 659048
rect 79078 644429 80078 658992
rect 79078 644373 79200 644429
rect 79256 644373 79500 644429
rect 79556 644373 79800 644429
rect 79856 644373 80078 644429
rect 79078 644229 80078 644373
rect 79078 644173 79200 644229
rect 79256 644173 79500 644229
rect 79556 644173 79800 644229
rect 79856 644173 80078 644229
rect 79078 642622 80078 644173
rect 79078 642566 79300 642622
rect 79356 642566 79600 642622
rect 79656 642566 79900 642622
rect 79956 642566 80078 642622
rect 79078 635622 80078 642566
rect 79078 635566 79300 635622
rect 79356 635566 79600 635622
rect 79656 635566 79900 635622
rect 79956 635566 80078 635622
rect 79078 628622 80078 635566
rect 79078 628566 79300 628622
rect 79356 628566 79600 628622
rect 79656 628566 79900 628622
rect 79956 628566 80078 628622
rect 79078 618048 80078 628566
rect 79078 617992 79284 618048
rect 79340 617992 79584 618048
rect 79640 617992 79884 618048
rect 79940 617992 80078 618048
rect 79078 608429 80078 617992
rect 79078 608373 79200 608429
rect 79256 608373 79500 608429
rect 79556 608373 79800 608429
rect 79856 608373 80078 608429
rect 79078 608229 80078 608373
rect 79078 608173 79200 608229
rect 79256 608173 79500 608229
rect 79556 608173 79800 608229
rect 79856 608173 80078 608229
rect 79078 601622 80078 608173
rect 79078 601566 79300 601622
rect 79356 601566 79600 601622
rect 79656 601566 79900 601622
rect 79956 601566 80078 601622
rect 79078 594622 80078 601566
rect 79078 594566 79300 594622
rect 79356 594566 79600 594622
rect 79656 594566 79900 594622
rect 79956 594566 80078 594622
rect 79078 587622 80078 594566
rect 79078 587566 79300 587622
rect 79356 587566 79600 587622
rect 79656 587566 79900 587622
rect 79956 587566 80078 587622
rect 79078 577048 80078 587566
rect 79078 576992 79284 577048
rect 79340 576992 79584 577048
rect 79640 576992 79884 577048
rect 79940 576992 80078 577048
rect 79078 572429 80078 576992
rect 79078 572373 79200 572429
rect 79256 572373 79500 572429
rect 79556 572373 79800 572429
rect 79856 572373 80078 572429
rect 79078 572229 80078 572373
rect 79078 572173 79200 572229
rect 79256 572173 79500 572229
rect 79556 572173 79800 572229
rect 79856 572173 80078 572229
rect 79078 560622 80078 572173
rect 79078 560566 79300 560622
rect 79356 560566 79600 560622
rect 79656 560566 79900 560622
rect 79956 560566 80078 560622
rect 79078 553622 80078 560566
rect 79078 553566 79300 553622
rect 79356 553566 79600 553622
rect 79656 553566 79900 553622
rect 79956 553566 80078 553622
rect 79078 546622 80078 553566
rect 79078 546566 79300 546622
rect 79356 546566 79600 546622
rect 79656 546566 79900 546622
rect 79956 546566 80078 546622
rect 79078 536429 80078 546566
rect 79078 536373 79200 536429
rect 79256 536373 79500 536429
rect 79556 536373 79800 536429
rect 79856 536373 80078 536429
rect 79078 536229 80078 536373
rect 79078 536173 79200 536229
rect 79256 536173 79500 536229
rect 79556 536173 79800 536229
rect 79856 536173 80078 536229
rect 79078 536048 80078 536173
rect 79078 535992 79284 536048
rect 79340 535992 79584 536048
rect 79640 535992 79884 536048
rect 79940 535992 80078 536048
rect 79078 519622 80078 535992
rect 79078 519566 79300 519622
rect 79356 519566 79600 519622
rect 79656 519566 79900 519622
rect 79956 519566 80078 519622
rect 79078 512622 80078 519566
rect 79078 512566 79300 512622
rect 79356 512566 79600 512622
rect 79656 512566 79900 512622
rect 79956 512566 80078 512622
rect 79078 505622 80078 512566
rect 79078 505566 79300 505622
rect 79356 505566 79600 505622
rect 79656 505566 79900 505622
rect 79956 505566 80078 505622
rect 79078 500429 80078 505566
rect 79078 500373 79200 500429
rect 79256 500373 79500 500429
rect 79556 500373 79800 500429
rect 79856 500373 80078 500429
rect 79078 500229 80078 500373
rect 79078 500173 79200 500229
rect 79256 500173 79500 500229
rect 79556 500173 79800 500229
rect 79856 500173 80078 500229
rect 79078 433670 80078 500173
rect 79078 433614 79208 433670
rect 79264 433614 79332 433670
rect 79388 433614 79456 433670
rect 79512 433614 79580 433670
rect 79636 433614 79704 433670
rect 79760 433614 79828 433670
rect 79884 433614 79952 433670
rect 80008 433614 80078 433670
rect 79078 433546 80078 433614
rect 79078 433490 79208 433546
rect 79264 433490 79332 433546
rect 79388 433490 79456 433546
rect 79512 433490 79580 433546
rect 79636 433490 79704 433546
rect 79760 433490 79828 433546
rect 79884 433490 79952 433546
rect 80008 433490 80078 433546
rect 79078 433422 80078 433490
rect 79078 433366 79208 433422
rect 79264 433366 79332 433422
rect 79388 433366 79456 433422
rect 79512 433366 79580 433422
rect 79636 433366 79704 433422
rect 79760 433366 79828 433422
rect 79884 433366 79952 433422
rect 80008 433366 80078 433422
rect 79078 433298 80078 433366
rect 79078 433242 79208 433298
rect 79264 433242 79332 433298
rect 79388 433242 79456 433298
rect 79512 433242 79580 433298
rect 79636 433242 79704 433298
rect 79760 433242 79828 433298
rect 79884 433242 79952 433298
rect 80008 433242 80078 433298
rect 79078 433174 80078 433242
rect 79078 433118 79208 433174
rect 79264 433118 79332 433174
rect 79388 433118 79456 433174
rect 79512 433118 79580 433174
rect 79636 433118 79704 433174
rect 79760 433118 79828 433174
rect 79884 433118 79952 433174
rect 80008 433118 80078 433174
rect 79078 433050 80078 433118
rect 79078 432994 79208 433050
rect 79264 432994 79332 433050
rect 79388 432994 79456 433050
rect 79512 432994 79580 433050
rect 79636 432994 79704 433050
rect 79760 432994 79828 433050
rect 79884 432994 79952 433050
rect 80008 432994 80078 433050
rect 79078 432926 80078 432994
rect 79078 432870 79208 432926
rect 79264 432870 79332 432926
rect 79388 432870 79456 432926
rect 79512 432870 79580 432926
rect 79636 432870 79704 432926
rect 79760 432870 79828 432926
rect 79884 432870 79952 432926
rect 80008 432870 80078 432926
rect 79078 432802 80078 432870
rect 79078 432746 79208 432802
rect 79264 432746 79332 432802
rect 79388 432746 79456 432802
rect 79512 432746 79580 432802
rect 79636 432746 79704 432802
rect 79760 432746 79828 432802
rect 79884 432746 79952 432802
rect 80008 432746 80078 432802
rect 79078 432678 80078 432746
rect 79078 432622 79208 432678
rect 79264 432622 79332 432678
rect 79388 432622 79456 432678
rect 79512 432622 79580 432678
rect 79636 432622 79704 432678
rect 79760 432622 79828 432678
rect 79884 432622 79952 432678
rect 80008 432622 80078 432678
rect 79078 432554 80078 432622
rect 79078 432498 79208 432554
rect 79264 432498 79332 432554
rect 79388 432498 79456 432554
rect 79512 432498 79580 432554
rect 79636 432498 79704 432554
rect 79760 432498 79828 432554
rect 79884 432498 79952 432554
rect 80008 432498 80078 432554
rect 79078 432430 80078 432498
rect 79078 432374 79208 432430
rect 79264 432374 79332 432430
rect 79388 432374 79456 432430
rect 79512 432374 79580 432430
rect 79636 432374 79704 432430
rect 79760 432374 79828 432430
rect 79884 432374 79952 432430
rect 80008 432374 80078 432430
rect 79078 432306 80078 432374
rect 79078 432250 79208 432306
rect 79264 432250 79332 432306
rect 79388 432250 79456 432306
rect 79512 432250 79580 432306
rect 79636 432250 79704 432306
rect 79760 432250 79828 432306
rect 79884 432250 79952 432306
rect 80008 432250 80078 432306
rect 79078 432182 80078 432250
rect 79078 432126 79208 432182
rect 79264 432126 79332 432182
rect 79388 432126 79456 432182
rect 79512 432126 79580 432182
rect 79636 432126 79704 432182
rect 79760 432126 79828 432182
rect 79884 432126 79952 432182
rect 80008 432126 80078 432182
rect 79078 432058 80078 432126
rect 79078 432002 79208 432058
rect 79264 432002 79332 432058
rect 79388 432002 79456 432058
rect 79512 432002 79580 432058
rect 79636 432002 79704 432058
rect 79760 432002 79828 432058
rect 79884 432002 79952 432058
rect 80008 432002 80078 432058
rect 79078 431934 80078 432002
rect 79078 431878 79208 431934
rect 79264 431878 79332 431934
rect 79388 431878 79456 431934
rect 79512 431878 79580 431934
rect 79636 431878 79704 431934
rect 79760 431878 79828 431934
rect 79884 431878 79952 431934
rect 80008 431878 80078 431934
rect 79078 431190 80078 431878
rect 79078 431134 79208 431190
rect 79264 431134 79332 431190
rect 79388 431134 79456 431190
rect 79512 431134 79580 431190
rect 79636 431134 79704 431190
rect 79760 431134 79828 431190
rect 79884 431134 79952 431190
rect 80008 431134 80078 431190
rect 79078 431066 80078 431134
rect 79078 431010 79208 431066
rect 79264 431010 79332 431066
rect 79388 431010 79456 431066
rect 79512 431010 79580 431066
rect 79636 431010 79704 431066
rect 79760 431010 79828 431066
rect 79884 431010 79952 431066
rect 80008 431010 80078 431066
rect 79078 430942 80078 431010
rect 79078 430886 79208 430942
rect 79264 430886 79332 430942
rect 79388 430886 79456 430942
rect 79512 430886 79580 430942
rect 79636 430886 79704 430942
rect 79760 430886 79828 430942
rect 79884 430886 79952 430942
rect 80008 430886 80078 430942
rect 79078 430818 80078 430886
rect 79078 430762 79208 430818
rect 79264 430762 79332 430818
rect 79388 430762 79456 430818
rect 79512 430762 79580 430818
rect 79636 430762 79704 430818
rect 79760 430762 79828 430818
rect 79884 430762 79952 430818
rect 80008 430762 80078 430818
rect 79078 430694 80078 430762
rect 79078 430638 79208 430694
rect 79264 430638 79332 430694
rect 79388 430638 79456 430694
rect 79512 430638 79580 430694
rect 79636 430638 79704 430694
rect 79760 430638 79828 430694
rect 79884 430638 79952 430694
rect 80008 430638 80078 430694
rect 79078 430570 80078 430638
rect 79078 430514 79208 430570
rect 79264 430514 79332 430570
rect 79388 430514 79456 430570
rect 79512 430514 79580 430570
rect 79636 430514 79704 430570
rect 79760 430514 79828 430570
rect 79884 430514 79952 430570
rect 80008 430514 80078 430570
rect 79078 430446 80078 430514
rect 79078 430390 79208 430446
rect 79264 430390 79332 430446
rect 79388 430390 79456 430446
rect 79512 430390 79580 430446
rect 79636 430390 79704 430446
rect 79760 430390 79828 430446
rect 79884 430390 79952 430446
rect 80008 430390 80078 430446
rect 79078 430322 80078 430390
rect 79078 430266 79208 430322
rect 79264 430266 79332 430322
rect 79388 430266 79456 430322
rect 79512 430266 79580 430322
rect 79636 430266 79704 430322
rect 79760 430266 79828 430322
rect 79884 430266 79952 430322
rect 80008 430266 80078 430322
rect 79078 430198 80078 430266
rect 79078 430142 79208 430198
rect 79264 430142 79332 430198
rect 79388 430142 79456 430198
rect 79512 430142 79580 430198
rect 79636 430142 79704 430198
rect 79760 430142 79828 430198
rect 79884 430142 79952 430198
rect 80008 430142 80078 430198
rect 79078 430074 80078 430142
rect 79078 430018 79208 430074
rect 79264 430018 79332 430074
rect 79388 430018 79456 430074
rect 79512 430018 79580 430074
rect 79636 430018 79704 430074
rect 79760 430018 79828 430074
rect 79884 430018 79952 430074
rect 80008 430018 80078 430074
rect 79078 429950 80078 430018
rect 79078 429894 79208 429950
rect 79264 429894 79332 429950
rect 79388 429894 79456 429950
rect 79512 429894 79580 429950
rect 79636 429894 79704 429950
rect 79760 429894 79828 429950
rect 79884 429894 79952 429950
rect 80008 429894 80078 429950
rect 79078 429826 80078 429894
rect 79078 429770 79208 429826
rect 79264 429770 79332 429826
rect 79388 429770 79456 429826
rect 79512 429770 79580 429826
rect 79636 429770 79704 429826
rect 79760 429770 79828 429826
rect 79884 429770 79952 429826
rect 80008 429770 80078 429826
rect 79078 429702 80078 429770
rect 79078 429646 79208 429702
rect 79264 429646 79332 429702
rect 79388 429646 79456 429702
rect 79512 429646 79580 429702
rect 79636 429646 79704 429702
rect 79760 429646 79828 429702
rect 79884 429646 79952 429702
rect 80008 429646 80078 429702
rect 79078 429578 80078 429646
rect 79078 429522 79208 429578
rect 79264 429522 79332 429578
rect 79388 429522 79456 429578
rect 79512 429522 79580 429578
rect 79636 429522 79704 429578
rect 79760 429522 79828 429578
rect 79884 429522 79952 429578
rect 80008 429522 80078 429578
rect 79078 429454 80078 429522
rect 79078 429398 79208 429454
rect 79264 429398 79332 429454
rect 79388 429398 79456 429454
rect 79512 429398 79580 429454
rect 79636 429398 79704 429454
rect 79760 429398 79828 429454
rect 79884 429398 79952 429454
rect 80008 429398 80078 429454
rect 79078 429330 80078 429398
rect 79078 429274 79208 429330
rect 79264 429274 79332 429330
rect 79388 429274 79456 429330
rect 79512 429274 79580 429330
rect 79636 429274 79704 429330
rect 79760 429274 79828 429330
rect 79884 429274 79952 429330
rect 80008 429274 80078 429330
rect 79078 428820 80078 429274
rect 79078 428764 79208 428820
rect 79264 428764 79332 428820
rect 79388 428764 79456 428820
rect 79512 428764 79580 428820
rect 79636 428764 79704 428820
rect 79760 428764 79828 428820
rect 79884 428764 79952 428820
rect 80008 428764 80078 428820
rect 79078 428696 80078 428764
rect 79078 428640 79208 428696
rect 79264 428640 79332 428696
rect 79388 428640 79456 428696
rect 79512 428640 79580 428696
rect 79636 428640 79704 428696
rect 79760 428640 79828 428696
rect 79884 428640 79952 428696
rect 80008 428640 80078 428696
rect 79078 428572 80078 428640
rect 79078 428516 79208 428572
rect 79264 428516 79332 428572
rect 79388 428516 79456 428572
rect 79512 428516 79580 428572
rect 79636 428516 79704 428572
rect 79760 428516 79828 428572
rect 79884 428516 79952 428572
rect 80008 428516 80078 428572
rect 79078 428448 80078 428516
rect 79078 428392 79208 428448
rect 79264 428392 79332 428448
rect 79388 428392 79456 428448
rect 79512 428392 79580 428448
rect 79636 428392 79704 428448
rect 79760 428392 79828 428448
rect 79884 428392 79952 428448
rect 80008 428392 80078 428448
rect 79078 428324 80078 428392
rect 79078 428268 79208 428324
rect 79264 428268 79332 428324
rect 79388 428268 79456 428324
rect 79512 428268 79580 428324
rect 79636 428268 79704 428324
rect 79760 428268 79828 428324
rect 79884 428268 79952 428324
rect 80008 428268 80078 428324
rect 79078 428200 80078 428268
rect 79078 428144 79208 428200
rect 79264 428144 79332 428200
rect 79388 428144 79456 428200
rect 79512 428144 79580 428200
rect 79636 428144 79704 428200
rect 79760 428144 79828 428200
rect 79884 428144 79952 428200
rect 80008 428144 80078 428200
rect 79078 428076 80078 428144
rect 79078 428020 79208 428076
rect 79264 428020 79332 428076
rect 79388 428020 79456 428076
rect 79512 428020 79580 428076
rect 79636 428020 79704 428076
rect 79760 428020 79828 428076
rect 79884 428020 79952 428076
rect 80008 428020 80078 428076
rect 79078 427952 80078 428020
rect 79078 427896 79208 427952
rect 79264 427896 79332 427952
rect 79388 427896 79456 427952
rect 79512 427896 79580 427952
rect 79636 427896 79704 427952
rect 79760 427896 79828 427952
rect 79884 427896 79952 427952
rect 80008 427896 80078 427952
rect 79078 427828 80078 427896
rect 79078 427772 79208 427828
rect 79264 427772 79332 427828
rect 79388 427772 79456 427828
rect 79512 427772 79580 427828
rect 79636 427772 79704 427828
rect 79760 427772 79828 427828
rect 79884 427772 79952 427828
rect 80008 427772 80078 427828
rect 79078 427704 80078 427772
rect 79078 427648 79208 427704
rect 79264 427648 79332 427704
rect 79388 427648 79456 427704
rect 79512 427648 79580 427704
rect 79636 427648 79704 427704
rect 79760 427648 79828 427704
rect 79884 427648 79952 427704
rect 80008 427648 80078 427704
rect 79078 427580 80078 427648
rect 79078 427524 79208 427580
rect 79264 427524 79332 427580
rect 79388 427524 79456 427580
rect 79512 427524 79580 427580
rect 79636 427524 79704 427580
rect 79760 427524 79828 427580
rect 79884 427524 79952 427580
rect 80008 427524 80078 427580
rect 79078 427456 80078 427524
rect 79078 427400 79208 427456
rect 79264 427400 79332 427456
rect 79388 427400 79456 427456
rect 79512 427400 79580 427456
rect 79636 427400 79704 427456
rect 79760 427400 79828 427456
rect 79884 427400 79952 427456
rect 80008 427400 80078 427456
rect 79078 427332 80078 427400
rect 79078 427276 79208 427332
rect 79264 427276 79332 427332
rect 79388 427276 79456 427332
rect 79512 427276 79580 427332
rect 79636 427276 79704 427332
rect 79760 427276 79828 427332
rect 79884 427276 79952 427332
rect 80008 427276 80078 427332
rect 79078 427208 80078 427276
rect 79078 427152 79208 427208
rect 79264 427152 79332 427208
rect 79388 427152 79456 427208
rect 79512 427152 79580 427208
rect 79636 427152 79704 427208
rect 79760 427152 79828 427208
rect 79884 427152 79952 427208
rect 80008 427152 80078 427208
rect 79078 427084 80078 427152
rect 79078 427028 79208 427084
rect 79264 427028 79332 427084
rect 79388 427028 79456 427084
rect 79512 427028 79580 427084
rect 79636 427028 79704 427084
rect 79760 427028 79828 427084
rect 79884 427028 79952 427084
rect 80008 427028 80078 427084
rect 79078 426960 80078 427028
rect 79078 426904 79208 426960
rect 79264 426904 79332 426960
rect 79388 426904 79456 426960
rect 79512 426904 79580 426960
rect 79636 426904 79704 426960
rect 79760 426904 79828 426960
rect 79884 426904 79952 426960
rect 80008 426904 80078 426960
rect 79078 426114 80078 426904
rect 79078 426058 79208 426114
rect 79264 426058 79332 426114
rect 79388 426058 79456 426114
rect 79512 426058 79580 426114
rect 79636 426058 79704 426114
rect 79760 426058 79828 426114
rect 79884 426058 79952 426114
rect 80008 426058 80078 426114
rect 79078 425990 80078 426058
rect 79078 425934 79208 425990
rect 79264 425934 79332 425990
rect 79388 425934 79456 425990
rect 79512 425934 79580 425990
rect 79636 425934 79704 425990
rect 79760 425934 79828 425990
rect 79884 425934 79952 425990
rect 80008 425934 80078 425990
rect 79078 425866 80078 425934
rect 79078 425810 79208 425866
rect 79264 425810 79332 425866
rect 79388 425810 79456 425866
rect 79512 425810 79580 425866
rect 79636 425810 79704 425866
rect 79760 425810 79828 425866
rect 79884 425810 79952 425866
rect 80008 425810 80078 425866
rect 79078 425742 80078 425810
rect 79078 425686 79208 425742
rect 79264 425686 79332 425742
rect 79388 425686 79456 425742
rect 79512 425686 79580 425742
rect 79636 425686 79704 425742
rect 79760 425686 79828 425742
rect 79884 425686 79952 425742
rect 80008 425686 80078 425742
rect 79078 425618 80078 425686
rect 79078 425562 79208 425618
rect 79264 425562 79332 425618
rect 79388 425562 79456 425618
rect 79512 425562 79580 425618
rect 79636 425562 79704 425618
rect 79760 425562 79828 425618
rect 79884 425562 79952 425618
rect 80008 425562 80078 425618
rect 79078 425494 80078 425562
rect 79078 425438 79208 425494
rect 79264 425438 79332 425494
rect 79388 425438 79456 425494
rect 79512 425438 79580 425494
rect 79636 425438 79704 425494
rect 79760 425438 79828 425494
rect 79884 425438 79952 425494
rect 80008 425438 80078 425494
rect 79078 425370 80078 425438
rect 79078 425314 79208 425370
rect 79264 425314 79332 425370
rect 79388 425314 79456 425370
rect 79512 425314 79580 425370
rect 79636 425314 79704 425370
rect 79760 425314 79828 425370
rect 79884 425314 79952 425370
rect 80008 425314 80078 425370
rect 79078 425246 80078 425314
rect 79078 425190 79208 425246
rect 79264 425190 79332 425246
rect 79388 425190 79456 425246
rect 79512 425190 79580 425246
rect 79636 425190 79704 425246
rect 79760 425190 79828 425246
rect 79884 425190 79952 425246
rect 80008 425190 80078 425246
rect 79078 425122 80078 425190
rect 79078 425066 79208 425122
rect 79264 425066 79332 425122
rect 79388 425066 79456 425122
rect 79512 425066 79580 425122
rect 79636 425066 79704 425122
rect 79760 425066 79828 425122
rect 79884 425066 79952 425122
rect 80008 425066 80078 425122
rect 79078 424998 80078 425066
rect 79078 424942 79208 424998
rect 79264 424942 79332 424998
rect 79388 424942 79456 424998
rect 79512 424942 79580 424998
rect 79636 424942 79704 424998
rect 79760 424942 79828 424998
rect 79884 424942 79952 424998
rect 80008 424942 80078 424998
rect 79078 424874 80078 424942
rect 79078 424818 79208 424874
rect 79264 424818 79332 424874
rect 79388 424818 79456 424874
rect 79512 424818 79580 424874
rect 79636 424818 79704 424874
rect 79760 424818 79828 424874
rect 79884 424818 79952 424874
rect 80008 424818 80078 424874
rect 79078 424750 80078 424818
rect 79078 424694 79208 424750
rect 79264 424694 79332 424750
rect 79388 424694 79456 424750
rect 79512 424694 79580 424750
rect 79636 424694 79704 424750
rect 79760 424694 79828 424750
rect 79884 424694 79952 424750
rect 80008 424694 80078 424750
rect 79078 424626 80078 424694
rect 79078 424570 79208 424626
rect 79264 424570 79332 424626
rect 79388 424570 79456 424626
rect 79512 424570 79580 424626
rect 79636 424570 79704 424626
rect 79760 424570 79828 424626
rect 79884 424570 79952 424626
rect 80008 424570 80078 424626
rect 79078 424502 80078 424570
rect 79078 424446 79208 424502
rect 79264 424446 79332 424502
rect 79388 424446 79456 424502
rect 79512 424446 79580 424502
rect 79636 424446 79704 424502
rect 79760 424446 79828 424502
rect 79884 424446 79952 424502
rect 80008 424446 80078 424502
rect 79078 424378 80078 424446
rect 79078 424322 79208 424378
rect 79264 424322 79332 424378
rect 79388 424322 79456 424378
rect 79512 424322 79580 424378
rect 79636 424322 79704 424378
rect 79760 424322 79828 424378
rect 79884 424322 79952 424378
rect 80008 424322 80078 424378
rect 79078 424254 80078 424322
rect 79078 424198 79208 424254
rect 79264 424198 79332 424254
rect 79388 424198 79456 424254
rect 79512 424198 79580 424254
rect 79636 424198 79704 424254
rect 79760 424198 79828 424254
rect 79884 424198 79952 424254
rect 80008 424198 80078 424254
rect 79078 423744 80078 424198
rect 79078 423688 79208 423744
rect 79264 423688 79332 423744
rect 79388 423688 79456 423744
rect 79512 423688 79580 423744
rect 79636 423688 79704 423744
rect 79760 423688 79828 423744
rect 79884 423688 79952 423744
rect 80008 423688 80078 423744
rect 79078 423620 80078 423688
rect 79078 423564 79208 423620
rect 79264 423564 79332 423620
rect 79388 423564 79456 423620
rect 79512 423564 79580 423620
rect 79636 423564 79704 423620
rect 79760 423564 79828 423620
rect 79884 423564 79952 423620
rect 80008 423564 80078 423620
rect 79078 423496 80078 423564
rect 79078 423440 79208 423496
rect 79264 423440 79332 423496
rect 79388 423440 79456 423496
rect 79512 423440 79580 423496
rect 79636 423440 79704 423496
rect 79760 423440 79828 423496
rect 79884 423440 79952 423496
rect 80008 423440 80078 423496
rect 79078 423372 80078 423440
rect 79078 423316 79208 423372
rect 79264 423316 79332 423372
rect 79388 423316 79456 423372
rect 79512 423316 79580 423372
rect 79636 423316 79704 423372
rect 79760 423316 79828 423372
rect 79884 423316 79952 423372
rect 80008 423316 80078 423372
rect 79078 423248 80078 423316
rect 79078 423192 79208 423248
rect 79264 423192 79332 423248
rect 79388 423192 79456 423248
rect 79512 423192 79580 423248
rect 79636 423192 79704 423248
rect 79760 423192 79828 423248
rect 79884 423192 79952 423248
rect 80008 423192 80078 423248
rect 79078 423124 80078 423192
rect 79078 423068 79208 423124
rect 79264 423068 79332 423124
rect 79388 423068 79456 423124
rect 79512 423068 79580 423124
rect 79636 423068 79704 423124
rect 79760 423068 79828 423124
rect 79884 423068 79952 423124
rect 80008 423068 80078 423124
rect 79078 423000 80078 423068
rect 79078 422944 79208 423000
rect 79264 422944 79332 423000
rect 79388 422944 79456 423000
rect 79512 422944 79580 423000
rect 79636 422944 79704 423000
rect 79760 422944 79828 423000
rect 79884 422944 79952 423000
rect 80008 422944 80078 423000
rect 79078 422876 80078 422944
rect 79078 422820 79208 422876
rect 79264 422820 79332 422876
rect 79388 422820 79456 422876
rect 79512 422820 79580 422876
rect 79636 422820 79704 422876
rect 79760 422820 79828 422876
rect 79884 422820 79952 422876
rect 80008 422820 80078 422876
rect 79078 422752 80078 422820
rect 79078 422696 79208 422752
rect 79264 422696 79332 422752
rect 79388 422696 79456 422752
rect 79512 422696 79580 422752
rect 79636 422696 79704 422752
rect 79760 422696 79828 422752
rect 79884 422696 79952 422752
rect 80008 422696 80078 422752
rect 79078 422628 80078 422696
rect 79078 422572 79208 422628
rect 79264 422572 79332 422628
rect 79388 422572 79456 422628
rect 79512 422572 79580 422628
rect 79636 422572 79704 422628
rect 79760 422572 79828 422628
rect 79884 422572 79952 422628
rect 80008 422572 80078 422628
rect 79078 422504 80078 422572
rect 79078 422448 79208 422504
rect 79264 422448 79332 422504
rect 79388 422448 79456 422504
rect 79512 422448 79580 422504
rect 79636 422448 79704 422504
rect 79760 422448 79828 422504
rect 79884 422448 79952 422504
rect 80008 422448 80078 422504
rect 79078 422380 80078 422448
rect 79078 422324 79208 422380
rect 79264 422324 79332 422380
rect 79388 422324 79456 422380
rect 79512 422324 79580 422380
rect 79636 422324 79704 422380
rect 79760 422324 79828 422380
rect 79884 422324 79952 422380
rect 80008 422324 80078 422380
rect 79078 422256 80078 422324
rect 79078 422200 79208 422256
rect 79264 422200 79332 422256
rect 79388 422200 79456 422256
rect 79512 422200 79580 422256
rect 79636 422200 79704 422256
rect 79760 422200 79828 422256
rect 79884 422200 79952 422256
rect 80008 422200 80078 422256
rect 79078 422132 80078 422200
rect 79078 422076 79208 422132
rect 79264 422076 79332 422132
rect 79388 422076 79456 422132
rect 79512 422076 79580 422132
rect 79636 422076 79704 422132
rect 79760 422076 79828 422132
rect 79884 422076 79952 422132
rect 80008 422076 80078 422132
rect 79078 422008 80078 422076
rect 79078 421952 79208 422008
rect 79264 421952 79332 422008
rect 79388 421952 79456 422008
rect 79512 421952 79580 422008
rect 79636 421952 79704 422008
rect 79760 421952 79828 422008
rect 79884 421952 79952 422008
rect 80008 421952 80078 422008
rect 79078 421884 80078 421952
rect 79078 421828 79208 421884
rect 79264 421828 79332 421884
rect 79388 421828 79456 421884
rect 79512 421828 79580 421884
rect 79636 421828 79704 421884
rect 79760 421828 79828 421884
rect 79884 421828 79952 421884
rect 80008 421828 80078 421884
rect 79078 421140 80078 421828
rect 79078 421084 79208 421140
rect 79264 421084 79332 421140
rect 79388 421084 79456 421140
rect 79512 421084 79580 421140
rect 79636 421084 79704 421140
rect 79760 421084 79828 421140
rect 79884 421084 79952 421140
rect 80008 421084 80078 421140
rect 79078 421016 80078 421084
rect 79078 420960 79208 421016
rect 79264 420960 79332 421016
rect 79388 420960 79456 421016
rect 79512 420960 79580 421016
rect 79636 420960 79704 421016
rect 79760 420960 79828 421016
rect 79884 420960 79952 421016
rect 80008 420960 80078 421016
rect 79078 420892 80078 420960
rect 79078 420836 79208 420892
rect 79264 420836 79332 420892
rect 79388 420836 79456 420892
rect 79512 420836 79580 420892
rect 79636 420836 79704 420892
rect 79760 420836 79828 420892
rect 79884 420836 79952 420892
rect 80008 420836 80078 420892
rect 79078 420768 80078 420836
rect 79078 420712 79208 420768
rect 79264 420712 79332 420768
rect 79388 420712 79456 420768
rect 79512 420712 79580 420768
rect 79636 420712 79704 420768
rect 79760 420712 79828 420768
rect 79884 420712 79952 420768
rect 80008 420712 80078 420768
rect 79078 420644 80078 420712
rect 79078 420588 79208 420644
rect 79264 420588 79332 420644
rect 79388 420588 79456 420644
rect 79512 420588 79580 420644
rect 79636 420588 79704 420644
rect 79760 420588 79828 420644
rect 79884 420588 79952 420644
rect 80008 420588 80078 420644
rect 79078 420520 80078 420588
rect 79078 420464 79208 420520
rect 79264 420464 79332 420520
rect 79388 420464 79456 420520
rect 79512 420464 79580 420520
rect 79636 420464 79704 420520
rect 79760 420464 79828 420520
rect 79884 420464 79952 420520
rect 80008 420464 80078 420520
rect 79078 420396 80078 420464
rect 79078 420340 79208 420396
rect 79264 420340 79332 420396
rect 79388 420340 79456 420396
rect 79512 420340 79580 420396
rect 79636 420340 79704 420396
rect 79760 420340 79828 420396
rect 79884 420340 79952 420396
rect 80008 420340 80078 420396
rect 79078 420272 80078 420340
rect 79078 420216 79208 420272
rect 79264 420216 79332 420272
rect 79388 420216 79456 420272
rect 79512 420216 79580 420272
rect 79636 420216 79704 420272
rect 79760 420216 79828 420272
rect 79884 420216 79952 420272
rect 80008 420216 80078 420272
rect 79078 420148 80078 420216
rect 79078 420092 79208 420148
rect 79264 420092 79332 420148
rect 79388 420092 79456 420148
rect 79512 420092 79580 420148
rect 79636 420092 79704 420148
rect 79760 420092 79828 420148
rect 79884 420092 79952 420148
rect 80008 420092 80078 420148
rect 79078 420024 80078 420092
rect 79078 419968 79208 420024
rect 79264 419968 79332 420024
rect 79388 419968 79456 420024
rect 79512 419968 79580 420024
rect 79636 419968 79704 420024
rect 79760 419968 79828 420024
rect 79884 419968 79952 420024
rect 80008 419968 80078 420024
rect 79078 419900 80078 419968
rect 79078 419844 79208 419900
rect 79264 419844 79332 419900
rect 79388 419844 79456 419900
rect 79512 419844 79580 419900
rect 79636 419844 79704 419900
rect 79760 419844 79828 419900
rect 79884 419844 79952 419900
rect 80008 419844 80078 419900
rect 79078 419776 80078 419844
rect 79078 419720 79208 419776
rect 79264 419720 79332 419776
rect 79388 419720 79456 419776
rect 79512 419720 79580 419776
rect 79636 419720 79704 419776
rect 79760 419720 79828 419776
rect 79884 419720 79952 419776
rect 80008 419720 80078 419776
rect 79078 419652 80078 419720
rect 79078 419596 79208 419652
rect 79264 419596 79332 419652
rect 79388 419596 79456 419652
rect 79512 419596 79580 419652
rect 79636 419596 79704 419652
rect 79760 419596 79828 419652
rect 79884 419596 79952 419652
rect 80008 419596 80078 419652
rect 79078 419528 80078 419596
rect 79078 419472 79208 419528
rect 79264 419472 79332 419528
rect 79388 419472 79456 419528
rect 79512 419472 79580 419528
rect 79636 419472 79704 419528
rect 79760 419472 79828 419528
rect 79884 419472 79952 419528
rect 80008 419472 80078 419528
rect 79078 419404 80078 419472
rect 79078 419348 79208 419404
rect 79264 419348 79332 419404
rect 79388 419348 79456 419404
rect 79512 419348 79580 419404
rect 79636 419348 79704 419404
rect 79760 419348 79828 419404
rect 79884 419348 79952 419404
rect 80008 419348 80078 419404
rect 79078 413048 80078 419348
rect 79078 412992 79284 413048
rect 79340 412992 79584 413048
rect 79640 412992 79884 413048
rect 79940 412992 80078 413048
rect 79078 396622 80078 412992
rect 79078 396566 79300 396622
rect 79356 396566 79600 396622
rect 79656 396566 79900 396622
rect 79956 396566 80078 396622
rect 79078 392429 80078 396566
rect 79078 392373 79200 392429
rect 79256 392373 79500 392429
rect 79556 392373 79800 392429
rect 79856 392373 80078 392429
rect 79078 392229 80078 392373
rect 79078 392173 79200 392229
rect 79256 392173 79500 392229
rect 79556 392173 79800 392229
rect 79856 392173 80078 392229
rect 79078 389622 80078 392173
rect 79078 389566 79300 389622
rect 79356 389566 79600 389622
rect 79656 389566 79900 389622
rect 79956 389566 80078 389622
rect 79078 382622 80078 389566
rect 79078 382566 79300 382622
rect 79356 382566 79600 382622
rect 79656 382566 79900 382622
rect 79956 382566 80078 382622
rect 79078 372048 80078 382566
rect 79078 371992 79284 372048
rect 79340 371992 79584 372048
rect 79640 371992 79884 372048
rect 79940 371992 80078 372048
rect 79078 356429 80078 371992
rect 79078 356373 79200 356429
rect 79256 356373 79500 356429
rect 79556 356373 79800 356429
rect 79856 356373 80078 356429
rect 79078 356229 80078 356373
rect 79078 356173 79200 356229
rect 79256 356173 79500 356229
rect 79556 356173 79800 356229
rect 79856 356173 80078 356229
rect 79078 355622 80078 356173
rect 79078 355566 79300 355622
rect 79356 355566 79600 355622
rect 79656 355566 79900 355622
rect 79956 355566 80078 355622
rect 79078 348622 80078 355566
rect 79078 348566 79300 348622
rect 79356 348566 79600 348622
rect 79656 348566 79900 348622
rect 79956 348566 80078 348622
rect 79078 341622 80078 348566
rect 79078 341566 79300 341622
rect 79356 341566 79600 341622
rect 79656 341566 79900 341622
rect 79956 341566 80078 341622
rect 79078 331040 80078 341566
rect 697922 922434 698922 939992
rect 697922 922378 698044 922434
rect 698100 922378 698344 922434
rect 698400 922378 698644 922434
rect 698700 922378 698922 922434
rect 697922 915434 698922 922378
rect 697922 915378 698044 915434
rect 698100 915378 698344 915434
rect 698400 915378 698644 915434
rect 698700 915378 698922 915434
rect 697922 908434 698922 915378
rect 697922 908378 698044 908434
rect 698100 908378 698344 908434
rect 698400 908378 698644 908434
rect 698700 908378 698922 908434
rect 697922 896429 698922 908378
rect 697922 896373 698144 896429
rect 698200 896373 698444 896429
rect 698500 896373 698744 896429
rect 698800 896373 698922 896429
rect 697922 896229 698922 896373
rect 697922 896173 698144 896229
rect 698200 896173 698444 896229
rect 698500 896173 698744 896229
rect 698800 896173 698922 896229
rect 697922 892008 698922 896173
rect 697922 891952 698060 892008
rect 698116 891952 698360 892008
rect 698416 891952 698660 892008
rect 698716 891952 698922 892008
rect 697922 860429 698922 891952
rect 697922 860373 698144 860429
rect 698200 860373 698444 860429
rect 698500 860373 698744 860429
rect 698800 860373 698922 860429
rect 697922 860229 698922 860373
rect 697922 860173 698144 860229
rect 698200 860173 698444 860229
rect 698500 860173 698744 860229
rect 698800 860173 698922 860229
rect 697922 836434 698922 860173
rect 697922 836378 698044 836434
rect 698100 836378 698344 836434
rect 698400 836378 698644 836434
rect 698700 836378 698922 836434
rect 697922 829434 698922 836378
rect 697922 829378 698044 829434
rect 698100 829378 698344 829434
rect 698400 829378 698644 829434
rect 698700 829378 698922 829434
rect 697922 824429 698922 829378
rect 697922 824373 698144 824429
rect 698200 824373 698444 824429
rect 698500 824373 698744 824429
rect 698800 824373 698922 824429
rect 697922 824229 698922 824373
rect 697922 824173 698144 824229
rect 698200 824173 698444 824229
rect 698500 824173 698744 824229
rect 698800 824173 698922 824229
rect 697922 822434 698922 824173
rect 697922 822378 698044 822434
rect 698100 822378 698344 822434
rect 698400 822378 698644 822434
rect 698700 822378 698922 822434
rect 697922 806008 698922 822378
rect 697922 805952 698060 806008
rect 698116 805952 698360 806008
rect 698416 805952 698660 806008
rect 698716 805952 698922 806008
rect 697922 752429 698922 805952
rect 697922 752373 698144 752429
rect 698200 752373 698444 752429
rect 698500 752373 698744 752429
rect 698800 752373 698922 752429
rect 697922 752229 698922 752373
rect 697922 752173 698144 752229
rect 698200 752173 698444 752229
rect 698500 752173 698744 752229
rect 698800 752173 698922 752229
rect 697922 750434 698922 752173
rect 697922 750378 698044 750434
rect 698100 750378 698344 750434
rect 698400 750378 698644 750434
rect 698700 750378 698922 750434
rect 697922 743434 698922 750378
rect 697922 743378 698044 743434
rect 698100 743378 698344 743434
rect 698400 743378 698644 743434
rect 698700 743378 698922 743434
rect 697922 736434 698922 743378
rect 697922 736378 698044 736434
rect 698100 736378 698344 736434
rect 698400 736378 698644 736434
rect 698700 736378 698922 736434
rect 697922 720008 698922 736378
rect 697922 719952 698060 720008
rect 698116 719952 698360 720008
rect 698416 719952 698660 720008
rect 698716 719952 698922 720008
rect 697922 716429 698922 719952
rect 697922 716373 698144 716429
rect 698200 716373 698444 716429
rect 698500 716373 698744 716429
rect 698800 716373 698922 716429
rect 697922 716229 698922 716373
rect 697922 716173 698144 716229
rect 698200 716173 698444 716229
rect 698500 716173 698744 716229
rect 698800 716173 698922 716229
rect 697922 707434 698922 716173
rect 697922 707378 698044 707434
rect 698100 707378 698344 707434
rect 698400 707378 698644 707434
rect 698700 707378 698922 707434
rect 697922 700434 698922 707378
rect 697922 700378 698044 700434
rect 698100 700378 698344 700434
rect 698400 700378 698644 700434
rect 698700 700378 698922 700434
rect 697922 693434 698922 700378
rect 697922 693378 698044 693434
rect 698100 693378 698344 693434
rect 698400 693378 698644 693434
rect 698700 693378 698922 693434
rect 697922 680429 698922 693378
rect 697922 680373 698144 680429
rect 698200 680373 698444 680429
rect 698500 680373 698744 680429
rect 698800 680373 698922 680429
rect 697922 680229 698922 680373
rect 697922 680173 698144 680229
rect 698200 680173 698444 680229
rect 698500 680173 698744 680229
rect 698800 680173 698922 680229
rect 697922 677008 698922 680173
rect 697922 676952 698060 677008
rect 698116 676952 698360 677008
rect 698416 676952 698660 677008
rect 698716 676952 698922 677008
rect 697922 664434 698922 676952
rect 697922 664378 698044 664434
rect 698100 664378 698344 664434
rect 698400 664378 698644 664434
rect 698700 664378 698922 664434
rect 697922 657434 698922 664378
rect 697922 657378 698044 657434
rect 698100 657378 698344 657434
rect 698400 657378 698644 657434
rect 698700 657378 698922 657434
rect 697922 650434 698922 657378
rect 697922 650378 698044 650434
rect 698100 650378 698344 650434
rect 698400 650378 698644 650434
rect 698700 650378 698922 650434
rect 697922 644429 698922 650378
rect 697922 644373 698144 644429
rect 698200 644373 698444 644429
rect 698500 644373 698744 644429
rect 698800 644373 698922 644429
rect 697922 644229 698922 644373
rect 697922 644173 698144 644229
rect 698200 644173 698444 644229
rect 698500 644173 698744 644229
rect 698800 644173 698922 644229
rect 697922 634008 698922 644173
rect 697922 633952 698060 634008
rect 698116 633952 698360 634008
rect 698416 633952 698660 634008
rect 698716 633952 698922 634008
rect 697922 621434 698922 633952
rect 697922 621378 698044 621434
rect 698100 621378 698344 621434
rect 698400 621378 698644 621434
rect 698700 621378 698922 621434
rect 697922 614434 698922 621378
rect 697922 614378 698044 614434
rect 698100 614378 698344 614434
rect 698400 614378 698644 614434
rect 698700 614378 698922 614434
rect 697922 608429 698922 614378
rect 697922 608373 698144 608429
rect 698200 608373 698444 608429
rect 698500 608373 698744 608429
rect 698800 608373 698922 608429
rect 697922 608229 698922 608373
rect 697922 608173 698144 608229
rect 698200 608173 698444 608229
rect 698500 608173 698744 608229
rect 698800 608173 698922 608229
rect 697922 607434 698922 608173
rect 697922 607378 698044 607434
rect 698100 607378 698344 607434
rect 698400 607378 698644 607434
rect 698700 607378 698922 607434
rect 697922 591008 698922 607378
rect 697922 590952 698060 591008
rect 698116 590952 698360 591008
rect 698416 590952 698660 591008
rect 698716 590952 698922 591008
rect 697922 578434 698922 590952
rect 697922 578378 698044 578434
rect 698100 578378 698344 578434
rect 698400 578378 698644 578434
rect 698700 578378 698922 578434
rect 697922 572429 698922 578378
rect 697922 572373 698144 572429
rect 698200 572373 698444 572429
rect 698500 572373 698744 572429
rect 698800 572373 698922 572429
rect 697922 572229 698922 572373
rect 697922 572173 698144 572229
rect 698200 572173 698444 572229
rect 698500 572173 698744 572229
rect 698800 572173 698922 572229
rect 697922 571434 698922 572173
rect 697922 571378 698044 571434
rect 698100 571378 698344 571434
rect 698400 571378 698644 571434
rect 698700 571378 698922 571434
rect 697922 564434 698922 571378
rect 697922 564378 698044 564434
rect 698100 564378 698344 564434
rect 698400 564378 698644 564434
rect 698700 564378 698922 564434
rect 697922 548008 698922 564378
rect 697922 547952 698060 548008
rect 698116 547952 698360 548008
rect 698416 547952 698660 548008
rect 698716 547952 698922 548008
rect 697922 536429 698922 547952
rect 697922 536373 698144 536429
rect 698200 536373 698444 536429
rect 698500 536373 698744 536429
rect 698800 536373 698922 536429
rect 697922 536229 698922 536373
rect 697922 536173 698144 536229
rect 698200 536173 698444 536229
rect 698500 536173 698744 536229
rect 698800 536173 698922 536229
rect 697922 535434 698922 536173
rect 697922 535378 698044 535434
rect 698100 535378 698344 535434
rect 698400 535378 698644 535434
rect 698700 535378 698922 535434
rect 697922 528434 698922 535378
rect 697922 528378 698044 528434
rect 698100 528378 698344 528434
rect 698400 528378 698644 528434
rect 698700 528378 698922 528434
rect 697922 521434 698922 528378
rect 697922 521378 698044 521434
rect 698100 521378 698344 521434
rect 698400 521378 698644 521434
rect 698700 521378 698922 521434
rect 697922 505008 698922 521378
rect 697922 504952 698060 505008
rect 698116 504952 698360 505008
rect 698416 504952 698660 505008
rect 698716 504952 698922 505008
rect 697922 500429 698922 504952
rect 697922 500373 698144 500429
rect 698200 500373 698444 500429
rect 698500 500373 698744 500429
rect 698800 500373 698922 500429
rect 697922 500229 698922 500373
rect 697922 500173 698144 500229
rect 698200 500173 698444 500229
rect 698500 500173 698744 500229
rect 698800 500173 698922 500229
rect 697922 464429 698922 500173
rect 697922 464373 698144 464429
rect 698200 464373 698444 464429
rect 698500 464373 698744 464429
rect 698800 464373 698922 464429
rect 697922 464229 698922 464373
rect 697922 464173 698144 464229
rect 698200 464173 698444 464229
rect 698500 464173 698744 464229
rect 698800 464173 698922 464229
rect 697922 453652 698922 464173
rect 697922 453596 697992 453652
rect 698048 453596 698116 453652
rect 698172 453596 698240 453652
rect 698296 453596 698364 453652
rect 698420 453596 698488 453652
rect 698544 453596 698612 453652
rect 698668 453596 698736 453652
rect 698792 453596 698922 453652
rect 697922 453528 698922 453596
rect 697922 453472 697992 453528
rect 698048 453472 698116 453528
rect 698172 453472 698240 453528
rect 698296 453472 698364 453528
rect 698420 453472 698488 453528
rect 698544 453472 698612 453528
rect 698668 453472 698736 453528
rect 698792 453472 698922 453528
rect 697922 453404 698922 453472
rect 697922 453348 697992 453404
rect 698048 453348 698116 453404
rect 698172 453348 698240 453404
rect 698296 453348 698364 453404
rect 698420 453348 698488 453404
rect 698544 453348 698612 453404
rect 698668 453348 698736 453404
rect 698792 453348 698922 453404
rect 697922 453280 698922 453348
rect 697922 453224 697992 453280
rect 698048 453224 698116 453280
rect 698172 453224 698240 453280
rect 698296 453224 698364 453280
rect 698420 453224 698488 453280
rect 698544 453224 698612 453280
rect 698668 453224 698736 453280
rect 698792 453224 698922 453280
rect 697922 453156 698922 453224
rect 697922 453100 697992 453156
rect 698048 453100 698116 453156
rect 698172 453100 698240 453156
rect 698296 453100 698364 453156
rect 698420 453100 698488 453156
rect 698544 453100 698612 453156
rect 698668 453100 698736 453156
rect 698792 453100 698922 453156
rect 697922 453032 698922 453100
rect 697922 452976 697992 453032
rect 698048 452976 698116 453032
rect 698172 452976 698240 453032
rect 698296 452976 698364 453032
rect 698420 452976 698488 453032
rect 698544 452976 698612 453032
rect 698668 452976 698736 453032
rect 698792 452976 698922 453032
rect 697922 452908 698922 452976
rect 697922 452852 697992 452908
rect 698048 452852 698116 452908
rect 698172 452852 698240 452908
rect 698296 452852 698364 452908
rect 698420 452852 698488 452908
rect 698544 452852 698612 452908
rect 698668 452852 698736 452908
rect 698792 452852 698922 452908
rect 697922 452784 698922 452852
rect 697922 452728 697992 452784
rect 698048 452728 698116 452784
rect 698172 452728 698240 452784
rect 698296 452728 698364 452784
rect 698420 452728 698488 452784
rect 698544 452728 698612 452784
rect 698668 452728 698736 452784
rect 698792 452728 698922 452784
rect 697922 452660 698922 452728
rect 697922 452604 697992 452660
rect 698048 452604 698116 452660
rect 698172 452604 698240 452660
rect 698296 452604 698364 452660
rect 698420 452604 698488 452660
rect 698544 452604 698612 452660
rect 698668 452604 698736 452660
rect 698792 452604 698922 452660
rect 697922 452536 698922 452604
rect 697922 452480 697992 452536
rect 698048 452480 698116 452536
rect 698172 452480 698240 452536
rect 698296 452480 698364 452536
rect 698420 452480 698488 452536
rect 698544 452480 698612 452536
rect 698668 452480 698736 452536
rect 698792 452480 698922 452536
rect 697922 452412 698922 452480
rect 697922 452356 697992 452412
rect 698048 452356 698116 452412
rect 698172 452356 698240 452412
rect 698296 452356 698364 452412
rect 698420 452356 698488 452412
rect 698544 452356 698612 452412
rect 698668 452356 698736 452412
rect 698792 452356 698922 452412
rect 697922 452288 698922 452356
rect 697922 452232 697992 452288
rect 698048 452232 698116 452288
rect 698172 452232 698240 452288
rect 698296 452232 698364 452288
rect 698420 452232 698488 452288
rect 698544 452232 698612 452288
rect 698668 452232 698736 452288
rect 698792 452232 698922 452288
rect 697922 452164 698922 452232
rect 697922 452108 697992 452164
rect 698048 452108 698116 452164
rect 698172 452108 698240 452164
rect 698296 452108 698364 452164
rect 698420 452108 698488 452164
rect 698544 452108 698612 452164
rect 698668 452108 698736 452164
rect 698792 452108 698922 452164
rect 697922 452040 698922 452108
rect 697922 451984 697992 452040
rect 698048 451984 698116 452040
rect 698172 451984 698240 452040
rect 698296 451984 698364 452040
rect 698420 451984 698488 452040
rect 698544 451984 698612 452040
rect 698668 451984 698736 452040
rect 698792 451984 698922 452040
rect 697922 451916 698922 451984
rect 697922 451860 697992 451916
rect 698048 451860 698116 451916
rect 698172 451860 698240 451916
rect 698296 451860 698364 451916
rect 698420 451860 698488 451916
rect 698544 451860 698612 451916
rect 698668 451860 698736 451916
rect 698792 451860 698922 451916
rect 697922 451172 698922 451860
rect 697922 451116 697992 451172
rect 698048 451116 698116 451172
rect 698172 451116 698240 451172
rect 698296 451116 698364 451172
rect 698420 451116 698488 451172
rect 698544 451116 698612 451172
rect 698668 451116 698736 451172
rect 698792 451116 698922 451172
rect 697922 451048 698922 451116
rect 697922 450992 697992 451048
rect 698048 450992 698116 451048
rect 698172 450992 698240 451048
rect 698296 450992 698364 451048
rect 698420 450992 698488 451048
rect 698544 450992 698612 451048
rect 698668 450992 698736 451048
rect 698792 450992 698922 451048
rect 697922 450924 698922 450992
rect 697922 450868 697992 450924
rect 698048 450868 698116 450924
rect 698172 450868 698240 450924
rect 698296 450868 698364 450924
rect 698420 450868 698488 450924
rect 698544 450868 698612 450924
rect 698668 450868 698736 450924
rect 698792 450868 698922 450924
rect 697922 450800 698922 450868
rect 697922 450744 697992 450800
rect 698048 450744 698116 450800
rect 698172 450744 698240 450800
rect 698296 450744 698364 450800
rect 698420 450744 698488 450800
rect 698544 450744 698612 450800
rect 698668 450744 698736 450800
rect 698792 450744 698922 450800
rect 697922 450676 698922 450744
rect 697922 450620 697992 450676
rect 698048 450620 698116 450676
rect 698172 450620 698240 450676
rect 698296 450620 698364 450676
rect 698420 450620 698488 450676
rect 698544 450620 698612 450676
rect 698668 450620 698736 450676
rect 698792 450620 698922 450676
rect 697922 450552 698922 450620
rect 697922 450496 697992 450552
rect 698048 450496 698116 450552
rect 698172 450496 698240 450552
rect 698296 450496 698364 450552
rect 698420 450496 698488 450552
rect 698544 450496 698612 450552
rect 698668 450496 698736 450552
rect 698792 450496 698922 450552
rect 697922 450428 698922 450496
rect 697922 450372 697992 450428
rect 698048 450372 698116 450428
rect 698172 450372 698240 450428
rect 698296 450372 698364 450428
rect 698420 450372 698488 450428
rect 698544 450372 698612 450428
rect 698668 450372 698736 450428
rect 698792 450372 698922 450428
rect 697922 450304 698922 450372
rect 697922 450248 697992 450304
rect 698048 450248 698116 450304
rect 698172 450248 698240 450304
rect 698296 450248 698364 450304
rect 698420 450248 698488 450304
rect 698544 450248 698612 450304
rect 698668 450248 698736 450304
rect 698792 450248 698922 450304
rect 697922 450180 698922 450248
rect 697922 450124 697992 450180
rect 698048 450124 698116 450180
rect 698172 450124 698240 450180
rect 698296 450124 698364 450180
rect 698420 450124 698488 450180
rect 698544 450124 698612 450180
rect 698668 450124 698736 450180
rect 698792 450124 698922 450180
rect 697922 450056 698922 450124
rect 697922 450000 697992 450056
rect 698048 450000 698116 450056
rect 698172 450000 698240 450056
rect 698296 450000 698364 450056
rect 698420 450000 698488 450056
rect 698544 450000 698612 450056
rect 698668 450000 698736 450056
rect 698792 450000 698922 450056
rect 697922 449932 698922 450000
rect 697922 449876 697992 449932
rect 698048 449876 698116 449932
rect 698172 449876 698240 449932
rect 698296 449876 698364 449932
rect 698420 449876 698488 449932
rect 698544 449876 698612 449932
rect 698668 449876 698736 449932
rect 698792 449876 698922 449932
rect 697922 449808 698922 449876
rect 697922 449752 697992 449808
rect 698048 449752 698116 449808
rect 698172 449752 698240 449808
rect 698296 449752 698364 449808
rect 698420 449752 698488 449808
rect 698544 449752 698612 449808
rect 698668 449752 698736 449808
rect 698792 449752 698922 449808
rect 697922 449684 698922 449752
rect 697922 449628 697992 449684
rect 698048 449628 698116 449684
rect 698172 449628 698240 449684
rect 698296 449628 698364 449684
rect 698420 449628 698488 449684
rect 698544 449628 698612 449684
rect 698668 449628 698736 449684
rect 698792 449628 698922 449684
rect 697922 449560 698922 449628
rect 697922 449504 697992 449560
rect 698048 449504 698116 449560
rect 698172 449504 698240 449560
rect 698296 449504 698364 449560
rect 698420 449504 698488 449560
rect 698544 449504 698612 449560
rect 698668 449504 698736 449560
rect 698792 449504 698922 449560
rect 697922 449436 698922 449504
rect 697922 449380 697992 449436
rect 698048 449380 698116 449436
rect 698172 449380 698240 449436
rect 698296 449380 698364 449436
rect 698420 449380 698488 449436
rect 698544 449380 698612 449436
rect 698668 449380 698736 449436
rect 698792 449380 698922 449436
rect 697922 449312 698922 449380
rect 697922 449256 697992 449312
rect 698048 449256 698116 449312
rect 698172 449256 698240 449312
rect 698296 449256 698364 449312
rect 698420 449256 698488 449312
rect 698544 449256 698612 449312
rect 698668 449256 698736 449312
rect 698792 449256 698922 449312
rect 697922 448802 698922 449256
rect 697922 448746 697992 448802
rect 698048 448746 698116 448802
rect 698172 448746 698240 448802
rect 698296 448746 698364 448802
rect 698420 448746 698488 448802
rect 698544 448746 698612 448802
rect 698668 448746 698736 448802
rect 698792 448746 698922 448802
rect 697922 448678 698922 448746
rect 697922 448622 697992 448678
rect 698048 448622 698116 448678
rect 698172 448622 698240 448678
rect 698296 448622 698364 448678
rect 698420 448622 698488 448678
rect 698544 448622 698612 448678
rect 698668 448622 698736 448678
rect 698792 448622 698922 448678
rect 697922 448554 698922 448622
rect 697922 448498 697992 448554
rect 698048 448498 698116 448554
rect 698172 448498 698240 448554
rect 698296 448498 698364 448554
rect 698420 448498 698488 448554
rect 698544 448498 698612 448554
rect 698668 448498 698736 448554
rect 698792 448498 698922 448554
rect 697922 448430 698922 448498
rect 697922 448374 697992 448430
rect 698048 448374 698116 448430
rect 698172 448374 698240 448430
rect 698296 448374 698364 448430
rect 698420 448374 698488 448430
rect 698544 448374 698612 448430
rect 698668 448374 698736 448430
rect 698792 448374 698922 448430
rect 697922 448306 698922 448374
rect 697922 448250 697992 448306
rect 698048 448250 698116 448306
rect 698172 448250 698240 448306
rect 698296 448250 698364 448306
rect 698420 448250 698488 448306
rect 698544 448250 698612 448306
rect 698668 448250 698736 448306
rect 698792 448250 698922 448306
rect 697922 448182 698922 448250
rect 697922 448126 697992 448182
rect 698048 448126 698116 448182
rect 698172 448126 698240 448182
rect 698296 448126 698364 448182
rect 698420 448126 698488 448182
rect 698544 448126 698612 448182
rect 698668 448126 698736 448182
rect 698792 448126 698922 448182
rect 697922 448058 698922 448126
rect 697922 448002 697992 448058
rect 698048 448002 698116 448058
rect 698172 448002 698240 448058
rect 698296 448002 698364 448058
rect 698420 448002 698488 448058
rect 698544 448002 698612 448058
rect 698668 448002 698736 448058
rect 698792 448002 698922 448058
rect 697922 447934 698922 448002
rect 697922 447878 697992 447934
rect 698048 447878 698116 447934
rect 698172 447878 698240 447934
rect 698296 447878 698364 447934
rect 698420 447878 698488 447934
rect 698544 447878 698612 447934
rect 698668 447878 698736 447934
rect 698792 447878 698922 447934
rect 697922 447810 698922 447878
rect 697922 447754 697992 447810
rect 698048 447754 698116 447810
rect 698172 447754 698240 447810
rect 698296 447754 698364 447810
rect 698420 447754 698488 447810
rect 698544 447754 698612 447810
rect 698668 447754 698736 447810
rect 698792 447754 698922 447810
rect 697922 447686 698922 447754
rect 697922 447630 697992 447686
rect 698048 447630 698116 447686
rect 698172 447630 698240 447686
rect 698296 447630 698364 447686
rect 698420 447630 698488 447686
rect 698544 447630 698612 447686
rect 698668 447630 698736 447686
rect 698792 447630 698922 447686
rect 697922 447562 698922 447630
rect 697922 447506 697992 447562
rect 698048 447506 698116 447562
rect 698172 447506 698240 447562
rect 698296 447506 698364 447562
rect 698420 447506 698488 447562
rect 698544 447506 698612 447562
rect 698668 447506 698736 447562
rect 698792 447506 698922 447562
rect 697922 447438 698922 447506
rect 697922 447382 697992 447438
rect 698048 447382 698116 447438
rect 698172 447382 698240 447438
rect 698296 447382 698364 447438
rect 698420 447382 698488 447438
rect 698544 447382 698612 447438
rect 698668 447382 698736 447438
rect 698792 447382 698922 447438
rect 697922 447314 698922 447382
rect 697922 447258 697992 447314
rect 698048 447258 698116 447314
rect 698172 447258 698240 447314
rect 698296 447258 698364 447314
rect 698420 447258 698488 447314
rect 698544 447258 698612 447314
rect 698668 447258 698736 447314
rect 698792 447258 698922 447314
rect 697922 447190 698922 447258
rect 697922 447134 697992 447190
rect 698048 447134 698116 447190
rect 698172 447134 698240 447190
rect 698296 447134 698364 447190
rect 698420 447134 698488 447190
rect 698544 447134 698612 447190
rect 698668 447134 698736 447190
rect 698792 447134 698922 447190
rect 697922 447066 698922 447134
rect 697922 447010 697992 447066
rect 698048 447010 698116 447066
rect 698172 447010 698240 447066
rect 698296 447010 698364 447066
rect 698420 447010 698488 447066
rect 698544 447010 698612 447066
rect 698668 447010 698736 447066
rect 698792 447010 698922 447066
rect 697922 446942 698922 447010
rect 697922 446886 697992 446942
rect 698048 446886 698116 446942
rect 698172 446886 698240 446942
rect 698296 446886 698364 446942
rect 698420 446886 698488 446942
rect 698544 446886 698612 446942
rect 698668 446886 698736 446942
rect 698792 446886 698922 446942
rect 697922 446096 698922 446886
rect 697922 446040 697992 446096
rect 698048 446040 698116 446096
rect 698172 446040 698240 446096
rect 698296 446040 698364 446096
rect 698420 446040 698488 446096
rect 698544 446040 698612 446096
rect 698668 446040 698736 446096
rect 698792 446040 698922 446096
rect 697922 445972 698922 446040
rect 697922 445916 697992 445972
rect 698048 445916 698116 445972
rect 698172 445916 698240 445972
rect 698296 445916 698364 445972
rect 698420 445916 698488 445972
rect 698544 445916 698612 445972
rect 698668 445916 698736 445972
rect 698792 445916 698922 445972
rect 697922 445848 698922 445916
rect 697922 445792 697992 445848
rect 698048 445792 698116 445848
rect 698172 445792 698240 445848
rect 698296 445792 698364 445848
rect 698420 445792 698488 445848
rect 698544 445792 698612 445848
rect 698668 445792 698736 445848
rect 698792 445792 698922 445848
rect 697922 445724 698922 445792
rect 697922 445668 697992 445724
rect 698048 445668 698116 445724
rect 698172 445668 698240 445724
rect 698296 445668 698364 445724
rect 698420 445668 698488 445724
rect 698544 445668 698612 445724
rect 698668 445668 698736 445724
rect 698792 445668 698922 445724
rect 697922 445600 698922 445668
rect 697922 445544 697992 445600
rect 698048 445544 698116 445600
rect 698172 445544 698240 445600
rect 698296 445544 698364 445600
rect 698420 445544 698488 445600
rect 698544 445544 698612 445600
rect 698668 445544 698736 445600
rect 698792 445544 698922 445600
rect 697922 445476 698922 445544
rect 697922 445420 697992 445476
rect 698048 445420 698116 445476
rect 698172 445420 698240 445476
rect 698296 445420 698364 445476
rect 698420 445420 698488 445476
rect 698544 445420 698612 445476
rect 698668 445420 698736 445476
rect 698792 445420 698922 445476
rect 697922 445352 698922 445420
rect 697922 445296 697992 445352
rect 698048 445296 698116 445352
rect 698172 445296 698240 445352
rect 698296 445296 698364 445352
rect 698420 445296 698488 445352
rect 698544 445296 698612 445352
rect 698668 445296 698736 445352
rect 698792 445296 698922 445352
rect 697922 445228 698922 445296
rect 697922 445172 697992 445228
rect 698048 445172 698116 445228
rect 698172 445172 698240 445228
rect 698296 445172 698364 445228
rect 698420 445172 698488 445228
rect 698544 445172 698612 445228
rect 698668 445172 698736 445228
rect 698792 445172 698922 445228
rect 697922 445104 698922 445172
rect 697922 445048 697992 445104
rect 698048 445048 698116 445104
rect 698172 445048 698240 445104
rect 698296 445048 698364 445104
rect 698420 445048 698488 445104
rect 698544 445048 698612 445104
rect 698668 445048 698736 445104
rect 698792 445048 698922 445104
rect 697922 444980 698922 445048
rect 697922 444924 697992 444980
rect 698048 444924 698116 444980
rect 698172 444924 698240 444980
rect 698296 444924 698364 444980
rect 698420 444924 698488 444980
rect 698544 444924 698612 444980
rect 698668 444924 698736 444980
rect 698792 444924 698922 444980
rect 697922 444856 698922 444924
rect 697922 444800 697992 444856
rect 698048 444800 698116 444856
rect 698172 444800 698240 444856
rect 698296 444800 698364 444856
rect 698420 444800 698488 444856
rect 698544 444800 698612 444856
rect 698668 444800 698736 444856
rect 698792 444800 698922 444856
rect 697922 444732 698922 444800
rect 697922 444676 697992 444732
rect 698048 444676 698116 444732
rect 698172 444676 698240 444732
rect 698296 444676 698364 444732
rect 698420 444676 698488 444732
rect 698544 444676 698612 444732
rect 698668 444676 698736 444732
rect 698792 444676 698922 444732
rect 697922 444608 698922 444676
rect 697922 444552 697992 444608
rect 698048 444552 698116 444608
rect 698172 444552 698240 444608
rect 698296 444552 698364 444608
rect 698420 444552 698488 444608
rect 698544 444552 698612 444608
rect 698668 444552 698736 444608
rect 698792 444552 698922 444608
rect 697922 444484 698922 444552
rect 697922 444428 697992 444484
rect 698048 444428 698116 444484
rect 698172 444428 698240 444484
rect 698296 444428 698364 444484
rect 698420 444428 698488 444484
rect 698544 444428 698612 444484
rect 698668 444428 698736 444484
rect 698792 444428 698922 444484
rect 697922 444360 698922 444428
rect 697922 444304 697992 444360
rect 698048 444304 698116 444360
rect 698172 444304 698240 444360
rect 698296 444304 698364 444360
rect 698420 444304 698488 444360
rect 698544 444304 698612 444360
rect 698668 444304 698736 444360
rect 698792 444304 698922 444360
rect 697922 444236 698922 444304
rect 697922 444180 697992 444236
rect 698048 444180 698116 444236
rect 698172 444180 698240 444236
rect 698296 444180 698364 444236
rect 698420 444180 698488 444236
rect 698544 444180 698612 444236
rect 698668 444180 698736 444236
rect 698792 444180 698922 444236
rect 697922 443726 698922 444180
rect 697922 443670 697992 443726
rect 698048 443670 698116 443726
rect 698172 443670 698240 443726
rect 698296 443670 698364 443726
rect 698420 443670 698488 443726
rect 698544 443670 698612 443726
rect 698668 443670 698736 443726
rect 698792 443670 698922 443726
rect 697922 443602 698922 443670
rect 697922 443546 697992 443602
rect 698048 443546 698116 443602
rect 698172 443546 698240 443602
rect 698296 443546 698364 443602
rect 698420 443546 698488 443602
rect 698544 443546 698612 443602
rect 698668 443546 698736 443602
rect 698792 443546 698922 443602
rect 697922 443478 698922 443546
rect 697922 443422 697992 443478
rect 698048 443422 698116 443478
rect 698172 443422 698240 443478
rect 698296 443422 698364 443478
rect 698420 443422 698488 443478
rect 698544 443422 698612 443478
rect 698668 443422 698736 443478
rect 698792 443422 698922 443478
rect 697922 443354 698922 443422
rect 697922 443298 697992 443354
rect 698048 443298 698116 443354
rect 698172 443298 698240 443354
rect 698296 443298 698364 443354
rect 698420 443298 698488 443354
rect 698544 443298 698612 443354
rect 698668 443298 698736 443354
rect 698792 443298 698922 443354
rect 697922 443230 698922 443298
rect 697922 443174 697992 443230
rect 698048 443174 698116 443230
rect 698172 443174 698240 443230
rect 698296 443174 698364 443230
rect 698420 443174 698488 443230
rect 698544 443174 698612 443230
rect 698668 443174 698736 443230
rect 698792 443174 698922 443230
rect 697922 443106 698922 443174
rect 697922 443050 697992 443106
rect 698048 443050 698116 443106
rect 698172 443050 698240 443106
rect 698296 443050 698364 443106
rect 698420 443050 698488 443106
rect 698544 443050 698612 443106
rect 698668 443050 698736 443106
rect 698792 443050 698922 443106
rect 697922 442982 698922 443050
rect 697922 442926 697992 442982
rect 698048 442926 698116 442982
rect 698172 442926 698240 442982
rect 698296 442926 698364 442982
rect 698420 442926 698488 442982
rect 698544 442926 698612 442982
rect 698668 442926 698736 442982
rect 698792 442926 698922 442982
rect 697922 442858 698922 442926
rect 697922 442802 697992 442858
rect 698048 442802 698116 442858
rect 698172 442802 698240 442858
rect 698296 442802 698364 442858
rect 698420 442802 698488 442858
rect 698544 442802 698612 442858
rect 698668 442802 698736 442858
rect 698792 442802 698922 442858
rect 697922 442734 698922 442802
rect 697922 442678 697992 442734
rect 698048 442678 698116 442734
rect 698172 442678 698240 442734
rect 698296 442678 698364 442734
rect 698420 442678 698488 442734
rect 698544 442678 698612 442734
rect 698668 442678 698736 442734
rect 698792 442678 698922 442734
rect 697922 442610 698922 442678
rect 697922 442554 697992 442610
rect 698048 442554 698116 442610
rect 698172 442554 698240 442610
rect 698296 442554 698364 442610
rect 698420 442554 698488 442610
rect 698544 442554 698612 442610
rect 698668 442554 698736 442610
rect 698792 442554 698922 442610
rect 697922 442486 698922 442554
rect 697922 442430 697992 442486
rect 698048 442430 698116 442486
rect 698172 442430 698240 442486
rect 698296 442430 698364 442486
rect 698420 442430 698488 442486
rect 698544 442430 698612 442486
rect 698668 442430 698736 442486
rect 698792 442430 698922 442486
rect 697922 442362 698922 442430
rect 697922 442306 697992 442362
rect 698048 442306 698116 442362
rect 698172 442306 698240 442362
rect 698296 442306 698364 442362
rect 698420 442306 698488 442362
rect 698544 442306 698612 442362
rect 698668 442306 698736 442362
rect 698792 442306 698922 442362
rect 697922 442238 698922 442306
rect 697922 442182 697992 442238
rect 698048 442182 698116 442238
rect 698172 442182 698240 442238
rect 698296 442182 698364 442238
rect 698420 442182 698488 442238
rect 698544 442182 698612 442238
rect 698668 442182 698736 442238
rect 698792 442182 698922 442238
rect 697922 442114 698922 442182
rect 697922 442058 697992 442114
rect 698048 442058 698116 442114
rect 698172 442058 698240 442114
rect 698296 442058 698364 442114
rect 698420 442058 698488 442114
rect 698544 442058 698612 442114
rect 698668 442058 698736 442114
rect 698792 442058 698922 442114
rect 697922 441990 698922 442058
rect 697922 441934 697992 441990
rect 698048 441934 698116 441990
rect 698172 441934 698240 441990
rect 698296 441934 698364 441990
rect 698420 441934 698488 441990
rect 698544 441934 698612 441990
rect 698668 441934 698736 441990
rect 698792 441934 698922 441990
rect 697922 441866 698922 441934
rect 697922 441810 697992 441866
rect 698048 441810 698116 441866
rect 698172 441810 698240 441866
rect 698296 441810 698364 441866
rect 698420 441810 698488 441866
rect 698544 441810 698612 441866
rect 698668 441810 698736 441866
rect 698792 441810 698922 441866
rect 697922 441122 698922 441810
rect 697922 441066 697992 441122
rect 698048 441066 698116 441122
rect 698172 441066 698240 441122
rect 698296 441066 698364 441122
rect 698420 441066 698488 441122
rect 698544 441066 698612 441122
rect 698668 441066 698736 441122
rect 698792 441066 698922 441122
rect 697922 440998 698922 441066
rect 697922 440942 697992 440998
rect 698048 440942 698116 440998
rect 698172 440942 698240 440998
rect 698296 440942 698364 440998
rect 698420 440942 698488 440998
rect 698544 440942 698612 440998
rect 698668 440942 698736 440998
rect 698792 440942 698922 440998
rect 697922 440874 698922 440942
rect 697922 440818 697992 440874
rect 698048 440818 698116 440874
rect 698172 440818 698240 440874
rect 698296 440818 698364 440874
rect 698420 440818 698488 440874
rect 698544 440818 698612 440874
rect 698668 440818 698736 440874
rect 698792 440818 698922 440874
rect 697922 440750 698922 440818
rect 697922 440694 697992 440750
rect 698048 440694 698116 440750
rect 698172 440694 698240 440750
rect 698296 440694 698364 440750
rect 698420 440694 698488 440750
rect 698544 440694 698612 440750
rect 698668 440694 698736 440750
rect 698792 440694 698922 440750
rect 697922 440626 698922 440694
rect 697922 440570 697992 440626
rect 698048 440570 698116 440626
rect 698172 440570 698240 440626
rect 698296 440570 698364 440626
rect 698420 440570 698488 440626
rect 698544 440570 698612 440626
rect 698668 440570 698736 440626
rect 698792 440570 698922 440626
rect 697922 440502 698922 440570
rect 697922 440446 697992 440502
rect 698048 440446 698116 440502
rect 698172 440446 698240 440502
rect 698296 440446 698364 440502
rect 698420 440446 698488 440502
rect 698544 440446 698612 440502
rect 698668 440446 698736 440502
rect 698792 440446 698922 440502
rect 697922 440378 698922 440446
rect 697922 440322 697992 440378
rect 698048 440322 698116 440378
rect 698172 440322 698240 440378
rect 698296 440322 698364 440378
rect 698420 440322 698488 440378
rect 698544 440322 698612 440378
rect 698668 440322 698736 440378
rect 698792 440322 698922 440378
rect 697922 440254 698922 440322
rect 697922 440198 697992 440254
rect 698048 440198 698116 440254
rect 698172 440198 698240 440254
rect 698296 440198 698364 440254
rect 698420 440198 698488 440254
rect 698544 440198 698612 440254
rect 698668 440198 698736 440254
rect 698792 440198 698922 440254
rect 697922 440130 698922 440198
rect 697922 440074 697992 440130
rect 698048 440074 698116 440130
rect 698172 440074 698240 440130
rect 698296 440074 698364 440130
rect 698420 440074 698488 440130
rect 698544 440074 698612 440130
rect 698668 440074 698736 440130
rect 698792 440074 698922 440130
rect 697922 440006 698922 440074
rect 697922 439950 697992 440006
rect 698048 439950 698116 440006
rect 698172 439950 698240 440006
rect 698296 439950 698364 440006
rect 698420 439950 698488 440006
rect 698544 439950 698612 440006
rect 698668 439950 698736 440006
rect 698792 439950 698922 440006
rect 697922 439882 698922 439950
rect 697922 439826 697992 439882
rect 698048 439826 698116 439882
rect 698172 439826 698240 439882
rect 698296 439826 698364 439882
rect 698420 439826 698488 439882
rect 698544 439826 698612 439882
rect 698668 439826 698736 439882
rect 698792 439826 698922 439882
rect 697922 439758 698922 439826
rect 697922 439702 697992 439758
rect 698048 439702 698116 439758
rect 698172 439702 698240 439758
rect 698296 439702 698364 439758
rect 698420 439702 698488 439758
rect 698544 439702 698612 439758
rect 698668 439702 698736 439758
rect 698792 439702 698922 439758
rect 697922 439634 698922 439702
rect 697922 439578 697992 439634
rect 698048 439578 698116 439634
rect 698172 439578 698240 439634
rect 698296 439578 698364 439634
rect 698420 439578 698488 439634
rect 698544 439578 698612 439634
rect 698668 439578 698736 439634
rect 698792 439578 698922 439634
rect 697922 439510 698922 439578
rect 697922 439454 697992 439510
rect 698048 439454 698116 439510
rect 698172 439454 698240 439510
rect 698296 439454 698364 439510
rect 698420 439454 698488 439510
rect 698544 439454 698612 439510
rect 698668 439454 698736 439510
rect 698792 439454 698922 439510
rect 697922 439386 698922 439454
rect 697922 439330 697992 439386
rect 698048 439330 698116 439386
rect 698172 439330 698240 439386
rect 698296 439330 698364 439386
rect 698420 439330 698488 439386
rect 698544 439330 698612 439386
rect 698668 439330 698736 439386
rect 698792 439330 698922 439386
rect 697922 428429 698922 439330
rect 697922 428373 698144 428429
rect 698200 428373 698444 428429
rect 698500 428373 698744 428429
rect 698800 428373 698922 428429
rect 697922 428229 698922 428373
rect 697922 428173 698144 428229
rect 698200 428173 698444 428229
rect 698500 428173 698744 428229
rect 698800 428173 698922 428229
rect 697922 410652 698922 428173
rect 697922 410596 697992 410652
rect 698048 410596 698116 410652
rect 698172 410596 698240 410652
rect 698296 410596 698364 410652
rect 698420 410596 698488 410652
rect 698544 410596 698612 410652
rect 698668 410596 698736 410652
rect 698792 410596 698922 410652
rect 697922 410528 698922 410596
rect 697922 410472 697992 410528
rect 698048 410472 698116 410528
rect 698172 410472 698240 410528
rect 698296 410472 698364 410528
rect 698420 410472 698488 410528
rect 698544 410472 698612 410528
rect 698668 410472 698736 410528
rect 698792 410472 698922 410528
rect 697922 410404 698922 410472
rect 697922 410348 697992 410404
rect 698048 410348 698116 410404
rect 698172 410348 698240 410404
rect 698296 410348 698364 410404
rect 698420 410348 698488 410404
rect 698544 410348 698612 410404
rect 698668 410348 698736 410404
rect 698792 410348 698922 410404
rect 697922 410280 698922 410348
rect 697922 410224 697992 410280
rect 698048 410224 698116 410280
rect 698172 410224 698240 410280
rect 698296 410224 698364 410280
rect 698420 410224 698488 410280
rect 698544 410224 698612 410280
rect 698668 410224 698736 410280
rect 698792 410224 698922 410280
rect 697922 410156 698922 410224
rect 697922 410100 697992 410156
rect 698048 410100 698116 410156
rect 698172 410100 698240 410156
rect 698296 410100 698364 410156
rect 698420 410100 698488 410156
rect 698544 410100 698612 410156
rect 698668 410100 698736 410156
rect 698792 410100 698922 410156
rect 697922 410032 698922 410100
rect 697922 409976 697992 410032
rect 698048 409976 698116 410032
rect 698172 409976 698240 410032
rect 698296 409976 698364 410032
rect 698420 409976 698488 410032
rect 698544 409976 698612 410032
rect 698668 409976 698736 410032
rect 698792 409976 698922 410032
rect 697922 409908 698922 409976
rect 697922 409852 697992 409908
rect 698048 409852 698116 409908
rect 698172 409852 698240 409908
rect 698296 409852 698364 409908
rect 698420 409852 698488 409908
rect 698544 409852 698612 409908
rect 698668 409852 698736 409908
rect 698792 409852 698922 409908
rect 697922 409784 698922 409852
rect 697922 409728 697992 409784
rect 698048 409728 698116 409784
rect 698172 409728 698240 409784
rect 698296 409728 698364 409784
rect 698420 409728 698488 409784
rect 698544 409728 698612 409784
rect 698668 409728 698736 409784
rect 698792 409728 698922 409784
rect 697922 409660 698922 409728
rect 697922 409604 697992 409660
rect 698048 409604 698116 409660
rect 698172 409604 698240 409660
rect 698296 409604 698364 409660
rect 698420 409604 698488 409660
rect 698544 409604 698612 409660
rect 698668 409604 698736 409660
rect 698792 409604 698922 409660
rect 697922 409536 698922 409604
rect 697922 409480 697992 409536
rect 698048 409480 698116 409536
rect 698172 409480 698240 409536
rect 698296 409480 698364 409536
rect 698420 409480 698488 409536
rect 698544 409480 698612 409536
rect 698668 409480 698736 409536
rect 698792 409480 698922 409536
rect 697922 409412 698922 409480
rect 697922 409356 697992 409412
rect 698048 409356 698116 409412
rect 698172 409356 698240 409412
rect 698296 409356 698364 409412
rect 698420 409356 698488 409412
rect 698544 409356 698612 409412
rect 698668 409356 698736 409412
rect 698792 409356 698922 409412
rect 697922 409288 698922 409356
rect 697922 409232 697992 409288
rect 698048 409232 698116 409288
rect 698172 409232 698240 409288
rect 698296 409232 698364 409288
rect 698420 409232 698488 409288
rect 698544 409232 698612 409288
rect 698668 409232 698736 409288
rect 698792 409232 698922 409288
rect 697922 409164 698922 409232
rect 697922 409108 697992 409164
rect 698048 409108 698116 409164
rect 698172 409108 698240 409164
rect 698296 409108 698364 409164
rect 698420 409108 698488 409164
rect 698544 409108 698612 409164
rect 698668 409108 698736 409164
rect 698792 409108 698922 409164
rect 697922 409040 698922 409108
rect 697922 408984 697992 409040
rect 698048 408984 698116 409040
rect 698172 408984 698240 409040
rect 698296 408984 698364 409040
rect 698420 408984 698488 409040
rect 698544 408984 698612 409040
rect 698668 408984 698736 409040
rect 698792 408984 698922 409040
rect 697922 408916 698922 408984
rect 697922 408860 697992 408916
rect 698048 408860 698116 408916
rect 698172 408860 698240 408916
rect 698296 408860 698364 408916
rect 698420 408860 698488 408916
rect 698544 408860 698612 408916
rect 698668 408860 698736 408916
rect 698792 408860 698922 408916
rect 697922 408172 698922 408860
rect 697922 408116 697992 408172
rect 698048 408116 698116 408172
rect 698172 408116 698240 408172
rect 698296 408116 698364 408172
rect 698420 408116 698488 408172
rect 698544 408116 698612 408172
rect 698668 408116 698736 408172
rect 698792 408116 698922 408172
rect 697922 408048 698922 408116
rect 697922 407992 697992 408048
rect 698048 407992 698116 408048
rect 698172 407992 698240 408048
rect 698296 407992 698364 408048
rect 698420 407992 698488 408048
rect 698544 407992 698612 408048
rect 698668 407992 698736 408048
rect 698792 407992 698922 408048
rect 697922 407924 698922 407992
rect 697922 407868 697992 407924
rect 698048 407868 698116 407924
rect 698172 407868 698240 407924
rect 698296 407868 698364 407924
rect 698420 407868 698488 407924
rect 698544 407868 698612 407924
rect 698668 407868 698736 407924
rect 698792 407868 698922 407924
rect 697922 407800 698922 407868
rect 697922 407744 697992 407800
rect 698048 407744 698116 407800
rect 698172 407744 698240 407800
rect 698296 407744 698364 407800
rect 698420 407744 698488 407800
rect 698544 407744 698612 407800
rect 698668 407744 698736 407800
rect 698792 407744 698922 407800
rect 697922 407676 698922 407744
rect 697922 407620 697992 407676
rect 698048 407620 698116 407676
rect 698172 407620 698240 407676
rect 698296 407620 698364 407676
rect 698420 407620 698488 407676
rect 698544 407620 698612 407676
rect 698668 407620 698736 407676
rect 698792 407620 698922 407676
rect 697922 407552 698922 407620
rect 697922 407496 697992 407552
rect 698048 407496 698116 407552
rect 698172 407496 698240 407552
rect 698296 407496 698364 407552
rect 698420 407496 698488 407552
rect 698544 407496 698612 407552
rect 698668 407496 698736 407552
rect 698792 407496 698922 407552
rect 697922 407428 698922 407496
rect 697922 407372 697992 407428
rect 698048 407372 698116 407428
rect 698172 407372 698240 407428
rect 698296 407372 698364 407428
rect 698420 407372 698488 407428
rect 698544 407372 698612 407428
rect 698668 407372 698736 407428
rect 698792 407372 698922 407428
rect 697922 407304 698922 407372
rect 697922 407248 697992 407304
rect 698048 407248 698116 407304
rect 698172 407248 698240 407304
rect 698296 407248 698364 407304
rect 698420 407248 698488 407304
rect 698544 407248 698612 407304
rect 698668 407248 698736 407304
rect 698792 407248 698922 407304
rect 697922 407180 698922 407248
rect 697922 407124 697992 407180
rect 698048 407124 698116 407180
rect 698172 407124 698240 407180
rect 698296 407124 698364 407180
rect 698420 407124 698488 407180
rect 698544 407124 698612 407180
rect 698668 407124 698736 407180
rect 698792 407124 698922 407180
rect 697922 407056 698922 407124
rect 697922 407000 697992 407056
rect 698048 407000 698116 407056
rect 698172 407000 698240 407056
rect 698296 407000 698364 407056
rect 698420 407000 698488 407056
rect 698544 407000 698612 407056
rect 698668 407000 698736 407056
rect 698792 407000 698922 407056
rect 697922 406932 698922 407000
rect 697922 406876 697992 406932
rect 698048 406876 698116 406932
rect 698172 406876 698240 406932
rect 698296 406876 698364 406932
rect 698420 406876 698488 406932
rect 698544 406876 698612 406932
rect 698668 406876 698736 406932
rect 698792 406876 698922 406932
rect 697922 406808 698922 406876
rect 697922 406752 697992 406808
rect 698048 406752 698116 406808
rect 698172 406752 698240 406808
rect 698296 406752 698364 406808
rect 698420 406752 698488 406808
rect 698544 406752 698612 406808
rect 698668 406752 698736 406808
rect 698792 406752 698922 406808
rect 697922 406684 698922 406752
rect 697922 406628 697992 406684
rect 698048 406628 698116 406684
rect 698172 406628 698240 406684
rect 698296 406628 698364 406684
rect 698420 406628 698488 406684
rect 698544 406628 698612 406684
rect 698668 406628 698736 406684
rect 698792 406628 698922 406684
rect 697922 406560 698922 406628
rect 697922 406504 697992 406560
rect 698048 406504 698116 406560
rect 698172 406504 698240 406560
rect 698296 406504 698364 406560
rect 698420 406504 698488 406560
rect 698544 406504 698612 406560
rect 698668 406504 698736 406560
rect 698792 406504 698922 406560
rect 697922 406436 698922 406504
rect 697922 406380 697992 406436
rect 698048 406380 698116 406436
rect 698172 406380 698240 406436
rect 698296 406380 698364 406436
rect 698420 406380 698488 406436
rect 698544 406380 698612 406436
rect 698668 406380 698736 406436
rect 698792 406380 698922 406436
rect 697922 406312 698922 406380
rect 697922 406256 697992 406312
rect 698048 406256 698116 406312
rect 698172 406256 698240 406312
rect 698296 406256 698364 406312
rect 698420 406256 698488 406312
rect 698544 406256 698612 406312
rect 698668 406256 698736 406312
rect 698792 406256 698922 406312
rect 697922 405802 698922 406256
rect 697922 405746 697992 405802
rect 698048 405746 698116 405802
rect 698172 405746 698240 405802
rect 698296 405746 698364 405802
rect 698420 405746 698488 405802
rect 698544 405746 698612 405802
rect 698668 405746 698736 405802
rect 698792 405746 698922 405802
rect 697922 405678 698922 405746
rect 697922 405622 697992 405678
rect 698048 405622 698116 405678
rect 698172 405622 698240 405678
rect 698296 405622 698364 405678
rect 698420 405622 698488 405678
rect 698544 405622 698612 405678
rect 698668 405622 698736 405678
rect 698792 405622 698922 405678
rect 697922 405554 698922 405622
rect 697922 405498 697992 405554
rect 698048 405498 698116 405554
rect 698172 405498 698240 405554
rect 698296 405498 698364 405554
rect 698420 405498 698488 405554
rect 698544 405498 698612 405554
rect 698668 405498 698736 405554
rect 698792 405498 698922 405554
rect 697922 405430 698922 405498
rect 697922 405374 697992 405430
rect 698048 405374 698116 405430
rect 698172 405374 698240 405430
rect 698296 405374 698364 405430
rect 698420 405374 698488 405430
rect 698544 405374 698612 405430
rect 698668 405374 698736 405430
rect 698792 405374 698922 405430
rect 697922 405306 698922 405374
rect 697922 405250 697992 405306
rect 698048 405250 698116 405306
rect 698172 405250 698240 405306
rect 698296 405250 698364 405306
rect 698420 405250 698488 405306
rect 698544 405250 698612 405306
rect 698668 405250 698736 405306
rect 698792 405250 698922 405306
rect 697922 405182 698922 405250
rect 697922 405126 697992 405182
rect 698048 405126 698116 405182
rect 698172 405126 698240 405182
rect 698296 405126 698364 405182
rect 698420 405126 698488 405182
rect 698544 405126 698612 405182
rect 698668 405126 698736 405182
rect 698792 405126 698922 405182
rect 697922 405058 698922 405126
rect 697922 405002 697992 405058
rect 698048 405002 698116 405058
rect 698172 405002 698240 405058
rect 698296 405002 698364 405058
rect 698420 405002 698488 405058
rect 698544 405002 698612 405058
rect 698668 405002 698736 405058
rect 698792 405002 698922 405058
rect 697922 404934 698922 405002
rect 697922 404878 697992 404934
rect 698048 404878 698116 404934
rect 698172 404878 698240 404934
rect 698296 404878 698364 404934
rect 698420 404878 698488 404934
rect 698544 404878 698612 404934
rect 698668 404878 698736 404934
rect 698792 404878 698922 404934
rect 697922 404810 698922 404878
rect 697922 404754 697992 404810
rect 698048 404754 698116 404810
rect 698172 404754 698240 404810
rect 698296 404754 698364 404810
rect 698420 404754 698488 404810
rect 698544 404754 698612 404810
rect 698668 404754 698736 404810
rect 698792 404754 698922 404810
rect 697922 404686 698922 404754
rect 697922 404630 697992 404686
rect 698048 404630 698116 404686
rect 698172 404630 698240 404686
rect 698296 404630 698364 404686
rect 698420 404630 698488 404686
rect 698544 404630 698612 404686
rect 698668 404630 698736 404686
rect 698792 404630 698922 404686
rect 697922 404562 698922 404630
rect 697922 404506 697992 404562
rect 698048 404506 698116 404562
rect 698172 404506 698240 404562
rect 698296 404506 698364 404562
rect 698420 404506 698488 404562
rect 698544 404506 698612 404562
rect 698668 404506 698736 404562
rect 698792 404506 698922 404562
rect 697922 404438 698922 404506
rect 697922 404382 697992 404438
rect 698048 404382 698116 404438
rect 698172 404382 698240 404438
rect 698296 404382 698364 404438
rect 698420 404382 698488 404438
rect 698544 404382 698612 404438
rect 698668 404382 698736 404438
rect 698792 404382 698922 404438
rect 697922 404314 698922 404382
rect 697922 404258 697992 404314
rect 698048 404258 698116 404314
rect 698172 404258 698240 404314
rect 698296 404258 698364 404314
rect 698420 404258 698488 404314
rect 698544 404258 698612 404314
rect 698668 404258 698736 404314
rect 698792 404258 698922 404314
rect 697922 404190 698922 404258
rect 697922 404134 697992 404190
rect 698048 404134 698116 404190
rect 698172 404134 698240 404190
rect 698296 404134 698364 404190
rect 698420 404134 698488 404190
rect 698544 404134 698612 404190
rect 698668 404134 698736 404190
rect 698792 404134 698922 404190
rect 697922 404066 698922 404134
rect 697922 404010 697992 404066
rect 698048 404010 698116 404066
rect 698172 404010 698240 404066
rect 698296 404010 698364 404066
rect 698420 404010 698488 404066
rect 698544 404010 698612 404066
rect 698668 404010 698736 404066
rect 698792 404010 698922 404066
rect 697922 403942 698922 404010
rect 697922 403886 697992 403942
rect 698048 403886 698116 403942
rect 698172 403886 698240 403942
rect 698296 403886 698364 403942
rect 698420 403886 698488 403942
rect 698544 403886 698612 403942
rect 698668 403886 698736 403942
rect 698792 403886 698922 403942
rect 697922 403096 698922 403886
rect 697922 403040 697992 403096
rect 698048 403040 698116 403096
rect 698172 403040 698240 403096
rect 698296 403040 698364 403096
rect 698420 403040 698488 403096
rect 698544 403040 698612 403096
rect 698668 403040 698736 403096
rect 698792 403040 698922 403096
rect 697922 402972 698922 403040
rect 697922 402916 697992 402972
rect 698048 402916 698116 402972
rect 698172 402916 698240 402972
rect 698296 402916 698364 402972
rect 698420 402916 698488 402972
rect 698544 402916 698612 402972
rect 698668 402916 698736 402972
rect 698792 402916 698922 402972
rect 697922 402848 698922 402916
rect 697922 402792 697992 402848
rect 698048 402792 698116 402848
rect 698172 402792 698240 402848
rect 698296 402792 698364 402848
rect 698420 402792 698488 402848
rect 698544 402792 698612 402848
rect 698668 402792 698736 402848
rect 698792 402792 698922 402848
rect 697922 402724 698922 402792
rect 697922 402668 697992 402724
rect 698048 402668 698116 402724
rect 698172 402668 698240 402724
rect 698296 402668 698364 402724
rect 698420 402668 698488 402724
rect 698544 402668 698612 402724
rect 698668 402668 698736 402724
rect 698792 402668 698922 402724
rect 697922 402600 698922 402668
rect 697922 402544 697992 402600
rect 698048 402544 698116 402600
rect 698172 402544 698240 402600
rect 698296 402544 698364 402600
rect 698420 402544 698488 402600
rect 698544 402544 698612 402600
rect 698668 402544 698736 402600
rect 698792 402544 698922 402600
rect 697922 402476 698922 402544
rect 697922 402420 697992 402476
rect 698048 402420 698116 402476
rect 698172 402420 698240 402476
rect 698296 402420 698364 402476
rect 698420 402420 698488 402476
rect 698544 402420 698612 402476
rect 698668 402420 698736 402476
rect 698792 402420 698922 402476
rect 697922 402352 698922 402420
rect 697922 402296 697992 402352
rect 698048 402296 698116 402352
rect 698172 402296 698240 402352
rect 698296 402296 698364 402352
rect 698420 402296 698488 402352
rect 698544 402296 698612 402352
rect 698668 402296 698736 402352
rect 698792 402296 698922 402352
rect 697922 402228 698922 402296
rect 697922 402172 697992 402228
rect 698048 402172 698116 402228
rect 698172 402172 698240 402228
rect 698296 402172 698364 402228
rect 698420 402172 698488 402228
rect 698544 402172 698612 402228
rect 698668 402172 698736 402228
rect 698792 402172 698922 402228
rect 697922 402104 698922 402172
rect 697922 402048 697992 402104
rect 698048 402048 698116 402104
rect 698172 402048 698240 402104
rect 698296 402048 698364 402104
rect 698420 402048 698488 402104
rect 698544 402048 698612 402104
rect 698668 402048 698736 402104
rect 698792 402048 698922 402104
rect 697922 401980 698922 402048
rect 697922 401924 697992 401980
rect 698048 401924 698116 401980
rect 698172 401924 698240 401980
rect 698296 401924 698364 401980
rect 698420 401924 698488 401980
rect 698544 401924 698612 401980
rect 698668 401924 698736 401980
rect 698792 401924 698922 401980
rect 697922 401856 698922 401924
rect 697922 401800 697992 401856
rect 698048 401800 698116 401856
rect 698172 401800 698240 401856
rect 698296 401800 698364 401856
rect 698420 401800 698488 401856
rect 698544 401800 698612 401856
rect 698668 401800 698736 401856
rect 698792 401800 698922 401856
rect 697922 401732 698922 401800
rect 697922 401676 697992 401732
rect 698048 401676 698116 401732
rect 698172 401676 698240 401732
rect 698296 401676 698364 401732
rect 698420 401676 698488 401732
rect 698544 401676 698612 401732
rect 698668 401676 698736 401732
rect 698792 401676 698922 401732
rect 697922 401608 698922 401676
rect 697922 401552 697992 401608
rect 698048 401552 698116 401608
rect 698172 401552 698240 401608
rect 698296 401552 698364 401608
rect 698420 401552 698488 401608
rect 698544 401552 698612 401608
rect 698668 401552 698736 401608
rect 698792 401552 698922 401608
rect 697922 401484 698922 401552
rect 697922 401428 697992 401484
rect 698048 401428 698116 401484
rect 698172 401428 698240 401484
rect 698296 401428 698364 401484
rect 698420 401428 698488 401484
rect 698544 401428 698612 401484
rect 698668 401428 698736 401484
rect 698792 401428 698922 401484
rect 697922 401360 698922 401428
rect 697922 401304 697992 401360
rect 698048 401304 698116 401360
rect 698172 401304 698240 401360
rect 698296 401304 698364 401360
rect 698420 401304 698488 401360
rect 698544 401304 698612 401360
rect 698668 401304 698736 401360
rect 698792 401304 698922 401360
rect 697922 401236 698922 401304
rect 697922 401180 697992 401236
rect 698048 401180 698116 401236
rect 698172 401180 698240 401236
rect 698296 401180 698364 401236
rect 698420 401180 698488 401236
rect 698544 401180 698612 401236
rect 698668 401180 698736 401236
rect 698792 401180 698922 401236
rect 697922 400726 698922 401180
rect 697922 400670 697992 400726
rect 698048 400670 698116 400726
rect 698172 400670 698240 400726
rect 698296 400670 698364 400726
rect 698420 400670 698488 400726
rect 698544 400670 698612 400726
rect 698668 400670 698736 400726
rect 698792 400670 698922 400726
rect 697922 400602 698922 400670
rect 697922 400546 697992 400602
rect 698048 400546 698116 400602
rect 698172 400546 698240 400602
rect 698296 400546 698364 400602
rect 698420 400546 698488 400602
rect 698544 400546 698612 400602
rect 698668 400546 698736 400602
rect 698792 400546 698922 400602
rect 697922 400478 698922 400546
rect 697922 400422 697992 400478
rect 698048 400422 698116 400478
rect 698172 400422 698240 400478
rect 698296 400422 698364 400478
rect 698420 400422 698488 400478
rect 698544 400422 698612 400478
rect 698668 400422 698736 400478
rect 698792 400422 698922 400478
rect 697922 400354 698922 400422
rect 697922 400298 697992 400354
rect 698048 400298 698116 400354
rect 698172 400298 698240 400354
rect 698296 400298 698364 400354
rect 698420 400298 698488 400354
rect 698544 400298 698612 400354
rect 698668 400298 698736 400354
rect 698792 400298 698922 400354
rect 697922 400230 698922 400298
rect 697922 400174 697992 400230
rect 698048 400174 698116 400230
rect 698172 400174 698240 400230
rect 698296 400174 698364 400230
rect 698420 400174 698488 400230
rect 698544 400174 698612 400230
rect 698668 400174 698736 400230
rect 698792 400174 698922 400230
rect 697922 400106 698922 400174
rect 697922 400050 697992 400106
rect 698048 400050 698116 400106
rect 698172 400050 698240 400106
rect 698296 400050 698364 400106
rect 698420 400050 698488 400106
rect 698544 400050 698612 400106
rect 698668 400050 698736 400106
rect 698792 400050 698922 400106
rect 697922 399982 698922 400050
rect 697922 399926 697992 399982
rect 698048 399926 698116 399982
rect 698172 399926 698240 399982
rect 698296 399926 698364 399982
rect 698420 399926 698488 399982
rect 698544 399926 698612 399982
rect 698668 399926 698736 399982
rect 698792 399926 698922 399982
rect 697922 399858 698922 399926
rect 697922 399802 697992 399858
rect 698048 399802 698116 399858
rect 698172 399802 698240 399858
rect 698296 399802 698364 399858
rect 698420 399802 698488 399858
rect 698544 399802 698612 399858
rect 698668 399802 698736 399858
rect 698792 399802 698922 399858
rect 697922 399734 698922 399802
rect 697922 399678 697992 399734
rect 698048 399678 698116 399734
rect 698172 399678 698240 399734
rect 698296 399678 698364 399734
rect 698420 399678 698488 399734
rect 698544 399678 698612 399734
rect 698668 399678 698736 399734
rect 698792 399678 698922 399734
rect 697922 399610 698922 399678
rect 697922 399554 697992 399610
rect 698048 399554 698116 399610
rect 698172 399554 698240 399610
rect 698296 399554 698364 399610
rect 698420 399554 698488 399610
rect 698544 399554 698612 399610
rect 698668 399554 698736 399610
rect 698792 399554 698922 399610
rect 697922 399486 698922 399554
rect 697922 399430 697992 399486
rect 698048 399430 698116 399486
rect 698172 399430 698240 399486
rect 698296 399430 698364 399486
rect 698420 399430 698488 399486
rect 698544 399430 698612 399486
rect 698668 399430 698736 399486
rect 698792 399430 698922 399486
rect 697922 399362 698922 399430
rect 697922 399306 697992 399362
rect 698048 399306 698116 399362
rect 698172 399306 698240 399362
rect 698296 399306 698364 399362
rect 698420 399306 698488 399362
rect 698544 399306 698612 399362
rect 698668 399306 698736 399362
rect 698792 399306 698922 399362
rect 697922 399238 698922 399306
rect 697922 399182 697992 399238
rect 698048 399182 698116 399238
rect 698172 399182 698240 399238
rect 698296 399182 698364 399238
rect 698420 399182 698488 399238
rect 698544 399182 698612 399238
rect 698668 399182 698736 399238
rect 698792 399182 698922 399238
rect 697922 399114 698922 399182
rect 697922 399058 697992 399114
rect 698048 399058 698116 399114
rect 698172 399058 698240 399114
rect 698296 399058 698364 399114
rect 698420 399058 698488 399114
rect 698544 399058 698612 399114
rect 698668 399058 698736 399114
rect 698792 399058 698922 399114
rect 697922 398990 698922 399058
rect 697922 398934 697992 398990
rect 698048 398934 698116 398990
rect 698172 398934 698240 398990
rect 698296 398934 698364 398990
rect 698420 398934 698488 398990
rect 698544 398934 698612 398990
rect 698668 398934 698736 398990
rect 698792 398934 698922 398990
rect 697922 398866 698922 398934
rect 697922 398810 697992 398866
rect 698048 398810 698116 398866
rect 698172 398810 698240 398866
rect 698296 398810 698364 398866
rect 698420 398810 698488 398866
rect 698544 398810 698612 398866
rect 698668 398810 698736 398866
rect 698792 398810 698922 398866
rect 697922 398122 698922 398810
rect 697922 398066 697992 398122
rect 698048 398066 698116 398122
rect 698172 398066 698240 398122
rect 698296 398066 698364 398122
rect 698420 398066 698488 398122
rect 698544 398066 698612 398122
rect 698668 398066 698736 398122
rect 698792 398066 698922 398122
rect 697922 397998 698922 398066
rect 697922 397942 697992 397998
rect 698048 397942 698116 397998
rect 698172 397942 698240 397998
rect 698296 397942 698364 397998
rect 698420 397942 698488 397998
rect 698544 397942 698612 397998
rect 698668 397942 698736 397998
rect 698792 397942 698922 397998
rect 697922 397874 698922 397942
rect 697922 397818 697992 397874
rect 698048 397818 698116 397874
rect 698172 397818 698240 397874
rect 698296 397818 698364 397874
rect 698420 397818 698488 397874
rect 698544 397818 698612 397874
rect 698668 397818 698736 397874
rect 698792 397818 698922 397874
rect 697922 397750 698922 397818
rect 697922 397694 697992 397750
rect 698048 397694 698116 397750
rect 698172 397694 698240 397750
rect 698296 397694 698364 397750
rect 698420 397694 698488 397750
rect 698544 397694 698612 397750
rect 698668 397694 698736 397750
rect 698792 397694 698922 397750
rect 697922 397626 698922 397694
rect 697922 397570 697992 397626
rect 698048 397570 698116 397626
rect 698172 397570 698240 397626
rect 698296 397570 698364 397626
rect 698420 397570 698488 397626
rect 698544 397570 698612 397626
rect 698668 397570 698736 397626
rect 698792 397570 698922 397626
rect 697922 397502 698922 397570
rect 697922 397446 697992 397502
rect 698048 397446 698116 397502
rect 698172 397446 698240 397502
rect 698296 397446 698364 397502
rect 698420 397446 698488 397502
rect 698544 397446 698612 397502
rect 698668 397446 698736 397502
rect 698792 397446 698922 397502
rect 697922 397378 698922 397446
rect 697922 397322 697992 397378
rect 698048 397322 698116 397378
rect 698172 397322 698240 397378
rect 698296 397322 698364 397378
rect 698420 397322 698488 397378
rect 698544 397322 698612 397378
rect 698668 397322 698736 397378
rect 698792 397322 698922 397378
rect 697922 397254 698922 397322
rect 697922 397198 697992 397254
rect 698048 397198 698116 397254
rect 698172 397198 698240 397254
rect 698296 397198 698364 397254
rect 698420 397198 698488 397254
rect 698544 397198 698612 397254
rect 698668 397198 698736 397254
rect 698792 397198 698922 397254
rect 697922 397130 698922 397198
rect 697922 397074 697992 397130
rect 698048 397074 698116 397130
rect 698172 397074 698240 397130
rect 698296 397074 698364 397130
rect 698420 397074 698488 397130
rect 698544 397074 698612 397130
rect 698668 397074 698736 397130
rect 698792 397074 698922 397130
rect 697922 397006 698922 397074
rect 697922 396950 697992 397006
rect 698048 396950 698116 397006
rect 698172 396950 698240 397006
rect 698296 396950 698364 397006
rect 698420 396950 698488 397006
rect 698544 396950 698612 397006
rect 698668 396950 698736 397006
rect 698792 396950 698922 397006
rect 697922 396882 698922 396950
rect 697922 396826 697992 396882
rect 698048 396826 698116 396882
rect 698172 396826 698240 396882
rect 698296 396826 698364 396882
rect 698420 396826 698488 396882
rect 698544 396826 698612 396882
rect 698668 396826 698736 396882
rect 698792 396826 698922 396882
rect 697922 396758 698922 396826
rect 697922 396702 697992 396758
rect 698048 396702 698116 396758
rect 698172 396702 698240 396758
rect 698296 396702 698364 396758
rect 698420 396702 698488 396758
rect 698544 396702 698612 396758
rect 698668 396702 698736 396758
rect 698792 396702 698922 396758
rect 697922 396634 698922 396702
rect 697922 396578 697992 396634
rect 698048 396578 698116 396634
rect 698172 396578 698240 396634
rect 698296 396578 698364 396634
rect 698420 396578 698488 396634
rect 698544 396578 698612 396634
rect 698668 396578 698736 396634
rect 698792 396578 698922 396634
rect 697922 396510 698922 396578
rect 697922 396454 697992 396510
rect 698048 396454 698116 396510
rect 698172 396454 698240 396510
rect 698296 396454 698364 396510
rect 698420 396454 698488 396510
rect 698544 396454 698612 396510
rect 698668 396454 698736 396510
rect 698792 396454 698922 396510
rect 697922 396386 698922 396454
rect 697922 396330 697992 396386
rect 698048 396330 698116 396386
rect 698172 396330 698240 396386
rect 698296 396330 698364 396386
rect 698420 396330 698488 396386
rect 698544 396330 698612 396386
rect 698668 396330 698736 396386
rect 698792 396330 698922 396386
rect 697922 392429 698922 396330
rect 697922 392373 698144 392429
rect 698200 392373 698444 392429
rect 698500 392373 698744 392429
rect 698800 392373 698922 392429
rect 697922 392229 698922 392373
rect 697922 392173 698144 392229
rect 698200 392173 698444 392229
rect 698500 392173 698744 392229
rect 698800 392173 698922 392229
rect 697922 363434 698922 392173
rect 697922 363378 698044 363434
rect 698100 363378 698344 363434
rect 698400 363378 698644 363434
rect 698700 363378 698922 363434
rect 697922 356429 698922 363378
rect 697922 356373 698144 356429
rect 698200 356373 698444 356429
rect 698500 356373 698744 356429
rect 698800 356373 698922 356429
rect 697922 356229 698922 356373
rect 697922 356173 698144 356229
rect 698200 356173 698444 356229
rect 698500 356173 698744 356229
rect 698800 356173 698922 356229
rect 697922 349434 698922 356173
rect 697922 349378 698044 349434
rect 698100 349378 698344 349434
rect 698400 349378 698644 349434
rect 698700 349378 698922 349434
rect 79078 330984 79208 331040
rect 79264 330984 79332 331040
rect 79388 330984 79456 331040
rect 79512 330984 79580 331040
rect 79636 330984 79704 331040
rect 79760 330984 79828 331040
rect 79884 330984 79952 331040
rect 80008 330984 80078 331040
rect 79078 330916 80078 330984
rect 79078 330860 79208 330916
rect 79264 330860 79332 330916
rect 79388 330860 79456 330916
rect 79512 330860 79580 330916
rect 79636 330860 79704 330916
rect 79760 330860 79828 330916
rect 79884 330860 79952 330916
rect 80008 330860 80078 330916
rect 79078 330792 80078 330860
rect 79078 330736 79208 330792
rect 79264 330736 79332 330792
rect 79388 330736 79456 330792
rect 79512 330736 79580 330792
rect 79636 330736 79704 330792
rect 79760 330736 79828 330792
rect 79884 330736 79952 330792
rect 80008 330736 80078 330792
rect 79078 330668 80078 330736
rect 79078 330612 79208 330668
rect 79264 330612 79332 330668
rect 79388 330612 79456 330668
rect 79512 330612 79580 330668
rect 79636 330612 79704 330668
rect 79760 330612 79828 330668
rect 79884 330612 79952 330668
rect 80008 330612 80078 330668
rect 79078 330544 80078 330612
rect 79078 330488 79208 330544
rect 79264 330488 79332 330544
rect 79388 330488 79456 330544
rect 79512 330488 79580 330544
rect 79636 330488 79704 330544
rect 79760 330488 79828 330544
rect 79884 330488 79952 330544
rect 80008 330488 80078 330544
rect 79078 330420 80078 330488
rect 79078 330364 79208 330420
rect 79264 330364 79332 330420
rect 79388 330364 79456 330420
rect 79512 330364 79580 330420
rect 79636 330364 79704 330420
rect 79760 330364 79828 330420
rect 79884 330364 79952 330420
rect 80008 330364 80078 330420
rect 79078 330296 80078 330364
rect 79078 330240 79208 330296
rect 79264 330240 79332 330296
rect 79388 330240 79456 330296
rect 79512 330240 79580 330296
rect 79636 330240 79704 330296
rect 79760 330240 79828 330296
rect 79884 330240 79952 330296
rect 80008 330240 80078 330296
rect 79078 314622 80078 330240
rect 88006 329488 88626 334520
rect 106006 330888 106626 333560
rect 106006 330832 106207 330888
rect 106263 330832 106407 330888
rect 106463 330832 106626 330888
rect 106006 330588 106626 330832
rect 106006 330532 106207 330588
rect 106263 330532 106407 330588
rect 106463 330532 106626 330588
rect 106006 330288 106626 330532
rect 106006 330232 106207 330288
rect 106263 330232 106407 330288
rect 106463 330232 106626 330288
rect 106006 330110 106626 330232
rect 88006 329432 88207 329488
rect 88263 329432 88407 329488
rect 88463 329432 88626 329488
rect 88006 329188 88626 329432
rect 88006 329132 88207 329188
rect 88263 329132 88407 329188
rect 88463 329132 88626 329188
rect 88006 328888 88626 329132
rect 88006 328832 88207 328888
rect 88263 328832 88407 328888
rect 88463 328832 88626 328888
rect 88006 328710 88626 328832
rect 124006 329488 124626 334520
rect 142006 330888 142626 333560
rect 142006 330832 142207 330888
rect 142263 330832 142407 330888
rect 142463 330832 142626 330888
rect 142006 330588 142626 330832
rect 142006 330532 142207 330588
rect 142263 330532 142407 330588
rect 142463 330532 142626 330588
rect 142006 330288 142626 330532
rect 142006 330232 142207 330288
rect 142263 330232 142407 330288
rect 142463 330232 142626 330288
rect 142006 330110 142626 330232
rect 158108 331040 158728 331110
rect 158108 330984 158178 331040
rect 158234 330984 158302 331040
rect 158358 330984 158426 331040
rect 158482 330984 158550 331040
rect 158606 330984 158728 331040
rect 158108 330916 158728 330984
rect 158108 330860 158178 330916
rect 158234 330860 158302 330916
rect 158358 330860 158426 330916
rect 158482 330860 158550 330916
rect 158606 330860 158728 330916
rect 158108 330792 158728 330860
rect 158108 330736 158178 330792
rect 158234 330736 158302 330792
rect 158358 330736 158426 330792
rect 158482 330736 158550 330792
rect 158606 330736 158728 330792
rect 158108 330668 158728 330736
rect 158108 330612 158178 330668
rect 158234 330612 158302 330668
rect 158358 330612 158426 330668
rect 158482 330612 158550 330668
rect 158606 330612 158728 330668
rect 158108 330544 158728 330612
rect 158108 330488 158178 330544
rect 158234 330488 158302 330544
rect 158358 330488 158426 330544
rect 158482 330488 158550 330544
rect 158606 330488 158728 330544
rect 158108 330420 158728 330488
rect 158108 330364 158178 330420
rect 158234 330364 158302 330420
rect 158358 330364 158426 330420
rect 158482 330364 158550 330420
rect 158606 330364 158728 330420
rect 158108 330296 158728 330364
rect 158108 330240 158178 330296
rect 158234 330240 158302 330296
rect 158358 330240 158426 330296
rect 158482 330240 158550 330296
rect 158606 330240 158728 330296
rect 124006 329432 124207 329488
rect 124263 329432 124407 329488
rect 124463 329432 124626 329488
rect 124006 329188 124626 329432
rect 124006 329132 124207 329188
rect 124263 329132 124407 329188
rect 124463 329132 124626 329188
rect 124006 328888 124626 329132
rect 124006 328832 124207 328888
rect 124263 328832 124407 328888
rect 124463 328832 124626 328888
rect 124006 328710 124626 328832
rect 157088 329640 157708 329710
rect 157088 329584 157158 329640
rect 157214 329584 157282 329640
rect 157338 329584 157406 329640
rect 157462 329584 157530 329640
rect 157586 329584 157708 329640
rect 157088 329516 157708 329584
rect 157088 329460 157158 329516
rect 157214 329460 157282 329516
rect 157338 329460 157406 329516
rect 157462 329460 157530 329516
rect 157586 329460 157708 329516
rect 157088 329392 157708 329460
rect 157088 329336 157158 329392
rect 157214 329336 157282 329392
rect 157338 329336 157406 329392
rect 157462 329336 157530 329392
rect 157586 329336 157708 329392
rect 157088 329268 157708 329336
rect 157088 329212 157158 329268
rect 157214 329212 157282 329268
rect 157338 329212 157406 329268
rect 157462 329212 157530 329268
rect 157586 329212 157708 329268
rect 157088 329144 157708 329212
rect 157088 329088 157158 329144
rect 157214 329088 157282 329144
rect 157338 329088 157406 329144
rect 157462 329088 157530 329144
rect 157586 329088 157708 329144
rect 157088 329020 157708 329088
rect 157088 328964 157158 329020
rect 157214 328964 157282 329020
rect 157338 328964 157406 329020
rect 157462 328964 157530 329020
rect 157586 328964 157708 329020
rect 157088 328896 157708 328964
rect 157088 328840 157158 328896
rect 157214 328840 157282 328896
rect 157338 328840 157406 328896
rect 157462 328840 157530 328896
rect 157586 328840 157708 328896
rect 79078 314566 79300 314622
rect 79356 314566 79600 314622
rect 79656 314566 79900 314622
rect 79956 314566 80078 314622
rect 79078 307622 80078 314566
rect 157088 318424 157708 328840
rect 157088 318368 157210 318424
rect 157266 318368 157510 318424
rect 157566 318368 157708 318424
rect 157088 317026 157708 318368
rect 157088 316970 157210 317026
rect 157266 316970 157510 317026
rect 157566 316970 157708 317026
rect 157088 315628 157708 316970
rect 157088 315572 157210 315628
rect 157266 315572 157510 315628
rect 157566 315572 157708 315628
rect 79078 307566 79300 307622
rect 79356 307566 79600 307622
rect 79656 307566 79900 307622
rect 79956 307566 80078 307622
rect 79078 307186 80078 307566
rect 79078 307130 79208 307186
rect 79264 307130 79332 307186
rect 79388 307130 79456 307186
rect 79512 307130 79580 307186
rect 79636 307130 79704 307186
rect 79760 307130 79828 307186
rect 79884 307130 79952 307186
rect 80008 307130 80078 307186
rect 79078 307062 80078 307130
rect 79078 307006 79208 307062
rect 79264 307006 79332 307062
rect 79388 307006 79456 307062
rect 79512 307006 79580 307062
rect 79636 307006 79704 307062
rect 79760 307006 79828 307062
rect 79884 307006 79952 307062
rect 80008 307006 80078 307062
rect 79078 306938 80078 307006
rect 79078 306882 79208 306938
rect 79264 306882 79332 306938
rect 79388 306882 79456 306938
rect 79512 306882 79580 306938
rect 79636 306882 79704 306938
rect 79760 306882 79828 306938
rect 79884 306882 79952 306938
rect 80008 306882 80078 306938
rect 79078 306814 80078 306882
rect 79078 306758 79208 306814
rect 79264 306758 79332 306814
rect 79388 306758 79456 306814
rect 79512 306758 79580 306814
rect 79636 306758 79704 306814
rect 79760 306758 79828 306814
rect 79884 306758 79952 306814
rect 80008 306758 80078 306814
rect 79078 306690 80078 306758
rect 79078 306634 79208 306690
rect 79264 306634 79332 306690
rect 79388 306634 79456 306690
rect 79512 306634 79580 306690
rect 79636 306634 79704 306690
rect 79760 306634 79828 306690
rect 79884 306634 79952 306690
rect 80008 306634 80078 306690
rect 79078 306566 80078 306634
rect 79078 306510 79208 306566
rect 79264 306510 79332 306566
rect 79388 306510 79456 306566
rect 79512 306510 79580 306566
rect 79636 306510 79704 306566
rect 79760 306510 79828 306566
rect 79884 306510 79952 306566
rect 80008 306510 80078 306566
rect 79078 306442 80078 306510
rect 79078 306386 79208 306442
rect 79264 306386 79332 306442
rect 79388 306386 79456 306442
rect 79512 306386 79580 306442
rect 79636 306386 79704 306442
rect 79760 306386 79828 306442
rect 79884 306386 79952 306442
rect 80008 306386 80078 306442
rect 79078 300622 80078 306386
rect 114555 305786 114875 314284
rect 116150 307186 116470 314284
rect 116150 307130 116220 307186
rect 116276 307130 116344 307186
rect 116400 307130 116470 307186
rect 116150 307062 116470 307130
rect 116150 307006 116220 307062
rect 116276 307006 116344 307062
rect 116400 307006 116470 307062
rect 116150 306938 116470 307006
rect 116150 306882 116220 306938
rect 116276 306882 116344 306938
rect 116400 306882 116470 306938
rect 116150 306814 116470 306882
rect 116150 306758 116220 306814
rect 116276 306758 116344 306814
rect 116400 306758 116470 306814
rect 116150 306690 116470 306758
rect 116150 306634 116220 306690
rect 116276 306634 116344 306690
rect 116400 306634 116470 306690
rect 116150 306566 116470 306634
rect 116150 306510 116220 306566
rect 116276 306510 116344 306566
rect 116400 306510 116470 306566
rect 116150 306442 116470 306510
rect 116150 306386 116220 306442
rect 116276 306386 116344 306442
rect 116400 306386 116470 306442
rect 116150 306256 116470 306386
rect 114555 305730 114625 305786
rect 114681 305730 114749 305786
rect 114805 305730 114875 305786
rect 114555 305662 114875 305730
rect 114555 305606 114625 305662
rect 114681 305606 114749 305662
rect 114805 305606 114875 305662
rect 114555 305538 114875 305606
rect 114555 305482 114625 305538
rect 114681 305482 114749 305538
rect 114805 305482 114875 305538
rect 114555 305414 114875 305482
rect 114555 305358 114625 305414
rect 114681 305358 114749 305414
rect 114805 305358 114875 305414
rect 114555 305290 114875 305358
rect 114555 305234 114625 305290
rect 114681 305234 114749 305290
rect 114805 305234 114875 305290
rect 114555 305166 114875 305234
rect 114555 305110 114625 305166
rect 114681 305110 114749 305166
rect 114805 305110 114875 305166
rect 114555 305042 114875 305110
rect 114555 304986 114625 305042
rect 114681 304986 114749 305042
rect 114805 304986 114875 305042
rect 114555 304856 114875 304986
rect 117745 305786 118065 314284
rect 119340 307186 119660 314284
rect 119340 307130 119410 307186
rect 119466 307130 119534 307186
rect 119590 307130 119660 307186
rect 119340 307062 119660 307130
rect 119340 307006 119410 307062
rect 119466 307006 119534 307062
rect 119590 307006 119660 307062
rect 119340 306938 119660 307006
rect 119340 306882 119410 306938
rect 119466 306882 119534 306938
rect 119590 306882 119660 306938
rect 119340 306814 119660 306882
rect 119340 306758 119410 306814
rect 119466 306758 119534 306814
rect 119590 306758 119660 306814
rect 119340 306690 119660 306758
rect 119340 306634 119410 306690
rect 119466 306634 119534 306690
rect 119590 306634 119660 306690
rect 119340 306566 119660 306634
rect 119340 306510 119410 306566
rect 119466 306510 119534 306566
rect 119590 306510 119660 306566
rect 119340 306442 119660 306510
rect 119340 306386 119410 306442
rect 119466 306386 119534 306442
rect 119590 306386 119660 306442
rect 119340 306256 119660 306386
rect 117745 305730 117815 305786
rect 117871 305730 117939 305786
rect 117995 305730 118065 305786
rect 117745 305662 118065 305730
rect 117745 305606 117815 305662
rect 117871 305606 117939 305662
rect 117995 305606 118065 305662
rect 117745 305538 118065 305606
rect 117745 305482 117815 305538
rect 117871 305482 117939 305538
rect 117995 305482 118065 305538
rect 117745 305414 118065 305482
rect 117745 305358 117815 305414
rect 117871 305358 117939 305414
rect 117995 305358 118065 305414
rect 117745 305290 118065 305358
rect 117745 305234 117815 305290
rect 117871 305234 117939 305290
rect 117995 305234 118065 305290
rect 117745 305166 118065 305234
rect 117745 305110 117815 305166
rect 117871 305110 117939 305166
rect 117995 305110 118065 305166
rect 117745 305042 118065 305110
rect 117745 304986 117815 305042
rect 117871 304986 117939 305042
rect 117995 304986 118065 305042
rect 117745 304856 118065 304986
rect 120935 305786 121255 314284
rect 122530 307186 122850 314284
rect 122530 307130 122600 307186
rect 122656 307130 122724 307186
rect 122780 307130 122850 307186
rect 122530 307062 122850 307130
rect 122530 307006 122600 307062
rect 122656 307006 122724 307062
rect 122780 307006 122850 307062
rect 122530 306938 122850 307006
rect 122530 306882 122600 306938
rect 122656 306882 122724 306938
rect 122780 306882 122850 306938
rect 122530 306814 122850 306882
rect 122530 306758 122600 306814
rect 122656 306758 122724 306814
rect 122780 306758 122850 306814
rect 122530 306690 122850 306758
rect 122530 306634 122600 306690
rect 122656 306634 122724 306690
rect 122780 306634 122850 306690
rect 122530 306566 122850 306634
rect 122530 306510 122600 306566
rect 122656 306510 122724 306566
rect 122780 306510 122850 306566
rect 122530 306442 122850 306510
rect 122530 306386 122600 306442
rect 122656 306386 122724 306442
rect 122780 306386 122850 306442
rect 122530 306256 122850 306386
rect 120935 305730 121005 305786
rect 121061 305730 121129 305786
rect 121185 305730 121255 305786
rect 120935 305662 121255 305730
rect 120935 305606 121005 305662
rect 121061 305606 121129 305662
rect 121185 305606 121255 305662
rect 120935 305538 121255 305606
rect 120935 305482 121005 305538
rect 121061 305482 121129 305538
rect 121185 305482 121255 305538
rect 120935 305414 121255 305482
rect 120935 305358 121005 305414
rect 121061 305358 121129 305414
rect 121185 305358 121255 305414
rect 120935 305290 121255 305358
rect 120935 305234 121005 305290
rect 121061 305234 121129 305290
rect 121185 305234 121255 305290
rect 120935 305166 121255 305234
rect 120935 305110 121005 305166
rect 121061 305110 121129 305166
rect 121185 305110 121255 305166
rect 120935 305042 121255 305110
rect 120935 304986 121005 305042
rect 121061 304986 121129 305042
rect 121185 304986 121255 305042
rect 120935 304856 121255 304986
rect 124125 305786 124445 314284
rect 124125 305730 124195 305786
rect 124251 305730 124319 305786
rect 124375 305730 124445 305786
rect 124125 305662 124445 305730
rect 124125 305606 124195 305662
rect 124251 305606 124319 305662
rect 124375 305606 124445 305662
rect 124125 305538 124445 305606
rect 124125 305482 124195 305538
rect 124251 305482 124319 305538
rect 124375 305482 124445 305538
rect 124125 305414 124445 305482
rect 124125 305358 124195 305414
rect 124251 305358 124319 305414
rect 124375 305358 124445 305414
rect 124125 305290 124445 305358
rect 124125 305234 124195 305290
rect 124251 305234 124319 305290
rect 124375 305234 124445 305290
rect 124125 305166 124445 305234
rect 124125 305110 124195 305166
rect 124251 305110 124319 305166
rect 124375 305110 124445 305166
rect 124125 305042 124445 305110
rect 124125 304986 124195 305042
rect 124251 304986 124319 305042
rect 124375 304986 124445 305042
rect 124125 304856 124445 304986
rect 157088 314230 157708 315572
rect 157088 314174 157210 314230
rect 157266 314174 157510 314230
rect 157566 314174 157708 314230
rect 157088 305726 157708 314174
rect 158108 317725 158728 330240
rect 160006 329488 160626 334520
rect 178006 330888 178626 333560
rect 178006 330832 178207 330888
rect 178263 330832 178407 330888
rect 178463 330832 178626 330888
rect 178006 330588 178626 330832
rect 178006 330532 178207 330588
rect 178263 330532 178407 330588
rect 178463 330532 178626 330588
rect 178006 330288 178626 330532
rect 178006 330232 178207 330288
rect 178263 330232 178407 330288
rect 178463 330232 178626 330288
rect 178006 330110 178626 330232
rect 160006 329432 160207 329488
rect 160263 329432 160407 329488
rect 160463 329432 160626 329488
rect 160006 329188 160626 329432
rect 160006 329132 160207 329188
rect 160263 329132 160407 329188
rect 160463 329132 160626 329188
rect 160006 328888 160626 329132
rect 160006 328832 160207 328888
rect 160263 328832 160407 328888
rect 160463 328832 160626 328888
rect 160006 328710 160626 328832
rect 196006 329488 196626 334520
rect 214006 330888 214626 333560
rect 214006 330832 214207 330888
rect 214263 330832 214407 330888
rect 214463 330832 214626 330888
rect 214006 330588 214626 330832
rect 214006 330532 214207 330588
rect 214263 330532 214407 330588
rect 214463 330532 214626 330588
rect 214006 330288 214626 330532
rect 214006 330232 214207 330288
rect 214263 330232 214407 330288
rect 214463 330232 214626 330288
rect 214006 330110 214626 330232
rect 196006 329432 196207 329488
rect 196263 329432 196407 329488
rect 196463 329432 196626 329488
rect 196006 329188 196626 329432
rect 196006 329132 196207 329188
rect 196263 329132 196407 329188
rect 196463 329132 196626 329188
rect 196006 328888 196626 329132
rect 196006 328832 196207 328888
rect 196263 328832 196407 328888
rect 196463 328832 196626 328888
rect 196006 328710 196626 328832
rect 232006 329488 232626 334520
rect 250006 330888 250626 333560
rect 250006 330832 250207 330888
rect 250263 330832 250407 330888
rect 250463 330832 250626 330888
rect 250006 330588 250626 330832
rect 250006 330532 250207 330588
rect 250263 330532 250407 330588
rect 250463 330532 250626 330588
rect 250006 330288 250626 330532
rect 250006 330232 250207 330288
rect 250263 330232 250407 330288
rect 250463 330232 250626 330288
rect 250006 330110 250626 330232
rect 232006 329432 232207 329488
rect 232263 329432 232407 329488
rect 232463 329432 232626 329488
rect 232006 329188 232626 329432
rect 232006 329132 232207 329188
rect 232263 329132 232407 329188
rect 232463 329132 232626 329188
rect 232006 328888 232626 329132
rect 232006 328832 232207 328888
rect 232263 328832 232407 328888
rect 232463 328832 232626 328888
rect 232006 328710 232626 328832
rect 268006 329488 268626 334520
rect 286006 330888 286626 333560
rect 286006 330832 286207 330888
rect 286263 330832 286407 330888
rect 286463 330832 286626 330888
rect 286006 330588 286626 330832
rect 286006 330532 286207 330588
rect 286263 330532 286407 330588
rect 286463 330532 286626 330588
rect 286006 330288 286626 330532
rect 286006 330232 286207 330288
rect 286263 330232 286407 330288
rect 286463 330232 286626 330288
rect 286006 330110 286626 330232
rect 268006 329432 268207 329488
rect 268263 329432 268407 329488
rect 268463 329432 268626 329488
rect 268006 329188 268626 329432
rect 268006 329132 268207 329188
rect 268263 329132 268407 329188
rect 268463 329132 268626 329188
rect 268006 328888 268626 329132
rect 268006 328832 268207 328888
rect 268263 328832 268407 328888
rect 268463 328832 268626 328888
rect 268006 328710 268626 328832
rect 304006 329488 304626 334520
rect 322006 330888 322626 333560
rect 322006 330832 322207 330888
rect 322263 330832 322407 330888
rect 322463 330832 322626 330888
rect 322006 330588 322626 330832
rect 322006 330532 322207 330588
rect 322263 330532 322407 330588
rect 322463 330532 322626 330588
rect 322006 330288 322626 330532
rect 322006 330232 322207 330288
rect 322263 330232 322407 330288
rect 322463 330232 322626 330288
rect 322006 330110 322626 330232
rect 304006 329432 304207 329488
rect 304263 329432 304407 329488
rect 304463 329432 304626 329488
rect 304006 329188 304626 329432
rect 304006 329132 304207 329188
rect 304263 329132 304407 329188
rect 304463 329132 304626 329188
rect 304006 328888 304626 329132
rect 304006 328832 304207 328888
rect 304263 328832 304407 328888
rect 304463 328832 304626 328888
rect 304006 328710 304626 328832
rect 340006 329488 340626 334520
rect 358006 330888 358626 333560
rect 358006 330832 358207 330888
rect 358263 330832 358407 330888
rect 358463 330832 358626 330888
rect 358006 330588 358626 330832
rect 358006 330532 358207 330588
rect 358263 330532 358407 330588
rect 358463 330532 358626 330588
rect 358006 330288 358626 330532
rect 358006 330232 358207 330288
rect 358263 330232 358407 330288
rect 358463 330232 358626 330288
rect 358006 330110 358626 330232
rect 340006 329432 340207 329488
rect 340263 329432 340407 329488
rect 340463 329432 340626 329488
rect 340006 329188 340626 329432
rect 340006 329132 340207 329188
rect 340263 329132 340407 329188
rect 340463 329132 340626 329188
rect 340006 328888 340626 329132
rect 340006 328832 340207 328888
rect 340263 328832 340407 328888
rect 340463 328832 340626 328888
rect 340006 328710 340626 328832
rect 376006 329488 376626 334520
rect 376006 329432 376207 329488
rect 376263 329432 376407 329488
rect 376463 329432 376626 329488
rect 376006 329188 376626 329432
rect 376006 329132 376207 329188
rect 376263 329132 376407 329188
rect 376463 329132 376626 329188
rect 376006 328888 376626 329132
rect 376006 328832 376207 328888
rect 376263 328832 376407 328888
rect 376463 328832 376626 328888
rect 376006 328710 376626 328832
rect 381240 331040 381860 331110
rect 381240 330984 381310 331040
rect 381366 330984 381434 331040
rect 381490 330984 381558 331040
rect 381614 330984 381682 331040
rect 381738 330984 381860 331040
rect 381240 330916 381860 330984
rect 381240 330860 381310 330916
rect 381366 330860 381434 330916
rect 381490 330860 381558 330916
rect 381614 330860 381682 330916
rect 381738 330860 381860 330916
rect 381240 330792 381860 330860
rect 381240 330736 381310 330792
rect 381366 330736 381434 330792
rect 381490 330736 381558 330792
rect 381614 330736 381682 330792
rect 381738 330736 381860 330792
rect 381240 330668 381860 330736
rect 381240 330612 381310 330668
rect 381366 330612 381434 330668
rect 381490 330612 381558 330668
rect 381614 330612 381682 330668
rect 381738 330612 381860 330668
rect 381240 330544 381860 330612
rect 381240 330488 381310 330544
rect 381366 330488 381434 330544
rect 381490 330488 381558 330544
rect 381614 330488 381682 330544
rect 381738 330488 381860 330544
rect 381240 330420 381860 330488
rect 381240 330364 381310 330420
rect 381366 330364 381434 330420
rect 381490 330364 381558 330420
rect 381614 330364 381682 330420
rect 381738 330364 381860 330420
rect 381240 330296 381860 330364
rect 381240 330240 381310 330296
rect 381366 330240 381434 330296
rect 381490 330240 381558 330296
rect 381614 330240 381682 330296
rect 381738 330240 381860 330296
rect 158108 317669 158230 317725
rect 158286 317669 158530 317725
rect 158586 317669 158728 317725
rect 158108 316327 158728 317669
rect 158108 316271 158230 316327
rect 158286 316271 158530 316327
rect 158586 316271 158728 316327
rect 158108 314929 158728 316271
rect 158108 314873 158230 314929
rect 158286 314873 158530 314929
rect 158586 314873 158728 314929
rect 158108 307126 158728 314873
rect 158108 307070 158178 307126
rect 158234 307070 158302 307126
rect 158358 307070 158426 307126
rect 158482 307070 158550 307126
rect 158606 307070 158728 307126
rect 158108 307002 158728 307070
rect 158108 306946 158178 307002
rect 158234 306946 158302 307002
rect 158358 306946 158426 307002
rect 158482 306946 158550 307002
rect 158606 306946 158728 307002
rect 158108 306878 158728 306946
rect 158108 306822 158178 306878
rect 158234 306822 158302 306878
rect 158358 306822 158426 306878
rect 158482 306822 158550 306878
rect 158606 306822 158728 306878
rect 158108 306754 158728 306822
rect 158108 306698 158178 306754
rect 158234 306698 158302 306754
rect 158358 306698 158426 306754
rect 158482 306698 158550 306754
rect 158606 306698 158728 306754
rect 158108 306630 158728 306698
rect 158108 306574 158178 306630
rect 158234 306574 158302 306630
rect 158358 306574 158426 306630
rect 158482 306574 158550 306630
rect 158606 306574 158728 306630
rect 158108 306506 158728 306574
rect 158108 306450 158178 306506
rect 158234 306450 158302 306506
rect 158358 306450 158426 306506
rect 158482 306450 158550 306506
rect 158606 306450 158728 306506
rect 158108 306382 158728 306450
rect 158108 306326 158178 306382
rect 158234 306326 158302 306382
rect 158358 306326 158426 306382
rect 158482 306326 158550 306382
rect 158606 306326 158728 306382
rect 158108 306256 158728 306326
rect 381240 317727 381860 330240
rect 394006 330888 394626 333560
rect 394006 330832 394207 330888
rect 394263 330832 394407 330888
rect 394463 330832 394626 330888
rect 394006 330588 394626 330832
rect 394006 330532 394207 330588
rect 394263 330532 394407 330588
rect 394463 330532 394626 330588
rect 394006 330288 394626 330532
rect 394006 330232 394207 330288
rect 394263 330232 394407 330288
rect 394463 330232 394626 330288
rect 394006 330110 394626 330232
rect 381240 317671 381382 317727
rect 381438 317671 381682 317727
rect 381738 317671 381860 317727
rect 381240 316329 381860 317671
rect 381240 316273 381382 316329
rect 381438 316273 381682 316329
rect 381738 316273 381860 316329
rect 381240 314931 381860 316273
rect 381240 314875 381382 314931
rect 381438 314875 381682 314931
rect 381738 314875 381860 314931
rect 381240 307126 381860 314875
rect 381240 307070 381310 307126
rect 381366 307070 381434 307126
rect 381490 307070 381558 307126
rect 381614 307070 381682 307126
rect 381738 307070 381860 307126
rect 381240 307002 381860 307070
rect 381240 306946 381310 307002
rect 381366 306946 381434 307002
rect 381490 306946 381558 307002
rect 381614 306946 381682 307002
rect 381738 306946 381860 307002
rect 381240 306878 381860 306946
rect 381240 306822 381310 306878
rect 381366 306822 381434 306878
rect 381490 306822 381558 306878
rect 381614 306822 381682 306878
rect 381738 306822 381860 306878
rect 381240 306754 381860 306822
rect 381240 306698 381310 306754
rect 381366 306698 381434 306754
rect 381490 306698 381558 306754
rect 381614 306698 381682 306754
rect 381738 306698 381860 306754
rect 381240 306630 381860 306698
rect 381240 306574 381310 306630
rect 381366 306574 381434 306630
rect 381490 306574 381558 306630
rect 381614 306574 381682 306630
rect 381738 306574 381860 306630
rect 381240 306506 381860 306574
rect 381240 306450 381310 306506
rect 381366 306450 381434 306506
rect 381490 306450 381558 306506
rect 381614 306450 381682 306506
rect 381738 306450 381860 306506
rect 381240 306382 381860 306450
rect 381240 306326 381310 306382
rect 381366 306326 381434 306382
rect 381490 306326 381558 306382
rect 381614 306326 381682 306382
rect 381738 306326 381860 306382
rect 381240 306256 381860 306326
rect 382260 329640 382880 329710
rect 382260 329584 382330 329640
rect 382386 329584 382454 329640
rect 382510 329584 382578 329640
rect 382634 329584 382702 329640
rect 382758 329584 382880 329640
rect 382260 329516 382880 329584
rect 382260 329460 382330 329516
rect 382386 329460 382454 329516
rect 382510 329460 382578 329516
rect 382634 329460 382702 329516
rect 382758 329460 382880 329516
rect 382260 329392 382880 329460
rect 382260 329336 382330 329392
rect 382386 329336 382454 329392
rect 382510 329336 382578 329392
rect 382634 329336 382702 329392
rect 382758 329336 382880 329392
rect 382260 329268 382880 329336
rect 382260 329212 382330 329268
rect 382386 329212 382454 329268
rect 382510 329212 382578 329268
rect 382634 329212 382702 329268
rect 382758 329212 382880 329268
rect 382260 329144 382880 329212
rect 382260 329088 382330 329144
rect 382386 329088 382454 329144
rect 382510 329088 382578 329144
rect 382634 329088 382702 329144
rect 382758 329088 382880 329144
rect 382260 329020 382880 329088
rect 382260 328964 382330 329020
rect 382386 328964 382454 329020
rect 382510 328964 382578 329020
rect 382634 328964 382702 329020
rect 382758 328964 382880 329020
rect 382260 328896 382880 328964
rect 382260 328840 382330 328896
rect 382386 328840 382454 328896
rect 382510 328840 382578 328896
rect 382634 328840 382702 328896
rect 382758 328840 382880 328896
rect 382260 318426 382880 328840
rect 412006 329488 412626 334520
rect 430006 330888 430626 333560
rect 430006 330832 430207 330888
rect 430263 330832 430407 330888
rect 430463 330832 430626 330888
rect 430006 330588 430626 330832
rect 430006 330532 430207 330588
rect 430263 330532 430407 330588
rect 430463 330532 430626 330588
rect 430006 330288 430626 330532
rect 430006 330232 430207 330288
rect 430263 330232 430407 330288
rect 430463 330232 430626 330288
rect 430006 330110 430626 330232
rect 412006 329432 412207 329488
rect 412263 329432 412407 329488
rect 412463 329432 412626 329488
rect 412006 329188 412626 329432
rect 412006 329132 412207 329188
rect 412263 329132 412407 329188
rect 412463 329132 412626 329188
rect 412006 328888 412626 329132
rect 412006 328832 412207 328888
rect 412263 328832 412407 328888
rect 412463 328832 412626 328888
rect 412006 328710 412626 328832
rect 448006 329488 448626 334520
rect 466006 330888 466626 333560
rect 466006 330832 466207 330888
rect 466263 330832 466407 330888
rect 466463 330832 466626 330888
rect 466006 330588 466626 330832
rect 466006 330532 466207 330588
rect 466263 330532 466407 330588
rect 466463 330532 466626 330588
rect 466006 330288 466626 330532
rect 466006 330232 466207 330288
rect 466263 330232 466407 330288
rect 466463 330232 466626 330288
rect 466006 330110 466626 330232
rect 448006 329432 448207 329488
rect 448263 329432 448407 329488
rect 448463 329432 448626 329488
rect 448006 329188 448626 329432
rect 448006 329132 448207 329188
rect 448263 329132 448407 329188
rect 448463 329132 448626 329188
rect 448006 328888 448626 329132
rect 448006 328832 448207 328888
rect 448263 328832 448407 328888
rect 448463 328832 448626 328888
rect 448006 328710 448626 328832
rect 484006 329488 484626 334520
rect 502006 330888 502626 333560
rect 502006 330832 502207 330888
rect 502263 330832 502407 330888
rect 502463 330832 502626 330888
rect 502006 330588 502626 330832
rect 502006 330532 502207 330588
rect 502263 330532 502407 330588
rect 502463 330532 502626 330588
rect 502006 330288 502626 330532
rect 502006 330232 502207 330288
rect 502263 330232 502407 330288
rect 502463 330232 502626 330288
rect 502006 330110 502626 330232
rect 484006 329432 484207 329488
rect 484263 329432 484407 329488
rect 484463 329432 484626 329488
rect 484006 329188 484626 329432
rect 484006 329132 484207 329188
rect 484263 329132 484407 329188
rect 484463 329132 484626 329188
rect 484006 328888 484626 329132
rect 484006 328832 484207 328888
rect 484263 328832 484407 328888
rect 484463 328832 484626 328888
rect 484006 328710 484626 328832
rect 520006 329488 520626 334520
rect 538006 330888 538626 333560
rect 538006 330832 538207 330888
rect 538263 330832 538407 330888
rect 538463 330832 538626 330888
rect 538006 330588 538626 330832
rect 538006 330532 538207 330588
rect 538263 330532 538407 330588
rect 538463 330532 538626 330588
rect 538006 330288 538626 330532
rect 538006 330232 538207 330288
rect 538263 330232 538407 330288
rect 538463 330232 538626 330288
rect 538006 330110 538626 330232
rect 520006 329432 520207 329488
rect 520263 329432 520407 329488
rect 520463 329432 520626 329488
rect 520006 329188 520626 329432
rect 520006 329132 520207 329188
rect 520263 329132 520407 329188
rect 520463 329132 520626 329188
rect 520006 328888 520626 329132
rect 520006 328832 520207 328888
rect 520263 328832 520407 328888
rect 520463 328832 520626 328888
rect 520006 328710 520626 328832
rect 556006 329488 556626 334520
rect 574006 330888 574626 333560
rect 574006 330832 574207 330888
rect 574263 330832 574407 330888
rect 574463 330832 574626 330888
rect 574006 330588 574626 330832
rect 574006 330532 574207 330588
rect 574263 330532 574407 330588
rect 574463 330532 574626 330588
rect 574006 330288 574626 330532
rect 574006 330232 574207 330288
rect 574263 330232 574407 330288
rect 574463 330232 574626 330288
rect 574006 330110 574626 330232
rect 556006 329432 556207 329488
rect 556263 329432 556407 329488
rect 556463 329432 556626 329488
rect 556006 329188 556626 329432
rect 556006 329132 556207 329188
rect 556263 329132 556407 329188
rect 556463 329132 556626 329188
rect 556006 328888 556626 329132
rect 556006 328832 556207 328888
rect 556263 328832 556407 328888
rect 556463 328832 556626 328888
rect 556006 328710 556626 328832
rect 592006 329488 592626 334520
rect 610006 330888 610626 333560
rect 610006 330832 610207 330888
rect 610263 330832 610407 330888
rect 610463 330832 610626 330888
rect 610006 330588 610626 330832
rect 610006 330532 610207 330588
rect 610263 330532 610407 330588
rect 610463 330532 610626 330588
rect 610006 330288 610626 330532
rect 610006 330232 610207 330288
rect 610263 330232 610407 330288
rect 610463 330232 610626 330288
rect 610006 330110 610626 330232
rect 592006 329432 592207 329488
rect 592263 329432 592407 329488
rect 592463 329432 592626 329488
rect 592006 329188 592626 329432
rect 592006 329132 592207 329188
rect 592263 329132 592407 329188
rect 592463 329132 592626 329188
rect 592006 328888 592626 329132
rect 592006 328832 592207 328888
rect 592263 328832 592407 328888
rect 592463 328832 592626 328888
rect 592006 328710 592626 328832
rect 628006 329488 628626 334520
rect 646006 330888 646626 333560
rect 646006 330832 646207 330888
rect 646263 330832 646407 330888
rect 646463 330832 646626 330888
rect 646006 330588 646626 330832
rect 646006 330532 646207 330588
rect 646263 330532 646407 330588
rect 646463 330532 646626 330588
rect 646006 330288 646626 330532
rect 646006 330232 646207 330288
rect 646263 330232 646407 330288
rect 646463 330232 646626 330288
rect 646006 330110 646626 330232
rect 628006 329432 628207 329488
rect 628263 329432 628407 329488
rect 628463 329432 628626 329488
rect 628006 329188 628626 329432
rect 628006 329132 628207 329188
rect 628263 329132 628407 329188
rect 628463 329132 628626 329188
rect 628006 328888 628626 329132
rect 628006 328832 628207 328888
rect 628263 328832 628407 328888
rect 628463 328832 628626 328888
rect 628006 328710 628626 328832
rect 664006 329488 664626 334520
rect 682006 330888 682626 333560
rect 682006 330832 682207 330888
rect 682263 330832 682407 330888
rect 682463 330832 682626 330888
rect 682006 330588 682626 330832
rect 682006 330532 682207 330588
rect 682263 330532 682407 330588
rect 682463 330532 682626 330588
rect 682006 330288 682626 330532
rect 682006 330232 682207 330288
rect 682263 330232 682407 330288
rect 682463 330232 682626 330288
rect 682006 330110 682626 330232
rect 697922 333008 698922 349378
rect 697922 332952 698060 333008
rect 698116 332952 698360 333008
rect 698416 332952 698660 333008
rect 698716 332952 698922 333008
rect 697922 331040 698922 332952
rect 697922 330984 698052 331040
rect 698108 330984 698176 331040
rect 698232 330984 698300 331040
rect 698356 330984 698424 331040
rect 698480 330984 698548 331040
rect 698604 330984 698672 331040
rect 698728 330984 698796 331040
rect 698852 330984 698922 331040
rect 697922 330916 698922 330984
rect 697922 330860 698052 330916
rect 698108 330860 698176 330916
rect 698232 330860 698300 330916
rect 698356 330860 698424 330916
rect 698480 330860 698548 330916
rect 698604 330860 698672 330916
rect 698728 330860 698796 330916
rect 698852 330860 698922 330916
rect 697922 330792 698922 330860
rect 697922 330736 698052 330792
rect 698108 330736 698176 330792
rect 698232 330736 698300 330792
rect 698356 330736 698424 330792
rect 698480 330736 698548 330792
rect 698604 330736 698672 330792
rect 698728 330736 698796 330792
rect 698852 330736 698922 330792
rect 697922 330668 698922 330736
rect 697922 330612 698052 330668
rect 698108 330612 698176 330668
rect 698232 330612 698300 330668
rect 698356 330612 698424 330668
rect 698480 330612 698548 330668
rect 698604 330612 698672 330668
rect 698728 330612 698796 330668
rect 698852 330612 698922 330668
rect 697922 330544 698922 330612
rect 697922 330488 698052 330544
rect 698108 330488 698176 330544
rect 698232 330488 698300 330544
rect 698356 330488 698424 330544
rect 698480 330488 698548 330544
rect 698604 330488 698672 330544
rect 698728 330488 698796 330544
rect 698852 330488 698922 330544
rect 697922 330420 698922 330488
rect 697922 330364 698052 330420
rect 698108 330364 698176 330420
rect 698232 330364 698300 330420
rect 698356 330364 698424 330420
rect 698480 330364 698548 330420
rect 698604 330364 698672 330420
rect 698728 330364 698796 330420
rect 698852 330364 698922 330420
rect 697922 330296 698922 330364
rect 697922 330240 698052 330296
rect 698108 330240 698176 330296
rect 698232 330240 698300 330296
rect 698356 330240 698424 330296
rect 698480 330240 698548 330296
rect 698604 330240 698672 330296
rect 698728 330240 698796 330296
rect 698852 330240 698922 330296
rect 664006 329432 664207 329488
rect 664263 329432 664407 329488
rect 664463 329432 664626 329488
rect 664006 329188 664626 329432
rect 664006 329132 664207 329188
rect 664263 329132 664407 329188
rect 664463 329132 664626 329188
rect 664006 328888 664626 329132
rect 664006 328832 664207 328888
rect 664263 328832 664407 328888
rect 664463 328832 664626 328888
rect 664006 328710 664626 328832
rect 382260 318370 382402 318426
rect 382458 318370 382702 318426
rect 382758 318370 382880 318426
rect 382260 317028 382880 318370
rect 382260 316972 382402 317028
rect 382458 316972 382702 317028
rect 382758 316972 382880 317028
rect 382260 315630 382880 316972
rect 382260 315574 382402 315630
rect 382458 315574 382702 315630
rect 382758 315574 382880 315630
rect 382260 314232 382880 315574
rect 697922 320434 698922 330240
rect 697922 320378 698044 320434
rect 698100 320378 698344 320434
rect 698400 320378 698644 320434
rect 698700 320378 698922 320434
rect 382260 314176 382402 314232
rect 382458 314176 382702 314232
rect 382758 314176 382880 314232
rect 157088 305670 157158 305726
rect 157214 305670 157282 305726
rect 157338 305670 157406 305726
rect 157462 305670 157530 305726
rect 157586 305670 157708 305726
rect 157088 305602 157708 305670
rect 157088 305546 157158 305602
rect 157214 305546 157282 305602
rect 157338 305546 157406 305602
rect 157462 305546 157530 305602
rect 157586 305546 157708 305602
rect 157088 305478 157708 305546
rect 157088 305422 157158 305478
rect 157214 305422 157282 305478
rect 157338 305422 157406 305478
rect 157462 305422 157530 305478
rect 157586 305422 157708 305478
rect 157088 305354 157708 305422
rect 157088 305298 157158 305354
rect 157214 305298 157282 305354
rect 157338 305298 157406 305354
rect 157462 305298 157530 305354
rect 157586 305298 157708 305354
rect 157088 305230 157708 305298
rect 157088 305174 157158 305230
rect 157214 305174 157282 305230
rect 157338 305174 157406 305230
rect 157462 305174 157530 305230
rect 157586 305174 157708 305230
rect 157088 305106 157708 305174
rect 157088 305050 157158 305106
rect 157214 305050 157282 305106
rect 157338 305050 157406 305106
rect 157462 305050 157530 305106
rect 157586 305050 157708 305106
rect 157088 304982 157708 305050
rect 157088 304926 157158 304982
rect 157214 304926 157282 304982
rect 157338 304926 157406 304982
rect 157462 304926 157530 304982
rect 157586 304926 157708 304982
rect 157088 304856 157708 304926
rect 382260 305726 382880 314176
rect 382260 305670 382330 305726
rect 382386 305670 382454 305726
rect 382510 305670 382578 305726
rect 382634 305670 382702 305726
rect 382758 305670 382880 305726
rect 382260 305602 382880 305670
rect 382260 305546 382330 305602
rect 382386 305546 382454 305602
rect 382510 305546 382578 305602
rect 382634 305546 382702 305602
rect 382758 305546 382880 305602
rect 382260 305478 382880 305546
rect 382260 305422 382330 305478
rect 382386 305422 382454 305478
rect 382510 305422 382578 305478
rect 382634 305422 382702 305478
rect 382758 305422 382880 305478
rect 382260 305354 382880 305422
rect 382260 305298 382330 305354
rect 382386 305298 382454 305354
rect 382510 305298 382578 305354
rect 382634 305298 382702 305354
rect 382758 305298 382880 305354
rect 382260 305230 382880 305298
rect 382260 305174 382330 305230
rect 382386 305174 382454 305230
rect 382510 305174 382578 305230
rect 382634 305174 382702 305230
rect 382758 305174 382880 305230
rect 382260 305106 382880 305174
rect 382260 305050 382330 305106
rect 382386 305050 382454 305106
rect 382510 305050 382578 305106
rect 382634 305050 382702 305106
rect 382758 305050 382880 305106
rect 382260 304982 382880 305050
rect 382260 304926 382330 304982
rect 382386 304926 382454 304982
rect 382510 304926 382578 304982
rect 382634 304926 382702 304982
rect 382758 304926 382880 304982
rect 382260 304856 382880 304926
rect 388555 305786 388875 314284
rect 390150 307186 390470 314284
rect 390150 307130 390220 307186
rect 390276 307130 390344 307186
rect 390400 307130 390470 307186
rect 390150 307062 390470 307130
rect 390150 307006 390220 307062
rect 390276 307006 390344 307062
rect 390400 307006 390470 307062
rect 390150 306938 390470 307006
rect 390150 306882 390220 306938
rect 390276 306882 390344 306938
rect 390400 306882 390470 306938
rect 390150 306814 390470 306882
rect 390150 306758 390220 306814
rect 390276 306758 390344 306814
rect 390400 306758 390470 306814
rect 390150 306690 390470 306758
rect 390150 306634 390220 306690
rect 390276 306634 390344 306690
rect 390400 306634 390470 306690
rect 390150 306566 390470 306634
rect 390150 306510 390220 306566
rect 390276 306510 390344 306566
rect 390400 306510 390470 306566
rect 390150 306442 390470 306510
rect 390150 306386 390220 306442
rect 390276 306386 390344 306442
rect 390400 306386 390470 306442
rect 390150 306256 390470 306386
rect 388555 305730 388625 305786
rect 388681 305730 388749 305786
rect 388805 305730 388875 305786
rect 388555 305662 388875 305730
rect 388555 305606 388625 305662
rect 388681 305606 388749 305662
rect 388805 305606 388875 305662
rect 388555 305538 388875 305606
rect 388555 305482 388625 305538
rect 388681 305482 388749 305538
rect 388805 305482 388875 305538
rect 388555 305414 388875 305482
rect 388555 305358 388625 305414
rect 388681 305358 388749 305414
rect 388805 305358 388875 305414
rect 388555 305290 388875 305358
rect 388555 305234 388625 305290
rect 388681 305234 388749 305290
rect 388805 305234 388875 305290
rect 388555 305166 388875 305234
rect 388555 305110 388625 305166
rect 388681 305110 388749 305166
rect 388805 305110 388875 305166
rect 388555 305042 388875 305110
rect 388555 304986 388625 305042
rect 388681 304986 388749 305042
rect 388805 304986 388875 305042
rect 388555 304856 388875 304986
rect 391745 305786 392065 314284
rect 393340 307186 393660 314284
rect 393340 307130 393410 307186
rect 393466 307130 393534 307186
rect 393590 307130 393660 307186
rect 393340 307062 393660 307130
rect 393340 307006 393410 307062
rect 393466 307006 393534 307062
rect 393590 307006 393660 307062
rect 393340 306938 393660 307006
rect 393340 306882 393410 306938
rect 393466 306882 393534 306938
rect 393590 306882 393660 306938
rect 393340 306814 393660 306882
rect 393340 306758 393410 306814
rect 393466 306758 393534 306814
rect 393590 306758 393660 306814
rect 393340 306690 393660 306758
rect 393340 306634 393410 306690
rect 393466 306634 393534 306690
rect 393590 306634 393660 306690
rect 393340 306566 393660 306634
rect 393340 306510 393410 306566
rect 393466 306510 393534 306566
rect 393590 306510 393660 306566
rect 393340 306442 393660 306510
rect 393340 306386 393410 306442
rect 393466 306386 393534 306442
rect 393590 306386 393660 306442
rect 393340 306256 393660 306386
rect 391745 305730 391815 305786
rect 391871 305730 391939 305786
rect 391995 305730 392065 305786
rect 391745 305662 392065 305730
rect 391745 305606 391815 305662
rect 391871 305606 391939 305662
rect 391995 305606 392065 305662
rect 391745 305538 392065 305606
rect 391745 305482 391815 305538
rect 391871 305482 391939 305538
rect 391995 305482 392065 305538
rect 391745 305414 392065 305482
rect 391745 305358 391815 305414
rect 391871 305358 391939 305414
rect 391995 305358 392065 305414
rect 391745 305290 392065 305358
rect 391745 305234 391815 305290
rect 391871 305234 391939 305290
rect 391995 305234 392065 305290
rect 391745 305166 392065 305234
rect 391745 305110 391815 305166
rect 391871 305110 391939 305166
rect 391995 305110 392065 305166
rect 391745 305042 392065 305110
rect 391745 304986 391815 305042
rect 391871 304986 391939 305042
rect 391995 304986 392065 305042
rect 391745 304856 392065 304986
rect 394935 305786 395255 314284
rect 396530 307186 396850 314284
rect 396530 307130 396600 307186
rect 396656 307130 396724 307186
rect 396780 307130 396850 307186
rect 396530 307062 396850 307130
rect 396530 307006 396600 307062
rect 396656 307006 396724 307062
rect 396780 307006 396850 307062
rect 396530 306938 396850 307006
rect 396530 306882 396600 306938
rect 396656 306882 396724 306938
rect 396780 306882 396850 306938
rect 396530 306814 396850 306882
rect 396530 306758 396600 306814
rect 396656 306758 396724 306814
rect 396780 306758 396850 306814
rect 396530 306690 396850 306758
rect 396530 306634 396600 306690
rect 396656 306634 396724 306690
rect 396780 306634 396850 306690
rect 396530 306566 396850 306634
rect 396530 306510 396600 306566
rect 396656 306510 396724 306566
rect 396780 306510 396850 306566
rect 396530 306442 396850 306510
rect 396530 306386 396600 306442
rect 396656 306386 396724 306442
rect 396780 306386 396850 306442
rect 396530 306256 396850 306386
rect 394935 305730 395005 305786
rect 395061 305730 395129 305786
rect 395185 305730 395255 305786
rect 394935 305662 395255 305730
rect 394935 305606 395005 305662
rect 395061 305606 395129 305662
rect 395185 305606 395255 305662
rect 394935 305538 395255 305606
rect 394935 305482 395005 305538
rect 395061 305482 395129 305538
rect 395185 305482 395255 305538
rect 394935 305414 395255 305482
rect 394935 305358 395005 305414
rect 395061 305358 395129 305414
rect 395185 305358 395255 305414
rect 394935 305290 395255 305358
rect 394935 305234 395005 305290
rect 395061 305234 395129 305290
rect 395185 305234 395255 305290
rect 394935 305166 395255 305234
rect 394935 305110 395005 305166
rect 395061 305110 395129 305166
rect 395185 305110 395255 305166
rect 394935 305042 395255 305110
rect 394935 304986 395005 305042
rect 395061 304986 395129 305042
rect 395185 304986 395255 305042
rect 394935 304856 395255 304986
rect 398125 305786 398445 314284
rect 398125 305730 398195 305786
rect 398251 305730 398319 305786
rect 398375 305730 398445 305786
rect 398125 305662 398445 305730
rect 398125 305606 398195 305662
rect 398251 305606 398319 305662
rect 398375 305606 398445 305662
rect 398125 305538 398445 305606
rect 398125 305482 398195 305538
rect 398251 305482 398319 305538
rect 398375 305482 398445 305538
rect 398125 305414 398445 305482
rect 398125 305358 398195 305414
rect 398251 305358 398319 305414
rect 398375 305358 398445 305414
rect 398125 305290 398445 305358
rect 398125 305234 398195 305290
rect 398251 305234 398319 305290
rect 398375 305234 398445 305290
rect 398125 305166 398445 305234
rect 398125 305110 398195 305166
rect 398251 305110 398319 305166
rect 398375 305110 398445 305166
rect 398125 305042 398445 305110
rect 398125 304986 398195 305042
rect 398251 304986 398319 305042
rect 398375 304986 398445 305042
rect 398125 304856 398445 304986
rect 488555 305786 488875 314284
rect 490150 307186 490470 314284
rect 490150 307130 490220 307186
rect 490276 307130 490344 307186
rect 490400 307130 490470 307186
rect 490150 307062 490470 307130
rect 490150 307006 490220 307062
rect 490276 307006 490344 307062
rect 490400 307006 490470 307062
rect 490150 306938 490470 307006
rect 490150 306882 490220 306938
rect 490276 306882 490344 306938
rect 490400 306882 490470 306938
rect 490150 306814 490470 306882
rect 490150 306758 490220 306814
rect 490276 306758 490344 306814
rect 490400 306758 490470 306814
rect 490150 306690 490470 306758
rect 490150 306634 490220 306690
rect 490276 306634 490344 306690
rect 490400 306634 490470 306690
rect 490150 306566 490470 306634
rect 490150 306510 490220 306566
rect 490276 306510 490344 306566
rect 490400 306510 490470 306566
rect 490150 306442 490470 306510
rect 490150 306386 490220 306442
rect 490276 306386 490344 306442
rect 490400 306386 490470 306442
rect 490150 306256 490470 306386
rect 488555 305730 488625 305786
rect 488681 305730 488749 305786
rect 488805 305730 488875 305786
rect 488555 305662 488875 305730
rect 488555 305606 488625 305662
rect 488681 305606 488749 305662
rect 488805 305606 488875 305662
rect 488555 305538 488875 305606
rect 488555 305482 488625 305538
rect 488681 305482 488749 305538
rect 488805 305482 488875 305538
rect 488555 305414 488875 305482
rect 488555 305358 488625 305414
rect 488681 305358 488749 305414
rect 488805 305358 488875 305414
rect 488555 305290 488875 305358
rect 488555 305234 488625 305290
rect 488681 305234 488749 305290
rect 488805 305234 488875 305290
rect 488555 305166 488875 305234
rect 488555 305110 488625 305166
rect 488681 305110 488749 305166
rect 488805 305110 488875 305166
rect 488555 305042 488875 305110
rect 488555 304986 488625 305042
rect 488681 304986 488749 305042
rect 488805 304986 488875 305042
rect 488555 304856 488875 304986
rect 491745 305786 492065 314284
rect 493340 307186 493660 314284
rect 493340 307130 493410 307186
rect 493466 307130 493534 307186
rect 493590 307130 493660 307186
rect 493340 307062 493660 307130
rect 493340 307006 493410 307062
rect 493466 307006 493534 307062
rect 493590 307006 493660 307062
rect 493340 306938 493660 307006
rect 493340 306882 493410 306938
rect 493466 306882 493534 306938
rect 493590 306882 493660 306938
rect 493340 306814 493660 306882
rect 493340 306758 493410 306814
rect 493466 306758 493534 306814
rect 493590 306758 493660 306814
rect 493340 306690 493660 306758
rect 493340 306634 493410 306690
rect 493466 306634 493534 306690
rect 493590 306634 493660 306690
rect 493340 306566 493660 306634
rect 493340 306510 493410 306566
rect 493466 306510 493534 306566
rect 493590 306510 493660 306566
rect 493340 306442 493660 306510
rect 493340 306386 493410 306442
rect 493466 306386 493534 306442
rect 493590 306386 493660 306442
rect 493340 306256 493660 306386
rect 491745 305730 491815 305786
rect 491871 305730 491939 305786
rect 491995 305730 492065 305786
rect 491745 305662 492065 305730
rect 491745 305606 491815 305662
rect 491871 305606 491939 305662
rect 491995 305606 492065 305662
rect 491745 305538 492065 305606
rect 491745 305482 491815 305538
rect 491871 305482 491939 305538
rect 491995 305482 492065 305538
rect 491745 305414 492065 305482
rect 491745 305358 491815 305414
rect 491871 305358 491939 305414
rect 491995 305358 492065 305414
rect 491745 305290 492065 305358
rect 491745 305234 491815 305290
rect 491871 305234 491939 305290
rect 491995 305234 492065 305290
rect 491745 305166 492065 305234
rect 491745 305110 491815 305166
rect 491871 305110 491939 305166
rect 491995 305110 492065 305166
rect 491745 305042 492065 305110
rect 491745 304986 491815 305042
rect 491871 304986 491939 305042
rect 491995 304986 492065 305042
rect 491745 304856 492065 304986
rect 494935 305786 495255 314284
rect 496530 307186 496850 314284
rect 496530 307130 496600 307186
rect 496656 307130 496724 307186
rect 496780 307130 496850 307186
rect 496530 307062 496850 307130
rect 496530 307006 496600 307062
rect 496656 307006 496724 307062
rect 496780 307006 496850 307062
rect 496530 306938 496850 307006
rect 496530 306882 496600 306938
rect 496656 306882 496724 306938
rect 496780 306882 496850 306938
rect 496530 306814 496850 306882
rect 496530 306758 496600 306814
rect 496656 306758 496724 306814
rect 496780 306758 496850 306814
rect 496530 306690 496850 306758
rect 496530 306634 496600 306690
rect 496656 306634 496724 306690
rect 496780 306634 496850 306690
rect 496530 306566 496850 306634
rect 496530 306510 496600 306566
rect 496656 306510 496724 306566
rect 496780 306510 496850 306566
rect 496530 306442 496850 306510
rect 496530 306386 496600 306442
rect 496656 306386 496724 306442
rect 496780 306386 496850 306442
rect 496530 306256 496850 306386
rect 494935 305730 495005 305786
rect 495061 305730 495129 305786
rect 495185 305730 495255 305786
rect 494935 305662 495255 305730
rect 494935 305606 495005 305662
rect 495061 305606 495129 305662
rect 495185 305606 495255 305662
rect 494935 305538 495255 305606
rect 494935 305482 495005 305538
rect 495061 305482 495129 305538
rect 495185 305482 495255 305538
rect 494935 305414 495255 305482
rect 494935 305358 495005 305414
rect 495061 305358 495129 305414
rect 495185 305358 495255 305414
rect 494935 305290 495255 305358
rect 494935 305234 495005 305290
rect 495061 305234 495129 305290
rect 495185 305234 495255 305290
rect 494935 305166 495255 305234
rect 494935 305110 495005 305166
rect 495061 305110 495129 305166
rect 495185 305110 495255 305166
rect 494935 305042 495255 305110
rect 494935 304986 495005 305042
rect 495061 304986 495129 305042
rect 495185 304986 495255 305042
rect 494935 304856 495255 304986
rect 498125 305786 498445 314284
rect 498125 305730 498195 305786
rect 498251 305730 498319 305786
rect 498375 305730 498445 305786
rect 498125 305662 498445 305730
rect 498125 305606 498195 305662
rect 498251 305606 498319 305662
rect 498375 305606 498445 305662
rect 498125 305538 498445 305606
rect 498125 305482 498195 305538
rect 498251 305482 498319 305538
rect 498375 305482 498445 305538
rect 498125 305414 498445 305482
rect 498125 305358 498195 305414
rect 498251 305358 498319 305414
rect 498375 305358 498445 305414
rect 498125 305290 498445 305358
rect 498125 305234 498195 305290
rect 498251 305234 498319 305290
rect 498375 305234 498445 305290
rect 498125 305166 498445 305234
rect 498125 305110 498195 305166
rect 498251 305110 498319 305166
rect 498375 305110 498445 305166
rect 498125 305042 498445 305110
rect 498125 304986 498195 305042
rect 498251 304986 498319 305042
rect 498375 304986 498445 305042
rect 498125 304856 498445 304986
rect 590840 307126 591840 307256
rect 590840 307070 590910 307126
rect 590966 307070 591034 307126
rect 591090 307070 591158 307126
rect 591214 307070 591282 307126
rect 591338 307070 591406 307126
rect 591462 307070 591530 307126
rect 591586 307070 591654 307126
rect 591710 307070 591840 307126
rect 590840 307002 591840 307070
rect 590840 306946 590910 307002
rect 590966 306946 591034 307002
rect 591090 306946 591158 307002
rect 591214 306946 591282 307002
rect 591338 306946 591406 307002
rect 591462 306946 591530 307002
rect 591586 306946 591654 307002
rect 591710 306946 591840 307002
rect 590840 306878 591840 306946
rect 590840 306822 590910 306878
rect 590966 306822 591034 306878
rect 591090 306822 591158 306878
rect 591214 306822 591282 306878
rect 591338 306822 591406 306878
rect 591462 306822 591530 306878
rect 591586 306822 591654 306878
rect 591710 306822 591840 306878
rect 590840 306754 591840 306822
rect 590840 306698 590910 306754
rect 590966 306698 591034 306754
rect 591090 306698 591158 306754
rect 591214 306698 591282 306754
rect 591338 306698 591406 306754
rect 591462 306698 591530 306754
rect 591586 306698 591654 306754
rect 591710 306698 591840 306754
rect 590840 306630 591840 306698
rect 590840 306574 590910 306630
rect 590966 306574 591034 306630
rect 591090 306574 591158 306630
rect 591214 306574 591282 306630
rect 591338 306574 591406 306630
rect 591462 306574 591530 306630
rect 591586 306574 591654 306630
rect 591710 306574 591840 306630
rect 590840 306506 591840 306574
rect 590840 306450 590910 306506
rect 590966 306450 591034 306506
rect 591090 306450 591158 306506
rect 591214 306450 591282 306506
rect 591338 306450 591406 306506
rect 591462 306450 591530 306506
rect 591586 306450 591654 306506
rect 591710 306450 591840 306506
rect 590840 306382 591840 306450
rect 590840 306326 590910 306382
rect 590966 306326 591034 306382
rect 591090 306326 591158 306382
rect 591214 306326 591282 306382
rect 591338 306326 591406 306382
rect 591462 306326 591530 306382
rect 591586 306326 591654 306382
rect 591710 306326 591840 306382
rect 79078 300566 79300 300622
rect 79356 300566 79600 300622
rect 79656 300566 79900 300622
rect 79956 300566 80078 300622
rect 79078 290048 80078 300566
rect 79078 289992 79284 290048
rect 79340 289992 79584 290048
rect 79640 289992 79884 290048
rect 79940 289992 80078 290048
rect 79078 283372 80078 289992
rect 79078 283316 79208 283372
rect 79264 283316 79332 283372
rect 79388 283316 79456 283372
rect 79512 283316 79580 283372
rect 79636 283316 79704 283372
rect 79760 283316 79828 283372
rect 79884 283316 79952 283372
rect 80008 283316 80078 283372
rect 79078 283248 80078 283316
rect 79078 283192 79208 283248
rect 79264 283192 79332 283248
rect 79388 283192 79456 283248
rect 79512 283192 79580 283248
rect 79636 283192 79704 283248
rect 79760 283192 79828 283248
rect 79884 283192 79952 283248
rect 80008 283192 80078 283248
rect 79078 283124 80078 283192
rect 79078 283068 79208 283124
rect 79264 283068 79332 283124
rect 79388 283068 79456 283124
rect 79512 283068 79580 283124
rect 79636 283068 79704 283124
rect 79760 283068 79828 283124
rect 79884 283068 79952 283124
rect 80008 283068 80078 283124
rect 79078 283000 80078 283068
rect 79078 282944 79208 283000
rect 79264 282944 79332 283000
rect 79388 282944 79456 283000
rect 79512 282944 79580 283000
rect 79636 282944 79704 283000
rect 79760 282944 79828 283000
rect 79884 282944 79952 283000
rect 80008 282944 80078 283000
rect 79078 282876 80078 282944
rect 79078 282820 79208 282876
rect 79264 282820 79332 282876
rect 79388 282820 79456 282876
rect 79512 282820 79580 282876
rect 79636 282820 79704 282876
rect 79760 282820 79828 282876
rect 79884 282820 79952 282876
rect 80008 282820 80078 282876
rect 79078 282752 80078 282820
rect 79078 282696 79208 282752
rect 79264 282696 79332 282752
rect 79388 282696 79456 282752
rect 79512 282696 79580 282752
rect 79636 282696 79704 282752
rect 79760 282696 79828 282752
rect 79884 282696 79952 282752
rect 80008 282696 80078 282752
rect 79078 282628 80078 282696
rect 79078 282572 79208 282628
rect 79264 282572 79332 282628
rect 79388 282572 79456 282628
rect 79512 282572 79580 282628
rect 79636 282572 79704 282628
rect 79760 282572 79828 282628
rect 79884 282572 79952 282628
rect 80008 282572 80078 282628
rect 79078 273622 80078 282572
rect 99224 283312 99544 283442
rect 99224 283256 99294 283312
rect 99350 283256 99418 283312
rect 99474 283256 99544 283312
rect 99224 283188 99544 283256
rect 99224 283132 99294 283188
rect 99350 283132 99418 283188
rect 99474 283132 99544 283188
rect 99224 283064 99544 283132
rect 99224 283008 99294 283064
rect 99350 283008 99418 283064
rect 99474 283008 99544 283064
rect 99224 282940 99544 283008
rect 99224 282884 99294 282940
rect 99350 282884 99418 282940
rect 99474 282884 99544 282940
rect 99224 282816 99544 282884
rect 99224 282760 99294 282816
rect 99350 282760 99418 282816
rect 99474 282760 99544 282816
rect 99224 282692 99544 282760
rect 99224 282636 99294 282692
rect 99350 282636 99418 282692
rect 99474 282636 99544 282692
rect 99224 282568 99544 282636
rect 99224 282512 99294 282568
rect 99350 282512 99418 282568
rect 99474 282512 99544 282568
rect 94224 281912 94544 282042
rect 94224 281856 94294 281912
rect 94350 281856 94418 281912
rect 94474 281856 94544 281912
rect 94224 281788 94544 281856
rect 94224 281732 94294 281788
rect 94350 281732 94418 281788
rect 94474 281732 94544 281788
rect 94224 281664 94544 281732
rect 94224 281608 94294 281664
rect 94350 281608 94418 281664
rect 94474 281608 94544 281664
rect 94224 281540 94544 281608
rect 94224 281484 94294 281540
rect 94350 281484 94418 281540
rect 94474 281484 94544 281540
rect 94224 281416 94544 281484
rect 94224 281360 94294 281416
rect 94350 281360 94418 281416
rect 94474 281360 94544 281416
rect 94224 281292 94544 281360
rect 94224 281236 94294 281292
rect 94350 281236 94418 281292
rect 94474 281236 94544 281292
rect 94224 281168 94544 281236
rect 94224 281112 94294 281168
rect 94350 281112 94418 281168
rect 94474 281112 94544 281168
rect 94224 279368 94544 281112
rect 99224 279368 99544 282512
rect 109224 283312 109544 283442
rect 109224 283256 109294 283312
rect 109350 283256 109418 283312
rect 109474 283256 109544 283312
rect 109224 283188 109544 283256
rect 109224 283132 109294 283188
rect 109350 283132 109418 283188
rect 109474 283132 109544 283188
rect 109224 283064 109544 283132
rect 109224 283008 109294 283064
rect 109350 283008 109418 283064
rect 109474 283008 109544 283064
rect 109224 282940 109544 283008
rect 109224 282884 109294 282940
rect 109350 282884 109418 282940
rect 109474 282884 109544 282940
rect 109224 282816 109544 282884
rect 109224 282760 109294 282816
rect 109350 282760 109418 282816
rect 109474 282760 109544 282816
rect 109224 282692 109544 282760
rect 109224 282636 109294 282692
rect 109350 282636 109418 282692
rect 109474 282636 109544 282692
rect 109224 282568 109544 282636
rect 109224 282512 109294 282568
rect 109350 282512 109418 282568
rect 109474 282512 109544 282568
rect 104224 281912 104544 282042
rect 104224 281856 104294 281912
rect 104350 281856 104418 281912
rect 104474 281856 104544 281912
rect 104224 281788 104544 281856
rect 104224 281732 104294 281788
rect 104350 281732 104418 281788
rect 104474 281732 104544 281788
rect 104224 281664 104544 281732
rect 104224 281608 104294 281664
rect 104350 281608 104418 281664
rect 104474 281608 104544 281664
rect 104224 281540 104544 281608
rect 104224 281484 104294 281540
rect 104350 281484 104418 281540
rect 104474 281484 104544 281540
rect 104224 281416 104544 281484
rect 104224 281360 104294 281416
rect 104350 281360 104418 281416
rect 104474 281360 104544 281416
rect 104224 281292 104544 281360
rect 104224 281236 104294 281292
rect 104350 281236 104418 281292
rect 104474 281236 104544 281292
rect 104224 281168 104544 281236
rect 104224 281112 104294 281168
rect 104350 281112 104418 281168
rect 104474 281112 104544 281168
rect 104224 279368 104544 281112
rect 109224 279368 109544 282512
rect 119224 283312 119544 283442
rect 119224 283256 119294 283312
rect 119350 283256 119418 283312
rect 119474 283256 119544 283312
rect 119224 283188 119544 283256
rect 119224 283132 119294 283188
rect 119350 283132 119418 283188
rect 119474 283132 119544 283188
rect 119224 283064 119544 283132
rect 119224 283008 119294 283064
rect 119350 283008 119418 283064
rect 119474 283008 119544 283064
rect 119224 282940 119544 283008
rect 119224 282884 119294 282940
rect 119350 282884 119418 282940
rect 119474 282884 119544 282940
rect 119224 282816 119544 282884
rect 119224 282760 119294 282816
rect 119350 282760 119418 282816
rect 119474 282760 119544 282816
rect 119224 282692 119544 282760
rect 119224 282636 119294 282692
rect 119350 282636 119418 282692
rect 119474 282636 119544 282692
rect 119224 282568 119544 282636
rect 119224 282512 119294 282568
rect 119350 282512 119418 282568
rect 119474 282512 119544 282568
rect 114224 281912 114544 282042
rect 114224 281856 114294 281912
rect 114350 281856 114418 281912
rect 114474 281856 114544 281912
rect 114224 281788 114544 281856
rect 114224 281732 114294 281788
rect 114350 281732 114418 281788
rect 114474 281732 114544 281788
rect 114224 281664 114544 281732
rect 114224 281608 114294 281664
rect 114350 281608 114418 281664
rect 114474 281608 114544 281664
rect 114224 281540 114544 281608
rect 114224 281484 114294 281540
rect 114350 281484 114418 281540
rect 114474 281484 114544 281540
rect 114224 281416 114544 281484
rect 114224 281360 114294 281416
rect 114350 281360 114418 281416
rect 114474 281360 114544 281416
rect 114224 281292 114544 281360
rect 114224 281236 114294 281292
rect 114350 281236 114418 281292
rect 114474 281236 114544 281292
rect 114224 281168 114544 281236
rect 114224 281112 114294 281168
rect 114350 281112 114418 281168
rect 114474 281112 114544 281168
rect 114224 279368 114544 281112
rect 119224 279368 119544 282512
rect 129224 283312 129544 283442
rect 129224 283256 129294 283312
rect 129350 283256 129418 283312
rect 129474 283256 129544 283312
rect 129224 283188 129544 283256
rect 129224 283132 129294 283188
rect 129350 283132 129418 283188
rect 129474 283132 129544 283188
rect 129224 283064 129544 283132
rect 129224 283008 129294 283064
rect 129350 283008 129418 283064
rect 129474 283008 129544 283064
rect 129224 282940 129544 283008
rect 129224 282884 129294 282940
rect 129350 282884 129418 282940
rect 129474 282884 129544 282940
rect 129224 282816 129544 282884
rect 129224 282760 129294 282816
rect 129350 282760 129418 282816
rect 129474 282760 129544 282816
rect 129224 282692 129544 282760
rect 129224 282636 129294 282692
rect 129350 282636 129418 282692
rect 129474 282636 129544 282692
rect 129224 282568 129544 282636
rect 129224 282512 129294 282568
rect 129350 282512 129418 282568
rect 129474 282512 129544 282568
rect 124224 281912 124544 282042
rect 124224 281856 124294 281912
rect 124350 281856 124418 281912
rect 124474 281856 124544 281912
rect 124224 281788 124544 281856
rect 124224 281732 124294 281788
rect 124350 281732 124418 281788
rect 124474 281732 124544 281788
rect 124224 281664 124544 281732
rect 124224 281608 124294 281664
rect 124350 281608 124418 281664
rect 124474 281608 124544 281664
rect 124224 281540 124544 281608
rect 124224 281484 124294 281540
rect 124350 281484 124418 281540
rect 124474 281484 124544 281540
rect 124224 281416 124544 281484
rect 124224 281360 124294 281416
rect 124350 281360 124418 281416
rect 124474 281360 124544 281416
rect 124224 281292 124544 281360
rect 124224 281236 124294 281292
rect 124350 281236 124418 281292
rect 124474 281236 124544 281292
rect 124224 281168 124544 281236
rect 124224 281112 124294 281168
rect 124350 281112 124418 281168
rect 124474 281112 124544 281168
rect 124224 279368 124544 281112
rect 129224 279368 129544 282512
rect 139224 283312 139544 283442
rect 139224 283256 139294 283312
rect 139350 283256 139418 283312
rect 139474 283256 139544 283312
rect 139224 283188 139544 283256
rect 139224 283132 139294 283188
rect 139350 283132 139418 283188
rect 139474 283132 139544 283188
rect 139224 283064 139544 283132
rect 139224 283008 139294 283064
rect 139350 283008 139418 283064
rect 139474 283008 139544 283064
rect 139224 282940 139544 283008
rect 139224 282884 139294 282940
rect 139350 282884 139418 282940
rect 139474 282884 139544 282940
rect 139224 282816 139544 282884
rect 139224 282760 139294 282816
rect 139350 282760 139418 282816
rect 139474 282760 139544 282816
rect 139224 282692 139544 282760
rect 139224 282636 139294 282692
rect 139350 282636 139418 282692
rect 139474 282636 139544 282692
rect 139224 282568 139544 282636
rect 139224 282512 139294 282568
rect 139350 282512 139418 282568
rect 139474 282512 139544 282568
rect 134224 281912 134544 282042
rect 134224 281856 134294 281912
rect 134350 281856 134418 281912
rect 134474 281856 134544 281912
rect 134224 281788 134544 281856
rect 134224 281732 134294 281788
rect 134350 281732 134418 281788
rect 134474 281732 134544 281788
rect 134224 281664 134544 281732
rect 134224 281608 134294 281664
rect 134350 281608 134418 281664
rect 134474 281608 134544 281664
rect 134224 281540 134544 281608
rect 134224 281484 134294 281540
rect 134350 281484 134418 281540
rect 134474 281484 134544 281540
rect 134224 281416 134544 281484
rect 134224 281360 134294 281416
rect 134350 281360 134418 281416
rect 134474 281360 134544 281416
rect 134224 281292 134544 281360
rect 134224 281236 134294 281292
rect 134350 281236 134418 281292
rect 134474 281236 134544 281292
rect 134224 281168 134544 281236
rect 134224 281112 134294 281168
rect 134350 281112 134418 281168
rect 134474 281112 134544 281168
rect 134224 279368 134544 281112
rect 139224 279368 139544 282512
rect 149224 283312 149544 283442
rect 149224 283256 149294 283312
rect 149350 283256 149418 283312
rect 149474 283256 149544 283312
rect 149224 283188 149544 283256
rect 149224 283132 149294 283188
rect 149350 283132 149418 283188
rect 149474 283132 149544 283188
rect 149224 283064 149544 283132
rect 149224 283008 149294 283064
rect 149350 283008 149418 283064
rect 149474 283008 149544 283064
rect 149224 282940 149544 283008
rect 149224 282884 149294 282940
rect 149350 282884 149418 282940
rect 149474 282884 149544 282940
rect 149224 282816 149544 282884
rect 149224 282760 149294 282816
rect 149350 282760 149418 282816
rect 149474 282760 149544 282816
rect 149224 282692 149544 282760
rect 149224 282636 149294 282692
rect 149350 282636 149418 282692
rect 149474 282636 149544 282692
rect 149224 282568 149544 282636
rect 149224 282512 149294 282568
rect 149350 282512 149418 282568
rect 149474 282512 149544 282568
rect 144224 281912 144544 282042
rect 144224 281856 144294 281912
rect 144350 281856 144418 281912
rect 144474 281856 144544 281912
rect 144224 281788 144544 281856
rect 144224 281732 144294 281788
rect 144350 281732 144418 281788
rect 144474 281732 144544 281788
rect 144224 281664 144544 281732
rect 144224 281608 144294 281664
rect 144350 281608 144418 281664
rect 144474 281608 144544 281664
rect 144224 281540 144544 281608
rect 144224 281484 144294 281540
rect 144350 281484 144418 281540
rect 144474 281484 144544 281540
rect 144224 281416 144544 281484
rect 144224 281360 144294 281416
rect 144350 281360 144418 281416
rect 144474 281360 144544 281416
rect 144224 281292 144544 281360
rect 144224 281236 144294 281292
rect 144350 281236 144418 281292
rect 144474 281236 144544 281292
rect 144224 281168 144544 281236
rect 144224 281112 144294 281168
rect 144350 281112 144418 281168
rect 144474 281112 144544 281168
rect 144224 279368 144544 281112
rect 149224 279368 149544 282512
rect 159224 283312 159544 283442
rect 159224 283256 159294 283312
rect 159350 283256 159418 283312
rect 159474 283256 159544 283312
rect 159224 283188 159544 283256
rect 159224 283132 159294 283188
rect 159350 283132 159418 283188
rect 159474 283132 159544 283188
rect 159224 283064 159544 283132
rect 159224 283008 159294 283064
rect 159350 283008 159418 283064
rect 159474 283008 159544 283064
rect 159224 282940 159544 283008
rect 159224 282884 159294 282940
rect 159350 282884 159418 282940
rect 159474 282884 159544 282940
rect 159224 282816 159544 282884
rect 159224 282760 159294 282816
rect 159350 282760 159418 282816
rect 159474 282760 159544 282816
rect 159224 282692 159544 282760
rect 159224 282636 159294 282692
rect 159350 282636 159418 282692
rect 159474 282636 159544 282692
rect 159224 282568 159544 282636
rect 159224 282512 159294 282568
rect 159350 282512 159418 282568
rect 159474 282512 159544 282568
rect 154224 281912 154544 282042
rect 154224 281856 154294 281912
rect 154350 281856 154418 281912
rect 154474 281856 154544 281912
rect 154224 281788 154544 281856
rect 154224 281732 154294 281788
rect 154350 281732 154418 281788
rect 154474 281732 154544 281788
rect 154224 281664 154544 281732
rect 154224 281608 154294 281664
rect 154350 281608 154418 281664
rect 154474 281608 154544 281664
rect 154224 281540 154544 281608
rect 154224 281484 154294 281540
rect 154350 281484 154418 281540
rect 154474 281484 154544 281540
rect 154224 281416 154544 281484
rect 154224 281360 154294 281416
rect 154350 281360 154418 281416
rect 154474 281360 154544 281416
rect 154224 281292 154544 281360
rect 154224 281236 154294 281292
rect 154350 281236 154418 281292
rect 154474 281236 154544 281292
rect 154224 281168 154544 281236
rect 154224 281112 154294 281168
rect 154350 281112 154418 281168
rect 154474 281112 154544 281168
rect 154224 279368 154544 281112
rect 159224 279368 159544 282512
rect 169224 283312 169544 283442
rect 169224 283256 169294 283312
rect 169350 283256 169418 283312
rect 169474 283256 169544 283312
rect 169224 283188 169544 283256
rect 169224 283132 169294 283188
rect 169350 283132 169418 283188
rect 169474 283132 169544 283188
rect 169224 283064 169544 283132
rect 169224 283008 169294 283064
rect 169350 283008 169418 283064
rect 169474 283008 169544 283064
rect 169224 282940 169544 283008
rect 169224 282884 169294 282940
rect 169350 282884 169418 282940
rect 169474 282884 169544 282940
rect 169224 282816 169544 282884
rect 169224 282760 169294 282816
rect 169350 282760 169418 282816
rect 169474 282760 169544 282816
rect 169224 282692 169544 282760
rect 169224 282636 169294 282692
rect 169350 282636 169418 282692
rect 169474 282636 169544 282692
rect 169224 282568 169544 282636
rect 169224 282512 169294 282568
rect 169350 282512 169418 282568
rect 169474 282512 169544 282568
rect 164224 281912 164544 282042
rect 164224 281856 164294 281912
rect 164350 281856 164418 281912
rect 164474 281856 164544 281912
rect 164224 281788 164544 281856
rect 164224 281732 164294 281788
rect 164350 281732 164418 281788
rect 164474 281732 164544 281788
rect 164224 281664 164544 281732
rect 164224 281608 164294 281664
rect 164350 281608 164418 281664
rect 164474 281608 164544 281664
rect 164224 281540 164544 281608
rect 164224 281484 164294 281540
rect 164350 281484 164418 281540
rect 164474 281484 164544 281540
rect 164224 281416 164544 281484
rect 164224 281360 164294 281416
rect 164350 281360 164418 281416
rect 164474 281360 164544 281416
rect 164224 281292 164544 281360
rect 164224 281236 164294 281292
rect 164350 281236 164418 281292
rect 164474 281236 164544 281292
rect 164224 281168 164544 281236
rect 164224 281112 164294 281168
rect 164350 281112 164418 281168
rect 164474 281112 164544 281168
rect 164224 279368 164544 281112
rect 169224 279368 169544 282512
rect 179224 283312 179544 283442
rect 179224 283256 179294 283312
rect 179350 283256 179418 283312
rect 179474 283256 179544 283312
rect 179224 283188 179544 283256
rect 179224 283132 179294 283188
rect 179350 283132 179418 283188
rect 179474 283132 179544 283188
rect 179224 283064 179544 283132
rect 179224 283008 179294 283064
rect 179350 283008 179418 283064
rect 179474 283008 179544 283064
rect 179224 282940 179544 283008
rect 179224 282884 179294 282940
rect 179350 282884 179418 282940
rect 179474 282884 179544 282940
rect 179224 282816 179544 282884
rect 179224 282760 179294 282816
rect 179350 282760 179418 282816
rect 179474 282760 179544 282816
rect 179224 282692 179544 282760
rect 179224 282636 179294 282692
rect 179350 282636 179418 282692
rect 179474 282636 179544 282692
rect 179224 282568 179544 282636
rect 179224 282512 179294 282568
rect 179350 282512 179418 282568
rect 179474 282512 179544 282568
rect 174224 281912 174544 282042
rect 174224 281856 174294 281912
rect 174350 281856 174418 281912
rect 174474 281856 174544 281912
rect 174224 281788 174544 281856
rect 174224 281732 174294 281788
rect 174350 281732 174418 281788
rect 174474 281732 174544 281788
rect 174224 281664 174544 281732
rect 174224 281608 174294 281664
rect 174350 281608 174418 281664
rect 174474 281608 174544 281664
rect 174224 281540 174544 281608
rect 174224 281484 174294 281540
rect 174350 281484 174418 281540
rect 174474 281484 174544 281540
rect 174224 281416 174544 281484
rect 174224 281360 174294 281416
rect 174350 281360 174418 281416
rect 174474 281360 174544 281416
rect 174224 281292 174544 281360
rect 174224 281236 174294 281292
rect 174350 281236 174418 281292
rect 174474 281236 174544 281292
rect 174224 281168 174544 281236
rect 174224 281112 174294 281168
rect 174350 281112 174418 281168
rect 174474 281112 174544 281168
rect 174224 279368 174544 281112
rect 179224 279368 179544 282512
rect 189224 283312 189544 283442
rect 189224 283256 189294 283312
rect 189350 283256 189418 283312
rect 189474 283256 189544 283312
rect 189224 283188 189544 283256
rect 189224 283132 189294 283188
rect 189350 283132 189418 283188
rect 189474 283132 189544 283188
rect 189224 283064 189544 283132
rect 189224 283008 189294 283064
rect 189350 283008 189418 283064
rect 189474 283008 189544 283064
rect 189224 282940 189544 283008
rect 189224 282884 189294 282940
rect 189350 282884 189418 282940
rect 189474 282884 189544 282940
rect 189224 282816 189544 282884
rect 189224 282760 189294 282816
rect 189350 282760 189418 282816
rect 189474 282760 189544 282816
rect 189224 282692 189544 282760
rect 189224 282636 189294 282692
rect 189350 282636 189418 282692
rect 189474 282636 189544 282692
rect 189224 282568 189544 282636
rect 189224 282512 189294 282568
rect 189350 282512 189418 282568
rect 189474 282512 189544 282568
rect 184224 281912 184544 282042
rect 184224 281856 184294 281912
rect 184350 281856 184418 281912
rect 184474 281856 184544 281912
rect 184224 281788 184544 281856
rect 184224 281732 184294 281788
rect 184350 281732 184418 281788
rect 184474 281732 184544 281788
rect 184224 281664 184544 281732
rect 184224 281608 184294 281664
rect 184350 281608 184418 281664
rect 184474 281608 184544 281664
rect 184224 281540 184544 281608
rect 184224 281484 184294 281540
rect 184350 281484 184418 281540
rect 184474 281484 184544 281540
rect 184224 281416 184544 281484
rect 184224 281360 184294 281416
rect 184350 281360 184418 281416
rect 184474 281360 184544 281416
rect 184224 281292 184544 281360
rect 184224 281236 184294 281292
rect 184350 281236 184418 281292
rect 184474 281236 184544 281292
rect 184224 281168 184544 281236
rect 184224 281112 184294 281168
rect 184350 281112 184418 281168
rect 184474 281112 184544 281168
rect 184224 279368 184544 281112
rect 189224 279368 189544 282512
rect 199224 283312 199544 283442
rect 199224 283256 199294 283312
rect 199350 283256 199418 283312
rect 199474 283256 199544 283312
rect 199224 283188 199544 283256
rect 199224 283132 199294 283188
rect 199350 283132 199418 283188
rect 199474 283132 199544 283188
rect 199224 283064 199544 283132
rect 199224 283008 199294 283064
rect 199350 283008 199418 283064
rect 199474 283008 199544 283064
rect 199224 282940 199544 283008
rect 199224 282884 199294 282940
rect 199350 282884 199418 282940
rect 199474 282884 199544 282940
rect 199224 282816 199544 282884
rect 199224 282760 199294 282816
rect 199350 282760 199418 282816
rect 199474 282760 199544 282816
rect 199224 282692 199544 282760
rect 199224 282636 199294 282692
rect 199350 282636 199418 282692
rect 199474 282636 199544 282692
rect 199224 282568 199544 282636
rect 199224 282512 199294 282568
rect 199350 282512 199418 282568
rect 199474 282512 199544 282568
rect 194224 281912 194544 282042
rect 194224 281856 194294 281912
rect 194350 281856 194418 281912
rect 194474 281856 194544 281912
rect 194224 281788 194544 281856
rect 194224 281732 194294 281788
rect 194350 281732 194418 281788
rect 194474 281732 194544 281788
rect 194224 281664 194544 281732
rect 194224 281608 194294 281664
rect 194350 281608 194418 281664
rect 194474 281608 194544 281664
rect 194224 281540 194544 281608
rect 194224 281484 194294 281540
rect 194350 281484 194418 281540
rect 194474 281484 194544 281540
rect 194224 281416 194544 281484
rect 194224 281360 194294 281416
rect 194350 281360 194418 281416
rect 194474 281360 194544 281416
rect 194224 281292 194544 281360
rect 194224 281236 194294 281292
rect 194350 281236 194418 281292
rect 194474 281236 194544 281292
rect 194224 281168 194544 281236
rect 194224 281112 194294 281168
rect 194350 281112 194418 281168
rect 194474 281112 194544 281168
rect 194224 279368 194544 281112
rect 199224 279368 199544 282512
rect 209224 283312 209544 283442
rect 209224 283256 209294 283312
rect 209350 283256 209418 283312
rect 209474 283256 209544 283312
rect 209224 283188 209544 283256
rect 209224 283132 209294 283188
rect 209350 283132 209418 283188
rect 209474 283132 209544 283188
rect 209224 283064 209544 283132
rect 209224 283008 209294 283064
rect 209350 283008 209418 283064
rect 209474 283008 209544 283064
rect 209224 282940 209544 283008
rect 209224 282884 209294 282940
rect 209350 282884 209418 282940
rect 209474 282884 209544 282940
rect 209224 282816 209544 282884
rect 209224 282760 209294 282816
rect 209350 282760 209418 282816
rect 209474 282760 209544 282816
rect 209224 282692 209544 282760
rect 209224 282636 209294 282692
rect 209350 282636 209418 282692
rect 209474 282636 209544 282692
rect 209224 282568 209544 282636
rect 209224 282512 209294 282568
rect 209350 282512 209418 282568
rect 209474 282512 209544 282568
rect 204224 281912 204544 282042
rect 204224 281856 204294 281912
rect 204350 281856 204418 281912
rect 204474 281856 204544 281912
rect 204224 281788 204544 281856
rect 204224 281732 204294 281788
rect 204350 281732 204418 281788
rect 204474 281732 204544 281788
rect 204224 281664 204544 281732
rect 204224 281608 204294 281664
rect 204350 281608 204418 281664
rect 204474 281608 204544 281664
rect 204224 281540 204544 281608
rect 204224 281484 204294 281540
rect 204350 281484 204418 281540
rect 204474 281484 204544 281540
rect 204224 281416 204544 281484
rect 204224 281360 204294 281416
rect 204350 281360 204418 281416
rect 204474 281360 204544 281416
rect 204224 281292 204544 281360
rect 204224 281236 204294 281292
rect 204350 281236 204418 281292
rect 204474 281236 204544 281292
rect 204224 281168 204544 281236
rect 204224 281112 204294 281168
rect 204350 281112 204418 281168
rect 204474 281112 204544 281168
rect 204224 279368 204544 281112
rect 209224 279368 209544 282512
rect 219224 283312 219544 283442
rect 219224 283256 219294 283312
rect 219350 283256 219418 283312
rect 219474 283256 219544 283312
rect 219224 283188 219544 283256
rect 219224 283132 219294 283188
rect 219350 283132 219418 283188
rect 219474 283132 219544 283188
rect 219224 283064 219544 283132
rect 219224 283008 219294 283064
rect 219350 283008 219418 283064
rect 219474 283008 219544 283064
rect 219224 282940 219544 283008
rect 219224 282884 219294 282940
rect 219350 282884 219418 282940
rect 219474 282884 219544 282940
rect 219224 282816 219544 282884
rect 219224 282760 219294 282816
rect 219350 282760 219418 282816
rect 219474 282760 219544 282816
rect 219224 282692 219544 282760
rect 219224 282636 219294 282692
rect 219350 282636 219418 282692
rect 219474 282636 219544 282692
rect 219224 282568 219544 282636
rect 219224 282512 219294 282568
rect 219350 282512 219418 282568
rect 219474 282512 219544 282568
rect 214224 281912 214544 282042
rect 214224 281856 214294 281912
rect 214350 281856 214418 281912
rect 214474 281856 214544 281912
rect 214224 281788 214544 281856
rect 214224 281732 214294 281788
rect 214350 281732 214418 281788
rect 214474 281732 214544 281788
rect 214224 281664 214544 281732
rect 214224 281608 214294 281664
rect 214350 281608 214418 281664
rect 214474 281608 214544 281664
rect 214224 281540 214544 281608
rect 214224 281484 214294 281540
rect 214350 281484 214418 281540
rect 214474 281484 214544 281540
rect 214224 281416 214544 281484
rect 214224 281360 214294 281416
rect 214350 281360 214418 281416
rect 214474 281360 214544 281416
rect 214224 281292 214544 281360
rect 214224 281236 214294 281292
rect 214350 281236 214418 281292
rect 214474 281236 214544 281292
rect 214224 281168 214544 281236
rect 214224 281112 214294 281168
rect 214350 281112 214418 281168
rect 214474 281112 214544 281168
rect 214224 279368 214544 281112
rect 219224 279368 219544 282512
rect 229224 283312 229544 283442
rect 229224 283256 229294 283312
rect 229350 283256 229418 283312
rect 229474 283256 229544 283312
rect 229224 283188 229544 283256
rect 229224 283132 229294 283188
rect 229350 283132 229418 283188
rect 229474 283132 229544 283188
rect 229224 283064 229544 283132
rect 229224 283008 229294 283064
rect 229350 283008 229418 283064
rect 229474 283008 229544 283064
rect 229224 282940 229544 283008
rect 229224 282884 229294 282940
rect 229350 282884 229418 282940
rect 229474 282884 229544 282940
rect 229224 282816 229544 282884
rect 229224 282760 229294 282816
rect 229350 282760 229418 282816
rect 229474 282760 229544 282816
rect 229224 282692 229544 282760
rect 229224 282636 229294 282692
rect 229350 282636 229418 282692
rect 229474 282636 229544 282692
rect 229224 282568 229544 282636
rect 229224 282512 229294 282568
rect 229350 282512 229418 282568
rect 229474 282512 229544 282568
rect 224224 281912 224544 282042
rect 224224 281856 224294 281912
rect 224350 281856 224418 281912
rect 224474 281856 224544 281912
rect 224224 281788 224544 281856
rect 224224 281732 224294 281788
rect 224350 281732 224418 281788
rect 224474 281732 224544 281788
rect 224224 281664 224544 281732
rect 224224 281608 224294 281664
rect 224350 281608 224418 281664
rect 224474 281608 224544 281664
rect 224224 281540 224544 281608
rect 224224 281484 224294 281540
rect 224350 281484 224418 281540
rect 224474 281484 224544 281540
rect 224224 281416 224544 281484
rect 224224 281360 224294 281416
rect 224350 281360 224418 281416
rect 224474 281360 224544 281416
rect 224224 281292 224544 281360
rect 224224 281236 224294 281292
rect 224350 281236 224418 281292
rect 224474 281236 224544 281292
rect 224224 281168 224544 281236
rect 224224 281112 224294 281168
rect 224350 281112 224418 281168
rect 224474 281112 224544 281168
rect 224224 279368 224544 281112
rect 229224 279368 229544 282512
rect 239224 283312 239544 283442
rect 239224 283256 239294 283312
rect 239350 283256 239418 283312
rect 239474 283256 239544 283312
rect 239224 283188 239544 283256
rect 239224 283132 239294 283188
rect 239350 283132 239418 283188
rect 239474 283132 239544 283188
rect 239224 283064 239544 283132
rect 239224 283008 239294 283064
rect 239350 283008 239418 283064
rect 239474 283008 239544 283064
rect 239224 282940 239544 283008
rect 239224 282884 239294 282940
rect 239350 282884 239418 282940
rect 239474 282884 239544 282940
rect 239224 282816 239544 282884
rect 239224 282760 239294 282816
rect 239350 282760 239418 282816
rect 239474 282760 239544 282816
rect 239224 282692 239544 282760
rect 239224 282636 239294 282692
rect 239350 282636 239418 282692
rect 239474 282636 239544 282692
rect 239224 282568 239544 282636
rect 239224 282512 239294 282568
rect 239350 282512 239418 282568
rect 239474 282512 239544 282568
rect 234224 281912 234544 282042
rect 234224 281856 234294 281912
rect 234350 281856 234418 281912
rect 234474 281856 234544 281912
rect 234224 281788 234544 281856
rect 234224 281732 234294 281788
rect 234350 281732 234418 281788
rect 234474 281732 234544 281788
rect 234224 281664 234544 281732
rect 234224 281608 234294 281664
rect 234350 281608 234418 281664
rect 234474 281608 234544 281664
rect 234224 281540 234544 281608
rect 234224 281484 234294 281540
rect 234350 281484 234418 281540
rect 234474 281484 234544 281540
rect 234224 281416 234544 281484
rect 234224 281360 234294 281416
rect 234350 281360 234418 281416
rect 234474 281360 234544 281416
rect 234224 281292 234544 281360
rect 234224 281236 234294 281292
rect 234350 281236 234418 281292
rect 234474 281236 234544 281292
rect 234224 281168 234544 281236
rect 234224 281112 234294 281168
rect 234350 281112 234418 281168
rect 234474 281112 234544 281168
rect 234224 279368 234544 281112
rect 239224 279368 239544 282512
rect 249224 283312 249544 283442
rect 249224 283256 249294 283312
rect 249350 283256 249418 283312
rect 249474 283256 249544 283312
rect 249224 283188 249544 283256
rect 249224 283132 249294 283188
rect 249350 283132 249418 283188
rect 249474 283132 249544 283188
rect 249224 283064 249544 283132
rect 249224 283008 249294 283064
rect 249350 283008 249418 283064
rect 249474 283008 249544 283064
rect 249224 282940 249544 283008
rect 249224 282884 249294 282940
rect 249350 282884 249418 282940
rect 249474 282884 249544 282940
rect 249224 282816 249544 282884
rect 249224 282760 249294 282816
rect 249350 282760 249418 282816
rect 249474 282760 249544 282816
rect 249224 282692 249544 282760
rect 249224 282636 249294 282692
rect 249350 282636 249418 282692
rect 249474 282636 249544 282692
rect 249224 282568 249544 282636
rect 249224 282512 249294 282568
rect 249350 282512 249418 282568
rect 249474 282512 249544 282568
rect 244224 281912 244544 282042
rect 244224 281856 244294 281912
rect 244350 281856 244418 281912
rect 244474 281856 244544 281912
rect 244224 281788 244544 281856
rect 244224 281732 244294 281788
rect 244350 281732 244418 281788
rect 244474 281732 244544 281788
rect 244224 281664 244544 281732
rect 244224 281608 244294 281664
rect 244350 281608 244418 281664
rect 244474 281608 244544 281664
rect 244224 281540 244544 281608
rect 244224 281484 244294 281540
rect 244350 281484 244418 281540
rect 244474 281484 244544 281540
rect 244224 281416 244544 281484
rect 244224 281360 244294 281416
rect 244350 281360 244418 281416
rect 244474 281360 244544 281416
rect 244224 281292 244544 281360
rect 244224 281236 244294 281292
rect 244350 281236 244418 281292
rect 244474 281236 244544 281292
rect 244224 281168 244544 281236
rect 244224 281112 244294 281168
rect 244350 281112 244418 281168
rect 244474 281112 244544 281168
rect 244224 279368 244544 281112
rect 249224 279368 249544 282512
rect 259224 283312 259544 283442
rect 259224 283256 259294 283312
rect 259350 283256 259418 283312
rect 259474 283256 259544 283312
rect 259224 283188 259544 283256
rect 259224 283132 259294 283188
rect 259350 283132 259418 283188
rect 259474 283132 259544 283188
rect 259224 283064 259544 283132
rect 259224 283008 259294 283064
rect 259350 283008 259418 283064
rect 259474 283008 259544 283064
rect 259224 282940 259544 283008
rect 259224 282884 259294 282940
rect 259350 282884 259418 282940
rect 259474 282884 259544 282940
rect 259224 282816 259544 282884
rect 259224 282760 259294 282816
rect 259350 282760 259418 282816
rect 259474 282760 259544 282816
rect 259224 282692 259544 282760
rect 259224 282636 259294 282692
rect 259350 282636 259418 282692
rect 259474 282636 259544 282692
rect 259224 282568 259544 282636
rect 259224 282512 259294 282568
rect 259350 282512 259418 282568
rect 259474 282512 259544 282568
rect 254224 281912 254544 282042
rect 254224 281856 254294 281912
rect 254350 281856 254418 281912
rect 254474 281856 254544 281912
rect 254224 281788 254544 281856
rect 254224 281732 254294 281788
rect 254350 281732 254418 281788
rect 254474 281732 254544 281788
rect 254224 281664 254544 281732
rect 254224 281608 254294 281664
rect 254350 281608 254418 281664
rect 254474 281608 254544 281664
rect 254224 281540 254544 281608
rect 254224 281484 254294 281540
rect 254350 281484 254418 281540
rect 254474 281484 254544 281540
rect 254224 281416 254544 281484
rect 254224 281360 254294 281416
rect 254350 281360 254418 281416
rect 254474 281360 254544 281416
rect 254224 281292 254544 281360
rect 254224 281236 254294 281292
rect 254350 281236 254418 281292
rect 254474 281236 254544 281292
rect 254224 281168 254544 281236
rect 254224 281112 254294 281168
rect 254350 281112 254418 281168
rect 254474 281112 254544 281168
rect 254224 279368 254544 281112
rect 259224 279368 259544 282512
rect 269224 283312 269544 283442
rect 269224 283256 269294 283312
rect 269350 283256 269418 283312
rect 269474 283256 269544 283312
rect 269224 283188 269544 283256
rect 269224 283132 269294 283188
rect 269350 283132 269418 283188
rect 269474 283132 269544 283188
rect 269224 283064 269544 283132
rect 269224 283008 269294 283064
rect 269350 283008 269418 283064
rect 269474 283008 269544 283064
rect 269224 282940 269544 283008
rect 269224 282884 269294 282940
rect 269350 282884 269418 282940
rect 269474 282884 269544 282940
rect 269224 282816 269544 282884
rect 269224 282760 269294 282816
rect 269350 282760 269418 282816
rect 269474 282760 269544 282816
rect 269224 282692 269544 282760
rect 269224 282636 269294 282692
rect 269350 282636 269418 282692
rect 269474 282636 269544 282692
rect 269224 282568 269544 282636
rect 269224 282512 269294 282568
rect 269350 282512 269418 282568
rect 269474 282512 269544 282568
rect 264224 281912 264544 282042
rect 264224 281856 264294 281912
rect 264350 281856 264418 281912
rect 264474 281856 264544 281912
rect 264224 281788 264544 281856
rect 264224 281732 264294 281788
rect 264350 281732 264418 281788
rect 264474 281732 264544 281788
rect 264224 281664 264544 281732
rect 264224 281608 264294 281664
rect 264350 281608 264418 281664
rect 264474 281608 264544 281664
rect 264224 281540 264544 281608
rect 264224 281484 264294 281540
rect 264350 281484 264418 281540
rect 264474 281484 264544 281540
rect 264224 281416 264544 281484
rect 264224 281360 264294 281416
rect 264350 281360 264418 281416
rect 264474 281360 264544 281416
rect 264224 281292 264544 281360
rect 264224 281236 264294 281292
rect 264350 281236 264418 281292
rect 264474 281236 264544 281292
rect 264224 281168 264544 281236
rect 264224 281112 264294 281168
rect 264350 281112 264418 281168
rect 264474 281112 264544 281168
rect 264224 279368 264544 281112
rect 269224 279368 269544 282512
rect 279224 283312 279544 283442
rect 279224 283256 279294 283312
rect 279350 283256 279418 283312
rect 279474 283256 279544 283312
rect 279224 283188 279544 283256
rect 279224 283132 279294 283188
rect 279350 283132 279418 283188
rect 279474 283132 279544 283188
rect 279224 283064 279544 283132
rect 279224 283008 279294 283064
rect 279350 283008 279418 283064
rect 279474 283008 279544 283064
rect 279224 282940 279544 283008
rect 279224 282884 279294 282940
rect 279350 282884 279418 282940
rect 279474 282884 279544 282940
rect 279224 282816 279544 282884
rect 279224 282760 279294 282816
rect 279350 282760 279418 282816
rect 279474 282760 279544 282816
rect 279224 282692 279544 282760
rect 279224 282636 279294 282692
rect 279350 282636 279418 282692
rect 279474 282636 279544 282692
rect 279224 282568 279544 282636
rect 279224 282512 279294 282568
rect 279350 282512 279418 282568
rect 279474 282512 279544 282568
rect 274224 281912 274544 282042
rect 274224 281856 274294 281912
rect 274350 281856 274418 281912
rect 274474 281856 274544 281912
rect 274224 281788 274544 281856
rect 274224 281732 274294 281788
rect 274350 281732 274418 281788
rect 274474 281732 274544 281788
rect 274224 281664 274544 281732
rect 274224 281608 274294 281664
rect 274350 281608 274418 281664
rect 274474 281608 274544 281664
rect 274224 281540 274544 281608
rect 274224 281484 274294 281540
rect 274350 281484 274418 281540
rect 274474 281484 274544 281540
rect 274224 281416 274544 281484
rect 274224 281360 274294 281416
rect 274350 281360 274418 281416
rect 274474 281360 274544 281416
rect 274224 281292 274544 281360
rect 274224 281236 274294 281292
rect 274350 281236 274418 281292
rect 274474 281236 274544 281292
rect 274224 281168 274544 281236
rect 274224 281112 274294 281168
rect 274350 281112 274418 281168
rect 274474 281112 274544 281168
rect 274224 279368 274544 281112
rect 279224 279368 279544 282512
rect 289224 283312 289544 283442
rect 289224 283256 289294 283312
rect 289350 283256 289418 283312
rect 289474 283256 289544 283312
rect 289224 283188 289544 283256
rect 289224 283132 289294 283188
rect 289350 283132 289418 283188
rect 289474 283132 289544 283188
rect 289224 283064 289544 283132
rect 289224 283008 289294 283064
rect 289350 283008 289418 283064
rect 289474 283008 289544 283064
rect 289224 282940 289544 283008
rect 289224 282884 289294 282940
rect 289350 282884 289418 282940
rect 289474 282884 289544 282940
rect 289224 282816 289544 282884
rect 289224 282760 289294 282816
rect 289350 282760 289418 282816
rect 289474 282760 289544 282816
rect 289224 282692 289544 282760
rect 289224 282636 289294 282692
rect 289350 282636 289418 282692
rect 289474 282636 289544 282692
rect 289224 282568 289544 282636
rect 289224 282512 289294 282568
rect 289350 282512 289418 282568
rect 289474 282512 289544 282568
rect 284224 281912 284544 282042
rect 284224 281856 284294 281912
rect 284350 281856 284418 281912
rect 284474 281856 284544 281912
rect 284224 281788 284544 281856
rect 284224 281732 284294 281788
rect 284350 281732 284418 281788
rect 284474 281732 284544 281788
rect 284224 281664 284544 281732
rect 284224 281608 284294 281664
rect 284350 281608 284418 281664
rect 284474 281608 284544 281664
rect 284224 281540 284544 281608
rect 284224 281484 284294 281540
rect 284350 281484 284418 281540
rect 284474 281484 284544 281540
rect 284224 281416 284544 281484
rect 284224 281360 284294 281416
rect 284350 281360 284418 281416
rect 284474 281360 284544 281416
rect 284224 281292 284544 281360
rect 284224 281236 284294 281292
rect 284350 281236 284418 281292
rect 284474 281236 284544 281292
rect 284224 281168 284544 281236
rect 284224 281112 284294 281168
rect 284350 281112 284418 281168
rect 284474 281112 284544 281168
rect 284224 279368 284544 281112
rect 289224 279368 289544 282512
rect 299224 283312 299544 283442
rect 299224 283256 299294 283312
rect 299350 283256 299418 283312
rect 299474 283256 299544 283312
rect 299224 283188 299544 283256
rect 299224 283132 299294 283188
rect 299350 283132 299418 283188
rect 299474 283132 299544 283188
rect 299224 283064 299544 283132
rect 299224 283008 299294 283064
rect 299350 283008 299418 283064
rect 299474 283008 299544 283064
rect 299224 282940 299544 283008
rect 299224 282884 299294 282940
rect 299350 282884 299418 282940
rect 299474 282884 299544 282940
rect 299224 282816 299544 282884
rect 299224 282760 299294 282816
rect 299350 282760 299418 282816
rect 299474 282760 299544 282816
rect 299224 282692 299544 282760
rect 299224 282636 299294 282692
rect 299350 282636 299418 282692
rect 299474 282636 299544 282692
rect 299224 282568 299544 282636
rect 299224 282512 299294 282568
rect 299350 282512 299418 282568
rect 299474 282512 299544 282568
rect 294224 281912 294544 282042
rect 294224 281856 294294 281912
rect 294350 281856 294418 281912
rect 294474 281856 294544 281912
rect 294224 281788 294544 281856
rect 294224 281732 294294 281788
rect 294350 281732 294418 281788
rect 294474 281732 294544 281788
rect 294224 281664 294544 281732
rect 294224 281608 294294 281664
rect 294350 281608 294418 281664
rect 294474 281608 294544 281664
rect 294224 281540 294544 281608
rect 294224 281484 294294 281540
rect 294350 281484 294418 281540
rect 294474 281484 294544 281540
rect 294224 281416 294544 281484
rect 294224 281360 294294 281416
rect 294350 281360 294418 281416
rect 294474 281360 294544 281416
rect 294224 281292 294544 281360
rect 294224 281236 294294 281292
rect 294350 281236 294418 281292
rect 294474 281236 294544 281292
rect 294224 281168 294544 281236
rect 294224 281112 294294 281168
rect 294350 281112 294418 281168
rect 294474 281112 294544 281168
rect 294224 279368 294544 281112
rect 299224 279368 299544 282512
rect 309224 283312 309544 283442
rect 309224 283256 309294 283312
rect 309350 283256 309418 283312
rect 309474 283256 309544 283312
rect 309224 283188 309544 283256
rect 309224 283132 309294 283188
rect 309350 283132 309418 283188
rect 309474 283132 309544 283188
rect 309224 283064 309544 283132
rect 309224 283008 309294 283064
rect 309350 283008 309418 283064
rect 309474 283008 309544 283064
rect 309224 282940 309544 283008
rect 309224 282884 309294 282940
rect 309350 282884 309418 282940
rect 309474 282884 309544 282940
rect 309224 282816 309544 282884
rect 309224 282760 309294 282816
rect 309350 282760 309418 282816
rect 309474 282760 309544 282816
rect 309224 282692 309544 282760
rect 309224 282636 309294 282692
rect 309350 282636 309418 282692
rect 309474 282636 309544 282692
rect 309224 282568 309544 282636
rect 309224 282512 309294 282568
rect 309350 282512 309418 282568
rect 309474 282512 309544 282568
rect 304224 281912 304544 282042
rect 304224 281856 304294 281912
rect 304350 281856 304418 281912
rect 304474 281856 304544 281912
rect 304224 281788 304544 281856
rect 304224 281732 304294 281788
rect 304350 281732 304418 281788
rect 304474 281732 304544 281788
rect 304224 281664 304544 281732
rect 304224 281608 304294 281664
rect 304350 281608 304418 281664
rect 304474 281608 304544 281664
rect 304224 281540 304544 281608
rect 304224 281484 304294 281540
rect 304350 281484 304418 281540
rect 304474 281484 304544 281540
rect 304224 281416 304544 281484
rect 304224 281360 304294 281416
rect 304350 281360 304418 281416
rect 304474 281360 304544 281416
rect 304224 281292 304544 281360
rect 304224 281236 304294 281292
rect 304350 281236 304418 281292
rect 304474 281236 304544 281292
rect 304224 281168 304544 281236
rect 304224 281112 304294 281168
rect 304350 281112 304418 281168
rect 304474 281112 304544 281168
rect 304224 279368 304544 281112
rect 309224 279368 309544 282512
rect 319224 283312 319544 283442
rect 319224 283256 319294 283312
rect 319350 283256 319418 283312
rect 319474 283256 319544 283312
rect 319224 283188 319544 283256
rect 319224 283132 319294 283188
rect 319350 283132 319418 283188
rect 319474 283132 319544 283188
rect 319224 283064 319544 283132
rect 319224 283008 319294 283064
rect 319350 283008 319418 283064
rect 319474 283008 319544 283064
rect 319224 282940 319544 283008
rect 319224 282884 319294 282940
rect 319350 282884 319418 282940
rect 319474 282884 319544 282940
rect 319224 282816 319544 282884
rect 319224 282760 319294 282816
rect 319350 282760 319418 282816
rect 319474 282760 319544 282816
rect 319224 282692 319544 282760
rect 319224 282636 319294 282692
rect 319350 282636 319418 282692
rect 319474 282636 319544 282692
rect 319224 282568 319544 282636
rect 319224 282512 319294 282568
rect 319350 282512 319418 282568
rect 319474 282512 319544 282568
rect 314224 281912 314544 282042
rect 314224 281856 314294 281912
rect 314350 281856 314418 281912
rect 314474 281856 314544 281912
rect 314224 281788 314544 281856
rect 314224 281732 314294 281788
rect 314350 281732 314418 281788
rect 314474 281732 314544 281788
rect 314224 281664 314544 281732
rect 314224 281608 314294 281664
rect 314350 281608 314418 281664
rect 314474 281608 314544 281664
rect 314224 281540 314544 281608
rect 314224 281484 314294 281540
rect 314350 281484 314418 281540
rect 314474 281484 314544 281540
rect 314224 281416 314544 281484
rect 314224 281360 314294 281416
rect 314350 281360 314418 281416
rect 314474 281360 314544 281416
rect 314224 281292 314544 281360
rect 314224 281236 314294 281292
rect 314350 281236 314418 281292
rect 314474 281236 314544 281292
rect 314224 281168 314544 281236
rect 314224 281112 314294 281168
rect 314350 281112 314418 281168
rect 314474 281112 314544 281168
rect 314224 279368 314544 281112
rect 319224 279368 319544 282512
rect 329224 283312 329544 283442
rect 329224 283256 329294 283312
rect 329350 283256 329418 283312
rect 329474 283256 329544 283312
rect 329224 283188 329544 283256
rect 329224 283132 329294 283188
rect 329350 283132 329418 283188
rect 329474 283132 329544 283188
rect 329224 283064 329544 283132
rect 329224 283008 329294 283064
rect 329350 283008 329418 283064
rect 329474 283008 329544 283064
rect 329224 282940 329544 283008
rect 329224 282884 329294 282940
rect 329350 282884 329418 282940
rect 329474 282884 329544 282940
rect 329224 282816 329544 282884
rect 329224 282760 329294 282816
rect 329350 282760 329418 282816
rect 329474 282760 329544 282816
rect 329224 282692 329544 282760
rect 329224 282636 329294 282692
rect 329350 282636 329418 282692
rect 329474 282636 329544 282692
rect 329224 282568 329544 282636
rect 329224 282512 329294 282568
rect 329350 282512 329418 282568
rect 329474 282512 329544 282568
rect 324224 281912 324544 282042
rect 324224 281856 324294 281912
rect 324350 281856 324418 281912
rect 324474 281856 324544 281912
rect 324224 281788 324544 281856
rect 324224 281732 324294 281788
rect 324350 281732 324418 281788
rect 324474 281732 324544 281788
rect 324224 281664 324544 281732
rect 324224 281608 324294 281664
rect 324350 281608 324418 281664
rect 324474 281608 324544 281664
rect 324224 281540 324544 281608
rect 324224 281484 324294 281540
rect 324350 281484 324418 281540
rect 324474 281484 324544 281540
rect 324224 281416 324544 281484
rect 324224 281360 324294 281416
rect 324350 281360 324418 281416
rect 324474 281360 324544 281416
rect 324224 281292 324544 281360
rect 324224 281236 324294 281292
rect 324350 281236 324418 281292
rect 324474 281236 324544 281292
rect 324224 281168 324544 281236
rect 324224 281112 324294 281168
rect 324350 281112 324418 281168
rect 324474 281112 324544 281168
rect 324224 279368 324544 281112
rect 329224 279368 329544 282512
rect 339224 283312 339544 283442
rect 339224 283256 339294 283312
rect 339350 283256 339418 283312
rect 339474 283256 339544 283312
rect 339224 283188 339544 283256
rect 339224 283132 339294 283188
rect 339350 283132 339418 283188
rect 339474 283132 339544 283188
rect 339224 283064 339544 283132
rect 339224 283008 339294 283064
rect 339350 283008 339418 283064
rect 339474 283008 339544 283064
rect 339224 282940 339544 283008
rect 339224 282884 339294 282940
rect 339350 282884 339418 282940
rect 339474 282884 339544 282940
rect 339224 282816 339544 282884
rect 339224 282760 339294 282816
rect 339350 282760 339418 282816
rect 339474 282760 339544 282816
rect 339224 282692 339544 282760
rect 339224 282636 339294 282692
rect 339350 282636 339418 282692
rect 339474 282636 339544 282692
rect 339224 282568 339544 282636
rect 339224 282512 339294 282568
rect 339350 282512 339418 282568
rect 339474 282512 339544 282568
rect 334224 281912 334544 282042
rect 334224 281856 334294 281912
rect 334350 281856 334418 281912
rect 334474 281856 334544 281912
rect 334224 281788 334544 281856
rect 334224 281732 334294 281788
rect 334350 281732 334418 281788
rect 334474 281732 334544 281788
rect 334224 281664 334544 281732
rect 334224 281608 334294 281664
rect 334350 281608 334418 281664
rect 334474 281608 334544 281664
rect 334224 281540 334544 281608
rect 334224 281484 334294 281540
rect 334350 281484 334418 281540
rect 334474 281484 334544 281540
rect 334224 281416 334544 281484
rect 334224 281360 334294 281416
rect 334350 281360 334418 281416
rect 334474 281360 334544 281416
rect 334224 281292 334544 281360
rect 334224 281236 334294 281292
rect 334350 281236 334418 281292
rect 334474 281236 334544 281292
rect 334224 281168 334544 281236
rect 334224 281112 334294 281168
rect 334350 281112 334418 281168
rect 334474 281112 334544 281168
rect 334224 279368 334544 281112
rect 339224 279368 339544 282512
rect 349224 283312 349544 283442
rect 349224 283256 349294 283312
rect 349350 283256 349418 283312
rect 349474 283256 349544 283312
rect 349224 283188 349544 283256
rect 349224 283132 349294 283188
rect 349350 283132 349418 283188
rect 349474 283132 349544 283188
rect 349224 283064 349544 283132
rect 349224 283008 349294 283064
rect 349350 283008 349418 283064
rect 349474 283008 349544 283064
rect 349224 282940 349544 283008
rect 349224 282884 349294 282940
rect 349350 282884 349418 282940
rect 349474 282884 349544 282940
rect 349224 282816 349544 282884
rect 349224 282760 349294 282816
rect 349350 282760 349418 282816
rect 349474 282760 349544 282816
rect 349224 282692 349544 282760
rect 349224 282636 349294 282692
rect 349350 282636 349418 282692
rect 349474 282636 349544 282692
rect 349224 282568 349544 282636
rect 349224 282512 349294 282568
rect 349350 282512 349418 282568
rect 349474 282512 349544 282568
rect 344224 281912 344544 282042
rect 344224 281856 344294 281912
rect 344350 281856 344418 281912
rect 344474 281856 344544 281912
rect 344224 281788 344544 281856
rect 344224 281732 344294 281788
rect 344350 281732 344418 281788
rect 344474 281732 344544 281788
rect 344224 281664 344544 281732
rect 344224 281608 344294 281664
rect 344350 281608 344418 281664
rect 344474 281608 344544 281664
rect 344224 281540 344544 281608
rect 344224 281484 344294 281540
rect 344350 281484 344418 281540
rect 344474 281484 344544 281540
rect 344224 281416 344544 281484
rect 344224 281360 344294 281416
rect 344350 281360 344418 281416
rect 344474 281360 344544 281416
rect 344224 281292 344544 281360
rect 344224 281236 344294 281292
rect 344350 281236 344418 281292
rect 344474 281236 344544 281292
rect 344224 281168 344544 281236
rect 344224 281112 344294 281168
rect 344350 281112 344418 281168
rect 344474 281112 344544 281168
rect 344224 279368 344544 281112
rect 349224 279368 349544 282512
rect 359224 283312 359544 283442
rect 359224 283256 359294 283312
rect 359350 283256 359418 283312
rect 359474 283256 359544 283312
rect 359224 283188 359544 283256
rect 359224 283132 359294 283188
rect 359350 283132 359418 283188
rect 359474 283132 359544 283188
rect 359224 283064 359544 283132
rect 359224 283008 359294 283064
rect 359350 283008 359418 283064
rect 359474 283008 359544 283064
rect 359224 282940 359544 283008
rect 359224 282884 359294 282940
rect 359350 282884 359418 282940
rect 359474 282884 359544 282940
rect 359224 282816 359544 282884
rect 359224 282760 359294 282816
rect 359350 282760 359418 282816
rect 359474 282760 359544 282816
rect 359224 282692 359544 282760
rect 359224 282636 359294 282692
rect 359350 282636 359418 282692
rect 359474 282636 359544 282692
rect 359224 282568 359544 282636
rect 359224 282512 359294 282568
rect 359350 282512 359418 282568
rect 359474 282512 359544 282568
rect 354224 281912 354544 282042
rect 354224 281856 354294 281912
rect 354350 281856 354418 281912
rect 354474 281856 354544 281912
rect 354224 281788 354544 281856
rect 354224 281732 354294 281788
rect 354350 281732 354418 281788
rect 354474 281732 354544 281788
rect 354224 281664 354544 281732
rect 354224 281608 354294 281664
rect 354350 281608 354418 281664
rect 354474 281608 354544 281664
rect 354224 281540 354544 281608
rect 354224 281484 354294 281540
rect 354350 281484 354418 281540
rect 354474 281484 354544 281540
rect 354224 281416 354544 281484
rect 354224 281360 354294 281416
rect 354350 281360 354418 281416
rect 354474 281360 354544 281416
rect 354224 281292 354544 281360
rect 354224 281236 354294 281292
rect 354350 281236 354418 281292
rect 354474 281236 354544 281292
rect 354224 281168 354544 281236
rect 354224 281112 354294 281168
rect 354350 281112 354418 281168
rect 354474 281112 354544 281168
rect 354224 279368 354544 281112
rect 359224 279368 359544 282512
rect 369224 283312 369544 283442
rect 369224 283256 369294 283312
rect 369350 283256 369418 283312
rect 369474 283256 369544 283312
rect 369224 283188 369544 283256
rect 369224 283132 369294 283188
rect 369350 283132 369418 283188
rect 369474 283132 369544 283188
rect 369224 283064 369544 283132
rect 369224 283008 369294 283064
rect 369350 283008 369418 283064
rect 369474 283008 369544 283064
rect 369224 282940 369544 283008
rect 369224 282884 369294 282940
rect 369350 282884 369418 282940
rect 369474 282884 369544 282940
rect 369224 282816 369544 282884
rect 369224 282760 369294 282816
rect 369350 282760 369418 282816
rect 369474 282760 369544 282816
rect 369224 282692 369544 282760
rect 369224 282636 369294 282692
rect 369350 282636 369418 282692
rect 369474 282636 369544 282692
rect 369224 282568 369544 282636
rect 369224 282512 369294 282568
rect 369350 282512 369418 282568
rect 369474 282512 369544 282568
rect 364224 281912 364544 282042
rect 364224 281856 364294 281912
rect 364350 281856 364418 281912
rect 364474 281856 364544 281912
rect 364224 281788 364544 281856
rect 364224 281732 364294 281788
rect 364350 281732 364418 281788
rect 364474 281732 364544 281788
rect 364224 281664 364544 281732
rect 364224 281608 364294 281664
rect 364350 281608 364418 281664
rect 364474 281608 364544 281664
rect 364224 281540 364544 281608
rect 364224 281484 364294 281540
rect 364350 281484 364418 281540
rect 364474 281484 364544 281540
rect 364224 281416 364544 281484
rect 364224 281360 364294 281416
rect 364350 281360 364418 281416
rect 364474 281360 364544 281416
rect 364224 281292 364544 281360
rect 364224 281236 364294 281292
rect 364350 281236 364418 281292
rect 364474 281236 364544 281292
rect 364224 281168 364544 281236
rect 364224 281112 364294 281168
rect 364350 281112 364418 281168
rect 364474 281112 364544 281168
rect 364224 279368 364544 281112
rect 369224 279368 369544 282512
rect 379224 283312 379544 283442
rect 379224 283256 379294 283312
rect 379350 283256 379418 283312
rect 379474 283256 379544 283312
rect 379224 283188 379544 283256
rect 379224 283132 379294 283188
rect 379350 283132 379418 283188
rect 379474 283132 379544 283188
rect 379224 283064 379544 283132
rect 379224 283008 379294 283064
rect 379350 283008 379418 283064
rect 379474 283008 379544 283064
rect 379224 282940 379544 283008
rect 379224 282884 379294 282940
rect 379350 282884 379418 282940
rect 379474 282884 379544 282940
rect 379224 282816 379544 282884
rect 379224 282760 379294 282816
rect 379350 282760 379418 282816
rect 379474 282760 379544 282816
rect 379224 282692 379544 282760
rect 379224 282636 379294 282692
rect 379350 282636 379418 282692
rect 379474 282636 379544 282692
rect 379224 282568 379544 282636
rect 379224 282512 379294 282568
rect 379350 282512 379418 282568
rect 379474 282512 379544 282568
rect 374224 281912 374544 282042
rect 374224 281856 374294 281912
rect 374350 281856 374418 281912
rect 374474 281856 374544 281912
rect 374224 281788 374544 281856
rect 374224 281732 374294 281788
rect 374350 281732 374418 281788
rect 374474 281732 374544 281788
rect 374224 281664 374544 281732
rect 374224 281608 374294 281664
rect 374350 281608 374418 281664
rect 374474 281608 374544 281664
rect 374224 281540 374544 281608
rect 374224 281484 374294 281540
rect 374350 281484 374418 281540
rect 374474 281484 374544 281540
rect 374224 281416 374544 281484
rect 374224 281360 374294 281416
rect 374350 281360 374418 281416
rect 374474 281360 374544 281416
rect 374224 281292 374544 281360
rect 374224 281236 374294 281292
rect 374350 281236 374418 281292
rect 374474 281236 374544 281292
rect 374224 281168 374544 281236
rect 374224 281112 374294 281168
rect 374350 281112 374418 281168
rect 374474 281112 374544 281168
rect 374224 279368 374544 281112
rect 379224 279368 379544 282512
rect 389224 283312 389544 283442
rect 389224 283256 389294 283312
rect 389350 283256 389418 283312
rect 389474 283256 389544 283312
rect 389224 283188 389544 283256
rect 389224 283132 389294 283188
rect 389350 283132 389418 283188
rect 389474 283132 389544 283188
rect 389224 283064 389544 283132
rect 389224 283008 389294 283064
rect 389350 283008 389418 283064
rect 389474 283008 389544 283064
rect 389224 282940 389544 283008
rect 389224 282884 389294 282940
rect 389350 282884 389418 282940
rect 389474 282884 389544 282940
rect 389224 282816 389544 282884
rect 389224 282760 389294 282816
rect 389350 282760 389418 282816
rect 389474 282760 389544 282816
rect 389224 282692 389544 282760
rect 389224 282636 389294 282692
rect 389350 282636 389418 282692
rect 389474 282636 389544 282692
rect 389224 282568 389544 282636
rect 389224 282512 389294 282568
rect 389350 282512 389418 282568
rect 389474 282512 389544 282568
rect 384224 281912 384544 282042
rect 384224 281856 384294 281912
rect 384350 281856 384418 281912
rect 384474 281856 384544 281912
rect 384224 281788 384544 281856
rect 384224 281732 384294 281788
rect 384350 281732 384418 281788
rect 384474 281732 384544 281788
rect 384224 281664 384544 281732
rect 384224 281608 384294 281664
rect 384350 281608 384418 281664
rect 384474 281608 384544 281664
rect 384224 281540 384544 281608
rect 384224 281484 384294 281540
rect 384350 281484 384418 281540
rect 384474 281484 384544 281540
rect 384224 281416 384544 281484
rect 384224 281360 384294 281416
rect 384350 281360 384418 281416
rect 384474 281360 384544 281416
rect 384224 281292 384544 281360
rect 384224 281236 384294 281292
rect 384350 281236 384418 281292
rect 384474 281236 384544 281292
rect 384224 281168 384544 281236
rect 384224 281112 384294 281168
rect 384350 281112 384418 281168
rect 384474 281112 384544 281168
rect 384224 279368 384544 281112
rect 389224 279368 389544 282512
rect 399224 283312 399544 283442
rect 399224 283256 399294 283312
rect 399350 283256 399418 283312
rect 399474 283256 399544 283312
rect 399224 283188 399544 283256
rect 399224 283132 399294 283188
rect 399350 283132 399418 283188
rect 399474 283132 399544 283188
rect 399224 283064 399544 283132
rect 399224 283008 399294 283064
rect 399350 283008 399418 283064
rect 399474 283008 399544 283064
rect 399224 282940 399544 283008
rect 399224 282884 399294 282940
rect 399350 282884 399418 282940
rect 399474 282884 399544 282940
rect 399224 282816 399544 282884
rect 399224 282760 399294 282816
rect 399350 282760 399418 282816
rect 399474 282760 399544 282816
rect 399224 282692 399544 282760
rect 399224 282636 399294 282692
rect 399350 282636 399418 282692
rect 399474 282636 399544 282692
rect 399224 282568 399544 282636
rect 399224 282512 399294 282568
rect 399350 282512 399418 282568
rect 399474 282512 399544 282568
rect 394224 281912 394544 282042
rect 394224 281856 394294 281912
rect 394350 281856 394418 281912
rect 394474 281856 394544 281912
rect 394224 281788 394544 281856
rect 394224 281732 394294 281788
rect 394350 281732 394418 281788
rect 394474 281732 394544 281788
rect 394224 281664 394544 281732
rect 394224 281608 394294 281664
rect 394350 281608 394418 281664
rect 394474 281608 394544 281664
rect 394224 281540 394544 281608
rect 394224 281484 394294 281540
rect 394350 281484 394418 281540
rect 394474 281484 394544 281540
rect 394224 281416 394544 281484
rect 394224 281360 394294 281416
rect 394350 281360 394418 281416
rect 394474 281360 394544 281416
rect 394224 281292 394544 281360
rect 394224 281236 394294 281292
rect 394350 281236 394418 281292
rect 394474 281236 394544 281292
rect 394224 281168 394544 281236
rect 394224 281112 394294 281168
rect 394350 281112 394418 281168
rect 394474 281112 394544 281168
rect 394224 279368 394544 281112
rect 399224 279368 399544 282512
rect 409224 283312 409544 283442
rect 409224 283256 409294 283312
rect 409350 283256 409418 283312
rect 409474 283256 409544 283312
rect 409224 283188 409544 283256
rect 409224 283132 409294 283188
rect 409350 283132 409418 283188
rect 409474 283132 409544 283188
rect 409224 283064 409544 283132
rect 409224 283008 409294 283064
rect 409350 283008 409418 283064
rect 409474 283008 409544 283064
rect 409224 282940 409544 283008
rect 409224 282884 409294 282940
rect 409350 282884 409418 282940
rect 409474 282884 409544 282940
rect 409224 282816 409544 282884
rect 409224 282760 409294 282816
rect 409350 282760 409418 282816
rect 409474 282760 409544 282816
rect 409224 282692 409544 282760
rect 409224 282636 409294 282692
rect 409350 282636 409418 282692
rect 409474 282636 409544 282692
rect 409224 282568 409544 282636
rect 409224 282512 409294 282568
rect 409350 282512 409418 282568
rect 409474 282512 409544 282568
rect 404224 281912 404544 282042
rect 404224 281856 404294 281912
rect 404350 281856 404418 281912
rect 404474 281856 404544 281912
rect 404224 281788 404544 281856
rect 404224 281732 404294 281788
rect 404350 281732 404418 281788
rect 404474 281732 404544 281788
rect 404224 281664 404544 281732
rect 404224 281608 404294 281664
rect 404350 281608 404418 281664
rect 404474 281608 404544 281664
rect 404224 281540 404544 281608
rect 404224 281484 404294 281540
rect 404350 281484 404418 281540
rect 404474 281484 404544 281540
rect 404224 281416 404544 281484
rect 404224 281360 404294 281416
rect 404350 281360 404418 281416
rect 404474 281360 404544 281416
rect 404224 281292 404544 281360
rect 404224 281236 404294 281292
rect 404350 281236 404418 281292
rect 404474 281236 404544 281292
rect 404224 281168 404544 281236
rect 404224 281112 404294 281168
rect 404350 281112 404418 281168
rect 404474 281112 404544 281168
rect 404224 279368 404544 281112
rect 409224 279368 409544 282512
rect 419224 283312 419544 283442
rect 419224 283256 419294 283312
rect 419350 283256 419418 283312
rect 419474 283256 419544 283312
rect 419224 283188 419544 283256
rect 419224 283132 419294 283188
rect 419350 283132 419418 283188
rect 419474 283132 419544 283188
rect 419224 283064 419544 283132
rect 419224 283008 419294 283064
rect 419350 283008 419418 283064
rect 419474 283008 419544 283064
rect 419224 282940 419544 283008
rect 419224 282884 419294 282940
rect 419350 282884 419418 282940
rect 419474 282884 419544 282940
rect 419224 282816 419544 282884
rect 419224 282760 419294 282816
rect 419350 282760 419418 282816
rect 419474 282760 419544 282816
rect 419224 282692 419544 282760
rect 419224 282636 419294 282692
rect 419350 282636 419418 282692
rect 419474 282636 419544 282692
rect 419224 282568 419544 282636
rect 419224 282512 419294 282568
rect 419350 282512 419418 282568
rect 419474 282512 419544 282568
rect 414224 281912 414544 282042
rect 414224 281856 414294 281912
rect 414350 281856 414418 281912
rect 414474 281856 414544 281912
rect 414224 281788 414544 281856
rect 414224 281732 414294 281788
rect 414350 281732 414418 281788
rect 414474 281732 414544 281788
rect 414224 281664 414544 281732
rect 414224 281608 414294 281664
rect 414350 281608 414418 281664
rect 414474 281608 414544 281664
rect 414224 281540 414544 281608
rect 414224 281484 414294 281540
rect 414350 281484 414418 281540
rect 414474 281484 414544 281540
rect 414224 281416 414544 281484
rect 414224 281360 414294 281416
rect 414350 281360 414418 281416
rect 414474 281360 414544 281416
rect 414224 281292 414544 281360
rect 414224 281236 414294 281292
rect 414350 281236 414418 281292
rect 414474 281236 414544 281292
rect 414224 281168 414544 281236
rect 414224 281112 414294 281168
rect 414350 281112 414418 281168
rect 414474 281112 414544 281168
rect 414224 279368 414544 281112
rect 419224 279368 419544 282512
rect 429224 283312 429544 283442
rect 429224 283256 429294 283312
rect 429350 283256 429418 283312
rect 429474 283256 429544 283312
rect 429224 283188 429544 283256
rect 429224 283132 429294 283188
rect 429350 283132 429418 283188
rect 429474 283132 429544 283188
rect 429224 283064 429544 283132
rect 429224 283008 429294 283064
rect 429350 283008 429418 283064
rect 429474 283008 429544 283064
rect 429224 282940 429544 283008
rect 429224 282884 429294 282940
rect 429350 282884 429418 282940
rect 429474 282884 429544 282940
rect 429224 282816 429544 282884
rect 429224 282760 429294 282816
rect 429350 282760 429418 282816
rect 429474 282760 429544 282816
rect 429224 282692 429544 282760
rect 429224 282636 429294 282692
rect 429350 282636 429418 282692
rect 429474 282636 429544 282692
rect 429224 282568 429544 282636
rect 429224 282512 429294 282568
rect 429350 282512 429418 282568
rect 429474 282512 429544 282568
rect 424224 281912 424544 282042
rect 424224 281856 424294 281912
rect 424350 281856 424418 281912
rect 424474 281856 424544 281912
rect 424224 281788 424544 281856
rect 424224 281732 424294 281788
rect 424350 281732 424418 281788
rect 424474 281732 424544 281788
rect 424224 281664 424544 281732
rect 424224 281608 424294 281664
rect 424350 281608 424418 281664
rect 424474 281608 424544 281664
rect 424224 281540 424544 281608
rect 424224 281484 424294 281540
rect 424350 281484 424418 281540
rect 424474 281484 424544 281540
rect 424224 281416 424544 281484
rect 424224 281360 424294 281416
rect 424350 281360 424418 281416
rect 424474 281360 424544 281416
rect 424224 281292 424544 281360
rect 424224 281236 424294 281292
rect 424350 281236 424418 281292
rect 424474 281236 424544 281292
rect 424224 281168 424544 281236
rect 424224 281112 424294 281168
rect 424350 281112 424418 281168
rect 424474 281112 424544 281168
rect 424224 279368 424544 281112
rect 429224 279368 429544 282512
rect 439224 283312 439544 283442
rect 439224 283256 439294 283312
rect 439350 283256 439418 283312
rect 439474 283256 439544 283312
rect 439224 283188 439544 283256
rect 439224 283132 439294 283188
rect 439350 283132 439418 283188
rect 439474 283132 439544 283188
rect 439224 283064 439544 283132
rect 439224 283008 439294 283064
rect 439350 283008 439418 283064
rect 439474 283008 439544 283064
rect 439224 282940 439544 283008
rect 439224 282884 439294 282940
rect 439350 282884 439418 282940
rect 439474 282884 439544 282940
rect 439224 282816 439544 282884
rect 439224 282760 439294 282816
rect 439350 282760 439418 282816
rect 439474 282760 439544 282816
rect 439224 282692 439544 282760
rect 439224 282636 439294 282692
rect 439350 282636 439418 282692
rect 439474 282636 439544 282692
rect 439224 282568 439544 282636
rect 439224 282512 439294 282568
rect 439350 282512 439418 282568
rect 439474 282512 439544 282568
rect 434224 281912 434544 282042
rect 434224 281856 434294 281912
rect 434350 281856 434418 281912
rect 434474 281856 434544 281912
rect 434224 281788 434544 281856
rect 434224 281732 434294 281788
rect 434350 281732 434418 281788
rect 434474 281732 434544 281788
rect 434224 281664 434544 281732
rect 434224 281608 434294 281664
rect 434350 281608 434418 281664
rect 434474 281608 434544 281664
rect 434224 281540 434544 281608
rect 434224 281484 434294 281540
rect 434350 281484 434418 281540
rect 434474 281484 434544 281540
rect 434224 281416 434544 281484
rect 434224 281360 434294 281416
rect 434350 281360 434418 281416
rect 434474 281360 434544 281416
rect 434224 281292 434544 281360
rect 434224 281236 434294 281292
rect 434350 281236 434418 281292
rect 434474 281236 434544 281292
rect 434224 281168 434544 281236
rect 434224 281112 434294 281168
rect 434350 281112 434418 281168
rect 434474 281112 434544 281168
rect 434224 279368 434544 281112
rect 439224 279368 439544 282512
rect 449224 283312 449544 283442
rect 449224 283256 449294 283312
rect 449350 283256 449418 283312
rect 449474 283256 449544 283312
rect 449224 283188 449544 283256
rect 449224 283132 449294 283188
rect 449350 283132 449418 283188
rect 449474 283132 449544 283188
rect 449224 283064 449544 283132
rect 449224 283008 449294 283064
rect 449350 283008 449418 283064
rect 449474 283008 449544 283064
rect 449224 282940 449544 283008
rect 449224 282884 449294 282940
rect 449350 282884 449418 282940
rect 449474 282884 449544 282940
rect 449224 282816 449544 282884
rect 449224 282760 449294 282816
rect 449350 282760 449418 282816
rect 449474 282760 449544 282816
rect 449224 282692 449544 282760
rect 449224 282636 449294 282692
rect 449350 282636 449418 282692
rect 449474 282636 449544 282692
rect 449224 282568 449544 282636
rect 449224 282512 449294 282568
rect 449350 282512 449418 282568
rect 449474 282512 449544 282568
rect 444224 281912 444544 282042
rect 444224 281856 444294 281912
rect 444350 281856 444418 281912
rect 444474 281856 444544 281912
rect 444224 281788 444544 281856
rect 444224 281732 444294 281788
rect 444350 281732 444418 281788
rect 444474 281732 444544 281788
rect 444224 281664 444544 281732
rect 444224 281608 444294 281664
rect 444350 281608 444418 281664
rect 444474 281608 444544 281664
rect 444224 281540 444544 281608
rect 444224 281484 444294 281540
rect 444350 281484 444418 281540
rect 444474 281484 444544 281540
rect 444224 281416 444544 281484
rect 444224 281360 444294 281416
rect 444350 281360 444418 281416
rect 444474 281360 444544 281416
rect 444224 281292 444544 281360
rect 444224 281236 444294 281292
rect 444350 281236 444418 281292
rect 444474 281236 444544 281292
rect 444224 281168 444544 281236
rect 444224 281112 444294 281168
rect 444350 281112 444418 281168
rect 444474 281112 444544 281168
rect 444224 279368 444544 281112
rect 449224 279368 449544 282512
rect 459224 283312 459544 283442
rect 459224 283256 459294 283312
rect 459350 283256 459418 283312
rect 459474 283256 459544 283312
rect 459224 283188 459544 283256
rect 459224 283132 459294 283188
rect 459350 283132 459418 283188
rect 459474 283132 459544 283188
rect 459224 283064 459544 283132
rect 459224 283008 459294 283064
rect 459350 283008 459418 283064
rect 459474 283008 459544 283064
rect 459224 282940 459544 283008
rect 459224 282884 459294 282940
rect 459350 282884 459418 282940
rect 459474 282884 459544 282940
rect 459224 282816 459544 282884
rect 459224 282760 459294 282816
rect 459350 282760 459418 282816
rect 459474 282760 459544 282816
rect 459224 282692 459544 282760
rect 459224 282636 459294 282692
rect 459350 282636 459418 282692
rect 459474 282636 459544 282692
rect 459224 282568 459544 282636
rect 459224 282512 459294 282568
rect 459350 282512 459418 282568
rect 459474 282512 459544 282568
rect 454224 281912 454544 282042
rect 454224 281856 454294 281912
rect 454350 281856 454418 281912
rect 454474 281856 454544 281912
rect 454224 281788 454544 281856
rect 454224 281732 454294 281788
rect 454350 281732 454418 281788
rect 454474 281732 454544 281788
rect 454224 281664 454544 281732
rect 454224 281608 454294 281664
rect 454350 281608 454418 281664
rect 454474 281608 454544 281664
rect 454224 281540 454544 281608
rect 454224 281484 454294 281540
rect 454350 281484 454418 281540
rect 454474 281484 454544 281540
rect 454224 281416 454544 281484
rect 454224 281360 454294 281416
rect 454350 281360 454418 281416
rect 454474 281360 454544 281416
rect 454224 281292 454544 281360
rect 454224 281236 454294 281292
rect 454350 281236 454418 281292
rect 454474 281236 454544 281292
rect 454224 281168 454544 281236
rect 454224 281112 454294 281168
rect 454350 281112 454418 281168
rect 454474 281112 454544 281168
rect 454224 279368 454544 281112
rect 459224 279368 459544 282512
rect 469224 283312 469544 283442
rect 469224 283256 469294 283312
rect 469350 283256 469418 283312
rect 469474 283256 469544 283312
rect 469224 283188 469544 283256
rect 469224 283132 469294 283188
rect 469350 283132 469418 283188
rect 469474 283132 469544 283188
rect 469224 283064 469544 283132
rect 469224 283008 469294 283064
rect 469350 283008 469418 283064
rect 469474 283008 469544 283064
rect 469224 282940 469544 283008
rect 469224 282884 469294 282940
rect 469350 282884 469418 282940
rect 469474 282884 469544 282940
rect 469224 282816 469544 282884
rect 469224 282760 469294 282816
rect 469350 282760 469418 282816
rect 469474 282760 469544 282816
rect 469224 282692 469544 282760
rect 469224 282636 469294 282692
rect 469350 282636 469418 282692
rect 469474 282636 469544 282692
rect 469224 282568 469544 282636
rect 469224 282512 469294 282568
rect 469350 282512 469418 282568
rect 469474 282512 469544 282568
rect 464224 281912 464544 282042
rect 464224 281856 464294 281912
rect 464350 281856 464418 281912
rect 464474 281856 464544 281912
rect 464224 281788 464544 281856
rect 464224 281732 464294 281788
rect 464350 281732 464418 281788
rect 464474 281732 464544 281788
rect 464224 281664 464544 281732
rect 464224 281608 464294 281664
rect 464350 281608 464418 281664
rect 464474 281608 464544 281664
rect 464224 281540 464544 281608
rect 464224 281484 464294 281540
rect 464350 281484 464418 281540
rect 464474 281484 464544 281540
rect 464224 281416 464544 281484
rect 464224 281360 464294 281416
rect 464350 281360 464418 281416
rect 464474 281360 464544 281416
rect 464224 281292 464544 281360
rect 464224 281236 464294 281292
rect 464350 281236 464418 281292
rect 464474 281236 464544 281292
rect 464224 281168 464544 281236
rect 464224 281112 464294 281168
rect 464350 281112 464418 281168
rect 464474 281112 464544 281168
rect 464224 279368 464544 281112
rect 469224 279368 469544 282512
rect 479224 283312 479544 283442
rect 479224 283256 479294 283312
rect 479350 283256 479418 283312
rect 479474 283256 479544 283312
rect 479224 283188 479544 283256
rect 479224 283132 479294 283188
rect 479350 283132 479418 283188
rect 479474 283132 479544 283188
rect 479224 283064 479544 283132
rect 479224 283008 479294 283064
rect 479350 283008 479418 283064
rect 479474 283008 479544 283064
rect 479224 282940 479544 283008
rect 479224 282884 479294 282940
rect 479350 282884 479418 282940
rect 479474 282884 479544 282940
rect 479224 282816 479544 282884
rect 479224 282760 479294 282816
rect 479350 282760 479418 282816
rect 479474 282760 479544 282816
rect 479224 282692 479544 282760
rect 479224 282636 479294 282692
rect 479350 282636 479418 282692
rect 479474 282636 479544 282692
rect 479224 282568 479544 282636
rect 479224 282512 479294 282568
rect 479350 282512 479418 282568
rect 479474 282512 479544 282568
rect 474224 281912 474544 282042
rect 474224 281856 474294 281912
rect 474350 281856 474418 281912
rect 474474 281856 474544 281912
rect 474224 281788 474544 281856
rect 474224 281732 474294 281788
rect 474350 281732 474418 281788
rect 474474 281732 474544 281788
rect 474224 281664 474544 281732
rect 474224 281608 474294 281664
rect 474350 281608 474418 281664
rect 474474 281608 474544 281664
rect 474224 281540 474544 281608
rect 474224 281484 474294 281540
rect 474350 281484 474418 281540
rect 474474 281484 474544 281540
rect 474224 281416 474544 281484
rect 474224 281360 474294 281416
rect 474350 281360 474418 281416
rect 474474 281360 474544 281416
rect 474224 281292 474544 281360
rect 474224 281236 474294 281292
rect 474350 281236 474418 281292
rect 474474 281236 474544 281292
rect 474224 281168 474544 281236
rect 474224 281112 474294 281168
rect 474350 281112 474418 281168
rect 474474 281112 474544 281168
rect 474224 279368 474544 281112
rect 479224 279368 479544 282512
rect 489224 283312 489544 283442
rect 489224 283256 489294 283312
rect 489350 283256 489418 283312
rect 489474 283256 489544 283312
rect 489224 283188 489544 283256
rect 489224 283132 489294 283188
rect 489350 283132 489418 283188
rect 489474 283132 489544 283188
rect 489224 283064 489544 283132
rect 489224 283008 489294 283064
rect 489350 283008 489418 283064
rect 489474 283008 489544 283064
rect 489224 282940 489544 283008
rect 489224 282884 489294 282940
rect 489350 282884 489418 282940
rect 489474 282884 489544 282940
rect 489224 282816 489544 282884
rect 489224 282760 489294 282816
rect 489350 282760 489418 282816
rect 489474 282760 489544 282816
rect 489224 282692 489544 282760
rect 489224 282636 489294 282692
rect 489350 282636 489418 282692
rect 489474 282636 489544 282692
rect 489224 282568 489544 282636
rect 489224 282512 489294 282568
rect 489350 282512 489418 282568
rect 489474 282512 489544 282568
rect 484224 281912 484544 282042
rect 484224 281856 484294 281912
rect 484350 281856 484418 281912
rect 484474 281856 484544 281912
rect 484224 281788 484544 281856
rect 484224 281732 484294 281788
rect 484350 281732 484418 281788
rect 484474 281732 484544 281788
rect 484224 281664 484544 281732
rect 484224 281608 484294 281664
rect 484350 281608 484418 281664
rect 484474 281608 484544 281664
rect 484224 281540 484544 281608
rect 484224 281484 484294 281540
rect 484350 281484 484418 281540
rect 484474 281484 484544 281540
rect 484224 281416 484544 281484
rect 484224 281360 484294 281416
rect 484350 281360 484418 281416
rect 484474 281360 484544 281416
rect 484224 281292 484544 281360
rect 484224 281236 484294 281292
rect 484350 281236 484418 281292
rect 484474 281236 484544 281292
rect 484224 281168 484544 281236
rect 484224 281112 484294 281168
rect 484350 281112 484418 281168
rect 484474 281112 484544 281168
rect 484224 279368 484544 281112
rect 489224 279368 489544 282512
rect 499224 283312 499544 283442
rect 499224 283256 499294 283312
rect 499350 283256 499418 283312
rect 499474 283256 499544 283312
rect 499224 283188 499544 283256
rect 499224 283132 499294 283188
rect 499350 283132 499418 283188
rect 499474 283132 499544 283188
rect 499224 283064 499544 283132
rect 499224 283008 499294 283064
rect 499350 283008 499418 283064
rect 499474 283008 499544 283064
rect 499224 282940 499544 283008
rect 499224 282884 499294 282940
rect 499350 282884 499418 282940
rect 499474 282884 499544 282940
rect 499224 282816 499544 282884
rect 499224 282760 499294 282816
rect 499350 282760 499418 282816
rect 499474 282760 499544 282816
rect 499224 282692 499544 282760
rect 499224 282636 499294 282692
rect 499350 282636 499418 282692
rect 499474 282636 499544 282692
rect 499224 282568 499544 282636
rect 499224 282512 499294 282568
rect 499350 282512 499418 282568
rect 499474 282512 499544 282568
rect 494224 281912 494544 282042
rect 494224 281856 494294 281912
rect 494350 281856 494418 281912
rect 494474 281856 494544 281912
rect 494224 281788 494544 281856
rect 494224 281732 494294 281788
rect 494350 281732 494418 281788
rect 494474 281732 494544 281788
rect 494224 281664 494544 281732
rect 494224 281608 494294 281664
rect 494350 281608 494418 281664
rect 494474 281608 494544 281664
rect 494224 281540 494544 281608
rect 494224 281484 494294 281540
rect 494350 281484 494418 281540
rect 494474 281484 494544 281540
rect 494224 281416 494544 281484
rect 494224 281360 494294 281416
rect 494350 281360 494418 281416
rect 494474 281360 494544 281416
rect 494224 281292 494544 281360
rect 494224 281236 494294 281292
rect 494350 281236 494418 281292
rect 494474 281236 494544 281292
rect 494224 281168 494544 281236
rect 494224 281112 494294 281168
rect 494350 281112 494418 281168
rect 494474 281112 494544 281168
rect 494224 279368 494544 281112
rect 499224 279368 499544 282512
rect 509224 283312 509544 283442
rect 509224 283256 509294 283312
rect 509350 283256 509418 283312
rect 509474 283256 509544 283312
rect 509224 283188 509544 283256
rect 509224 283132 509294 283188
rect 509350 283132 509418 283188
rect 509474 283132 509544 283188
rect 509224 283064 509544 283132
rect 509224 283008 509294 283064
rect 509350 283008 509418 283064
rect 509474 283008 509544 283064
rect 509224 282940 509544 283008
rect 509224 282884 509294 282940
rect 509350 282884 509418 282940
rect 509474 282884 509544 282940
rect 509224 282816 509544 282884
rect 509224 282760 509294 282816
rect 509350 282760 509418 282816
rect 509474 282760 509544 282816
rect 509224 282692 509544 282760
rect 509224 282636 509294 282692
rect 509350 282636 509418 282692
rect 509474 282636 509544 282692
rect 509224 282568 509544 282636
rect 509224 282512 509294 282568
rect 509350 282512 509418 282568
rect 509474 282512 509544 282568
rect 504224 281912 504544 282042
rect 504224 281856 504294 281912
rect 504350 281856 504418 281912
rect 504474 281856 504544 281912
rect 504224 281788 504544 281856
rect 504224 281732 504294 281788
rect 504350 281732 504418 281788
rect 504474 281732 504544 281788
rect 504224 281664 504544 281732
rect 504224 281608 504294 281664
rect 504350 281608 504418 281664
rect 504474 281608 504544 281664
rect 504224 281540 504544 281608
rect 504224 281484 504294 281540
rect 504350 281484 504418 281540
rect 504474 281484 504544 281540
rect 504224 281416 504544 281484
rect 504224 281360 504294 281416
rect 504350 281360 504418 281416
rect 504474 281360 504544 281416
rect 504224 281292 504544 281360
rect 504224 281236 504294 281292
rect 504350 281236 504418 281292
rect 504474 281236 504544 281292
rect 504224 281168 504544 281236
rect 504224 281112 504294 281168
rect 504350 281112 504418 281168
rect 504474 281112 504544 281168
rect 504224 279368 504544 281112
rect 509224 279368 509544 282512
rect 519224 283312 519544 283442
rect 519224 283256 519294 283312
rect 519350 283256 519418 283312
rect 519474 283256 519544 283312
rect 519224 283188 519544 283256
rect 519224 283132 519294 283188
rect 519350 283132 519418 283188
rect 519474 283132 519544 283188
rect 519224 283064 519544 283132
rect 519224 283008 519294 283064
rect 519350 283008 519418 283064
rect 519474 283008 519544 283064
rect 519224 282940 519544 283008
rect 519224 282884 519294 282940
rect 519350 282884 519418 282940
rect 519474 282884 519544 282940
rect 519224 282816 519544 282884
rect 519224 282760 519294 282816
rect 519350 282760 519418 282816
rect 519474 282760 519544 282816
rect 519224 282692 519544 282760
rect 519224 282636 519294 282692
rect 519350 282636 519418 282692
rect 519474 282636 519544 282692
rect 519224 282568 519544 282636
rect 519224 282512 519294 282568
rect 519350 282512 519418 282568
rect 519474 282512 519544 282568
rect 514224 281912 514544 282042
rect 514224 281856 514294 281912
rect 514350 281856 514418 281912
rect 514474 281856 514544 281912
rect 514224 281788 514544 281856
rect 514224 281732 514294 281788
rect 514350 281732 514418 281788
rect 514474 281732 514544 281788
rect 514224 281664 514544 281732
rect 514224 281608 514294 281664
rect 514350 281608 514418 281664
rect 514474 281608 514544 281664
rect 514224 281540 514544 281608
rect 514224 281484 514294 281540
rect 514350 281484 514418 281540
rect 514474 281484 514544 281540
rect 514224 281416 514544 281484
rect 514224 281360 514294 281416
rect 514350 281360 514418 281416
rect 514474 281360 514544 281416
rect 514224 281292 514544 281360
rect 514224 281236 514294 281292
rect 514350 281236 514418 281292
rect 514474 281236 514544 281292
rect 514224 281168 514544 281236
rect 514224 281112 514294 281168
rect 514350 281112 514418 281168
rect 514474 281112 514544 281168
rect 514224 279368 514544 281112
rect 519224 279368 519544 282512
rect 529224 283312 529544 283442
rect 529224 283256 529294 283312
rect 529350 283256 529418 283312
rect 529474 283256 529544 283312
rect 529224 283188 529544 283256
rect 529224 283132 529294 283188
rect 529350 283132 529418 283188
rect 529474 283132 529544 283188
rect 529224 283064 529544 283132
rect 529224 283008 529294 283064
rect 529350 283008 529418 283064
rect 529474 283008 529544 283064
rect 529224 282940 529544 283008
rect 529224 282884 529294 282940
rect 529350 282884 529418 282940
rect 529474 282884 529544 282940
rect 529224 282816 529544 282884
rect 529224 282760 529294 282816
rect 529350 282760 529418 282816
rect 529474 282760 529544 282816
rect 529224 282692 529544 282760
rect 529224 282636 529294 282692
rect 529350 282636 529418 282692
rect 529474 282636 529544 282692
rect 529224 282568 529544 282636
rect 529224 282512 529294 282568
rect 529350 282512 529418 282568
rect 529474 282512 529544 282568
rect 524224 281912 524544 282042
rect 524224 281856 524294 281912
rect 524350 281856 524418 281912
rect 524474 281856 524544 281912
rect 524224 281788 524544 281856
rect 524224 281732 524294 281788
rect 524350 281732 524418 281788
rect 524474 281732 524544 281788
rect 524224 281664 524544 281732
rect 524224 281608 524294 281664
rect 524350 281608 524418 281664
rect 524474 281608 524544 281664
rect 524224 281540 524544 281608
rect 524224 281484 524294 281540
rect 524350 281484 524418 281540
rect 524474 281484 524544 281540
rect 524224 281416 524544 281484
rect 524224 281360 524294 281416
rect 524350 281360 524418 281416
rect 524474 281360 524544 281416
rect 524224 281292 524544 281360
rect 524224 281236 524294 281292
rect 524350 281236 524418 281292
rect 524474 281236 524544 281292
rect 524224 281168 524544 281236
rect 524224 281112 524294 281168
rect 524350 281112 524418 281168
rect 524474 281112 524544 281168
rect 524224 279368 524544 281112
rect 529224 279368 529544 282512
rect 539224 283312 539544 283442
rect 539224 283256 539294 283312
rect 539350 283256 539418 283312
rect 539474 283256 539544 283312
rect 539224 283188 539544 283256
rect 539224 283132 539294 283188
rect 539350 283132 539418 283188
rect 539474 283132 539544 283188
rect 539224 283064 539544 283132
rect 539224 283008 539294 283064
rect 539350 283008 539418 283064
rect 539474 283008 539544 283064
rect 539224 282940 539544 283008
rect 539224 282884 539294 282940
rect 539350 282884 539418 282940
rect 539474 282884 539544 282940
rect 539224 282816 539544 282884
rect 539224 282760 539294 282816
rect 539350 282760 539418 282816
rect 539474 282760 539544 282816
rect 539224 282692 539544 282760
rect 539224 282636 539294 282692
rect 539350 282636 539418 282692
rect 539474 282636 539544 282692
rect 539224 282568 539544 282636
rect 539224 282512 539294 282568
rect 539350 282512 539418 282568
rect 539474 282512 539544 282568
rect 534224 281912 534544 282042
rect 534224 281856 534294 281912
rect 534350 281856 534418 281912
rect 534474 281856 534544 281912
rect 534224 281788 534544 281856
rect 534224 281732 534294 281788
rect 534350 281732 534418 281788
rect 534474 281732 534544 281788
rect 534224 281664 534544 281732
rect 534224 281608 534294 281664
rect 534350 281608 534418 281664
rect 534474 281608 534544 281664
rect 534224 281540 534544 281608
rect 534224 281484 534294 281540
rect 534350 281484 534418 281540
rect 534474 281484 534544 281540
rect 534224 281416 534544 281484
rect 534224 281360 534294 281416
rect 534350 281360 534418 281416
rect 534474 281360 534544 281416
rect 534224 281292 534544 281360
rect 534224 281236 534294 281292
rect 534350 281236 534418 281292
rect 534474 281236 534544 281292
rect 534224 281168 534544 281236
rect 534224 281112 534294 281168
rect 534350 281112 534418 281168
rect 534474 281112 534544 281168
rect 534224 279368 534544 281112
rect 539224 279368 539544 282512
rect 549224 283312 549544 283442
rect 549224 283256 549294 283312
rect 549350 283256 549418 283312
rect 549474 283256 549544 283312
rect 549224 283188 549544 283256
rect 549224 283132 549294 283188
rect 549350 283132 549418 283188
rect 549474 283132 549544 283188
rect 549224 283064 549544 283132
rect 549224 283008 549294 283064
rect 549350 283008 549418 283064
rect 549474 283008 549544 283064
rect 549224 282940 549544 283008
rect 549224 282884 549294 282940
rect 549350 282884 549418 282940
rect 549474 282884 549544 282940
rect 549224 282816 549544 282884
rect 549224 282760 549294 282816
rect 549350 282760 549418 282816
rect 549474 282760 549544 282816
rect 549224 282692 549544 282760
rect 549224 282636 549294 282692
rect 549350 282636 549418 282692
rect 549474 282636 549544 282692
rect 549224 282568 549544 282636
rect 549224 282512 549294 282568
rect 549350 282512 549418 282568
rect 549474 282512 549544 282568
rect 544224 281912 544544 282042
rect 544224 281856 544294 281912
rect 544350 281856 544418 281912
rect 544474 281856 544544 281912
rect 544224 281788 544544 281856
rect 544224 281732 544294 281788
rect 544350 281732 544418 281788
rect 544474 281732 544544 281788
rect 544224 281664 544544 281732
rect 544224 281608 544294 281664
rect 544350 281608 544418 281664
rect 544474 281608 544544 281664
rect 544224 281540 544544 281608
rect 544224 281484 544294 281540
rect 544350 281484 544418 281540
rect 544474 281484 544544 281540
rect 544224 281416 544544 281484
rect 544224 281360 544294 281416
rect 544350 281360 544418 281416
rect 544474 281360 544544 281416
rect 544224 281292 544544 281360
rect 544224 281236 544294 281292
rect 544350 281236 544418 281292
rect 544474 281236 544544 281292
rect 544224 281168 544544 281236
rect 544224 281112 544294 281168
rect 544350 281112 544418 281168
rect 544474 281112 544544 281168
rect 544224 279368 544544 281112
rect 549224 279368 549544 282512
rect 590840 283372 591840 306326
rect 590840 283316 590970 283372
rect 591026 283316 591094 283372
rect 591150 283316 591218 283372
rect 591274 283316 591342 283372
rect 591398 283316 591466 283372
rect 591522 283316 591590 283372
rect 591646 283316 591714 283372
rect 591770 283316 591840 283372
rect 590840 283248 591840 283316
rect 590840 283192 590970 283248
rect 591026 283192 591094 283248
rect 591150 283192 591218 283248
rect 591274 283192 591342 283248
rect 591398 283192 591466 283248
rect 591522 283192 591590 283248
rect 591646 283192 591714 283248
rect 591770 283192 591840 283248
rect 590840 283124 591840 283192
rect 590840 283068 590970 283124
rect 591026 283068 591094 283124
rect 591150 283068 591218 283124
rect 591274 283068 591342 283124
rect 591398 283068 591466 283124
rect 591522 283068 591590 283124
rect 591646 283068 591714 283124
rect 591770 283068 591840 283124
rect 590840 283000 591840 283068
rect 590840 282944 590970 283000
rect 591026 282944 591094 283000
rect 591150 282944 591218 283000
rect 591274 282944 591342 283000
rect 591398 282944 591466 283000
rect 591522 282944 591590 283000
rect 591646 282944 591714 283000
rect 591770 282944 591840 283000
rect 590840 282876 591840 282944
rect 590840 282820 590970 282876
rect 591026 282820 591094 282876
rect 591150 282820 591218 282876
rect 591274 282820 591342 282876
rect 591398 282820 591466 282876
rect 591522 282820 591590 282876
rect 591646 282820 591714 282876
rect 591770 282820 591840 282876
rect 590840 282752 591840 282820
rect 590840 282696 590970 282752
rect 591026 282696 591094 282752
rect 591150 282696 591218 282752
rect 591274 282696 591342 282752
rect 591398 282696 591466 282752
rect 591522 282696 591590 282752
rect 591646 282696 591714 282752
rect 591770 282696 591840 282752
rect 590840 282628 591840 282696
rect 590840 282572 590970 282628
rect 591026 282572 591094 282628
rect 591150 282572 591218 282628
rect 591274 282572 591342 282628
rect 591398 282572 591466 282628
rect 591522 282572 591590 282628
rect 591646 282572 591714 282628
rect 591770 282572 591840 282628
rect 554224 281912 554544 282042
rect 554224 281856 554294 281912
rect 554350 281856 554418 281912
rect 554474 281856 554544 281912
rect 554224 281788 554544 281856
rect 554224 281732 554294 281788
rect 554350 281732 554418 281788
rect 554474 281732 554544 281788
rect 554224 281664 554544 281732
rect 554224 281608 554294 281664
rect 554350 281608 554418 281664
rect 554474 281608 554544 281664
rect 554224 281540 554544 281608
rect 554224 281484 554294 281540
rect 554350 281484 554418 281540
rect 554474 281484 554544 281540
rect 554224 281416 554544 281484
rect 554224 281360 554294 281416
rect 554350 281360 554418 281416
rect 554474 281360 554544 281416
rect 554224 281292 554544 281360
rect 554224 281236 554294 281292
rect 554350 281236 554418 281292
rect 554474 281236 554544 281292
rect 554224 281168 554544 281236
rect 554224 281112 554294 281168
rect 554350 281112 554418 281168
rect 554474 281112 554544 281168
rect 554224 279368 554544 281112
rect 79078 273566 79300 273622
rect 79356 273566 79600 273622
rect 79656 273566 79900 273622
rect 79956 273566 80078 273622
rect 79078 266622 80078 273566
rect 79078 266566 79300 266622
rect 79356 266566 79600 266622
rect 79656 266566 79900 266622
rect 79956 266566 80078 266622
rect 79078 259622 80078 266566
rect 79078 259566 79300 259622
rect 79356 259566 79600 259622
rect 79656 259566 79900 259622
rect 79956 259566 80078 259622
rect 79078 255372 80078 259566
rect 79078 255316 79148 255372
rect 79204 255316 79272 255372
rect 79328 255316 79396 255372
rect 79452 255316 79520 255372
rect 79576 255316 79644 255372
rect 79700 255316 79768 255372
rect 79824 255316 79892 255372
rect 79948 255316 80078 255372
rect 79078 255248 80078 255316
rect 79078 255192 79148 255248
rect 79204 255192 79272 255248
rect 79328 255192 79396 255248
rect 79452 255192 79520 255248
rect 79576 255192 79644 255248
rect 79700 255192 79768 255248
rect 79824 255192 79892 255248
rect 79948 255192 80078 255248
rect 79078 249048 80078 255192
rect 79078 248992 79284 249048
rect 79340 248992 79584 249048
rect 79640 248992 79884 249048
rect 79940 248992 80078 249048
rect 79078 232622 80078 248992
rect 79078 232566 79300 232622
rect 79356 232566 79600 232622
rect 79656 232566 79900 232622
rect 79956 232566 80078 232622
rect 79078 229372 80078 232566
rect 79078 229316 79148 229372
rect 79204 229316 79272 229372
rect 79328 229316 79396 229372
rect 79452 229316 79520 229372
rect 79576 229316 79644 229372
rect 79700 229316 79768 229372
rect 79824 229316 79892 229372
rect 79948 229316 80078 229372
rect 79078 229248 80078 229316
rect 79078 229192 79148 229248
rect 79204 229192 79272 229248
rect 79328 229192 79396 229248
rect 79452 229192 79520 229248
rect 79576 229192 79644 229248
rect 79700 229192 79768 229248
rect 79824 229192 79892 229248
rect 79948 229192 80078 229248
rect 79078 225622 80078 229192
rect 79078 225566 79300 225622
rect 79356 225566 79600 225622
rect 79656 225566 79900 225622
rect 79956 225566 80078 225622
rect 79078 218622 80078 225566
rect 79078 218566 79300 218622
rect 79356 218566 79600 218622
rect 79656 218566 79900 218622
rect 79956 218566 80078 218622
rect 79078 208048 80078 218566
rect 79078 207992 79284 208048
rect 79340 207992 79584 208048
rect 79640 207992 79884 208048
rect 79940 207992 80078 208048
rect 79078 203372 80078 207992
rect 79078 203316 79148 203372
rect 79204 203316 79272 203372
rect 79328 203316 79396 203372
rect 79452 203316 79520 203372
rect 79576 203316 79644 203372
rect 79700 203316 79768 203372
rect 79824 203316 79892 203372
rect 79948 203316 80078 203372
rect 79078 203248 80078 203316
rect 79078 203192 79148 203248
rect 79204 203192 79272 203248
rect 79328 203192 79396 203248
rect 79452 203192 79520 203248
rect 79576 203192 79644 203248
rect 79700 203192 79768 203248
rect 79824 203192 79892 203248
rect 79948 203192 80078 203248
rect 79078 191622 80078 203192
rect 79078 191566 79300 191622
rect 79356 191566 79600 191622
rect 79656 191566 79900 191622
rect 79956 191566 80078 191622
rect 79078 184622 80078 191566
rect 79078 184566 79300 184622
rect 79356 184566 79600 184622
rect 79656 184566 79900 184622
rect 79956 184566 80078 184622
rect 79078 177622 80078 184566
rect 79078 177566 79300 177622
rect 79356 177566 79600 177622
rect 79656 177566 79900 177622
rect 79956 177566 80078 177622
rect 79078 177372 80078 177566
rect 79078 177316 79148 177372
rect 79204 177316 79272 177372
rect 79328 177316 79396 177372
rect 79452 177316 79520 177372
rect 79576 177316 79644 177372
rect 79700 177316 79768 177372
rect 79824 177316 79892 177372
rect 79948 177316 80078 177372
rect 79078 177248 80078 177316
rect 79078 177192 79148 177248
rect 79204 177192 79272 177248
rect 79328 177192 79396 177248
rect 79452 177192 79520 177248
rect 79576 177192 79644 177248
rect 79700 177192 79768 177248
rect 79824 177192 79892 177248
rect 79948 177192 80078 177248
rect 79078 151372 80078 177192
rect 79078 151316 79148 151372
rect 79204 151316 79272 151372
rect 79328 151316 79396 151372
rect 79452 151316 79520 151372
rect 79576 151316 79644 151372
rect 79700 151316 79768 151372
rect 79824 151316 79892 151372
rect 79948 151316 80078 151372
rect 79078 151248 80078 151316
rect 79078 151192 79148 151248
rect 79204 151192 79272 151248
rect 79328 151192 79396 151248
rect 79452 151192 79520 151248
rect 79576 151192 79644 151248
rect 79700 151192 79768 151248
rect 79824 151192 79892 151248
rect 79948 151192 80078 151248
rect 79078 125372 80078 151192
rect 79078 125316 79148 125372
rect 79204 125316 79272 125372
rect 79328 125316 79396 125372
rect 79452 125316 79520 125372
rect 79576 125316 79644 125372
rect 79700 125316 79768 125372
rect 79824 125316 79892 125372
rect 79948 125316 80078 125372
rect 79078 125248 80078 125316
rect 79078 125192 79148 125248
rect 79204 125192 79272 125248
rect 79328 125192 79396 125248
rect 79452 125192 79520 125248
rect 79576 125192 79644 125248
rect 79700 125192 79768 125248
rect 79824 125192 79892 125248
rect 79948 125192 80078 125248
rect 79078 99372 80078 125192
rect 79078 99316 79148 99372
rect 79204 99316 79272 99372
rect 79328 99316 79396 99372
rect 79452 99316 79520 99372
rect 79576 99316 79644 99372
rect 79700 99316 79768 99372
rect 79824 99316 79892 99372
rect 79948 99316 80078 99372
rect 79078 99248 80078 99316
rect 79078 99192 79148 99248
rect 79204 99192 79272 99248
rect 79328 99192 79396 99248
rect 79452 99192 79520 99248
rect 79576 99192 79644 99248
rect 79700 99192 79768 99248
rect 79824 99192 79892 99248
rect 79948 99192 80078 99248
rect 79078 80008 80078 99192
rect 590840 255372 591840 282572
rect 590840 255316 590970 255372
rect 591026 255316 591094 255372
rect 591150 255316 591218 255372
rect 591274 255316 591342 255372
rect 591398 255316 591466 255372
rect 591522 255316 591590 255372
rect 591646 255316 591714 255372
rect 591770 255316 591840 255372
rect 590840 255248 591840 255316
rect 590840 255192 590970 255248
rect 591026 255192 591094 255248
rect 591150 255192 591218 255248
rect 591274 255192 591342 255248
rect 591398 255192 591466 255248
rect 591522 255192 591590 255248
rect 591646 255192 591714 255248
rect 591770 255192 591840 255248
rect 590840 229372 591840 255192
rect 590840 229316 590970 229372
rect 591026 229316 591094 229372
rect 591150 229316 591218 229372
rect 591274 229316 591342 229372
rect 591398 229316 591466 229372
rect 591522 229316 591590 229372
rect 591646 229316 591714 229372
rect 591770 229316 591840 229372
rect 590840 229248 591840 229316
rect 590840 229192 590970 229248
rect 591026 229192 591094 229248
rect 591150 229192 591218 229248
rect 591274 229192 591342 229248
rect 591398 229192 591466 229248
rect 591522 229192 591590 229248
rect 591646 229192 591714 229248
rect 591770 229192 591840 229248
rect 590840 203372 591840 229192
rect 590840 203316 590970 203372
rect 591026 203316 591094 203372
rect 591150 203316 591218 203372
rect 591274 203316 591342 203372
rect 591398 203316 591466 203372
rect 591522 203316 591590 203372
rect 591646 203316 591714 203372
rect 591770 203316 591840 203372
rect 590840 203248 591840 203316
rect 590840 203192 590970 203248
rect 591026 203192 591094 203248
rect 591150 203192 591218 203248
rect 591274 203192 591342 203248
rect 591398 203192 591466 203248
rect 591522 203192 591590 203248
rect 591646 203192 591714 203248
rect 591770 203192 591840 203248
rect 590840 177372 591840 203192
rect 590840 177316 590970 177372
rect 591026 177316 591094 177372
rect 591150 177316 591218 177372
rect 591274 177316 591342 177372
rect 591398 177316 591466 177372
rect 591522 177316 591590 177372
rect 591646 177316 591714 177372
rect 591770 177316 591840 177372
rect 590840 177248 591840 177316
rect 590840 177192 590970 177248
rect 591026 177192 591094 177248
rect 591150 177192 591218 177248
rect 591274 177192 591342 177248
rect 591398 177192 591466 177248
rect 591522 177192 591590 177248
rect 591646 177192 591714 177248
rect 591770 177192 591840 177248
rect 590840 151372 591840 177192
rect 590840 151316 590970 151372
rect 591026 151316 591094 151372
rect 591150 151316 591218 151372
rect 591274 151316 591342 151372
rect 591398 151316 591466 151372
rect 591522 151316 591590 151372
rect 591646 151316 591714 151372
rect 591770 151316 591840 151372
rect 590840 151248 591840 151316
rect 590840 151192 590970 151248
rect 591026 151192 591094 151248
rect 591150 151192 591218 151248
rect 591274 151192 591342 151248
rect 591398 151192 591466 151248
rect 591522 151192 591590 151248
rect 591646 151192 591714 151248
rect 591770 151192 591840 151248
rect 590840 125372 591840 151192
rect 590840 125316 590970 125372
rect 591026 125316 591094 125372
rect 591150 125316 591218 125372
rect 591274 125316 591342 125372
rect 591398 125316 591466 125372
rect 591522 125316 591590 125372
rect 591646 125316 591714 125372
rect 591770 125316 591840 125372
rect 590840 125248 591840 125316
rect 590840 125192 590970 125248
rect 591026 125192 591094 125248
rect 591150 125192 591218 125248
rect 591274 125192 591342 125248
rect 591398 125192 591466 125248
rect 591522 125192 591590 125248
rect 591646 125192 591714 125248
rect 591770 125192 591840 125248
rect 590840 120137 591840 125192
rect 590840 120081 590959 120137
rect 591015 120081 591259 120137
rect 591315 120081 591559 120137
rect 591615 120081 591840 120137
rect 590840 117029 591840 120081
rect 590840 116973 590959 117029
rect 591015 116973 591259 117029
rect 591315 116973 591559 117029
rect 591615 116973 591840 117029
rect 590840 113921 591840 116973
rect 590840 113865 590959 113921
rect 591015 113865 591259 113921
rect 591315 113865 591559 113921
rect 591615 113865 591840 113921
rect 590840 99372 591840 113865
rect 590840 99316 590970 99372
rect 591026 99316 591094 99372
rect 591150 99316 591218 99372
rect 591274 99316 591342 99372
rect 591398 99316 591466 99372
rect 591522 99316 591590 99372
rect 591646 99316 591714 99372
rect 591770 99316 591840 99372
rect 590840 99248 591840 99316
rect 590840 99192 590970 99248
rect 591026 99192 591094 99248
rect 591150 99192 591218 99248
rect 591274 99192 591342 99248
rect 591398 99192 591466 99248
rect 591522 99192 591590 99248
rect 591646 99192 591714 99248
rect 591770 99192 591840 99248
rect 79078 79952 79208 80008
rect 79264 79952 79332 80008
rect 79388 79952 79456 80008
rect 79512 79952 79580 80008
rect 79636 79952 79704 80008
rect 79760 79952 79828 80008
rect 79884 79952 79952 80008
rect 80008 79952 80078 80008
rect 79078 79884 80078 79952
rect 79078 79828 79208 79884
rect 79264 79828 79332 79884
rect 79388 79828 79456 79884
rect 79512 79828 79580 79884
rect 79636 79828 79704 79884
rect 79760 79828 79828 79884
rect 79884 79828 79952 79884
rect 80008 79828 80078 79884
rect 79078 79760 80078 79828
rect 79078 79704 79208 79760
rect 79264 79704 79332 79760
rect 79388 79704 79456 79760
rect 79512 79704 79580 79760
rect 79636 79704 79704 79760
rect 79760 79704 79828 79760
rect 79884 79704 79952 79760
rect 80008 79704 80078 79760
rect 79078 79636 80078 79704
rect 79078 79580 79208 79636
rect 79264 79580 79332 79636
rect 79388 79580 79456 79636
rect 79512 79580 79580 79636
rect 79636 79580 79704 79636
rect 79760 79580 79828 79636
rect 79884 79580 79952 79636
rect 80008 79580 80078 79636
rect 79078 79512 80078 79580
rect 79078 79456 79208 79512
rect 79264 79456 79332 79512
rect 79388 79456 79456 79512
rect 79512 79456 79580 79512
rect 79636 79456 79704 79512
rect 79760 79456 79828 79512
rect 79884 79456 79952 79512
rect 80008 79456 80078 79512
rect 79078 79388 80078 79456
rect 79078 79332 79208 79388
rect 79264 79332 79332 79388
rect 79388 79332 79456 79388
rect 79512 79332 79580 79388
rect 79636 79332 79704 79388
rect 79760 79332 79828 79388
rect 79884 79332 79952 79388
rect 80008 79332 80078 79388
rect 79078 79264 80078 79332
rect 79078 79208 79208 79264
rect 79264 79208 79332 79264
rect 79388 79208 79456 79264
rect 79512 79208 79580 79264
rect 79636 79208 79704 79264
rect 79760 79208 79828 79264
rect 79884 79208 79952 79264
rect 80008 79208 80078 79264
rect 79078 79078 80078 79208
rect 77678 78552 77808 78608
rect 77864 78552 77932 78608
rect 77988 78552 78056 78608
rect 78112 78552 78180 78608
rect 78236 78552 78304 78608
rect 78360 78552 78428 78608
rect 78484 78552 78552 78608
rect 78608 78552 78678 78608
rect 77678 78484 78678 78552
rect 77678 78428 77808 78484
rect 77864 78428 77932 78484
rect 77988 78428 78056 78484
rect 78112 78428 78180 78484
rect 78236 78428 78304 78484
rect 78360 78428 78428 78484
rect 78484 78428 78552 78484
rect 78608 78428 78678 78484
rect 77678 78360 78678 78428
rect 77678 78304 77808 78360
rect 77864 78304 77932 78360
rect 77988 78304 78056 78360
rect 78112 78304 78180 78360
rect 78236 78304 78304 78360
rect 78360 78304 78428 78360
rect 78484 78304 78552 78360
rect 78608 78304 78678 78360
rect 77678 78236 78678 78304
rect 77678 78180 77808 78236
rect 77864 78180 77932 78236
rect 77988 78180 78056 78236
rect 78112 78180 78180 78236
rect 78236 78180 78304 78236
rect 78360 78180 78428 78236
rect 78484 78180 78552 78236
rect 78608 78180 78678 78236
rect 77678 78112 78678 78180
rect 77678 78056 77808 78112
rect 77864 78056 77932 78112
rect 77988 78056 78056 78112
rect 78112 78056 78180 78112
rect 78236 78056 78304 78112
rect 78360 78056 78428 78112
rect 78484 78056 78552 78112
rect 78608 78056 78678 78112
rect 77678 77988 78678 78056
rect 77678 77932 77808 77988
rect 77864 77932 77932 77988
rect 77988 77932 78056 77988
rect 78112 77932 78180 77988
rect 78236 77932 78304 77988
rect 78360 77932 78428 77988
rect 78484 77932 78552 77988
rect 78608 77932 78678 77988
rect 77678 77864 78678 77932
rect 77678 77808 77808 77864
rect 77864 77808 77932 77864
rect 77988 77808 78056 77864
rect 78112 77808 78180 77864
rect 78236 77808 78304 77864
rect 78360 77808 78428 77864
rect 78484 77808 78552 77864
rect 78608 77808 78678 77864
rect 77678 77678 78678 77808
rect 94224 78608 94544 81752
rect 99224 80008 99544 81752
rect 99224 79952 99294 80008
rect 99350 79952 99418 80008
rect 99474 79952 99544 80008
rect 99224 79884 99544 79952
rect 99224 79828 99294 79884
rect 99350 79828 99418 79884
rect 99474 79828 99544 79884
rect 99224 79760 99544 79828
rect 99224 79704 99294 79760
rect 99350 79704 99418 79760
rect 99474 79704 99544 79760
rect 99224 79636 99544 79704
rect 99224 79580 99294 79636
rect 99350 79580 99418 79636
rect 99474 79580 99544 79636
rect 99224 79512 99544 79580
rect 99224 79456 99294 79512
rect 99350 79456 99418 79512
rect 99474 79456 99544 79512
rect 99224 79388 99544 79456
rect 99224 79332 99294 79388
rect 99350 79332 99418 79388
rect 99474 79332 99544 79388
rect 99224 79264 99544 79332
rect 99224 79208 99294 79264
rect 99350 79208 99418 79264
rect 99474 79208 99544 79264
rect 99224 79078 99544 79208
rect 94224 78552 94294 78608
rect 94350 78552 94418 78608
rect 94474 78552 94544 78608
rect 94224 78484 94544 78552
rect 94224 78428 94294 78484
rect 94350 78428 94418 78484
rect 94474 78428 94544 78484
rect 94224 78360 94544 78428
rect 94224 78304 94294 78360
rect 94350 78304 94418 78360
rect 94474 78304 94544 78360
rect 94224 78236 94544 78304
rect 94224 78180 94294 78236
rect 94350 78180 94418 78236
rect 94474 78180 94544 78236
rect 94224 78112 94544 78180
rect 94224 78056 94294 78112
rect 94350 78056 94418 78112
rect 94474 78056 94544 78112
rect 94224 77988 94544 78056
rect 94224 77932 94294 77988
rect 94350 77932 94418 77988
rect 94474 77932 94544 77988
rect 94224 77864 94544 77932
rect 94224 77808 94294 77864
rect 94350 77808 94418 77864
rect 94474 77808 94544 77864
rect 94224 77678 94544 77808
rect 104224 78608 104544 81752
rect 104224 78552 104294 78608
rect 104350 78552 104418 78608
rect 104474 78552 104544 78608
rect 104224 78484 104544 78552
rect 104224 78428 104294 78484
rect 104350 78428 104418 78484
rect 104474 78428 104544 78484
rect 104224 78360 104544 78428
rect 104224 78304 104294 78360
rect 104350 78304 104418 78360
rect 104474 78304 104544 78360
rect 104224 78236 104544 78304
rect 104224 78180 104294 78236
rect 104350 78180 104418 78236
rect 104474 78180 104544 78236
rect 104224 78112 104544 78180
rect 104224 78056 104294 78112
rect 104350 78056 104418 78112
rect 104474 78056 104544 78112
rect 104224 77988 104544 78056
rect 104224 77932 104294 77988
rect 104350 77932 104418 77988
rect 104474 77932 104544 77988
rect 104224 77864 104544 77932
rect 104224 77808 104294 77864
rect 104350 77808 104418 77864
rect 104474 77808 104544 77864
rect 104224 77678 104544 77808
rect 107272 80008 109172 80078
rect 107272 79952 107330 80008
rect 107386 79952 107454 80008
rect 107510 79952 107578 80008
rect 107634 79952 107702 80008
rect 107758 79952 107826 80008
rect 107882 79952 107950 80008
rect 108006 79952 108074 80008
rect 108130 79952 108198 80008
rect 108254 79952 108322 80008
rect 108378 79952 108446 80008
rect 108502 79952 108570 80008
rect 108626 79952 108694 80008
rect 108750 79952 108818 80008
rect 108874 79952 108942 80008
rect 108998 79952 109066 80008
rect 109122 79952 109172 80008
rect 107272 79884 109172 79952
rect 107272 79828 107330 79884
rect 107386 79828 107454 79884
rect 107510 79828 107578 79884
rect 107634 79828 107702 79884
rect 107758 79828 107826 79884
rect 107882 79828 107950 79884
rect 108006 79828 108074 79884
rect 108130 79828 108198 79884
rect 108254 79828 108322 79884
rect 108378 79828 108446 79884
rect 108502 79828 108570 79884
rect 108626 79828 108694 79884
rect 108750 79828 108818 79884
rect 108874 79828 108942 79884
rect 108998 79828 109066 79884
rect 109122 79828 109172 79884
rect 107272 79760 109172 79828
rect 107272 79704 107330 79760
rect 107386 79704 107454 79760
rect 107510 79704 107578 79760
rect 107634 79704 107702 79760
rect 107758 79704 107826 79760
rect 107882 79704 107950 79760
rect 108006 79704 108074 79760
rect 108130 79704 108198 79760
rect 108254 79704 108322 79760
rect 108378 79704 108446 79760
rect 108502 79704 108570 79760
rect 108626 79704 108694 79760
rect 108750 79704 108818 79760
rect 108874 79704 108942 79760
rect 108998 79704 109066 79760
rect 109122 79704 109172 79760
rect 107272 79636 109172 79704
rect 107272 79580 107330 79636
rect 107386 79580 107454 79636
rect 107510 79580 107578 79636
rect 107634 79580 107702 79636
rect 107758 79580 107826 79636
rect 107882 79580 107950 79636
rect 108006 79580 108074 79636
rect 108130 79580 108198 79636
rect 108254 79580 108322 79636
rect 108378 79580 108446 79636
rect 108502 79580 108570 79636
rect 108626 79580 108694 79636
rect 108750 79580 108818 79636
rect 108874 79580 108942 79636
rect 108998 79580 109066 79636
rect 109122 79580 109172 79636
rect 107272 79512 109172 79580
rect 107272 79456 107330 79512
rect 107386 79456 107454 79512
rect 107510 79456 107578 79512
rect 107634 79456 107702 79512
rect 107758 79456 107826 79512
rect 107882 79456 107950 79512
rect 108006 79456 108074 79512
rect 108130 79456 108198 79512
rect 108254 79456 108322 79512
rect 108378 79456 108446 79512
rect 108502 79456 108570 79512
rect 108626 79456 108694 79512
rect 108750 79456 108818 79512
rect 108874 79456 108942 79512
rect 108998 79456 109066 79512
rect 109122 79456 109172 79512
rect 107272 79388 109172 79456
rect 107272 79332 107330 79388
rect 107386 79332 107454 79388
rect 107510 79332 107578 79388
rect 107634 79332 107702 79388
rect 107758 79332 107826 79388
rect 107882 79332 107950 79388
rect 108006 79332 108074 79388
rect 108130 79332 108198 79388
rect 108254 79332 108322 79388
rect 108378 79332 108446 79388
rect 108502 79332 108570 79388
rect 108626 79332 108694 79388
rect 108750 79332 108818 79388
rect 108874 79332 108942 79388
rect 108998 79332 109066 79388
rect 109122 79332 109172 79388
rect 107272 79264 109172 79332
rect 107272 79208 107330 79264
rect 107386 79208 107454 79264
rect 107510 79208 107578 79264
rect 107634 79208 107702 79264
rect 107758 79208 107826 79264
rect 107882 79208 107950 79264
rect 108006 79208 108074 79264
rect 108130 79208 108198 79264
rect 108254 79208 108322 79264
rect 108378 79208 108446 79264
rect 108502 79208 108570 79264
rect 108626 79208 108694 79264
rect 108750 79208 108818 79264
rect 108874 79208 108942 79264
rect 108998 79208 109066 79264
rect 109122 79208 109172 79264
rect 107272 70130 109172 79208
rect 107272 70074 107342 70130
rect 107398 70074 107466 70130
rect 107522 70074 107590 70130
rect 107646 70074 107714 70130
rect 107770 70074 107838 70130
rect 107894 70074 107962 70130
rect 108018 70074 108086 70130
rect 108142 70074 108210 70130
rect 108266 70074 108334 70130
rect 108390 70074 108458 70130
rect 108514 70074 108582 70130
rect 108638 70074 108706 70130
rect 108762 70074 108830 70130
rect 108886 70074 108954 70130
rect 109010 70074 109078 70130
rect 109134 70074 109172 70130
rect 107272 70000 109172 70074
rect 109752 80008 111802 80078
rect 109752 79952 109810 80008
rect 109866 79952 109934 80008
rect 109990 79952 110058 80008
rect 110114 79952 110182 80008
rect 110238 79952 110306 80008
rect 110362 79952 110430 80008
rect 110486 79952 110554 80008
rect 110610 79952 110678 80008
rect 110734 79952 110802 80008
rect 110858 79952 110926 80008
rect 110982 79952 111050 80008
rect 111106 79952 111174 80008
rect 111230 79952 111298 80008
rect 111354 79952 111422 80008
rect 111478 79952 111546 80008
rect 111602 79952 111670 80008
rect 111726 79952 111802 80008
rect 109752 79884 111802 79952
rect 109752 79828 109810 79884
rect 109866 79828 109934 79884
rect 109990 79828 110058 79884
rect 110114 79828 110182 79884
rect 110238 79828 110306 79884
rect 110362 79828 110430 79884
rect 110486 79828 110554 79884
rect 110610 79828 110678 79884
rect 110734 79828 110802 79884
rect 110858 79828 110926 79884
rect 110982 79828 111050 79884
rect 111106 79828 111174 79884
rect 111230 79828 111298 79884
rect 111354 79828 111422 79884
rect 111478 79828 111546 79884
rect 111602 79828 111670 79884
rect 111726 79828 111802 79884
rect 109752 79760 111802 79828
rect 109752 79704 109810 79760
rect 109866 79704 109934 79760
rect 109990 79704 110058 79760
rect 110114 79704 110182 79760
rect 110238 79704 110306 79760
rect 110362 79704 110430 79760
rect 110486 79704 110554 79760
rect 110610 79704 110678 79760
rect 110734 79704 110802 79760
rect 110858 79704 110926 79760
rect 110982 79704 111050 79760
rect 111106 79704 111174 79760
rect 111230 79704 111298 79760
rect 111354 79704 111422 79760
rect 111478 79704 111546 79760
rect 111602 79704 111670 79760
rect 111726 79704 111802 79760
rect 109752 79636 111802 79704
rect 109752 79580 109810 79636
rect 109866 79580 109934 79636
rect 109990 79580 110058 79636
rect 110114 79580 110182 79636
rect 110238 79580 110306 79636
rect 110362 79580 110430 79636
rect 110486 79580 110554 79636
rect 110610 79580 110678 79636
rect 110734 79580 110802 79636
rect 110858 79580 110926 79636
rect 110982 79580 111050 79636
rect 111106 79580 111174 79636
rect 111230 79580 111298 79636
rect 111354 79580 111422 79636
rect 111478 79580 111546 79636
rect 111602 79580 111670 79636
rect 111726 79580 111802 79636
rect 109752 79512 111802 79580
rect 109752 79456 109810 79512
rect 109866 79456 109934 79512
rect 109990 79456 110058 79512
rect 110114 79456 110182 79512
rect 110238 79456 110306 79512
rect 110362 79456 110430 79512
rect 110486 79456 110554 79512
rect 110610 79456 110678 79512
rect 110734 79456 110802 79512
rect 110858 79456 110926 79512
rect 110982 79456 111050 79512
rect 111106 79456 111174 79512
rect 111230 79456 111298 79512
rect 111354 79456 111422 79512
rect 111478 79456 111546 79512
rect 111602 79456 111670 79512
rect 111726 79456 111802 79512
rect 109752 79388 111802 79456
rect 109752 79332 109810 79388
rect 109866 79332 109934 79388
rect 109990 79332 110058 79388
rect 110114 79332 110182 79388
rect 110238 79332 110306 79388
rect 110362 79332 110430 79388
rect 110486 79332 110554 79388
rect 110610 79332 110678 79388
rect 110734 79332 110802 79388
rect 110858 79332 110926 79388
rect 110982 79332 111050 79388
rect 111106 79332 111174 79388
rect 111230 79332 111298 79388
rect 111354 79332 111422 79388
rect 111478 79332 111546 79388
rect 111602 79332 111670 79388
rect 111726 79332 111802 79388
rect 109752 79264 111802 79332
rect 109752 79208 109810 79264
rect 109866 79208 109934 79264
rect 109990 79208 110058 79264
rect 110114 79208 110182 79264
rect 110238 79208 110306 79264
rect 110362 79208 110430 79264
rect 110486 79208 110554 79264
rect 110610 79208 110678 79264
rect 110734 79208 110802 79264
rect 110858 79208 110926 79264
rect 110982 79208 111050 79264
rect 111106 79208 111174 79264
rect 111230 79208 111298 79264
rect 111354 79208 111422 79264
rect 111478 79208 111546 79264
rect 111602 79208 111670 79264
rect 111726 79208 111802 79264
rect 109752 70130 111802 79208
rect 109752 70074 109822 70130
rect 109878 70074 109946 70130
rect 110002 70074 110070 70130
rect 110126 70074 110194 70130
rect 110250 70074 110318 70130
rect 110374 70074 110442 70130
rect 110498 70074 110566 70130
rect 110622 70074 110690 70130
rect 110746 70074 110814 70130
rect 110870 70074 110938 70130
rect 110994 70074 111062 70130
rect 111118 70074 111186 70130
rect 111242 70074 111310 70130
rect 111366 70074 111434 70130
rect 111490 70074 111558 70130
rect 111614 70074 111682 70130
rect 111738 70074 111802 70130
rect 109752 70000 111802 70074
rect 112122 80008 114172 80078
rect 112122 79952 112180 80008
rect 112236 79952 112304 80008
rect 112360 79952 112428 80008
rect 112484 79952 112552 80008
rect 112608 79952 112676 80008
rect 112732 79952 112800 80008
rect 112856 79952 112924 80008
rect 112980 79952 113048 80008
rect 113104 79952 113172 80008
rect 113228 79952 113296 80008
rect 113352 79952 113420 80008
rect 113476 79952 113544 80008
rect 113600 79952 113668 80008
rect 113724 79952 113792 80008
rect 113848 79952 113916 80008
rect 113972 79952 114040 80008
rect 114096 79952 114172 80008
rect 112122 79884 114172 79952
rect 112122 79828 112180 79884
rect 112236 79828 112304 79884
rect 112360 79828 112428 79884
rect 112484 79828 112552 79884
rect 112608 79828 112676 79884
rect 112732 79828 112800 79884
rect 112856 79828 112924 79884
rect 112980 79828 113048 79884
rect 113104 79828 113172 79884
rect 113228 79828 113296 79884
rect 113352 79828 113420 79884
rect 113476 79828 113544 79884
rect 113600 79828 113668 79884
rect 113724 79828 113792 79884
rect 113848 79828 113916 79884
rect 113972 79828 114040 79884
rect 114096 79828 114172 79884
rect 112122 79760 114172 79828
rect 112122 79704 112180 79760
rect 112236 79704 112304 79760
rect 112360 79704 112428 79760
rect 112484 79704 112552 79760
rect 112608 79704 112676 79760
rect 112732 79704 112800 79760
rect 112856 79704 112924 79760
rect 112980 79704 113048 79760
rect 113104 79704 113172 79760
rect 113228 79704 113296 79760
rect 113352 79704 113420 79760
rect 113476 79704 113544 79760
rect 113600 79704 113668 79760
rect 113724 79704 113792 79760
rect 113848 79704 113916 79760
rect 113972 79704 114040 79760
rect 114096 79704 114172 79760
rect 112122 79636 114172 79704
rect 112122 79580 112180 79636
rect 112236 79580 112304 79636
rect 112360 79580 112428 79636
rect 112484 79580 112552 79636
rect 112608 79580 112676 79636
rect 112732 79580 112800 79636
rect 112856 79580 112924 79636
rect 112980 79580 113048 79636
rect 113104 79580 113172 79636
rect 113228 79580 113296 79636
rect 113352 79580 113420 79636
rect 113476 79580 113544 79636
rect 113600 79580 113668 79636
rect 113724 79580 113792 79636
rect 113848 79580 113916 79636
rect 113972 79580 114040 79636
rect 114096 79580 114172 79636
rect 112122 79512 114172 79580
rect 112122 79456 112180 79512
rect 112236 79456 112304 79512
rect 112360 79456 112428 79512
rect 112484 79456 112552 79512
rect 112608 79456 112676 79512
rect 112732 79456 112800 79512
rect 112856 79456 112924 79512
rect 112980 79456 113048 79512
rect 113104 79456 113172 79512
rect 113228 79456 113296 79512
rect 113352 79456 113420 79512
rect 113476 79456 113544 79512
rect 113600 79456 113668 79512
rect 113724 79456 113792 79512
rect 113848 79456 113916 79512
rect 113972 79456 114040 79512
rect 114096 79456 114172 79512
rect 112122 79388 114172 79456
rect 112122 79332 112180 79388
rect 112236 79332 112304 79388
rect 112360 79332 112428 79388
rect 112484 79332 112552 79388
rect 112608 79332 112676 79388
rect 112732 79332 112800 79388
rect 112856 79332 112924 79388
rect 112980 79332 113048 79388
rect 113104 79332 113172 79388
rect 113228 79332 113296 79388
rect 113352 79332 113420 79388
rect 113476 79332 113544 79388
rect 113600 79332 113668 79388
rect 113724 79332 113792 79388
rect 113848 79332 113916 79388
rect 113972 79332 114040 79388
rect 114096 79332 114172 79388
rect 112122 79264 114172 79332
rect 112122 79208 112180 79264
rect 112236 79208 112304 79264
rect 112360 79208 112428 79264
rect 112484 79208 112552 79264
rect 112608 79208 112676 79264
rect 112732 79208 112800 79264
rect 112856 79208 112924 79264
rect 112980 79208 113048 79264
rect 113104 79208 113172 79264
rect 113228 79208 113296 79264
rect 113352 79208 113420 79264
rect 113476 79208 113544 79264
rect 113600 79208 113668 79264
rect 113724 79208 113792 79264
rect 113848 79208 113916 79264
rect 113972 79208 114040 79264
rect 114096 79208 114172 79264
rect 112122 70130 114172 79208
rect 112122 70074 112192 70130
rect 112248 70074 112316 70130
rect 112372 70074 112440 70130
rect 112496 70074 112564 70130
rect 112620 70074 112688 70130
rect 112744 70074 112812 70130
rect 112868 70074 112936 70130
rect 112992 70074 113060 70130
rect 113116 70074 113184 70130
rect 113240 70074 113308 70130
rect 113364 70074 113432 70130
rect 113488 70074 113556 70130
rect 113612 70074 113680 70130
rect 113736 70074 113804 70130
rect 113860 70074 113928 70130
rect 113984 70074 114052 70130
rect 114108 70074 114172 70130
rect 112122 70000 114172 70074
rect 114828 80008 116878 80078
rect 114828 79952 114886 80008
rect 114942 79952 115010 80008
rect 115066 79952 115134 80008
rect 115190 79952 115258 80008
rect 115314 79952 115382 80008
rect 115438 79952 115506 80008
rect 115562 79952 115630 80008
rect 115686 79952 115754 80008
rect 115810 79952 115878 80008
rect 115934 79952 116002 80008
rect 116058 79952 116126 80008
rect 116182 79952 116250 80008
rect 116306 79952 116374 80008
rect 116430 79952 116498 80008
rect 116554 79952 116622 80008
rect 116678 79952 116746 80008
rect 116802 79952 116878 80008
rect 114828 79884 116878 79952
rect 114828 79828 114886 79884
rect 114942 79828 115010 79884
rect 115066 79828 115134 79884
rect 115190 79828 115258 79884
rect 115314 79828 115382 79884
rect 115438 79828 115506 79884
rect 115562 79828 115630 79884
rect 115686 79828 115754 79884
rect 115810 79828 115878 79884
rect 115934 79828 116002 79884
rect 116058 79828 116126 79884
rect 116182 79828 116250 79884
rect 116306 79828 116374 79884
rect 116430 79828 116498 79884
rect 116554 79828 116622 79884
rect 116678 79828 116746 79884
rect 116802 79828 116878 79884
rect 114828 79760 116878 79828
rect 114828 79704 114886 79760
rect 114942 79704 115010 79760
rect 115066 79704 115134 79760
rect 115190 79704 115258 79760
rect 115314 79704 115382 79760
rect 115438 79704 115506 79760
rect 115562 79704 115630 79760
rect 115686 79704 115754 79760
rect 115810 79704 115878 79760
rect 115934 79704 116002 79760
rect 116058 79704 116126 79760
rect 116182 79704 116250 79760
rect 116306 79704 116374 79760
rect 116430 79704 116498 79760
rect 116554 79704 116622 79760
rect 116678 79704 116746 79760
rect 116802 79704 116878 79760
rect 114828 79636 116878 79704
rect 114828 79580 114886 79636
rect 114942 79580 115010 79636
rect 115066 79580 115134 79636
rect 115190 79580 115258 79636
rect 115314 79580 115382 79636
rect 115438 79580 115506 79636
rect 115562 79580 115630 79636
rect 115686 79580 115754 79636
rect 115810 79580 115878 79636
rect 115934 79580 116002 79636
rect 116058 79580 116126 79636
rect 116182 79580 116250 79636
rect 116306 79580 116374 79636
rect 116430 79580 116498 79636
rect 116554 79580 116622 79636
rect 116678 79580 116746 79636
rect 116802 79580 116878 79636
rect 114828 79512 116878 79580
rect 114828 79456 114886 79512
rect 114942 79456 115010 79512
rect 115066 79456 115134 79512
rect 115190 79456 115258 79512
rect 115314 79456 115382 79512
rect 115438 79456 115506 79512
rect 115562 79456 115630 79512
rect 115686 79456 115754 79512
rect 115810 79456 115878 79512
rect 115934 79456 116002 79512
rect 116058 79456 116126 79512
rect 116182 79456 116250 79512
rect 116306 79456 116374 79512
rect 116430 79456 116498 79512
rect 116554 79456 116622 79512
rect 116678 79456 116746 79512
rect 116802 79456 116878 79512
rect 114828 79388 116878 79456
rect 114828 79332 114886 79388
rect 114942 79332 115010 79388
rect 115066 79332 115134 79388
rect 115190 79332 115258 79388
rect 115314 79332 115382 79388
rect 115438 79332 115506 79388
rect 115562 79332 115630 79388
rect 115686 79332 115754 79388
rect 115810 79332 115878 79388
rect 115934 79332 116002 79388
rect 116058 79332 116126 79388
rect 116182 79332 116250 79388
rect 116306 79332 116374 79388
rect 116430 79332 116498 79388
rect 116554 79332 116622 79388
rect 116678 79332 116746 79388
rect 116802 79332 116878 79388
rect 114828 79264 116878 79332
rect 114828 79208 114886 79264
rect 114942 79208 115010 79264
rect 115066 79208 115134 79264
rect 115190 79208 115258 79264
rect 115314 79208 115382 79264
rect 115438 79208 115506 79264
rect 115562 79208 115630 79264
rect 115686 79208 115754 79264
rect 115810 79208 115878 79264
rect 115934 79208 116002 79264
rect 116058 79208 116126 79264
rect 116182 79208 116250 79264
rect 116306 79208 116374 79264
rect 116430 79208 116498 79264
rect 116554 79208 116622 79264
rect 116678 79208 116746 79264
rect 116802 79208 116878 79264
rect 114828 70130 116878 79208
rect 114828 70074 114892 70130
rect 114948 70074 115016 70130
rect 115072 70074 115140 70130
rect 115196 70074 115264 70130
rect 115320 70074 115388 70130
rect 115444 70074 115512 70130
rect 115568 70074 115636 70130
rect 115692 70074 115760 70130
rect 115816 70074 115884 70130
rect 115940 70074 116008 70130
rect 116064 70074 116132 70130
rect 116188 70074 116256 70130
rect 116312 70074 116380 70130
rect 116436 70074 116504 70130
rect 116560 70074 116628 70130
rect 116684 70074 116752 70130
rect 116808 70074 116878 70130
rect 114828 70000 116878 70074
rect 117198 80008 119248 80078
rect 117198 79952 117256 80008
rect 117312 79952 117380 80008
rect 117436 79952 117504 80008
rect 117560 79952 117628 80008
rect 117684 79952 117752 80008
rect 117808 79952 117876 80008
rect 117932 79952 118000 80008
rect 118056 79952 118124 80008
rect 118180 79952 118248 80008
rect 118304 79952 118372 80008
rect 118428 79952 118496 80008
rect 118552 79952 118620 80008
rect 118676 79952 118744 80008
rect 118800 79952 118868 80008
rect 118924 79952 118992 80008
rect 119048 79952 119116 80008
rect 119172 79952 119248 80008
rect 117198 79884 119248 79952
rect 117198 79828 117256 79884
rect 117312 79828 117380 79884
rect 117436 79828 117504 79884
rect 117560 79828 117628 79884
rect 117684 79828 117752 79884
rect 117808 79828 117876 79884
rect 117932 79828 118000 79884
rect 118056 79828 118124 79884
rect 118180 79828 118248 79884
rect 118304 79828 118372 79884
rect 118428 79828 118496 79884
rect 118552 79828 118620 79884
rect 118676 79828 118744 79884
rect 118800 79828 118868 79884
rect 118924 79828 118992 79884
rect 119048 79828 119116 79884
rect 119172 79828 119248 79884
rect 117198 79760 119248 79828
rect 117198 79704 117256 79760
rect 117312 79704 117380 79760
rect 117436 79704 117504 79760
rect 117560 79704 117628 79760
rect 117684 79704 117752 79760
rect 117808 79704 117876 79760
rect 117932 79704 118000 79760
rect 118056 79704 118124 79760
rect 118180 79704 118248 79760
rect 118304 79704 118372 79760
rect 118428 79704 118496 79760
rect 118552 79704 118620 79760
rect 118676 79704 118744 79760
rect 118800 79704 118868 79760
rect 118924 79704 118992 79760
rect 119048 79704 119116 79760
rect 119172 79704 119248 79760
rect 117198 79636 119248 79704
rect 117198 79580 117256 79636
rect 117312 79580 117380 79636
rect 117436 79580 117504 79636
rect 117560 79580 117628 79636
rect 117684 79580 117752 79636
rect 117808 79580 117876 79636
rect 117932 79580 118000 79636
rect 118056 79580 118124 79636
rect 118180 79580 118248 79636
rect 118304 79580 118372 79636
rect 118428 79580 118496 79636
rect 118552 79580 118620 79636
rect 118676 79580 118744 79636
rect 118800 79580 118868 79636
rect 118924 79580 118992 79636
rect 119048 79580 119116 79636
rect 119172 79580 119248 79636
rect 117198 79512 119248 79580
rect 117198 79456 117256 79512
rect 117312 79456 117380 79512
rect 117436 79456 117504 79512
rect 117560 79456 117628 79512
rect 117684 79456 117752 79512
rect 117808 79456 117876 79512
rect 117932 79456 118000 79512
rect 118056 79456 118124 79512
rect 118180 79456 118248 79512
rect 118304 79456 118372 79512
rect 118428 79456 118496 79512
rect 118552 79456 118620 79512
rect 118676 79456 118744 79512
rect 118800 79456 118868 79512
rect 118924 79456 118992 79512
rect 119048 79456 119116 79512
rect 119172 79456 119248 79512
rect 117198 79388 119248 79456
rect 117198 79332 117256 79388
rect 117312 79332 117380 79388
rect 117436 79332 117504 79388
rect 117560 79332 117628 79388
rect 117684 79332 117752 79388
rect 117808 79332 117876 79388
rect 117932 79332 118000 79388
rect 118056 79332 118124 79388
rect 118180 79332 118248 79388
rect 118304 79332 118372 79388
rect 118428 79332 118496 79388
rect 118552 79332 118620 79388
rect 118676 79332 118744 79388
rect 118800 79332 118868 79388
rect 118924 79332 118992 79388
rect 119048 79332 119116 79388
rect 119172 79332 119248 79388
rect 117198 79264 119248 79332
rect 117198 79208 117256 79264
rect 117312 79208 117380 79264
rect 117436 79208 117504 79264
rect 117560 79208 117628 79264
rect 117684 79208 117752 79264
rect 117808 79208 117876 79264
rect 117932 79208 118000 79264
rect 118056 79208 118124 79264
rect 118180 79208 118248 79264
rect 118304 79208 118372 79264
rect 118428 79208 118496 79264
rect 118552 79208 118620 79264
rect 118676 79208 118744 79264
rect 118800 79208 118868 79264
rect 118924 79208 118992 79264
rect 119048 79208 119116 79264
rect 119172 79208 119248 79264
rect 117198 70130 119248 79208
rect 117198 70074 117262 70130
rect 117318 70074 117386 70130
rect 117442 70074 117510 70130
rect 117566 70074 117634 70130
rect 117690 70074 117758 70130
rect 117814 70074 117882 70130
rect 117938 70074 118006 70130
rect 118062 70074 118130 70130
rect 118186 70074 118254 70130
rect 118310 70074 118378 70130
rect 118434 70074 118502 70130
rect 118558 70074 118626 70130
rect 118682 70074 118750 70130
rect 118806 70074 118874 70130
rect 118930 70074 118998 70130
rect 119054 70074 119122 70130
rect 119178 70074 119248 70130
rect 117198 70000 119248 70074
rect 119828 80008 121728 80078
rect 119828 79952 119860 80008
rect 119916 79952 119984 80008
rect 120040 79952 120108 80008
rect 120164 79952 120232 80008
rect 120288 79952 120356 80008
rect 120412 79952 120480 80008
rect 120536 79952 120604 80008
rect 120660 79952 120728 80008
rect 120784 79952 120852 80008
rect 120908 79952 120976 80008
rect 121032 79952 121100 80008
rect 121156 79952 121224 80008
rect 121280 79952 121348 80008
rect 121404 79952 121472 80008
rect 121528 79952 121596 80008
rect 121652 79952 121728 80008
rect 119828 79884 121728 79952
rect 119828 79828 119860 79884
rect 119916 79828 119984 79884
rect 120040 79828 120108 79884
rect 120164 79828 120232 79884
rect 120288 79828 120356 79884
rect 120412 79828 120480 79884
rect 120536 79828 120604 79884
rect 120660 79828 120728 79884
rect 120784 79828 120852 79884
rect 120908 79828 120976 79884
rect 121032 79828 121100 79884
rect 121156 79828 121224 79884
rect 121280 79828 121348 79884
rect 121404 79828 121472 79884
rect 121528 79828 121596 79884
rect 121652 79828 121728 79884
rect 119828 79760 121728 79828
rect 119828 79704 119860 79760
rect 119916 79704 119984 79760
rect 120040 79704 120108 79760
rect 120164 79704 120232 79760
rect 120288 79704 120356 79760
rect 120412 79704 120480 79760
rect 120536 79704 120604 79760
rect 120660 79704 120728 79760
rect 120784 79704 120852 79760
rect 120908 79704 120976 79760
rect 121032 79704 121100 79760
rect 121156 79704 121224 79760
rect 121280 79704 121348 79760
rect 121404 79704 121472 79760
rect 121528 79704 121596 79760
rect 121652 79704 121728 79760
rect 119828 79636 121728 79704
rect 119828 79580 119860 79636
rect 119916 79580 119984 79636
rect 120040 79580 120108 79636
rect 120164 79580 120232 79636
rect 120288 79580 120356 79636
rect 120412 79580 120480 79636
rect 120536 79580 120604 79636
rect 120660 79580 120728 79636
rect 120784 79580 120852 79636
rect 120908 79580 120976 79636
rect 121032 79580 121100 79636
rect 121156 79580 121224 79636
rect 121280 79580 121348 79636
rect 121404 79580 121472 79636
rect 121528 79580 121596 79636
rect 121652 79580 121728 79636
rect 119828 79512 121728 79580
rect 119828 79456 119860 79512
rect 119916 79456 119984 79512
rect 120040 79456 120108 79512
rect 120164 79456 120232 79512
rect 120288 79456 120356 79512
rect 120412 79456 120480 79512
rect 120536 79456 120604 79512
rect 120660 79456 120728 79512
rect 120784 79456 120852 79512
rect 120908 79456 120976 79512
rect 121032 79456 121100 79512
rect 121156 79456 121224 79512
rect 121280 79456 121348 79512
rect 121404 79456 121472 79512
rect 121528 79456 121596 79512
rect 121652 79456 121728 79512
rect 119828 79388 121728 79456
rect 119828 79332 119860 79388
rect 119916 79332 119984 79388
rect 120040 79332 120108 79388
rect 120164 79332 120232 79388
rect 120288 79332 120356 79388
rect 120412 79332 120480 79388
rect 120536 79332 120604 79388
rect 120660 79332 120728 79388
rect 120784 79332 120852 79388
rect 120908 79332 120976 79388
rect 121032 79332 121100 79388
rect 121156 79332 121224 79388
rect 121280 79332 121348 79388
rect 121404 79332 121472 79388
rect 121528 79332 121596 79388
rect 121652 79332 121728 79388
rect 119828 79264 121728 79332
rect 119828 79208 119860 79264
rect 119916 79208 119984 79264
rect 120040 79208 120108 79264
rect 120164 79208 120232 79264
rect 120288 79208 120356 79264
rect 120412 79208 120480 79264
rect 120536 79208 120604 79264
rect 120660 79208 120728 79264
rect 120784 79208 120852 79264
rect 120908 79208 120976 79264
rect 121032 79208 121100 79264
rect 121156 79208 121224 79264
rect 121280 79208 121348 79264
rect 121404 79208 121472 79264
rect 121528 79208 121596 79264
rect 121652 79208 121728 79264
rect 119828 70130 121728 79208
rect 124224 78608 124544 81752
rect 129224 80008 129544 81752
rect 129224 79952 129294 80008
rect 129350 79952 129418 80008
rect 129474 79952 129544 80008
rect 129224 79884 129544 79952
rect 129224 79828 129294 79884
rect 129350 79828 129418 79884
rect 129474 79828 129544 79884
rect 129224 79760 129544 79828
rect 129224 79704 129294 79760
rect 129350 79704 129418 79760
rect 129474 79704 129544 79760
rect 129224 79636 129544 79704
rect 129224 79580 129294 79636
rect 129350 79580 129418 79636
rect 129474 79580 129544 79636
rect 129224 79512 129544 79580
rect 129224 79456 129294 79512
rect 129350 79456 129418 79512
rect 129474 79456 129544 79512
rect 129224 79388 129544 79456
rect 129224 79332 129294 79388
rect 129350 79332 129418 79388
rect 129474 79332 129544 79388
rect 129224 79264 129544 79332
rect 129224 79208 129294 79264
rect 129350 79208 129418 79264
rect 129474 79208 129544 79264
rect 129224 79078 129544 79208
rect 124224 78552 124294 78608
rect 124350 78552 124418 78608
rect 124474 78552 124544 78608
rect 124224 78484 124544 78552
rect 124224 78428 124294 78484
rect 124350 78428 124418 78484
rect 124474 78428 124544 78484
rect 124224 78360 124544 78428
rect 124224 78304 124294 78360
rect 124350 78304 124418 78360
rect 124474 78304 124544 78360
rect 124224 78236 124544 78304
rect 124224 78180 124294 78236
rect 124350 78180 124418 78236
rect 124474 78180 124544 78236
rect 124224 78112 124544 78180
rect 124224 78056 124294 78112
rect 124350 78056 124418 78112
rect 124474 78056 124544 78112
rect 124224 77988 124544 78056
rect 124224 77932 124294 77988
rect 124350 77932 124418 77988
rect 124474 77932 124544 77988
rect 124224 77864 124544 77932
rect 124224 77808 124294 77864
rect 124350 77808 124418 77864
rect 124474 77808 124544 77864
rect 124224 77678 124544 77808
rect 134224 78608 134544 81752
rect 139224 80008 139544 81752
rect 139224 79952 139294 80008
rect 139350 79952 139418 80008
rect 139474 79952 139544 80008
rect 139224 79884 139544 79952
rect 139224 79828 139294 79884
rect 139350 79828 139418 79884
rect 139474 79828 139544 79884
rect 139224 79760 139544 79828
rect 139224 79704 139294 79760
rect 139350 79704 139418 79760
rect 139474 79704 139544 79760
rect 139224 79636 139544 79704
rect 139224 79580 139294 79636
rect 139350 79580 139418 79636
rect 139474 79580 139544 79636
rect 139224 79512 139544 79580
rect 139224 79456 139294 79512
rect 139350 79456 139418 79512
rect 139474 79456 139544 79512
rect 139224 79388 139544 79456
rect 139224 79332 139294 79388
rect 139350 79332 139418 79388
rect 139474 79332 139544 79388
rect 139224 79264 139544 79332
rect 139224 79208 139294 79264
rect 139350 79208 139418 79264
rect 139474 79208 139544 79264
rect 139224 79078 139544 79208
rect 134224 78552 134294 78608
rect 134350 78552 134418 78608
rect 134474 78552 134544 78608
rect 134224 78484 134544 78552
rect 134224 78428 134294 78484
rect 134350 78428 134418 78484
rect 134474 78428 134544 78484
rect 134224 78360 134544 78428
rect 134224 78304 134294 78360
rect 134350 78304 134418 78360
rect 134474 78304 134544 78360
rect 134224 78236 134544 78304
rect 134224 78180 134294 78236
rect 134350 78180 134418 78236
rect 134474 78180 134544 78236
rect 134224 78112 134544 78180
rect 134224 78056 134294 78112
rect 134350 78056 134418 78112
rect 134474 78056 134544 78112
rect 134224 77988 134544 78056
rect 134224 77932 134294 77988
rect 134350 77932 134418 77988
rect 134474 77932 134544 77988
rect 134224 77864 134544 77932
rect 134224 77808 134294 77864
rect 134350 77808 134418 77864
rect 134474 77808 134544 77864
rect 134224 77678 134544 77808
rect 144224 78608 144544 81752
rect 149224 80008 149544 81752
rect 149224 79952 149294 80008
rect 149350 79952 149418 80008
rect 149474 79952 149544 80008
rect 149224 79884 149544 79952
rect 149224 79828 149294 79884
rect 149350 79828 149418 79884
rect 149474 79828 149544 79884
rect 149224 79760 149544 79828
rect 149224 79704 149294 79760
rect 149350 79704 149418 79760
rect 149474 79704 149544 79760
rect 149224 79636 149544 79704
rect 149224 79580 149294 79636
rect 149350 79580 149418 79636
rect 149474 79580 149544 79636
rect 149224 79512 149544 79580
rect 149224 79456 149294 79512
rect 149350 79456 149418 79512
rect 149474 79456 149544 79512
rect 149224 79388 149544 79456
rect 149224 79332 149294 79388
rect 149350 79332 149418 79388
rect 149474 79332 149544 79388
rect 149224 79264 149544 79332
rect 149224 79208 149294 79264
rect 149350 79208 149418 79264
rect 149474 79208 149544 79264
rect 149224 79078 149544 79208
rect 144224 78552 144294 78608
rect 144350 78552 144418 78608
rect 144474 78552 144544 78608
rect 144224 78484 144544 78552
rect 144224 78428 144294 78484
rect 144350 78428 144418 78484
rect 144474 78428 144544 78484
rect 144224 78360 144544 78428
rect 144224 78304 144294 78360
rect 144350 78304 144418 78360
rect 144474 78304 144544 78360
rect 144224 78236 144544 78304
rect 144224 78180 144294 78236
rect 144350 78180 144418 78236
rect 144474 78180 144544 78236
rect 144224 78112 144544 78180
rect 144224 78056 144294 78112
rect 144350 78056 144418 78112
rect 144474 78056 144544 78112
rect 144224 77988 144544 78056
rect 144224 77932 144294 77988
rect 144350 77932 144418 77988
rect 144474 77932 144544 77988
rect 144224 77864 144544 77932
rect 144224 77808 144294 77864
rect 144350 77808 144418 77864
rect 144474 77808 144544 77864
rect 144224 77678 144544 77808
rect 154224 78608 154544 81752
rect 159224 80008 159544 81752
rect 159224 79952 159294 80008
rect 159350 79952 159418 80008
rect 159474 79952 159544 80008
rect 159224 79884 159544 79952
rect 159224 79828 159294 79884
rect 159350 79828 159418 79884
rect 159474 79828 159544 79884
rect 159224 79760 159544 79828
rect 159224 79704 159294 79760
rect 159350 79704 159418 79760
rect 159474 79704 159544 79760
rect 159224 79636 159544 79704
rect 159224 79580 159294 79636
rect 159350 79580 159418 79636
rect 159474 79580 159544 79636
rect 159224 79512 159544 79580
rect 159224 79456 159294 79512
rect 159350 79456 159418 79512
rect 159474 79456 159544 79512
rect 159224 79388 159544 79456
rect 159224 79332 159294 79388
rect 159350 79332 159418 79388
rect 159474 79332 159544 79388
rect 159224 79264 159544 79332
rect 159224 79208 159294 79264
rect 159350 79208 159418 79264
rect 159474 79208 159544 79264
rect 159224 79078 159544 79208
rect 154224 78552 154294 78608
rect 154350 78552 154418 78608
rect 154474 78552 154544 78608
rect 154224 78484 154544 78552
rect 154224 78428 154294 78484
rect 154350 78428 154418 78484
rect 154474 78428 154544 78484
rect 154224 78360 154544 78428
rect 154224 78304 154294 78360
rect 154350 78304 154418 78360
rect 154474 78304 154544 78360
rect 154224 78236 154544 78304
rect 154224 78180 154294 78236
rect 154350 78180 154418 78236
rect 154474 78180 154544 78236
rect 154224 78112 154544 78180
rect 154224 78056 154294 78112
rect 154350 78056 154418 78112
rect 154474 78056 154544 78112
rect 154224 77988 154544 78056
rect 154224 77932 154294 77988
rect 154350 77932 154418 77988
rect 154474 77932 154544 77988
rect 154224 77864 154544 77932
rect 154224 77808 154294 77864
rect 154350 77808 154418 77864
rect 154474 77808 154544 77864
rect 154224 77678 154544 77808
rect 164224 78608 164544 81752
rect 169224 80008 169544 81752
rect 169224 79952 169294 80008
rect 169350 79952 169418 80008
rect 169474 79952 169544 80008
rect 169224 79884 169544 79952
rect 169224 79828 169294 79884
rect 169350 79828 169418 79884
rect 169474 79828 169544 79884
rect 169224 79760 169544 79828
rect 169224 79704 169294 79760
rect 169350 79704 169418 79760
rect 169474 79704 169544 79760
rect 169224 79636 169544 79704
rect 169224 79580 169294 79636
rect 169350 79580 169418 79636
rect 169474 79580 169544 79636
rect 169224 79512 169544 79580
rect 169224 79456 169294 79512
rect 169350 79456 169418 79512
rect 169474 79456 169544 79512
rect 169224 79388 169544 79456
rect 169224 79332 169294 79388
rect 169350 79332 169418 79388
rect 169474 79332 169544 79388
rect 169224 79264 169544 79332
rect 169224 79208 169294 79264
rect 169350 79208 169418 79264
rect 169474 79208 169544 79264
rect 169224 79078 169544 79208
rect 164224 78552 164294 78608
rect 164350 78552 164418 78608
rect 164474 78552 164544 78608
rect 164224 78484 164544 78552
rect 164224 78428 164294 78484
rect 164350 78428 164418 78484
rect 164474 78428 164544 78484
rect 164224 78360 164544 78428
rect 164224 78304 164294 78360
rect 164350 78304 164418 78360
rect 164474 78304 164544 78360
rect 164224 78236 164544 78304
rect 164224 78180 164294 78236
rect 164350 78180 164418 78236
rect 164474 78180 164544 78236
rect 164224 78112 164544 78180
rect 164224 78056 164294 78112
rect 164350 78056 164418 78112
rect 164474 78056 164544 78112
rect 164224 77988 164544 78056
rect 164224 77932 164294 77988
rect 164350 77932 164418 77988
rect 164474 77932 164544 77988
rect 164224 77864 164544 77932
rect 164224 77808 164294 77864
rect 164350 77808 164418 77864
rect 164474 77808 164544 77864
rect 164224 77678 164544 77808
rect 174224 78608 174544 81752
rect 179224 80008 179544 81752
rect 179224 79952 179294 80008
rect 179350 79952 179418 80008
rect 179474 79952 179544 80008
rect 179224 79884 179544 79952
rect 179224 79828 179294 79884
rect 179350 79828 179418 79884
rect 179474 79828 179544 79884
rect 179224 79760 179544 79828
rect 179224 79704 179294 79760
rect 179350 79704 179418 79760
rect 179474 79704 179544 79760
rect 179224 79636 179544 79704
rect 179224 79580 179294 79636
rect 179350 79580 179418 79636
rect 179474 79580 179544 79636
rect 179224 79512 179544 79580
rect 179224 79456 179294 79512
rect 179350 79456 179418 79512
rect 179474 79456 179544 79512
rect 179224 79388 179544 79456
rect 179224 79332 179294 79388
rect 179350 79332 179418 79388
rect 179474 79332 179544 79388
rect 179224 79264 179544 79332
rect 179224 79208 179294 79264
rect 179350 79208 179418 79264
rect 179474 79208 179544 79264
rect 179224 79078 179544 79208
rect 174224 78552 174294 78608
rect 174350 78552 174418 78608
rect 174474 78552 174544 78608
rect 174224 78484 174544 78552
rect 174224 78428 174294 78484
rect 174350 78428 174418 78484
rect 174474 78428 174544 78484
rect 174224 78360 174544 78428
rect 174224 78304 174294 78360
rect 174350 78304 174418 78360
rect 174474 78304 174544 78360
rect 174224 78236 174544 78304
rect 174224 78180 174294 78236
rect 174350 78180 174418 78236
rect 174474 78180 174544 78236
rect 174224 78112 174544 78180
rect 174224 78056 174294 78112
rect 174350 78056 174418 78112
rect 174474 78056 174544 78112
rect 174224 77988 174544 78056
rect 174224 77932 174294 77988
rect 174350 77932 174418 77988
rect 174474 77932 174544 77988
rect 174224 77864 174544 77932
rect 174224 77808 174294 77864
rect 174350 77808 174418 77864
rect 174474 77808 174544 77864
rect 174224 77678 174544 77808
rect 184224 78608 184544 81752
rect 189224 80008 189544 81752
rect 189224 79952 189294 80008
rect 189350 79952 189418 80008
rect 189474 79952 189544 80008
rect 189224 79884 189544 79952
rect 189224 79828 189294 79884
rect 189350 79828 189418 79884
rect 189474 79828 189544 79884
rect 189224 79760 189544 79828
rect 189224 79704 189294 79760
rect 189350 79704 189418 79760
rect 189474 79704 189544 79760
rect 189224 79636 189544 79704
rect 189224 79580 189294 79636
rect 189350 79580 189418 79636
rect 189474 79580 189544 79636
rect 189224 79512 189544 79580
rect 189224 79456 189294 79512
rect 189350 79456 189418 79512
rect 189474 79456 189544 79512
rect 189224 79388 189544 79456
rect 189224 79332 189294 79388
rect 189350 79332 189418 79388
rect 189474 79332 189544 79388
rect 189224 79264 189544 79332
rect 189224 79208 189294 79264
rect 189350 79208 189418 79264
rect 189474 79208 189544 79264
rect 189224 79078 189544 79208
rect 184224 78552 184294 78608
rect 184350 78552 184418 78608
rect 184474 78552 184544 78608
rect 184224 78484 184544 78552
rect 184224 78428 184294 78484
rect 184350 78428 184418 78484
rect 184474 78428 184544 78484
rect 184224 78360 184544 78428
rect 184224 78304 184294 78360
rect 184350 78304 184418 78360
rect 184474 78304 184544 78360
rect 184224 78236 184544 78304
rect 184224 78180 184294 78236
rect 184350 78180 184418 78236
rect 184474 78180 184544 78236
rect 184224 78112 184544 78180
rect 184224 78056 184294 78112
rect 184350 78056 184418 78112
rect 184474 78056 184544 78112
rect 184224 77988 184544 78056
rect 184224 77932 184294 77988
rect 184350 77932 184418 77988
rect 184474 77932 184544 77988
rect 184224 77864 184544 77932
rect 184224 77808 184294 77864
rect 184350 77808 184418 77864
rect 184474 77808 184544 77864
rect 184224 77678 184544 77808
rect 194224 78608 194544 81752
rect 199224 80008 199544 81752
rect 199224 79952 199294 80008
rect 199350 79952 199418 80008
rect 199474 79952 199544 80008
rect 199224 79884 199544 79952
rect 199224 79828 199294 79884
rect 199350 79828 199418 79884
rect 199474 79828 199544 79884
rect 199224 79760 199544 79828
rect 199224 79704 199294 79760
rect 199350 79704 199418 79760
rect 199474 79704 199544 79760
rect 199224 79636 199544 79704
rect 199224 79580 199294 79636
rect 199350 79580 199418 79636
rect 199474 79580 199544 79636
rect 199224 79512 199544 79580
rect 199224 79456 199294 79512
rect 199350 79456 199418 79512
rect 199474 79456 199544 79512
rect 199224 79388 199544 79456
rect 199224 79332 199294 79388
rect 199350 79332 199418 79388
rect 199474 79332 199544 79388
rect 199224 79264 199544 79332
rect 199224 79208 199294 79264
rect 199350 79208 199418 79264
rect 199474 79208 199544 79264
rect 199224 79078 199544 79208
rect 194224 78552 194294 78608
rect 194350 78552 194418 78608
rect 194474 78552 194544 78608
rect 194224 78484 194544 78552
rect 194224 78428 194294 78484
rect 194350 78428 194418 78484
rect 194474 78428 194544 78484
rect 194224 78360 194544 78428
rect 194224 78304 194294 78360
rect 194350 78304 194418 78360
rect 194474 78304 194544 78360
rect 194224 78236 194544 78304
rect 194224 78180 194294 78236
rect 194350 78180 194418 78236
rect 194474 78180 194544 78236
rect 194224 78112 194544 78180
rect 194224 78056 194294 78112
rect 194350 78056 194418 78112
rect 194474 78056 194544 78112
rect 194224 77988 194544 78056
rect 194224 77932 194294 77988
rect 194350 77932 194418 77988
rect 194474 77932 194544 77988
rect 194224 77864 194544 77932
rect 194224 77808 194294 77864
rect 194350 77808 194418 77864
rect 194474 77808 194544 77864
rect 194224 77678 194544 77808
rect 204224 78608 204544 81752
rect 209224 80008 209544 81752
rect 209224 79952 209294 80008
rect 209350 79952 209418 80008
rect 209474 79952 209544 80008
rect 209224 79884 209544 79952
rect 209224 79828 209294 79884
rect 209350 79828 209418 79884
rect 209474 79828 209544 79884
rect 209224 79760 209544 79828
rect 209224 79704 209294 79760
rect 209350 79704 209418 79760
rect 209474 79704 209544 79760
rect 209224 79636 209544 79704
rect 209224 79580 209294 79636
rect 209350 79580 209418 79636
rect 209474 79580 209544 79636
rect 209224 79512 209544 79580
rect 209224 79456 209294 79512
rect 209350 79456 209418 79512
rect 209474 79456 209544 79512
rect 209224 79388 209544 79456
rect 209224 79332 209294 79388
rect 209350 79332 209418 79388
rect 209474 79332 209544 79388
rect 209224 79264 209544 79332
rect 209224 79208 209294 79264
rect 209350 79208 209418 79264
rect 209474 79208 209544 79264
rect 209224 79078 209544 79208
rect 204224 78552 204294 78608
rect 204350 78552 204418 78608
rect 204474 78552 204544 78608
rect 204224 78484 204544 78552
rect 204224 78428 204294 78484
rect 204350 78428 204418 78484
rect 204474 78428 204544 78484
rect 204224 78360 204544 78428
rect 204224 78304 204294 78360
rect 204350 78304 204418 78360
rect 204474 78304 204544 78360
rect 204224 78236 204544 78304
rect 204224 78180 204294 78236
rect 204350 78180 204418 78236
rect 204474 78180 204544 78236
rect 204224 78112 204544 78180
rect 204224 78056 204294 78112
rect 204350 78056 204418 78112
rect 204474 78056 204544 78112
rect 204224 77988 204544 78056
rect 204224 77932 204294 77988
rect 204350 77932 204418 77988
rect 204474 77932 204544 77988
rect 204224 77864 204544 77932
rect 204224 77808 204294 77864
rect 204350 77808 204418 77864
rect 204474 77808 204544 77864
rect 204224 77678 204544 77808
rect 214224 78608 214544 81752
rect 219224 80008 219544 81752
rect 219224 79952 219294 80008
rect 219350 79952 219418 80008
rect 219474 79952 219544 80008
rect 219224 79884 219544 79952
rect 219224 79828 219294 79884
rect 219350 79828 219418 79884
rect 219474 79828 219544 79884
rect 219224 79760 219544 79828
rect 219224 79704 219294 79760
rect 219350 79704 219418 79760
rect 219474 79704 219544 79760
rect 219224 79636 219544 79704
rect 219224 79580 219294 79636
rect 219350 79580 219418 79636
rect 219474 79580 219544 79636
rect 219224 79512 219544 79580
rect 219224 79456 219294 79512
rect 219350 79456 219418 79512
rect 219474 79456 219544 79512
rect 219224 79388 219544 79456
rect 219224 79332 219294 79388
rect 219350 79332 219418 79388
rect 219474 79332 219544 79388
rect 219224 79264 219544 79332
rect 219224 79208 219294 79264
rect 219350 79208 219418 79264
rect 219474 79208 219544 79264
rect 219224 79078 219544 79208
rect 214224 78552 214294 78608
rect 214350 78552 214418 78608
rect 214474 78552 214544 78608
rect 214224 78484 214544 78552
rect 214224 78428 214294 78484
rect 214350 78428 214418 78484
rect 214474 78428 214544 78484
rect 214224 78360 214544 78428
rect 214224 78304 214294 78360
rect 214350 78304 214418 78360
rect 214474 78304 214544 78360
rect 214224 78236 214544 78304
rect 214224 78180 214294 78236
rect 214350 78180 214418 78236
rect 214474 78180 214544 78236
rect 214224 78112 214544 78180
rect 214224 78056 214294 78112
rect 214350 78056 214418 78112
rect 214474 78056 214544 78112
rect 214224 77988 214544 78056
rect 214224 77932 214294 77988
rect 214350 77932 214418 77988
rect 214474 77932 214544 77988
rect 214224 77864 214544 77932
rect 214224 77808 214294 77864
rect 214350 77808 214418 77864
rect 214474 77808 214544 77864
rect 214224 77678 214544 77808
rect 224224 78608 224544 81752
rect 229224 80008 229544 81752
rect 229224 79952 229294 80008
rect 229350 79952 229418 80008
rect 229474 79952 229544 80008
rect 229224 79884 229544 79952
rect 229224 79828 229294 79884
rect 229350 79828 229418 79884
rect 229474 79828 229544 79884
rect 229224 79760 229544 79828
rect 229224 79704 229294 79760
rect 229350 79704 229418 79760
rect 229474 79704 229544 79760
rect 229224 79636 229544 79704
rect 229224 79580 229294 79636
rect 229350 79580 229418 79636
rect 229474 79580 229544 79636
rect 229224 79512 229544 79580
rect 229224 79456 229294 79512
rect 229350 79456 229418 79512
rect 229474 79456 229544 79512
rect 229224 79388 229544 79456
rect 229224 79332 229294 79388
rect 229350 79332 229418 79388
rect 229474 79332 229544 79388
rect 229224 79264 229544 79332
rect 229224 79208 229294 79264
rect 229350 79208 229418 79264
rect 229474 79208 229544 79264
rect 229224 79078 229544 79208
rect 224224 78552 224294 78608
rect 224350 78552 224418 78608
rect 224474 78552 224544 78608
rect 224224 78484 224544 78552
rect 224224 78428 224294 78484
rect 224350 78428 224418 78484
rect 224474 78428 224544 78484
rect 224224 78360 224544 78428
rect 224224 78304 224294 78360
rect 224350 78304 224418 78360
rect 224474 78304 224544 78360
rect 224224 78236 224544 78304
rect 224224 78180 224294 78236
rect 224350 78180 224418 78236
rect 224474 78180 224544 78236
rect 224224 78112 224544 78180
rect 224224 78056 224294 78112
rect 224350 78056 224418 78112
rect 224474 78056 224544 78112
rect 224224 77988 224544 78056
rect 224224 77932 224294 77988
rect 224350 77932 224418 77988
rect 224474 77932 224544 77988
rect 224224 77864 224544 77932
rect 224224 77808 224294 77864
rect 224350 77808 224418 77864
rect 224474 77808 224544 77864
rect 224224 77678 224544 77808
rect 234224 78608 234544 81752
rect 239224 80008 239544 81752
rect 239224 79952 239294 80008
rect 239350 79952 239418 80008
rect 239474 79952 239544 80008
rect 239224 79884 239544 79952
rect 239224 79828 239294 79884
rect 239350 79828 239418 79884
rect 239474 79828 239544 79884
rect 239224 79760 239544 79828
rect 239224 79704 239294 79760
rect 239350 79704 239418 79760
rect 239474 79704 239544 79760
rect 239224 79636 239544 79704
rect 239224 79580 239294 79636
rect 239350 79580 239418 79636
rect 239474 79580 239544 79636
rect 239224 79512 239544 79580
rect 239224 79456 239294 79512
rect 239350 79456 239418 79512
rect 239474 79456 239544 79512
rect 239224 79388 239544 79456
rect 239224 79332 239294 79388
rect 239350 79332 239418 79388
rect 239474 79332 239544 79388
rect 239224 79264 239544 79332
rect 239224 79208 239294 79264
rect 239350 79208 239418 79264
rect 239474 79208 239544 79264
rect 239224 79078 239544 79208
rect 234224 78552 234294 78608
rect 234350 78552 234418 78608
rect 234474 78552 234544 78608
rect 234224 78484 234544 78552
rect 234224 78428 234294 78484
rect 234350 78428 234418 78484
rect 234474 78428 234544 78484
rect 234224 78360 234544 78428
rect 234224 78304 234294 78360
rect 234350 78304 234418 78360
rect 234474 78304 234544 78360
rect 234224 78236 234544 78304
rect 234224 78180 234294 78236
rect 234350 78180 234418 78236
rect 234474 78180 234544 78236
rect 234224 78112 234544 78180
rect 234224 78056 234294 78112
rect 234350 78056 234418 78112
rect 234474 78056 234544 78112
rect 234224 77988 234544 78056
rect 234224 77932 234294 77988
rect 234350 77932 234418 77988
rect 234474 77932 234544 77988
rect 234224 77864 234544 77932
rect 234224 77808 234294 77864
rect 234350 77808 234418 77864
rect 234474 77808 234544 77864
rect 234224 77678 234544 77808
rect 244224 78608 244544 81752
rect 249224 80008 249544 81752
rect 249224 79952 249294 80008
rect 249350 79952 249418 80008
rect 249474 79952 249544 80008
rect 249224 79884 249544 79952
rect 249224 79828 249294 79884
rect 249350 79828 249418 79884
rect 249474 79828 249544 79884
rect 249224 79760 249544 79828
rect 249224 79704 249294 79760
rect 249350 79704 249418 79760
rect 249474 79704 249544 79760
rect 249224 79636 249544 79704
rect 249224 79580 249294 79636
rect 249350 79580 249418 79636
rect 249474 79580 249544 79636
rect 249224 79512 249544 79580
rect 249224 79456 249294 79512
rect 249350 79456 249418 79512
rect 249474 79456 249544 79512
rect 249224 79388 249544 79456
rect 249224 79332 249294 79388
rect 249350 79332 249418 79388
rect 249474 79332 249544 79388
rect 249224 79264 249544 79332
rect 249224 79208 249294 79264
rect 249350 79208 249418 79264
rect 249474 79208 249544 79264
rect 249224 79078 249544 79208
rect 244224 78552 244294 78608
rect 244350 78552 244418 78608
rect 244474 78552 244544 78608
rect 244224 78484 244544 78552
rect 244224 78428 244294 78484
rect 244350 78428 244418 78484
rect 244474 78428 244544 78484
rect 244224 78360 244544 78428
rect 244224 78304 244294 78360
rect 244350 78304 244418 78360
rect 244474 78304 244544 78360
rect 244224 78236 244544 78304
rect 244224 78180 244294 78236
rect 244350 78180 244418 78236
rect 244474 78180 244544 78236
rect 244224 78112 244544 78180
rect 244224 78056 244294 78112
rect 244350 78056 244418 78112
rect 244474 78056 244544 78112
rect 244224 77988 244544 78056
rect 244224 77932 244294 77988
rect 244350 77932 244418 77988
rect 244474 77932 244544 77988
rect 244224 77864 244544 77932
rect 244224 77808 244294 77864
rect 244350 77808 244418 77864
rect 244474 77808 244544 77864
rect 244224 77678 244544 77808
rect 254224 78608 254544 81752
rect 259224 80008 259544 81752
rect 259224 79952 259294 80008
rect 259350 79952 259418 80008
rect 259474 79952 259544 80008
rect 259224 79884 259544 79952
rect 259224 79828 259294 79884
rect 259350 79828 259418 79884
rect 259474 79828 259544 79884
rect 259224 79760 259544 79828
rect 259224 79704 259294 79760
rect 259350 79704 259418 79760
rect 259474 79704 259544 79760
rect 259224 79636 259544 79704
rect 259224 79580 259294 79636
rect 259350 79580 259418 79636
rect 259474 79580 259544 79636
rect 259224 79512 259544 79580
rect 259224 79456 259294 79512
rect 259350 79456 259418 79512
rect 259474 79456 259544 79512
rect 259224 79388 259544 79456
rect 259224 79332 259294 79388
rect 259350 79332 259418 79388
rect 259474 79332 259544 79388
rect 259224 79264 259544 79332
rect 259224 79208 259294 79264
rect 259350 79208 259418 79264
rect 259474 79208 259544 79264
rect 259224 79078 259544 79208
rect 254224 78552 254294 78608
rect 254350 78552 254418 78608
rect 254474 78552 254544 78608
rect 254224 78484 254544 78552
rect 254224 78428 254294 78484
rect 254350 78428 254418 78484
rect 254474 78428 254544 78484
rect 254224 78360 254544 78428
rect 254224 78304 254294 78360
rect 254350 78304 254418 78360
rect 254474 78304 254544 78360
rect 254224 78236 254544 78304
rect 254224 78180 254294 78236
rect 254350 78180 254418 78236
rect 254474 78180 254544 78236
rect 254224 78112 254544 78180
rect 254224 78056 254294 78112
rect 254350 78056 254418 78112
rect 254474 78056 254544 78112
rect 254224 77988 254544 78056
rect 254224 77932 254294 77988
rect 254350 77932 254418 77988
rect 254474 77932 254544 77988
rect 254224 77864 254544 77932
rect 254224 77808 254294 77864
rect 254350 77808 254418 77864
rect 254474 77808 254544 77864
rect 254224 77678 254544 77808
rect 264224 78608 264544 81752
rect 269224 80008 269544 81752
rect 269224 79952 269294 80008
rect 269350 79952 269418 80008
rect 269474 79952 269544 80008
rect 269224 79884 269544 79952
rect 269224 79828 269294 79884
rect 269350 79828 269418 79884
rect 269474 79828 269544 79884
rect 269224 79760 269544 79828
rect 269224 79704 269294 79760
rect 269350 79704 269418 79760
rect 269474 79704 269544 79760
rect 269224 79636 269544 79704
rect 269224 79580 269294 79636
rect 269350 79580 269418 79636
rect 269474 79580 269544 79636
rect 269224 79512 269544 79580
rect 269224 79456 269294 79512
rect 269350 79456 269418 79512
rect 269474 79456 269544 79512
rect 269224 79388 269544 79456
rect 269224 79332 269294 79388
rect 269350 79332 269418 79388
rect 269474 79332 269544 79388
rect 269224 79264 269544 79332
rect 269224 79208 269294 79264
rect 269350 79208 269418 79264
rect 269474 79208 269544 79264
rect 269224 79078 269544 79208
rect 272272 80008 274172 80078
rect 272272 79952 272330 80008
rect 272386 79952 272454 80008
rect 272510 79952 272578 80008
rect 272634 79952 272702 80008
rect 272758 79952 272826 80008
rect 272882 79952 272950 80008
rect 273006 79952 273074 80008
rect 273130 79952 273198 80008
rect 273254 79952 273322 80008
rect 273378 79952 273446 80008
rect 273502 79952 273570 80008
rect 273626 79952 273694 80008
rect 273750 79952 273818 80008
rect 273874 79952 273942 80008
rect 273998 79952 274066 80008
rect 274122 79952 274172 80008
rect 272272 79884 274172 79952
rect 272272 79828 272330 79884
rect 272386 79828 272454 79884
rect 272510 79828 272578 79884
rect 272634 79828 272702 79884
rect 272758 79828 272826 79884
rect 272882 79828 272950 79884
rect 273006 79828 273074 79884
rect 273130 79828 273198 79884
rect 273254 79828 273322 79884
rect 273378 79828 273446 79884
rect 273502 79828 273570 79884
rect 273626 79828 273694 79884
rect 273750 79828 273818 79884
rect 273874 79828 273942 79884
rect 273998 79828 274066 79884
rect 274122 79828 274172 79884
rect 272272 79760 274172 79828
rect 272272 79704 272330 79760
rect 272386 79704 272454 79760
rect 272510 79704 272578 79760
rect 272634 79704 272702 79760
rect 272758 79704 272826 79760
rect 272882 79704 272950 79760
rect 273006 79704 273074 79760
rect 273130 79704 273198 79760
rect 273254 79704 273322 79760
rect 273378 79704 273446 79760
rect 273502 79704 273570 79760
rect 273626 79704 273694 79760
rect 273750 79704 273818 79760
rect 273874 79704 273942 79760
rect 273998 79704 274066 79760
rect 274122 79704 274172 79760
rect 272272 79636 274172 79704
rect 272272 79580 272330 79636
rect 272386 79580 272454 79636
rect 272510 79580 272578 79636
rect 272634 79580 272702 79636
rect 272758 79580 272826 79636
rect 272882 79580 272950 79636
rect 273006 79580 273074 79636
rect 273130 79580 273198 79636
rect 273254 79580 273322 79636
rect 273378 79580 273446 79636
rect 273502 79580 273570 79636
rect 273626 79580 273694 79636
rect 273750 79580 273818 79636
rect 273874 79580 273942 79636
rect 273998 79580 274066 79636
rect 274122 79580 274172 79636
rect 272272 79512 274172 79580
rect 272272 79456 272330 79512
rect 272386 79456 272454 79512
rect 272510 79456 272578 79512
rect 272634 79456 272702 79512
rect 272758 79456 272826 79512
rect 272882 79456 272950 79512
rect 273006 79456 273074 79512
rect 273130 79456 273198 79512
rect 273254 79456 273322 79512
rect 273378 79456 273446 79512
rect 273502 79456 273570 79512
rect 273626 79456 273694 79512
rect 273750 79456 273818 79512
rect 273874 79456 273942 79512
rect 273998 79456 274066 79512
rect 274122 79456 274172 79512
rect 272272 79388 274172 79456
rect 272272 79332 272330 79388
rect 272386 79332 272454 79388
rect 272510 79332 272578 79388
rect 272634 79332 272702 79388
rect 272758 79332 272826 79388
rect 272882 79332 272950 79388
rect 273006 79332 273074 79388
rect 273130 79332 273198 79388
rect 273254 79332 273322 79388
rect 273378 79332 273446 79388
rect 273502 79332 273570 79388
rect 273626 79332 273694 79388
rect 273750 79332 273818 79388
rect 273874 79332 273942 79388
rect 273998 79332 274066 79388
rect 274122 79332 274172 79388
rect 272272 79264 274172 79332
rect 272272 79208 272330 79264
rect 272386 79208 272454 79264
rect 272510 79208 272578 79264
rect 272634 79208 272702 79264
rect 272758 79208 272826 79264
rect 272882 79208 272950 79264
rect 273006 79208 273074 79264
rect 273130 79208 273198 79264
rect 273254 79208 273322 79264
rect 273378 79208 273446 79264
rect 273502 79208 273570 79264
rect 273626 79208 273694 79264
rect 273750 79208 273818 79264
rect 273874 79208 273942 79264
rect 273998 79208 274066 79264
rect 274122 79208 274172 79264
rect 264224 78552 264294 78608
rect 264350 78552 264418 78608
rect 264474 78552 264544 78608
rect 264224 78484 264544 78552
rect 264224 78428 264294 78484
rect 264350 78428 264418 78484
rect 264474 78428 264544 78484
rect 264224 78360 264544 78428
rect 264224 78304 264294 78360
rect 264350 78304 264418 78360
rect 264474 78304 264544 78360
rect 264224 78236 264544 78304
rect 264224 78180 264294 78236
rect 264350 78180 264418 78236
rect 264474 78180 264544 78236
rect 264224 78112 264544 78180
rect 264224 78056 264294 78112
rect 264350 78056 264418 78112
rect 264474 78056 264544 78112
rect 264224 77988 264544 78056
rect 264224 77932 264294 77988
rect 264350 77932 264418 77988
rect 264474 77932 264544 77988
rect 264224 77864 264544 77932
rect 264224 77808 264294 77864
rect 264350 77808 264418 77864
rect 264474 77808 264544 77864
rect 264224 77678 264544 77808
rect 119828 70074 119866 70130
rect 119922 70074 119990 70130
rect 120046 70074 120114 70130
rect 120170 70074 120238 70130
rect 120294 70074 120362 70130
rect 120418 70074 120486 70130
rect 120542 70074 120610 70130
rect 120666 70074 120734 70130
rect 120790 70074 120858 70130
rect 120914 70074 120982 70130
rect 121038 70074 121106 70130
rect 121162 70074 121230 70130
rect 121286 70074 121354 70130
rect 121410 70074 121478 70130
rect 121534 70074 121602 70130
rect 121658 70074 121728 70130
rect 119828 70000 121728 70074
rect 272272 70130 274172 79208
rect 272272 70074 272342 70130
rect 272398 70074 272466 70130
rect 272522 70074 272590 70130
rect 272646 70074 272714 70130
rect 272770 70074 272838 70130
rect 272894 70074 272962 70130
rect 273018 70074 273086 70130
rect 273142 70074 273210 70130
rect 273266 70074 273334 70130
rect 273390 70074 273458 70130
rect 273514 70074 273582 70130
rect 273638 70074 273706 70130
rect 273762 70074 273830 70130
rect 273886 70074 273954 70130
rect 274010 70074 274078 70130
rect 274134 70074 274172 70130
rect 272272 70000 274172 70074
rect 274752 80008 276802 80078
rect 274752 79952 274810 80008
rect 274866 79952 274934 80008
rect 274990 79952 275058 80008
rect 275114 79952 275182 80008
rect 275238 79952 275306 80008
rect 275362 79952 275430 80008
rect 275486 79952 275554 80008
rect 275610 79952 275678 80008
rect 275734 79952 275802 80008
rect 275858 79952 275926 80008
rect 275982 79952 276050 80008
rect 276106 79952 276174 80008
rect 276230 79952 276298 80008
rect 276354 79952 276422 80008
rect 276478 79952 276546 80008
rect 276602 79952 276670 80008
rect 276726 79952 276802 80008
rect 274752 79884 276802 79952
rect 274752 79828 274810 79884
rect 274866 79828 274934 79884
rect 274990 79828 275058 79884
rect 275114 79828 275182 79884
rect 275238 79828 275306 79884
rect 275362 79828 275430 79884
rect 275486 79828 275554 79884
rect 275610 79828 275678 79884
rect 275734 79828 275802 79884
rect 275858 79828 275926 79884
rect 275982 79828 276050 79884
rect 276106 79828 276174 79884
rect 276230 79828 276298 79884
rect 276354 79828 276422 79884
rect 276478 79828 276546 79884
rect 276602 79828 276670 79884
rect 276726 79828 276802 79884
rect 274752 79760 276802 79828
rect 274752 79704 274810 79760
rect 274866 79704 274934 79760
rect 274990 79704 275058 79760
rect 275114 79704 275182 79760
rect 275238 79704 275306 79760
rect 275362 79704 275430 79760
rect 275486 79704 275554 79760
rect 275610 79704 275678 79760
rect 275734 79704 275802 79760
rect 275858 79704 275926 79760
rect 275982 79704 276050 79760
rect 276106 79704 276174 79760
rect 276230 79704 276298 79760
rect 276354 79704 276422 79760
rect 276478 79704 276546 79760
rect 276602 79704 276670 79760
rect 276726 79704 276802 79760
rect 274752 79636 276802 79704
rect 274752 79580 274810 79636
rect 274866 79580 274934 79636
rect 274990 79580 275058 79636
rect 275114 79580 275182 79636
rect 275238 79580 275306 79636
rect 275362 79580 275430 79636
rect 275486 79580 275554 79636
rect 275610 79580 275678 79636
rect 275734 79580 275802 79636
rect 275858 79580 275926 79636
rect 275982 79580 276050 79636
rect 276106 79580 276174 79636
rect 276230 79580 276298 79636
rect 276354 79580 276422 79636
rect 276478 79580 276546 79636
rect 276602 79580 276670 79636
rect 276726 79580 276802 79636
rect 274752 79512 276802 79580
rect 274752 79456 274810 79512
rect 274866 79456 274934 79512
rect 274990 79456 275058 79512
rect 275114 79456 275182 79512
rect 275238 79456 275306 79512
rect 275362 79456 275430 79512
rect 275486 79456 275554 79512
rect 275610 79456 275678 79512
rect 275734 79456 275802 79512
rect 275858 79456 275926 79512
rect 275982 79456 276050 79512
rect 276106 79456 276174 79512
rect 276230 79456 276298 79512
rect 276354 79456 276422 79512
rect 276478 79456 276546 79512
rect 276602 79456 276670 79512
rect 276726 79456 276802 79512
rect 274752 79388 276802 79456
rect 274752 79332 274810 79388
rect 274866 79332 274934 79388
rect 274990 79332 275058 79388
rect 275114 79332 275182 79388
rect 275238 79332 275306 79388
rect 275362 79332 275430 79388
rect 275486 79332 275554 79388
rect 275610 79332 275678 79388
rect 275734 79332 275802 79388
rect 275858 79332 275926 79388
rect 275982 79332 276050 79388
rect 276106 79332 276174 79388
rect 276230 79332 276298 79388
rect 276354 79332 276422 79388
rect 276478 79332 276546 79388
rect 276602 79332 276670 79388
rect 276726 79332 276802 79388
rect 274752 79264 276802 79332
rect 274752 79208 274810 79264
rect 274866 79208 274934 79264
rect 274990 79208 275058 79264
rect 275114 79208 275182 79264
rect 275238 79208 275306 79264
rect 275362 79208 275430 79264
rect 275486 79208 275554 79264
rect 275610 79208 275678 79264
rect 275734 79208 275802 79264
rect 275858 79208 275926 79264
rect 275982 79208 276050 79264
rect 276106 79208 276174 79264
rect 276230 79208 276298 79264
rect 276354 79208 276422 79264
rect 276478 79208 276546 79264
rect 276602 79208 276670 79264
rect 276726 79208 276802 79264
rect 274752 70130 276802 79208
rect 274752 70074 274822 70130
rect 274878 70074 274946 70130
rect 275002 70074 275070 70130
rect 275126 70074 275194 70130
rect 275250 70074 275318 70130
rect 275374 70074 275442 70130
rect 275498 70074 275566 70130
rect 275622 70074 275690 70130
rect 275746 70074 275814 70130
rect 275870 70074 275938 70130
rect 275994 70074 276062 70130
rect 276118 70074 276186 70130
rect 276242 70074 276310 70130
rect 276366 70074 276434 70130
rect 276490 70074 276558 70130
rect 276614 70074 276682 70130
rect 276738 70074 276802 70130
rect 274752 70000 276802 70074
rect 277122 80008 279172 80078
rect 277122 79952 277180 80008
rect 277236 79952 277304 80008
rect 277360 79952 277428 80008
rect 277484 79952 277552 80008
rect 277608 79952 277676 80008
rect 277732 79952 277800 80008
rect 277856 79952 277924 80008
rect 277980 79952 278048 80008
rect 278104 79952 278172 80008
rect 278228 79952 278296 80008
rect 278352 79952 278420 80008
rect 278476 79952 278544 80008
rect 278600 79952 278668 80008
rect 278724 79952 278792 80008
rect 278848 79952 278916 80008
rect 278972 79952 279040 80008
rect 279096 79952 279172 80008
rect 277122 79884 279172 79952
rect 277122 79828 277180 79884
rect 277236 79828 277304 79884
rect 277360 79828 277428 79884
rect 277484 79828 277552 79884
rect 277608 79828 277676 79884
rect 277732 79828 277800 79884
rect 277856 79828 277924 79884
rect 277980 79828 278048 79884
rect 278104 79828 278172 79884
rect 278228 79828 278296 79884
rect 278352 79828 278420 79884
rect 278476 79828 278544 79884
rect 278600 79828 278668 79884
rect 278724 79828 278792 79884
rect 278848 79828 278916 79884
rect 278972 79828 279040 79884
rect 279096 79828 279172 79884
rect 277122 79760 279172 79828
rect 277122 79704 277180 79760
rect 277236 79704 277304 79760
rect 277360 79704 277428 79760
rect 277484 79704 277552 79760
rect 277608 79704 277676 79760
rect 277732 79704 277800 79760
rect 277856 79704 277924 79760
rect 277980 79704 278048 79760
rect 278104 79704 278172 79760
rect 278228 79704 278296 79760
rect 278352 79704 278420 79760
rect 278476 79704 278544 79760
rect 278600 79704 278668 79760
rect 278724 79704 278792 79760
rect 278848 79704 278916 79760
rect 278972 79704 279040 79760
rect 279096 79704 279172 79760
rect 277122 79636 279172 79704
rect 277122 79580 277180 79636
rect 277236 79580 277304 79636
rect 277360 79580 277428 79636
rect 277484 79580 277552 79636
rect 277608 79580 277676 79636
rect 277732 79580 277800 79636
rect 277856 79580 277924 79636
rect 277980 79580 278048 79636
rect 278104 79580 278172 79636
rect 278228 79580 278296 79636
rect 278352 79580 278420 79636
rect 278476 79580 278544 79636
rect 278600 79580 278668 79636
rect 278724 79580 278792 79636
rect 278848 79580 278916 79636
rect 278972 79580 279040 79636
rect 279096 79580 279172 79636
rect 277122 79512 279172 79580
rect 277122 79456 277180 79512
rect 277236 79456 277304 79512
rect 277360 79456 277428 79512
rect 277484 79456 277552 79512
rect 277608 79456 277676 79512
rect 277732 79456 277800 79512
rect 277856 79456 277924 79512
rect 277980 79456 278048 79512
rect 278104 79456 278172 79512
rect 278228 79456 278296 79512
rect 278352 79456 278420 79512
rect 278476 79456 278544 79512
rect 278600 79456 278668 79512
rect 278724 79456 278792 79512
rect 278848 79456 278916 79512
rect 278972 79456 279040 79512
rect 279096 79456 279172 79512
rect 277122 79388 279172 79456
rect 277122 79332 277180 79388
rect 277236 79332 277304 79388
rect 277360 79332 277428 79388
rect 277484 79332 277552 79388
rect 277608 79332 277676 79388
rect 277732 79332 277800 79388
rect 277856 79332 277924 79388
rect 277980 79332 278048 79388
rect 278104 79332 278172 79388
rect 278228 79332 278296 79388
rect 278352 79332 278420 79388
rect 278476 79332 278544 79388
rect 278600 79332 278668 79388
rect 278724 79332 278792 79388
rect 278848 79332 278916 79388
rect 278972 79332 279040 79388
rect 279096 79332 279172 79388
rect 277122 79264 279172 79332
rect 277122 79208 277180 79264
rect 277236 79208 277304 79264
rect 277360 79208 277428 79264
rect 277484 79208 277552 79264
rect 277608 79208 277676 79264
rect 277732 79208 277800 79264
rect 277856 79208 277924 79264
rect 277980 79208 278048 79264
rect 278104 79208 278172 79264
rect 278228 79208 278296 79264
rect 278352 79208 278420 79264
rect 278476 79208 278544 79264
rect 278600 79208 278668 79264
rect 278724 79208 278792 79264
rect 278848 79208 278916 79264
rect 278972 79208 279040 79264
rect 279096 79208 279172 79264
rect 277122 70130 279172 79208
rect 277122 70074 277192 70130
rect 277248 70074 277316 70130
rect 277372 70074 277440 70130
rect 277496 70074 277564 70130
rect 277620 70074 277688 70130
rect 277744 70074 277812 70130
rect 277868 70074 277936 70130
rect 277992 70074 278060 70130
rect 278116 70074 278184 70130
rect 278240 70074 278308 70130
rect 278364 70074 278432 70130
rect 278488 70074 278556 70130
rect 278612 70074 278680 70130
rect 278736 70074 278804 70130
rect 278860 70074 278928 70130
rect 278984 70074 279052 70130
rect 279108 70074 279172 70130
rect 277122 70000 279172 70074
rect 279828 80008 281878 80078
rect 279828 79952 279886 80008
rect 279942 79952 280010 80008
rect 280066 79952 280134 80008
rect 280190 79952 280258 80008
rect 280314 79952 280382 80008
rect 280438 79952 280506 80008
rect 280562 79952 280630 80008
rect 280686 79952 280754 80008
rect 280810 79952 280878 80008
rect 280934 79952 281002 80008
rect 281058 79952 281126 80008
rect 281182 79952 281250 80008
rect 281306 79952 281374 80008
rect 281430 79952 281498 80008
rect 281554 79952 281622 80008
rect 281678 79952 281746 80008
rect 281802 79952 281878 80008
rect 279828 79884 281878 79952
rect 279828 79828 279886 79884
rect 279942 79828 280010 79884
rect 280066 79828 280134 79884
rect 280190 79828 280258 79884
rect 280314 79828 280382 79884
rect 280438 79828 280506 79884
rect 280562 79828 280630 79884
rect 280686 79828 280754 79884
rect 280810 79828 280878 79884
rect 280934 79828 281002 79884
rect 281058 79828 281126 79884
rect 281182 79828 281250 79884
rect 281306 79828 281374 79884
rect 281430 79828 281498 79884
rect 281554 79828 281622 79884
rect 281678 79828 281746 79884
rect 281802 79828 281878 79884
rect 279828 79760 281878 79828
rect 279828 79704 279886 79760
rect 279942 79704 280010 79760
rect 280066 79704 280134 79760
rect 280190 79704 280258 79760
rect 280314 79704 280382 79760
rect 280438 79704 280506 79760
rect 280562 79704 280630 79760
rect 280686 79704 280754 79760
rect 280810 79704 280878 79760
rect 280934 79704 281002 79760
rect 281058 79704 281126 79760
rect 281182 79704 281250 79760
rect 281306 79704 281374 79760
rect 281430 79704 281498 79760
rect 281554 79704 281622 79760
rect 281678 79704 281746 79760
rect 281802 79704 281878 79760
rect 279828 79636 281878 79704
rect 279828 79580 279886 79636
rect 279942 79580 280010 79636
rect 280066 79580 280134 79636
rect 280190 79580 280258 79636
rect 280314 79580 280382 79636
rect 280438 79580 280506 79636
rect 280562 79580 280630 79636
rect 280686 79580 280754 79636
rect 280810 79580 280878 79636
rect 280934 79580 281002 79636
rect 281058 79580 281126 79636
rect 281182 79580 281250 79636
rect 281306 79580 281374 79636
rect 281430 79580 281498 79636
rect 281554 79580 281622 79636
rect 281678 79580 281746 79636
rect 281802 79580 281878 79636
rect 279828 79512 281878 79580
rect 279828 79456 279886 79512
rect 279942 79456 280010 79512
rect 280066 79456 280134 79512
rect 280190 79456 280258 79512
rect 280314 79456 280382 79512
rect 280438 79456 280506 79512
rect 280562 79456 280630 79512
rect 280686 79456 280754 79512
rect 280810 79456 280878 79512
rect 280934 79456 281002 79512
rect 281058 79456 281126 79512
rect 281182 79456 281250 79512
rect 281306 79456 281374 79512
rect 281430 79456 281498 79512
rect 281554 79456 281622 79512
rect 281678 79456 281746 79512
rect 281802 79456 281878 79512
rect 279828 79388 281878 79456
rect 279828 79332 279886 79388
rect 279942 79332 280010 79388
rect 280066 79332 280134 79388
rect 280190 79332 280258 79388
rect 280314 79332 280382 79388
rect 280438 79332 280506 79388
rect 280562 79332 280630 79388
rect 280686 79332 280754 79388
rect 280810 79332 280878 79388
rect 280934 79332 281002 79388
rect 281058 79332 281126 79388
rect 281182 79332 281250 79388
rect 281306 79332 281374 79388
rect 281430 79332 281498 79388
rect 281554 79332 281622 79388
rect 281678 79332 281746 79388
rect 281802 79332 281878 79388
rect 279828 79264 281878 79332
rect 279828 79208 279886 79264
rect 279942 79208 280010 79264
rect 280066 79208 280134 79264
rect 280190 79208 280258 79264
rect 280314 79208 280382 79264
rect 280438 79208 280506 79264
rect 280562 79208 280630 79264
rect 280686 79208 280754 79264
rect 280810 79208 280878 79264
rect 280934 79208 281002 79264
rect 281058 79208 281126 79264
rect 281182 79208 281250 79264
rect 281306 79208 281374 79264
rect 281430 79208 281498 79264
rect 281554 79208 281622 79264
rect 281678 79208 281746 79264
rect 281802 79208 281878 79264
rect 279828 70130 281878 79208
rect 279828 70074 279892 70130
rect 279948 70074 280016 70130
rect 280072 70074 280140 70130
rect 280196 70074 280264 70130
rect 280320 70074 280388 70130
rect 280444 70074 280512 70130
rect 280568 70074 280636 70130
rect 280692 70074 280760 70130
rect 280816 70074 280884 70130
rect 280940 70074 281008 70130
rect 281064 70074 281132 70130
rect 281188 70074 281256 70130
rect 281312 70074 281380 70130
rect 281436 70074 281504 70130
rect 281560 70074 281628 70130
rect 281684 70074 281752 70130
rect 281808 70074 281878 70130
rect 279828 70000 281878 70074
rect 282198 80008 284248 80078
rect 282198 79952 282256 80008
rect 282312 79952 282380 80008
rect 282436 79952 282504 80008
rect 282560 79952 282628 80008
rect 282684 79952 282752 80008
rect 282808 79952 282876 80008
rect 282932 79952 283000 80008
rect 283056 79952 283124 80008
rect 283180 79952 283248 80008
rect 283304 79952 283372 80008
rect 283428 79952 283496 80008
rect 283552 79952 283620 80008
rect 283676 79952 283744 80008
rect 283800 79952 283868 80008
rect 283924 79952 283992 80008
rect 284048 79952 284116 80008
rect 284172 79952 284248 80008
rect 282198 79884 284248 79952
rect 282198 79828 282256 79884
rect 282312 79828 282380 79884
rect 282436 79828 282504 79884
rect 282560 79828 282628 79884
rect 282684 79828 282752 79884
rect 282808 79828 282876 79884
rect 282932 79828 283000 79884
rect 283056 79828 283124 79884
rect 283180 79828 283248 79884
rect 283304 79828 283372 79884
rect 283428 79828 283496 79884
rect 283552 79828 283620 79884
rect 283676 79828 283744 79884
rect 283800 79828 283868 79884
rect 283924 79828 283992 79884
rect 284048 79828 284116 79884
rect 284172 79828 284248 79884
rect 282198 79760 284248 79828
rect 282198 79704 282256 79760
rect 282312 79704 282380 79760
rect 282436 79704 282504 79760
rect 282560 79704 282628 79760
rect 282684 79704 282752 79760
rect 282808 79704 282876 79760
rect 282932 79704 283000 79760
rect 283056 79704 283124 79760
rect 283180 79704 283248 79760
rect 283304 79704 283372 79760
rect 283428 79704 283496 79760
rect 283552 79704 283620 79760
rect 283676 79704 283744 79760
rect 283800 79704 283868 79760
rect 283924 79704 283992 79760
rect 284048 79704 284116 79760
rect 284172 79704 284248 79760
rect 282198 79636 284248 79704
rect 282198 79580 282256 79636
rect 282312 79580 282380 79636
rect 282436 79580 282504 79636
rect 282560 79580 282628 79636
rect 282684 79580 282752 79636
rect 282808 79580 282876 79636
rect 282932 79580 283000 79636
rect 283056 79580 283124 79636
rect 283180 79580 283248 79636
rect 283304 79580 283372 79636
rect 283428 79580 283496 79636
rect 283552 79580 283620 79636
rect 283676 79580 283744 79636
rect 283800 79580 283868 79636
rect 283924 79580 283992 79636
rect 284048 79580 284116 79636
rect 284172 79580 284248 79636
rect 282198 79512 284248 79580
rect 282198 79456 282256 79512
rect 282312 79456 282380 79512
rect 282436 79456 282504 79512
rect 282560 79456 282628 79512
rect 282684 79456 282752 79512
rect 282808 79456 282876 79512
rect 282932 79456 283000 79512
rect 283056 79456 283124 79512
rect 283180 79456 283248 79512
rect 283304 79456 283372 79512
rect 283428 79456 283496 79512
rect 283552 79456 283620 79512
rect 283676 79456 283744 79512
rect 283800 79456 283868 79512
rect 283924 79456 283992 79512
rect 284048 79456 284116 79512
rect 284172 79456 284248 79512
rect 282198 79388 284248 79456
rect 282198 79332 282256 79388
rect 282312 79332 282380 79388
rect 282436 79332 282504 79388
rect 282560 79332 282628 79388
rect 282684 79332 282752 79388
rect 282808 79332 282876 79388
rect 282932 79332 283000 79388
rect 283056 79332 283124 79388
rect 283180 79332 283248 79388
rect 283304 79332 283372 79388
rect 283428 79332 283496 79388
rect 283552 79332 283620 79388
rect 283676 79332 283744 79388
rect 283800 79332 283868 79388
rect 283924 79332 283992 79388
rect 284048 79332 284116 79388
rect 284172 79332 284248 79388
rect 282198 79264 284248 79332
rect 282198 79208 282256 79264
rect 282312 79208 282380 79264
rect 282436 79208 282504 79264
rect 282560 79208 282628 79264
rect 282684 79208 282752 79264
rect 282808 79208 282876 79264
rect 282932 79208 283000 79264
rect 283056 79208 283124 79264
rect 283180 79208 283248 79264
rect 283304 79208 283372 79264
rect 283428 79208 283496 79264
rect 283552 79208 283620 79264
rect 283676 79208 283744 79264
rect 283800 79208 283868 79264
rect 283924 79208 283992 79264
rect 284048 79208 284116 79264
rect 284172 79208 284248 79264
rect 282198 70130 284248 79208
rect 282198 70074 282262 70130
rect 282318 70074 282386 70130
rect 282442 70074 282510 70130
rect 282566 70074 282634 70130
rect 282690 70074 282758 70130
rect 282814 70074 282882 70130
rect 282938 70074 283006 70130
rect 283062 70074 283130 70130
rect 283186 70074 283254 70130
rect 283310 70074 283378 70130
rect 283434 70074 283502 70130
rect 283558 70074 283626 70130
rect 283682 70074 283750 70130
rect 283806 70074 283874 70130
rect 283930 70074 283998 70130
rect 284054 70074 284122 70130
rect 284178 70074 284248 70130
rect 282198 70000 284248 70074
rect 284828 80008 286728 80078
rect 284828 79952 284860 80008
rect 284916 79952 284984 80008
rect 285040 79952 285108 80008
rect 285164 79952 285232 80008
rect 285288 79952 285356 80008
rect 285412 79952 285480 80008
rect 285536 79952 285604 80008
rect 285660 79952 285728 80008
rect 285784 79952 285852 80008
rect 285908 79952 285976 80008
rect 286032 79952 286100 80008
rect 286156 79952 286224 80008
rect 286280 79952 286348 80008
rect 286404 79952 286472 80008
rect 286528 79952 286596 80008
rect 286652 79952 286728 80008
rect 284828 79884 286728 79952
rect 284828 79828 284860 79884
rect 284916 79828 284984 79884
rect 285040 79828 285108 79884
rect 285164 79828 285232 79884
rect 285288 79828 285356 79884
rect 285412 79828 285480 79884
rect 285536 79828 285604 79884
rect 285660 79828 285728 79884
rect 285784 79828 285852 79884
rect 285908 79828 285976 79884
rect 286032 79828 286100 79884
rect 286156 79828 286224 79884
rect 286280 79828 286348 79884
rect 286404 79828 286472 79884
rect 286528 79828 286596 79884
rect 286652 79828 286728 79884
rect 284828 79760 286728 79828
rect 284828 79704 284860 79760
rect 284916 79704 284984 79760
rect 285040 79704 285108 79760
rect 285164 79704 285232 79760
rect 285288 79704 285356 79760
rect 285412 79704 285480 79760
rect 285536 79704 285604 79760
rect 285660 79704 285728 79760
rect 285784 79704 285852 79760
rect 285908 79704 285976 79760
rect 286032 79704 286100 79760
rect 286156 79704 286224 79760
rect 286280 79704 286348 79760
rect 286404 79704 286472 79760
rect 286528 79704 286596 79760
rect 286652 79704 286728 79760
rect 284828 79636 286728 79704
rect 284828 79580 284860 79636
rect 284916 79580 284984 79636
rect 285040 79580 285108 79636
rect 285164 79580 285232 79636
rect 285288 79580 285356 79636
rect 285412 79580 285480 79636
rect 285536 79580 285604 79636
rect 285660 79580 285728 79636
rect 285784 79580 285852 79636
rect 285908 79580 285976 79636
rect 286032 79580 286100 79636
rect 286156 79580 286224 79636
rect 286280 79580 286348 79636
rect 286404 79580 286472 79636
rect 286528 79580 286596 79636
rect 286652 79580 286728 79636
rect 284828 79512 286728 79580
rect 284828 79456 284860 79512
rect 284916 79456 284984 79512
rect 285040 79456 285108 79512
rect 285164 79456 285232 79512
rect 285288 79456 285356 79512
rect 285412 79456 285480 79512
rect 285536 79456 285604 79512
rect 285660 79456 285728 79512
rect 285784 79456 285852 79512
rect 285908 79456 285976 79512
rect 286032 79456 286100 79512
rect 286156 79456 286224 79512
rect 286280 79456 286348 79512
rect 286404 79456 286472 79512
rect 286528 79456 286596 79512
rect 286652 79456 286728 79512
rect 284828 79388 286728 79456
rect 284828 79332 284860 79388
rect 284916 79332 284984 79388
rect 285040 79332 285108 79388
rect 285164 79332 285232 79388
rect 285288 79332 285356 79388
rect 285412 79332 285480 79388
rect 285536 79332 285604 79388
rect 285660 79332 285728 79388
rect 285784 79332 285852 79388
rect 285908 79332 285976 79388
rect 286032 79332 286100 79388
rect 286156 79332 286224 79388
rect 286280 79332 286348 79388
rect 286404 79332 286472 79388
rect 286528 79332 286596 79388
rect 286652 79332 286728 79388
rect 284828 79264 286728 79332
rect 284828 79208 284860 79264
rect 284916 79208 284984 79264
rect 285040 79208 285108 79264
rect 285164 79208 285232 79264
rect 285288 79208 285356 79264
rect 285412 79208 285480 79264
rect 285536 79208 285604 79264
rect 285660 79208 285728 79264
rect 285784 79208 285852 79264
rect 285908 79208 285976 79264
rect 286032 79208 286100 79264
rect 286156 79208 286224 79264
rect 286280 79208 286348 79264
rect 286404 79208 286472 79264
rect 286528 79208 286596 79264
rect 286652 79208 286728 79264
rect 284828 70130 286728 79208
rect 289224 80008 289544 81752
rect 289224 79952 289294 80008
rect 289350 79952 289418 80008
rect 289474 79952 289544 80008
rect 289224 79884 289544 79952
rect 289224 79828 289294 79884
rect 289350 79828 289418 79884
rect 289474 79828 289544 79884
rect 289224 79760 289544 79828
rect 289224 79704 289294 79760
rect 289350 79704 289418 79760
rect 289474 79704 289544 79760
rect 289224 79636 289544 79704
rect 289224 79580 289294 79636
rect 289350 79580 289418 79636
rect 289474 79580 289544 79636
rect 289224 79512 289544 79580
rect 289224 79456 289294 79512
rect 289350 79456 289418 79512
rect 289474 79456 289544 79512
rect 289224 79388 289544 79456
rect 289224 79332 289294 79388
rect 289350 79332 289418 79388
rect 289474 79332 289544 79388
rect 289224 79264 289544 79332
rect 289224 79208 289294 79264
rect 289350 79208 289418 79264
rect 289474 79208 289544 79264
rect 289224 79078 289544 79208
rect 294224 78608 294544 81752
rect 299224 80008 299544 81752
rect 299224 79952 299294 80008
rect 299350 79952 299418 80008
rect 299474 79952 299544 80008
rect 299224 79884 299544 79952
rect 299224 79828 299294 79884
rect 299350 79828 299418 79884
rect 299474 79828 299544 79884
rect 299224 79760 299544 79828
rect 299224 79704 299294 79760
rect 299350 79704 299418 79760
rect 299474 79704 299544 79760
rect 299224 79636 299544 79704
rect 299224 79580 299294 79636
rect 299350 79580 299418 79636
rect 299474 79580 299544 79636
rect 299224 79512 299544 79580
rect 299224 79456 299294 79512
rect 299350 79456 299418 79512
rect 299474 79456 299544 79512
rect 299224 79388 299544 79456
rect 299224 79332 299294 79388
rect 299350 79332 299418 79388
rect 299474 79332 299544 79388
rect 299224 79264 299544 79332
rect 299224 79208 299294 79264
rect 299350 79208 299418 79264
rect 299474 79208 299544 79264
rect 299224 79078 299544 79208
rect 294224 78552 294294 78608
rect 294350 78552 294418 78608
rect 294474 78552 294544 78608
rect 294224 78484 294544 78552
rect 294224 78428 294294 78484
rect 294350 78428 294418 78484
rect 294474 78428 294544 78484
rect 294224 78360 294544 78428
rect 294224 78304 294294 78360
rect 294350 78304 294418 78360
rect 294474 78304 294544 78360
rect 294224 78236 294544 78304
rect 294224 78180 294294 78236
rect 294350 78180 294418 78236
rect 294474 78180 294544 78236
rect 294224 78112 294544 78180
rect 294224 78056 294294 78112
rect 294350 78056 294418 78112
rect 294474 78056 294544 78112
rect 294224 77988 294544 78056
rect 294224 77932 294294 77988
rect 294350 77932 294418 77988
rect 294474 77932 294544 77988
rect 294224 77864 294544 77932
rect 294224 77808 294294 77864
rect 294350 77808 294418 77864
rect 294474 77808 294544 77864
rect 294224 77678 294544 77808
rect 304224 78608 304544 81752
rect 309224 80008 309544 81752
rect 309224 79952 309294 80008
rect 309350 79952 309418 80008
rect 309474 79952 309544 80008
rect 309224 79884 309544 79952
rect 309224 79828 309294 79884
rect 309350 79828 309418 79884
rect 309474 79828 309544 79884
rect 309224 79760 309544 79828
rect 309224 79704 309294 79760
rect 309350 79704 309418 79760
rect 309474 79704 309544 79760
rect 309224 79636 309544 79704
rect 309224 79580 309294 79636
rect 309350 79580 309418 79636
rect 309474 79580 309544 79636
rect 309224 79512 309544 79580
rect 309224 79456 309294 79512
rect 309350 79456 309418 79512
rect 309474 79456 309544 79512
rect 309224 79388 309544 79456
rect 309224 79332 309294 79388
rect 309350 79332 309418 79388
rect 309474 79332 309544 79388
rect 309224 79264 309544 79332
rect 309224 79208 309294 79264
rect 309350 79208 309418 79264
rect 309474 79208 309544 79264
rect 309224 79078 309544 79208
rect 304224 78552 304294 78608
rect 304350 78552 304418 78608
rect 304474 78552 304544 78608
rect 304224 78484 304544 78552
rect 304224 78428 304294 78484
rect 304350 78428 304418 78484
rect 304474 78428 304544 78484
rect 304224 78360 304544 78428
rect 304224 78304 304294 78360
rect 304350 78304 304418 78360
rect 304474 78304 304544 78360
rect 304224 78236 304544 78304
rect 304224 78180 304294 78236
rect 304350 78180 304418 78236
rect 304474 78180 304544 78236
rect 304224 78112 304544 78180
rect 304224 78056 304294 78112
rect 304350 78056 304418 78112
rect 304474 78056 304544 78112
rect 304224 77988 304544 78056
rect 304224 77932 304294 77988
rect 304350 77932 304418 77988
rect 304474 77932 304544 77988
rect 304224 77864 304544 77932
rect 304224 77808 304294 77864
rect 304350 77808 304418 77864
rect 304474 77808 304544 77864
rect 304224 77678 304544 77808
rect 314224 78608 314544 81752
rect 319224 80008 319544 81752
rect 319224 79952 319294 80008
rect 319350 79952 319418 80008
rect 319474 79952 319544 80008
rect 319224 79884 319544 79952
rect 319224 79828 319294 79884
rect 319350 79828 319418 79884
rect 319474 79828 319544 79884
rect 319224 79760 319544 79828
rect 319224 79704 319294 79760
rect 319350 79704 319418 79760
rect 319474 79704 319544 79760
rect 319224 79636 319544 79704
rect 319224 79580 319294 79636
rect 319350 79580 319418 79636
rect 319474 79580 319544 79636
rect 319224 79512 319544 79580
rect 319224 79456 319294 79512
rect 319350 79456 319418 79512
rect 319474 79456 319544 79512
rect 319224 79388 319544 79456
rect 319224 79332 319294 79388
rect 319350 79332 319418 79388
rect 319474 79332 319544 79388
rect 319224 79264 319544 79332
rect 319224 79208 319294 79264
rect 319350 79208 319418 79264
rect 319474 79208 319544 79264
rect 319224 79078 319544 79208
rect 314224 78552 314294 78608
rect 314350 78552 314418 78608
rect 314474 78552 314544 78608
rect 314224 78484 314544 78552
rect 314224 78428 314294 78484
rect 314350 78428 314418 78484
rect 314474 78428 314544 78484
rect 314224 78360 314544 78428
rect 314224 78304 314294 78360
rect 314350 78304 314418 78360
rect 314474 78304 314544 78360
rect 314224 78236 314544 78304
rect 314224 78180 314294 78236
rect 314350 78180 314418 78236
rect 314474 78180 314544 78236
rect 314224 78112 314544 78180
rect 314224 78056 314294 78112
rect 314350 78056 314418 78112
rect 314474 78056 314544 78112
rect 314224 77988 314544 78056
rect 314224 77932 314294 77988
rect 314350 77932 314418 77988
rect 314474 77932 314544 77988
rect 314224 77864 314544 77932
rect 314224 77808 314294 77864
rect 314350 77808 314418 77864
rect 314474 77808 314544 77864
rect 314224 77678 314544 77808
rect 324224 78608 324544 81752
rect 329224 80008 329544 81752
rect 329224 79952 329294 80008
rect 329350 79952 329418 80008
rect 329474 79952 329544 80008
rect 329224 79884 329544 79952
rect 329224 79828 329294 79884
rect 329350 79828 329418 79884
rect 329474 79828 329544 79884
rect 329224 79760 329544 79828
rect 329224 79704 329294 79760
rect 329350 79704 329418 79760
rect 329474 79704 329544 79760
rect 329224 79636 329544 79704
rect 329224 79580 329294 79636
rect 329350 79580 329418 79636
rect 329474 79580 329544 79636
rect 329224 79512 329544 79580
rect 329224 79456 329294 79512
rect 329350 79456 329418 79512
rect 329474 79456 329544 79512
rect 329224 79388 329544 79456
rect 329224 79332 329294 79388
rect 329350 79332 329418 79388
rect 329474 79332 329544 79388
rect 329224 79264 329544 79332
rect 329224 79208 329294 79264
rect 329350 79208 329418 79264
rect 329474 79208 329544 79264
rect 329224 79078 329544 79208
rect 324224 78552 324294 78608
rect 324350 78552 324418 78608
rect 324474 78552 324544 78608
rect 324224 78484 324544 78552
rect 324224 78428 324294 78484
rect 324350 78428 324418 78484
rect 324474 78428 324544 78484
rect 324224 78360 324544 78428
rect 324224 78304 324294 78360
rect 324350 78304 324418 78360
rect 324474 78304 324544 78360
rect 324224 78236 324544 78304
rect 324224 78180 324294 78236
rect 324350 78180 324418 78236
rect 324474 78180 324544 78236
rect 324224 78112 324544 78180
rect 324224 78056 324294 78112
rect 324350 78056 324418 78112
rect 324474 78056 324544 78112
rect 324224 77988 324544 78056
rect 324224 77932 324294 77988
rect 324350 77932 324418 77988
rect 324474 77932 324544 77988
rect 324224 77864 324544 77932
rect 324224 77808 324294 77864
rect 324350 77808 324418 77864
rect 324474 77808 324544 77864
rect 324224 77678 324544 77808
rect 334224 78608 334544 81752
rect 339224 80008 339544 81752
rect 339224 79952 339294 80008
rect 339350 79952 339418 80008
rect 339474 79952 339544 80008
rect 339224 79884 339544 79952
rect 339224 79828 339294 79884
rect 339350 79828 339418 79884
rect 339474 79828 339544 79884
rect 339224 79760 339544 79828
rect 339224 79704 339294 79760
rect 339350 79704 339418 79760
rect 339474 79704 339544 79760
rect 339224 79636 339544 79704
rect 339224 79580 339294 79636
rect 339350 79580 339418 79636
rect 339474 79580 339544 79636
rect 339224 79512 339544 79580
rect 339224 79456 339294 79512
rect 339350 79456 339418 79512
rect 339474 79456 339544 79512
rect 339224 79388 339544 79456
rect 339224 79332 339294 79388
rect 339350 79332 339418 79388
rect 339474 79332 339544 79388
rect 339224 79264 339544 79332
rect 339224 79208 339294 79264
rect 339350 79208 339418 79264
rect 339474 79208 339544 79264
rect 339224 79078 339544 79208
rect 334224 78552 334294 78608
rect 334350 78552 334418 78608
rect 334474 78552 334544 78608
rect 334224 78484 334544 78552
rect 334224 78428 334294 78484
rect 334350 78428 334418 78484
rect 334474 78428 334544 78484
rect 334224 78360 334544 78428
rect 334224 78304 334294 78360
rect 334350 78304 334418 78360
rect 334474 78304 334544 78360
rect 334224 78236 334544 78304
rect 334224 78180 334294 78236
rect 334350 78180 334418 78236
rect 334474 78180 334544 78236
rect 334224 78112 334544 78180
rect 334224 78056 334294 78112
rect 334350 78056 334418 78112
rect 334474 78056 334544 78112
rect 334224 77988 334544 78056
rect 334224 77932 334294 77988
rect 334350 77932 334418 77988
rect 334474 77932 334544 77988
rect 334224 77864 334544 77932
rect 334224 77808 334294 77864
rect 334350 77808 334418 77864
rect 334474 77808 334544 77864
rect 334224 77678 334544 77808
rect 344224 78608 344544 81752
rect 349224 80008 349544 81752
rect 349224 79952 349294 80008
rect 349350 79952 349418 80008
rect 349474 79952 349544 80008
rect 349224 79884 349544 79952
rect 349224 79828 349294 79884
rect 349350 79828 349418 79884
rect 349474 79828 349544 79884
rect 349224 79760 349544 79828
rect 349224 79704 349294 79760
rect 349350 79704 349418 79760
rect 349474 79704 349544 79760
rect 349224 79636 349544 79704
rect 349224 79580 349294 79636
rect 349350 79580 349418 79636
rect 349474 79580 349544 79636
rect 349224 79512 349544 79580
rect 349224 79456 349294 79512
rect 349350 79456 349418 79512
rect 349474 79456 349544 79512
rect 349224 79388 349544 79456
rect 349224 79332 349294 79388
rect 349350 79332 349418 79388
rect 349474 79332 349544 79388
rect 349224 79264 349544 79332
rect 349224 79208 349294 79264
rect 349350 79208 349418 79264
rect 349474 79208 349544 79264
rect 349224 79078 349544 79208
rect 344224 78552 344294 78608
rect 344350 78552 344418 78608
rect 344474 78552 344544 78608
rect 344224 78484 344544 78552
rect 344224 78428 344294 78484
rect 344350 78428 344418 78484
rect 344474 78428 344544 78484
rect 344224 78360 344544 78428
rect 344224 78304 344294 78360
rect 344350 78304 344418 78360
rect 344474 78304 344544 78360
rect 344224 78236 344544 78304
rect 344224 78180 344294 78236
rect 344350 78180 344418 78236
rect 344474 78180 344544 78236
rect 344224 78112 344544 78180
rect 344224 78056 344294 78112
rect 344350 78056 344418 78112
rect 344474 78056 344544 78112
rect 344224 77988 344544 78056
rect 344224 77932 344294 77988
rect 344350 77932 344418 77988
rect 344474 77932 344544 77988
rect 344224 77864 344544 77932
rect 344224 77808 344294 77864
rect 344350 77808 344418 77864
rect 344474 77808 344544 77864
rect 344224 77678 344544 77808
rect 354224 78608 354544 81752
rect 359224 80008 359544 81752
rect 359224 79952 359294 80008
rect 359350 79952 359418 80008
rect 359474 79952 359544 80008
rect 359224 79884 359544 79952
rect 359224 79828 359294 79884
rect 359350 79828 359418 79884
rect 359474 79828 359544 79884
rect 359224 79760 359544 79828
rect 359224 79704 359294 79760
rect 359350 79704 359418 79760
rect 359474 79704 359544 79760
rect 359224 79636 359544 79704
rect 359224 79580 359294 79636
rect 359350 79580 359418 79636
rect 359474 79580 359544 79636
rect 359224 79512 359544 79580
rect 359224 79456 359294 79512
rect 359350 79456 359418 79512
rect 359474 79456 359544 79512
rect 359224 79388 359544 79456
rect 359224 79332 359294 79388
rect 359350 79332 359418 79388
rect 359474 79332 359544 79388
rect 359224 79264 359544 79332
rect 359224 79208 359294 79264
rect 359350 79208 359418 79264
rect 359474 79208 359544 79264
rect 359224 79078 359544 79208
rect 354224 78552 354294 78608
rect 354350 78552 354418 78608
rect 354474 78552 354544 78608
rect 354224 78484 354544 78552
rect 354224 78428 354294 78484
rect 354350 78428 354418 78484
rect 354474 78428 354544 78484
rect 354224 78360 354544 78428
rect 354224 78304 354294 78360
rect 354350 78304 354418 78360
rect 354474 78304 354544 78360
rect 354224 78236 354544 78304
rect 354224 78180 354294 78236
rect 354350 78180 354418 78236
rect 354474 78180 354544 78236
rect 354224 78112 354544 78180
rect 354224 78056 354294 78112
rect 354350 78056 354418 78112
rect 354474 78056 354544 78112
rect 354224 77988 354544 78056
rect 354224 77932 354294 77988
rect 354350 77932 354418 77988
rect 354474 77932 354544 77988
rect 354224 77864 354544 77932
rect 354224 77808 354294 77864
rect 354350 77808 354418 77864
rect 354474 77808 354544 77864
rect 354224 77678 354544 77808
rect 364224 78608 364544 81752
rect 369224 80008 369544 81752
rect 369224 79952 369294 80008
rect 369350 79952 369418 80008
rect 369474 79952 369544 80008
rect 369224 79884 369544 79952
rect 369224 79828 369294 79884
rect 369350 79828 369418 79884
rect 369474 79828 369544 79884
rect 369224 79760 369544 79828
rect 369224 79704 369294 79760
rect 369350 79704 369418 79760
rect 369474 79704 369544 79760
rect 369224 79636 369544 79704
rect 369224 79580 369294 79636
rect 369350 79580 369418 79636
rect 369474 79580 369544 79636
rect 369224 79512 369544 79580
rect 369224 79456 369294 79512
rect 369350 79456 369418 79512
rect 369474 79456 369544 79512
rect 369224 79388 369544 79456
rect 369224 79332 369294 79388
rect 369350 79332 369418 79388
rect 369474 79332 369544 79388
rect 369224 79264 369544 79332
rect 369224 79208 369294 79264
rect 369350 79208 369418 79264
rect 369474 79208 369544 79264
rect 369224 79078 369544 79208
rect 364224 78552 364294 78608
rect 364350 78552 364418 78608
rect 364474 78552 364544 78608
rect 364224 78484 364544 78552
rect 364224 78428 364294 78484
rect 364350 78428 364418 78484
rect 364474 78428 364544 78484
rect 364224 78360 364544 78428
rect 364224 78304 364294 78360
rect 364350 78304 364418 78360
rect 364474 78304 364544 78360
rect 364224 78236 364544 78304
rect 364224 78180 364294 78236
rect 364350 78180 364418 78236
rect 364474 78180 364544 78236
rect 364224 78112 364544 78180
rect 364224 78056 364294 78112
rect 364350 78056 364418 78112
rect 364474 78056 364544 78112
rect 364224 77988 364544 78056
rect 364224 77932 364294 77988
rect 364350 77932 364418 77988
rect 364474 77932 364544 77988
rect 364224 77864 364544 77932
rect 364224 77808 364294 77864
rect 364350 77808 364418 77864
rect 364474 77808 364544 77864
rect 364224 77678 364544 77808
rect 374224 78608 374544 81752
rect 379224 80008 379544 81752
rect 379224 79952 379294 80008
rect 379350 79952 379418 80008
rect 379474 79952 379544 80008
rect 379224 79884 379544 79952
rect 379224 79828 379294 79884
rect 379350 79828 379418 79884
rect 379474 79828 379544 79884
rect 379224 79760 379544 79828
rect 379224 79704 379294 79760
rect 379350 79704 379418 79760
rect 379474 79704 379544 79760
rect 379224 79636 379544 79704
rect 379224 79580 379294 79636
rect 379350 79580 379418 79636
rect 379474 79580 379544 79636
rect 379224 79512 379544 79580
rect 379224 79456 379294 79512
rect 379350 79456 379418 79512
rect 379474 79456 379544 79512
rect 379224 79388 379544 79456
rect 379224 79332 379294 79388
rect 379350 79332 379418 79388
rect 379474 79332 379544 79388
rect 379224 79264 379544 79332
rect 379224 79208 379294 79264
rect 379350 79208 379418 79264
rect 379474 79208 379544 79264
rect 379224 79078 379544 79208
rect 374224 78552 374294 78608
rect 374350 78552 374418 78608
rect 374474 78552 374544 78608
rect 374224 78484 374544 78552
rect 374224 78428 374294 78484
rect 374350 78428 374418 78484
rect 374474 78428 374544 78484
rect 374224 78360 374544 78428
rect 374224 78304 374294 78360
rect 374350 78304 374418 78360
rect 374474 78304 374544 78360
rect 374224 78236 374544 78304
rect 374224 78180 374294 78236
rect 374350 78180 374418 78236
rect 374474 78180 374544 78236
rect 374224 78112 374544 78180
rect 374224 78056 374294 78112
rect 374350 78056 374418 78112
rect 374474 78056 374544 78112
rect 374224 77988 374544 78056
rect 374224 77932 374294 77988
rect 374350 77932 374418 77988
rect 374474 77932 374544 77988
rect 374224 77864 374544 77932
rect 374224 77808 374294 77864
rect 374350 77808 374418 77864
rect 374474 77808 374544 77864
rect 374224 77678 374544 77808
rect 384224 78608 384544 81752
rect 389224 80008 389544 81752
rect 389224 79952 389294 80008
rect 389350 79952 389418 80008
rect 389474 79952 389544 80008
rect 389224 79884 389544 79952
rect 389224 79828 389294 79884
rect 389350 79828 389418 79884
rect 389474 79828 389544 79884
rect 389224 79760 389544 79828
rect 389224 79704 389294 79760
rect 389350 79704 389418 79760
rect 389474 79704 389544 79760
rect 389224 79636 389544 79704
rect 389224 79580 389294 79636
rect 389350 79580 389418 79636
rect 389474 79580 389544 79636
rect 389224 79512 389544 79580
rect 389224 79456 389294 79512
rect 389350 79456 389418 79512
rect 389474 79456 389544 79512
rect 389224 79388 389544 79456
rect 389224 79332 389294 79388
rect 389350 79332 389418 79388
rect 389474 79332 389544 79388
rect 389224 79264 389544 79332
rect 389224 79208 389294 79264
rect 389350 79208 389418 79264
rect 389474 79208 389544 79264
rect 389224 79078 389544 79208
rect 384224 78552 384294 78608
rect 384350 78552 384418 78608
rect 384474 78552 384544 78608
rect 384224 78484 384544 78552
rect 384224 78428 384294 78484
rect 384350 78428 384418 78484
rect 384474 78428 384544 78484
rect 384224 78360 384544 78428
rect 384224 78304 384294 78360
rect 384350 78304 384418 78360
rect 384474 78304 384544 78360
rect 384224 78236 384544 78304
rect 384224 78180 384294 78236
rect 384350 78180 384418 78236
rect 384474 78180 384544 78236
rect 384224 78112 384544 78180
rect 384224 78056 384294 78112
rect 384350 78056 384418 78112
rect 384474 78056 384544 78112
rect 384224 77988 384544 78056
rect 384224 77932 384294 77988
rect 384350 77932 384418 77988
rect 384474 77932 384544 77988
rect 384224 77864 384544 77932
rect 384224 77808 384294 77864
rect 384350 77808 384418 77864
rect 384474 77808 384544 77864
rect 384224 77678 384544 77808
rect 394224 78608 394544 81752
rect 399224 80008 399544 81752
rect 399224 79952 399294 80008
rect 399350 79952 399418 80008
rect 399474 79952 399544 80008
rect 399224 79884 399544 79952
rect 399224 79828 399294 79884
rect 399350 79828 399418 79884
rect 399474 79828 399544 79884
rect 399224 79760 399544 79828
rect 399224 79704 399294 79760
rect 399350 79704 399418 79760
rect 399474 79704 399544 79760
rect 399224 79636 399544 79704
rect 399224 79580 399294 79636
rect 399350 79580 399418 79636
rect 399474 79580 399544 79636
rect 399224 79512 399544 79580
rect 399224 79456 399294 79512
rect 399350 79456 399418 79512
rect 399474 79456 399544 79512
rect 399224 79388 399544 79456
rect 399224 79332 399294 79388
rect 399350 79332 399418 79388
rect 399474 79332 399544 79388
rect 399224 79264 399544 79332
rect 399224 79208 399294 79264
rect 399350 79208 399418 79264
rect 399474 79208 399544 79264
rect 399224 79078 399544 79208
rect 394224 78552 394294 78608
rect 394350 78552 394418 78608
rect 394474 78552 394544 78608
rect 394224 78484 394544 78552
rect 394224 78428 394294 78484
rect 394350 78428 394418 78484
rect 394474 78428 394544 78484
rect 394224 78360 394544 78428
rect 394224 78304 394294 78360
rect 394350 78304 394418 78360
rect 394474 78304 394544 78360
rect 394224 78236 394544 78304
rect 394224 78180 394294 78236
rect 394350 78180 394418 78236
rect 394474 78180 394544 78236
rect 394224 78112 394544 78180
rect 394224 78056 394294 78112
rect 394350 78056 394418 78112
rect 394474 78056 394544 78112
rect 394224 77988 394544 78056
rect 394224 77932 394294 77988
rect 394350 77932 394418 77988
rect 394474 77932 394544 77988
rect 394224 77864 394544 77932
rect 394224 77808 394294 77864
rect 394350 77808 394418 77864
rect 394474 77808 394544 77864
rect 394224 77678 394544 77808
rect 404224 78608 404544 81752
rect 409224 80008 409544 81752
rect 409224 79952 409294 80008
rect 409350 79952 409418 80008
rect 409474 79952 409544 80008
rect 409224 79884 409544 79952
rect 409224 79828 409294 79884
rect 409350 79828 409418 79884
rect 409474 79828 409544 79884
rect 409224 79760 409544 79828
rect 409224 79704 409294 79760
rect 409350 79704 409418 79760
rect 409474 79704 409544 79760
rect 409224 79636 409544 79704
rect 409224 79580 409294 79636
rect 409350 79580 409418 79636
rect 409474 79580 409544 79636
rect 409224 79512 409544 79580
rect 409224 79456 409294 79512
rect 409350 79456 409418 79512
rect 409474 79456 409544 79512
rect 409224 79388 409544 79456
rect 409224 79332 409294 79388
rect 409350 79332 409418 79388
rect 409474 79332 409544 79388
rect 409224 79264 409544 79332
rect 409224 79208 409294 79264
rect 409350 79208 409418 79264
rect 409474 79208 409544 79264
rect 409224 79078 409544 79208
rect 404224 78552 404294 78608
rect 404350 78552 404418 78608
rect 404474 78552 404544 78608
rect 404224 78484 404544 78552
rect 404224 78428 404294 78484
rect 404350 78428 404418 78484
rect 404474 78428 404544 78484
rect 404224 78360 404544 78428
rect 404224 78304 404294 78360
rect 404350 78304 404418 78360
rect 404474 78304 404544 78360
rect 404224 78236 404544 78304
rect 404224 78180 404294 78236
rect 404350 78180 404418 78236
rect 404474 78180 404544 78236
rect 404224 78112 404544 78180
rect 404224 78056 404294 78112
rect 404350 78056 404418 78112
rect 404474 78056 404544 78112
rect 404224 77988 404544 78056
rect 404224 77932 404294 77988
rect 404350 77932 404418 77988
rect 404474 77932 404544 77988
rect 404224 77864 404544 77932
rect 404224 77808 404294 77864
rect 404350 77808 404418 77864
rect 404474 77808 404544 77864
rect 404224 77678 404544 77808
rect 414224 78608 414544 81752
rect 419224 80008 419544 81752
rect 419224 79952 419294 80008
rect 419350 79952 419418 80008
rect 419474 79952 419544 80008
rect 419224 79884 419544 79952
rect 419224 79828 419294 79884
rect 419350 79828 419418 79884
rect 419474 79828 419544 79884
rect 419224 79760 419544 79828
rect 419224 79704 419294 79760
rect 419350 79704 419418 79760
rect 419474 79704 419544 79760
rect 419224 79636 419544 79704
rect 419224 79580 419294 79636
rect 419350 79580 419418 79636
rect 419474 79580 419544 79636
rect 419224 79512 419544 79580
rect 419224 79456 419294 79512
rect 419350 79456 419418 79512
rect 419474 79456 419544 79512
rect 419224 79388 419544 79456
rect 419224 79332 419294 79388
rect 419350 79332 419418 79388
rect 419474 79332 419544 79388
rect 419224 79264 419544 79332
rect 419224 79208 419294 79264
rect 419350 79208 419418 79264
rect 419474 79208 419544 79264
rect 419224 79078 419544 79208
rect 414224 78552 414294 78608
rect 414350 78552 414418 78608
rect 414474 78552 414544 78608
rect 414224 78484 414544 78552
rect 414224 78428 414294 78484
rect 414350 78428 414418 78484
rect 414474 78428 414544 78484
rect 414224 78360 414544 78428
rect 414224 78304 414294 78360
rect 414350 78304 414418 78360
rect 414474 78304 414544 78360
rect 414224 78236 414544 78304
rect 414224 78180 414294 78236
rect 414350 78180 414418 78236
rect 414474 78180 414544 78236
rect 414224 78112 414544 78180
rect 414224 78056 414294 78112
rect 414350 78056 414418 78112
rect 414474 78056 414544 78112
rect 414224 77988 414544 78056
rect 414224 77932 414294 77988
rect 414350 77932 414418 77988
rect 414474 77932 414544 77988
rect 414224 77864 414544 77932
rect 414224 77808 414294 77864
rect 414350 77808 414418 77864
rect 414474 77808 414544 77864
rect 414224 77678 414544 77808
rect 424224 78608 424544 81752
rect 429224 80008 429544 81752
rect 429224 79952 429294 80008
rect 429350 79952 429418 80008
rect 429474 79952 429544 80008
rect 429224 79884 429544 79952
rect 429224 79828 429294 79884
rect 429350 79828 429418 79884
rect 429474 79828 429544 79884
rect 429224 79760 429544 79828
rect 429224 79704 429294 79760
rect 429350 79704 429418 79760
rect 429474 79704 429544 79760
rect 429224 79636 429544 79704
rect 429224 79580 429294 79636
rect 429350 79580 429418 79636
rect 429474 79580 429544 79636
rect 429224 79512 429544 79580
rect 429224 79456 429294 79512
rect 429350 79456 429418 79512
rect 429474 79456 429544 79512
rect 429224 79388 429544 79456
rect 429224 79332 429294 79388
rect 429350 79332 429418 79388
rect 429474 79332 429544 79388
rect 429224 79264 429544 79332
rect 429224 79208 429294 79264
rect 429350 79208 429418 79264
rect 429474 79208 429544 79264
rect 429224 79078 429544 79208
rect 424224 78552 424294 78608
rect 424350 78552 424418 78608
rect 424474 78552 424544 78608
rect 424224 78484 424544 78552
rect 424224 78428 424294 78484
rect 424350 78428 424418 78484
rect 424474 78428 424544 78484
rect 424224 78360 424544 78428
rect 424224 78304 424294 78360
rect 424350 78304 424418 78360
rect 424474 78304 424544 78360
rect 424224 78236 424544 78304
rect 424224 78180 424294 78236
rect 424350 78180 424418 78236
rect 424474 78180 424544 78236
rect 424224 78112 424544 78180
rect 424224 78056 424294 78112
rect 424350 78056 424418 78112
rect 424474 78056 424544 78112
rect 424224 77988 424544 78056
rect 424224 77932 424294 77988
rect 424350 77932 424418 77988
rect 424474 77932 424544 77988
rect 424224 77864 424544 77932
rect 424224 77808 424294 77864
rect 424350 77808 424418 77864
rect 424474 77808 424544 77864
rect 424224 77678 424544 77808
rect 434224 78608 434544 81752
rect 439224 80008 439544 81752
rect 439224 79952 439294 80008
rect 439350 79952 439418 80008
rect 439474 79952 439544 80008
rect 439224 79884 439544 79952
rect 439224 79828 439294 79884
rect 439350 79828 439418 79884
rect 439474 79828 439544 79884
rect 439224 79760 439544 79828
rect 439224 79704 439294 79760
rect 439350 79704 439418 79760
rect 439474 79704 439544 79760
rect 439224 79636 439544 79704
rect 439224 79580 439294 79636
rect 439350 79580 439418 79636
rect 439474 79580 439544 79636
rect 439224 79512 439544 79580
rect 439224 79456 439294 79512
rect 439350 79456 439418 79512
rect 439474 79456 439544 79512
rect 439224 79388 439544 79456
rect 439224 79332 439294 79388
rect 439350 79332 439418 79388
rect 439474 79332 439544 79388
rect 439224 79264 439544 79332
rect 439224 79208 439294 79264
rect 439350 79208 439418 79264
rect 439474 79208 439544 79264
rect 439224 79078 439544 79208
rect 434224 78552 434294 78608
rect 434350 78552 434418 78608
rect 434474 78552 434544 78608
rect 434224 78484 434544 78552
rect 434224 78428 434294 78484
rect 434350 78428 434418 78484
rect 434474 78428 434544 78484
rect 434224 78360 434544 78428
rect 434224 78304 434294 78360
rect 434350 78304 434418 78360
rect 434474 78304 434544 78360
rect 434224 78236 434544 78304
rect 434224 78180 434294 78236
rect 434350 78180 434418 78236
rect 434474 78180 434544 78236
rect 434224 78112 434544 78180
rect 434224 78056 434294 78112
rect 434350 78056 434418 78112
rect 434474 78056 434544 78112
rect 434224 77988 434544 78056
rect 434224 77932 434294 77988
rect 434350 77932 434418 77988
rect 434474 77932 434544 77988
rect 434224 77864 434544 77932
rect 434224 77808 434294 77864
rect 434350 77808 434418 77864
rect 434474 77808 434544 77864
rect 434224 77678 434544 77808
rect 444224 78608 444544 81752
rect 449224 80008 449544 81752
rect 449224 79952 449294 80008
rect 449350 79952 449418 80008
rect 449474 79952 449544 80008
rect 449224 79884 449544 79952
rect 449224 79828 449294 79884
rect 449350 79828 449418 79884
rect 449474 79828 449544 79884
rect 449224 79760 449544 79828
rect 449224 79704 449294 79760
rect 449350 79704 449418 79760
rect 449474 79704 449544 79760
rect 449224 79636 449544 79704
rect 449224 79580 449294 79636
rect 449350 79580 449418 79636
rect 449474 79580 449544 79636
rect 449224 79512 449544 79580
rect 449224 79456 449294 79512
rect 449350 79456 449418 79512
rect 449474 79456 449544 79512
rect 449224 79388 449544 79456
rect 449224 79332 449294 79388
rect 449350 79332 449418 79388
rect 449474 79332 449544 79388
rect 449224 79264 449544 79332
rect 449224 79208 449294 79264
rect 449350 79208 449418 79264
rect 449474 79208 449544 79264
rect 449224 79078 449544 79208
rect 444224 78552 444294 78608
rect 444350 78552 444418 78608
rect 444474 78552 444544 78608
rect 444224 78484 444544 78552
rect 444224 78428 444294 78484
rect 444350 78428 444418 78484
rect 444474 78428 444544 78484
rect 444224 78360 444544 78428
rect 444224 78304 444294 78360
rect 444350 78304 444418 78360
rect 444474 78304 444544 78360
rect 444224 78236 444544 78304
rect 444224 78180 444294 78236
rect 444350 78180 444418 78236
rect 444474 78180 444544 78236
rect 444224 78112 444544 78180
rect 444224 78056 444294 78112
rect 444350 78056 444418 78112
rect 444474 78056 444544 78112
rect 444224 77988 444544 78056
rect 444224 77932 444294 77988
rect 444350 77932 444418 77988
rect 444474 77932 444544 77988
rect 444224 77864 444544 77932
rect 444224 77808 444294 77864
rect 444350 77808 444418 77864
rect 444474 77808 444544 77864
rect 444224 77678 444544 77808
rect 454224 78608 454544 81752
rect 459224 80008 459544 81752
rect 459224 79952 459294 80008
rect 459350 79952 459418 80008
rect 459474 79952 459544 80008
rect 459224 79884 459544 79952
rect 459224 79828 459294 79884
rect 459350 79828 459418 79884
rect 459474 79828 459544 79884
rect 459224 79760 459544 79828
rect 459224 79704 459294 79760
rect 459350 79704 459418 79760
rect 459474 79704 459544 79760
rect 459224 79636 459544 79704
rect 459224 79580 459294 79636
rect 459350 79580 459418 79636
rect 459474 79580 459544 79636
rect 459224 79512 459544 79580
rect 459224 79456 459294 79512
rect 459350 79456 459418 79512
rect 459474 79456 459544 79512
rect 459224 79388 459544 79456
rect 459224 79332 459294 79388
rect 459350 79332 459418 79388
rect 459474 79332 459544 79388
rect 459224 79264 459544 79332
rect 459224 79208 459294 79264
rect 459350 79208 459418 79264
rect 459474 79208 459544 79264
rect 459224 79078 459544 79208
rect 454224 78552 454294 78608
rect 454350 78552 454418 78608
rect 454474 78552 454544 78608
rect 454224 78484 454544 78552
rect 454224 78428 454294 78484
rect 454350 78428 454418 78484
rect 454474 78428 454544 78484
rect 454224 78360 454544 78428
rect 454224 78304 454294 78360
rect 454350 78304 454418 78360
rect 454474 78304 454544 78360
rect 454224 78236 454544 78304
rect 454224 78180 454294 78236
rect 454350 78180 454418 78236
rect 454474 78180 454544 78236
rect 454224 78112 454544 78180
rect 454224 78056 454294 78112
rect 454350 78056 454418 78112
rect 454474 78056 454544 78112
rect 454224 77988 454544 78056
rect 454224 77932 454294 77988
rect 454350 77932 454418 77988
rect 454474 77932 454544 77988
rect 454224 77864 454544 77932
rect 454224 77808 454294 77864
rect 454350 77808 454418 77864
rect 454474 77808 454544 77864
rect 454224 77678 454544 77808
rect 464224 78608 464544 81752
rect 469224 80008 469544 81752
rect 469224 79952 469294 80008
rect 469350 79952 469418 80008
rect 469474 79952 469544 80008
rect 469224 79884 469544 79952
rect 469224 79828 469294 79884
rect 469350 79828 469418 79884
rect 469474 79828 469544 79884
rect 469224 79760 469544 79828
rect 469224 79704 469294 79760
rect 469350 79704 469418 79760
rect 469474 79704 469544 79760
rect 469224 79636 469544 79704
rect 469224 79580 469294 79636
rect 469350 79580 469418 79636
rect 469474 79580 469544 79636
rect 469224 79512 469544 79580
rect 469224 79456 469294 79512
rect 469350 79456 469418 79512
rect 469474 79456 469544 79512
rect 469224 79388 469544 79456
rect 469224 79332 469294 79388
rect 469350 79332 469418 79388
rect 469474 79332 469544 79388
rect 469224 79264 469544 79332
rect 469224 79208 469294 79264
rect 469350 79208 469418 79264
rect 469474 79208 469544 79264
rect 469224 79078 469544 79208
rect 464224 78552 464294 78608
rect 464350 78552 464418 78608
rect 464474 78552 464544 78608
rect 464224 78484 464544 78552
rect 464224 78428 464294 78484
rect 464350 78428 464418 78484
rect 464474 78428 464544 78484
rect 464224 78360 464544 78428
rect 464224 78304 464294 78360
rect 464350 78304 464418 78360
rect 464474 78304 464544 78360
rect 464224 78236 464544 78304
rect 464224 78180 464294 78236
rect 464350 78180 464418 78236
rect 464474 78180 464544 78236
rect 464224 78112 464544 78180
rect 464224 78056 464294 78112
rect 464350 78056 464418 78112
rect 464474 78056 464544 78112
rect 464224 77988 464544 78056
rect 464224 77932 464294 77988
rect 464350 77932 464418 77988
rect 464474 77932 464544 77988
rect 464224 77864 464544 77932
rect 464224 77808 464294 77864
rect 464350 77808 464418 77864
rect 464474 77808 464544 77864
rect 464224 77678 464544 77808
rect 474224 78608 474544 81752
rect 479224 80008 479544 81752
rect 479224 79952 479294 80008
rect 479350 79952 479418 80008
rect 479474 79952 479544 80008
rect 479224 79884 479544 79952
rect 479224 79828 479294 79884
rect 479350 79828 479418 79884
rect 479474 79828 479544 79884
rect 479224 79760 479544 79828
rect 479224 79704 479294 79760
rect 479350 79704 479418 79760
rect 479474 79704 479544 79760
rect 479224 79636 479544 79704
rect 479224 79580 479294 79636
rect 479350 79580 479418 79636
rect 479474 79580 479544 79636
rect 479224 79512 479544 79580
rect 479224 79456 479294 79512
rect 479350 79456 479418 79512
rect 479474 79456 479544 79512
rect 479224 79388 479544 79456
rect 479224 79332 479294 79388
rect 479350 79332 479418 79388
rect 479474 79332 479544 79388
rect 479224 79264 479544 79332
rect 479224 79208 479294 79264
rect 479350 79208 479418 79264
rect 479474 79208 479544 79264
rect 479224 79078 479544 79208
rect 474224 78552 474294 78608
rect 474350 78552 474418 78608
rect 474474 78552 474544 78608
rect 474224 78484 474544 78552
rect 474224 78428 474294 78484
rect 474350 78428 474418 78484
rect 474474 78428 474544 78484
rect 474224 78360 474544 78428
rect 474224 78304 474294 78360
rect 474350 78304 474418 78360
rect 474474 78304 474544 78360
rect 474224 78236 474544 78304
rect 474224 78180 474294 78236
rect 474350 78180 474418 78236
rect 474474 78180 474544 78236
rect 474224 78112 474544 78180
rect 474224 78056 474294 78112
rect 474350 78056 474418 78112
rect 474474 78056 474544 78112
rect 474224 77988 474544 78056
rect 474224 77932 474294 77988
rect 474350 77932 474418 77988
rect 474474 77932 474544 77988
rect 474224 77864 474544 77932
rect 474224 77808 474294 77864
rect 474350 77808 474418 77864
rect 474474 77808 474544 77864
rect 474224 77678 474544 77808
rect 484224 78608 484544 81752
rect 489224 80008 489544 81752
rect 489224 79952 489294 80008
rect 489350 79952 489418 80008
rect 489474 79952 489544 80008
rect 489224 79884 489544 79952
rect 489224 79828 489294 79884
rect 489350 79828 489418 79884
rect 489474 79828 489544 79884
rect 489224 79760 489544 79828
rect 489224 79704 489294 79760
rect 489350 79704 489418 79760
rect 489474 79704 489544 79760
rect 489224 79636 489544 79704
rect 489224 79580 489294 79636
rect 489350 79580 489418 79636
rect 489474 79580 489544 79636
rect 489224 79512 489544 79580
rect 489224 79456 489294 79512
rect 489350 79456 489418 79512
rect 489474 79456 489544 79512
rect 489224 79388 489544 79456
rect 489224 79332 489294 79388
rect 489350 79332 489418 79388
rect 489474 79332 489544 79388
rect 489224 79264 489544 79332
rect 489224 79208 489294 79264
rect 489350 79208 489418 79264
rect 489474 79208 489544 79264
rect 489224 79078 489544 79208
rect 484224 78552 484294 78608
rect 484350 78552 484418 78608
rect 484474 78552 484544 78608
rect 484224 78484 484544 78552
rect 484224 78428 484294 78484
rect 484350 78428 484418 78484
rect 484474 78428 484544 78484
rect 484224 78360 484544 78428
rect 484224 78304 484294 78360
rect 484350 78304 484418 78360
rect 484474 78304 484544 78360
rect 484224 78236 484544 78304
rect 484224 78180 484294 78236
rect 484350 78180 484418 78236
rect 484474 78180 484544 78236
rect 484224 78112 484544 78180
rect 484224 78056 484294 78112
rect 484350 78056 484418 78112
rect 484474 78056 484544 78112
rect 484224 77988 484544 78056
rect 484224 77932 484294 77988
rect 484350 77932 484418 77988
rect 484474 77932 484544 77988
rect 484224 77864 484544 77932
rect 484224 77808 484294 77864
rect 484350 77808 484418 77864
rect 484474 77808 484544 77864
rect 484224 77678 484544 77808
rect 494224 78608 494544 81752
rect 499224 80008 499544 81752
rect 499224 79952 499294 80008
rect 499350 79952 499418 80008
rect 499474 79952 499544 80008
rect 499224 79884 499544 79952
rect 499224 79828 499294 79884
rect 499350 79828 499418 79884
rect 499474 79828 499544 79884
rect 499224 79760 499544 79828
rect 499224 79704 499294 79760
rect 499350 79704 499418 79760
rect 499474 79704 499544 79760
rect 499224 79636 499544 79704
rect 499224 79580 499294 79636
rect 499350 79580 499418 79636
rect 499474 79580 499544 79636
rect 499224 79512 499544 79580
rect 499224 79456 499294 79512
rect 499350 79456 499418 79512
rect 499474 79456 499544 79512
rect 499224 79388 499544 79456
rect 499224 79332 499294 79388
rect 499350 79332 499418 79388
rect 499474 79332 499544 79388
rect 499224 79264 499544 79332
rect 499224 79208 499294 79264
rect 499350 79208 499418 79264
rect 499474 79208 499544 79264
rect 499224 79078 499544 79208
rect 494224 78552 494294 78608
rect 494350 78552 494418 78608
rect 494474 78552 494544 78608
rect 494224 78484 494544 78552
rect 494224 78428 494294 78484
rect 494350 78428 494418 78484
rect 494474 78428 494544 78484
rect 494224 78360 494544 78428
rect 494224 78304 494294 78360
rect 494350 78304 494418 78360
rect 494474 78304 494544 78360
rect 494224 78236 494544 78304
rect 494224 78180 494294 78236
rect 494350 78180 494418 78236
rect 494474 78180 494544 78236
rect 494224 78112 494544 78180
rect 494224 78056 494294 78112
rect 494350 78056 494418 78112
rect 494474 78056 494544 78112
rect 494224 77988 494544 78056
rect 494224 77932 494294 77988
rect 494350 77932 494418 77988
rect 494474 77932 494544 77988
rect 494224 77864 494544 77932
rect 494224 77808 494294 77864
rect 494350 77808 494418 77864
rect 494474 77808 494544 77864
rect 494224 77678 494544 77808
rect 504224 78608 504544 81752
rect 509224 80008 509544 81752
rect 509224 79952 509294 80008
rect 509350 79952 509418 80008
rect 509474 79952 509544 80008
rect 509224 79884 509544 79952
rect 509224 79828 509294 79884
rect 509350 79828 509418 79884
rect 509474 79828 509544 79884
rect 509224 79760 509544 79828
rect 509224 79704 509294 79760
rect 509350 79704 509418 79760
rect 509474 79704 509544 79760
rect 509224 79636 509544 79704
rect 509224 79580 509294 79636
rect 509350 79580 509418 79636
rect 509474 79580 509544 79636
rect 509224 79512 509544 79580
rect 509224 79456 509294 79512
rect 509350 79456 509418 79512
rect 509474 79456 509544 79512
rect 509224 79388 509544 79456
rect 509224 79332 509294 79388
rect 509350 79332 509418 79388
rect 509474 79332 509544 79388
rect 509224 79264 509544 79332
rect 509224 79208 509294 79264
rect 509350 79208 509418 79264
rect 509474 79208 509544 79264
rect 509224 79078 509544 79208
rect 504224 78552 504294 78608
rect 504350 78552 504418 78608
rect 504474 78552 504544 78608
rect 504224 78484 504544 78552
rect 504224 78428 504294 78484
rect 504350 78428 504418 78484
rect 504474 78428 504544 78484
rect 504224 78360 504544 78428
rect 504224 78304 504294 78360
rect 504350 78304 504418 78360
rect 504474 78304 504544 78360
rect 504224 78236 504544 78304
rect 504224 78180 504294 78236
rect 504350 78180 504418 78236
rect 504474 78180 504544 78236
rect 504224 78112 504544 78180
rect 504224 78056 504294 78112
rect 504350 78056 504418 78112
rect 504474 78056 504544 78112
rect 504224 77988 504544 78056
rect 504224 77932 504294 77988
rect 504350 77932 504418 77988
rect 504474 77932 504544 77988
rect 504224 77864 504544 77932
rect 504224 77808 504294 77864
rect 504350 77808 504418 77864
rect 504474 77808 504544 77864
rect 504224 77678 504544 77808
rect 514224 78608 514544 81752
rect 519224 80008 519544 81752
rect 519224 79952 519294 80008
rect 519350 79952 519418 80008
rect 519474 79952 519544 80008
rect 519224 79884 519544 79952
rect 519224 79828 519294 79884
rect 519350 79828 519418 79884
rect 519474 79828 519544 79884
rect 519224 79760 519544 79828
rect 519224 79704 519294 79760
rect 519350 79704 519418 79760
rect 519474 79704 519544 79760
rect 519224 79636 519544 79704
rect 519224 79580 519294 79636
rect 519350 79580 519418 79636
rect 519474 79580 519544 79636
rect 519224 79512 519544 79580
rect 519224 79456 519294 79512
rect 519350 79456 519418 79512
rect 519474 79456 519544 79512
rect 519224 79388 519544 79456
rect 519224 79332 519294 79388
rect 519350 79332 519418 79388
rect 519474 79332 519544 79388
rect 519224 79264 519544 79332
rect 519224 79208 519294 79264
rect 519350 79208 519418 79264
rect 519474 79208 519544 79264
rect 519224 79078 519544 79208
rect 514224 78552 514294 78608
rect 514350 78552 514418 78608
rect 514474 78552 514544 78608
rect 514224 78484 514544 78552
rect 514224 78428 514294 78484
rect 514350 78428 514418 78484
rect 514474 78428 514544 78484
rect 514224 78360 514544 78428
rect 514224 78304 514294 78360
rect 514350 78304 514418 78360
rect 514474 78304 514544 78360
rect 514224 78236 514544 78304
rect 514224 78180 514294 78236
rect 514350 78180 514418 78236
rect 514474 78180 514544 78236
rect 514224 78112 514544 78180
rect 514224 78056 514294 78112
rect 514350 78056 514418 78112
rect 514474 78056 514544 78112
rect 514224 77988 514544 78056
rect 514224 77932 514294 77988
rect 514350 77932 514418 77988
rect 514474 77932 514544 77988
rect 514224 77864 514544 77932
rect 514224 77808 514294 77864
rect 514350 77808 514418 77864
rect 514474 77808 514544 77864
rect 514224 77678 514544 77808
rect 524224 78608 524544 81752
rect 529224 80008 529544 81752
rect 529224 79952 529294 80008
rect 529350 79952 529418 80008
rect 529474 79952 529544 80008
rect 529224 79884 529544 79952
rect 529224 79828 529294 79884
rect 529350 79828 529418 79884
rect 529474 79828 529544 79884
rect 529224 79760 529544 79828
rect 529224 79704 529294 79760
rect 529350 79704 529418 79760
rect 529474 79704 529544 79760
rect 529224 79636 529544 79704
rect 529224 79580 529294 79636
rect 529350 79580 529418 79636
rect 529474 79580 529544 79636
rect 529224 79512 529544 79580
rect 529224 79456 529294 79512
rect 529350 79456 529418 79512
rect 529474 79456 529544 79512
rect 529224 79388 529544 79456
rect 529224 79332 529294 79388
rect 529350 79332 529418 79388
rect 529474 79332 529544 79388
rect 529224 79264 529544 79332
rect 529224 79208 529294 79264
rect 529350 79208 529418 79264
rect 529474 79208 529544 79264
rect 529224 79078 529544 79208
rect 524224 78552 524294 78608
rect 524350 78552 524418 78608
rect 524474 78552 524544 78608
rect 524224 78484 524544 78552
rect 524224 78428 524294 78484
rect 524350 78428 524418 78484
rect 524474 78428 524544 78484
rect 524224 78360 524544 78428
rect 524224 78304 524294 78360
rect 524350 78304 524418 78360
rect 524474 78304 524544 78360
rect 524224 78236 524544 78304
rect 524224 78180 524294 78236
rect 524350 78180 524418 78236
rect 524474 78180 524544 78236
rect 524224 78112 524544 78180
rect 524224 78056 524294 78112
rect 524350 78056 524418 78112
rect 524474 78056 524544 78112
rect 524224 77988 524544 78056
rect 524224 77932 524294 77988
rect 524350 77932 524418 77988
rect 524474 77932 524544 77988
rect 524224 77864 524544 77932
rect 524224 77808 524294 77864
rect 524350 77808 524418 77864
rect 524474 77808 524544 77864
rect 524224 77678 524544 77808
rect 534224 78608 534544 81752
rect 539224 80008 539544 81752
rect 539224 79952 539294 80008
rect 539350 79952 539418 80008
rect 539474 79952 539544 80008
rect 539224 79884 539544 79952
rect 539224 79828 539294 79884
rect 539350 79828 539418 79884
rect 539474 79828 539544 79884
rect 539224 79760 539544 79828
rect 539224 79704 539294 79760
rect 539350 79704 539418 79760
rect 539474 79704 539544 79760
rect 539224 79636 539544 79704
rect 539224 79580 539294 79636
rect 539350 79580 539418 79636
rect 539474 79580 539544 79636
rect 539224 79512 539544 79580
rect 539224 79456 539294 79512
rect 539350 79456 539418 79512
rect 539474 79456 539544 79512
rect 539224 79388 539544 79456
rect 539224 79332 539294 79388
rect 539350 79332 539418 79388
rect 539474 79332 539544 79388
rect 539224 79264 539544 79332
rect 539224 79208 539294 79264
rect 539350 79208 539418 79264
rect 539474 79208 539544 79264
rect 539224 79078 539544 79208
rect 534224 78552 534294 78608
rect 534350 78552 534418 78608
rect 534474 78552 534544 78608
rect 534224 78484 534544 78552
rect 534224 78428 534294 78484
rect 534350 78428 534418 78484
rect 534474 78428 534544 78484
rect 534224 78360 534544 78428
rect 534224 78304 534294 78360
rect 534350 78304 534418 78360
rect 534474 78304 534544 78360
rect 534224 78236 534544 78304
rect 534224 78180 534294 78236
rect 534350 78180 534418 78236
rect 534474 78180 534544 78236
rect 534224 78112 534544 78180
rect 534224 78056 534294 78112
rect 534350 78056 534418 78112
rect 534474 78056 534544 78112
rect 534224 77988 534544 78056
rect 534224 77932 534294 77988
rect 534350 77932 534418 77988
rect 534474 77932 534544 77988
rect 534224 77864 534544 77932
rect 534224 77808 534294 77864
rect 534350 77808 534418 77864
rect 534474 77808 534544 77864
rect 534224 77678 534544 77808
rect 544224 78608 544544 81752
rect 549224 80008 549544 81752
rect 549224 79952 549294 80008
rect 549350 79952 549418 80008
rect 549474 79952 549544 80008
rect 549224 79884 549544 79952
rect 549224 79828 549294 79884
rect 549350 79828 549418 79884
rect 549474 79828 549544 79884
rect 549224 79760 549544 79828
rect 549224 79704 549294 79760
rect 549350 79704 549418 79760
rect 549474 79704 549544 79760
rect 549224 79636 549544 79704
rect 549224 79580 549294 79636
rect 549350 79580 549418 79636
rect 549474 79580 549544 79636
rect 549224 79512 549544 79580
rect 549224 79456 549294 79512
rect 549350 79456 549418 79512
rect 549474 79456 549544 79512
rect 549224 79388 549544 79456
rect 549224 79332 549294 79388
rect 549350 79332 549418 79388
rect 549474 79332 549544 79388
rect 549224 79264 549544 79332
rect 549224 79208 549294 79264
rect 549350 79208 549418 79264
rect 549474 79208 549544 79264
rect 549224 79078 549544 79208
rect 544224 78552 544294 78608
rect 544350 78552 544418 78608
rect 544474 78552 544544 78608
rect 544224 78484 544544 78552
rect 544224 78428 544294 78484
rect 544350 78428 544418 78484
rect 544474 78428 544544 78484
rect 544224 78360 544544 78428
rect 544224 78304 544294 78360
rect 544350 78304 544418 78360
rect 544474 78304 544544 78360
rect 544224 78236 544544 78304
rect 544224 78180 544294 78236
rect 544350 78180 544418 78236
rect 544474 78180 544544 78236
rect 544224 78112 544544 78180
rect 544224 78056 544294 78112
rect 544350 78056 544418 78112
rect 544474 78056 544544 78112
rect 544224 77988 544544 78056
rect 544224 77932 544294 77988
rect 544350 77932 544418 77988
rect 544474 77932 544544 77988
rect 544224 77864 544544 77932
rect 544224 77808 544294 77864
rect 544350 77808 544418 77864
rect 544474 77808 544544 77864
rect 544224 77678 544544 77808
rect 554224 78608 554544 81752
rect 590840 80008 591840 99192
rect 590840 79952 590970 80008
rect 591026 79952 591094 80008
rect 591150 79952 591218 80008
rect 591274 79952 591342 80008
rect 591398 79952 591466 80008
rect 591522 79952 591590 80008
rect 591646 79952 591714 80008
rect 591770 79952 591840 80008
rect 590840 79884 591840 79952
rect 590840 79828 590970 79884
rect 591026 79828 591094 79884
rect 591150 79828 591218 79884
rect 591274 79828 591342 79884
rect 591398 79828 591466 79884
rect 591522 79828 591590 79884
rect 591646 79828 591714 79884
rect 591770 79828 591840 79884
rect 590840 79760 591840 79828
rect 590840 79704 590970 79760
rect 591026 79704 591094 79760
rect 591150 79704 591218 79760
rect 591274 79704 591342 79760
rect 591398 79704 591466 79760
rect 591522 79704 591590 79760
rect 591646 79704 591714 79760
rect 591770 79704 591840 79760
rect 590840 79636 591840 79704
rect 590840 79580 590970 79636
rect 591026 79580 591094 79636
rect 591150 79580 591218 79636
rect 591274 79580 591342 79636
rect 591398 79580 591466 79636
rect 591522 79580 591590 79636
rect 591646 79580 591714 79636
rect 591770 79580 591840 79636
rect 590840 79512 591840 79580
rect 590840 79456 590970 79512
rect 591026 79456 591094 79512
rect 591150 79456 591218 79512
rect 591274 79456 591342 79512
rect 591398 79456 591466 79512
rect 591522 79456 591590 79512
rect 591646 79456 591714 79512
rect 591770 79456 591840 79512
rect 590840 79388 591840 79456
rect 590840 79332 590970 79388
rect 591026 79332 591094 79388
rect 591150 79332 591218 79388
rect 591274 79332 591342 79388
rect 591398 79332 591466 79388
rect 591522 79332 591590 79388
rect 591646 79332 591714 79388
rect 591770 79332 591840 79388
rect 590840 79264 591840 79332
rect 590840 79208 590970 79264
rect 591026 79208 591094 79264
rect 591150 79208 591218 79264
rect 591274 79208 591342 79264
rect 591398 79208 591466 79264
rect 591522 79208 591590 79264
rect 591646 79208 591714 79264
rect 591770 79208 591840 79264
rect 590840 79078 591840 79208
rect 592240 305726 593240 305856
rect 592240 305670 592310 305726
rect 592366 305670 592434 305726
rect 592490 305670 592558 305726
rect 592614 305670 592682 305726
rect 592738 305670 592806 305726
rect 592862 305670 592930 305726
rect 592986 305670 593054 305726
rect 593110 305670 593240 305726
rect 592240 305602 593240 305670
rect 592240 305546 592310 305602
rect 592366 305546 592434 305602
rect 592490 305546 592558 305602
rect 592614 305546 592682 305602
rect 592738 305546 592806 305602
rect 592862 305546 592930 305602
rect 592986 305546 593054 305602
rect 593110 305546 593240 305602
rect 592240 305478 593240 305546
rect 592240 305422 592310 305478
rect 592366 305422 592434 305478
rect 592490 305422 592558 305478
rect 592614 305422 592682 305478
rect 592738 305422 592806 305478
rect 592862 305422 592930 305478
rect 592986 305422 593054 305478
rect 593110 305422 593240 305478
rect 592240 305354 593240 305422
rect 592240 305298 592310 305354
rect 592366 305298 592434 305354
rect 592490 305298 592558 305354
rect 592614 305298 592682 305354
rect 592738 305298 592806 305354
rect 592862 305298 592930 305354
rect 592986 305298 593054 305354
rect 593110 305298 593240 305354
rect 592240 305230 593240 305298
rect 592240 305174 592310 305230
rect 592366 305174 592434 305230
rect 592490 305174 592558 305230
rect 592614 305174 592682 305230
rect 592738 305174 592806 305230
rect 592862 305174 592930 305230
rect 592986 305174 593054 305230
rect 593110 305174 593240 305230
rect 592240 305106 593240 305174
rect 592240 305050 592310 305106
rect 592366 305050 592434 305106
rect 592490 305050 592558 305106
rect 592614 305050 592682 305106
rect 592738 305050 592806 305106
rect 592862 305050 592930 305106
rect 592986 305050 593054 305106
rect 593110 305050 593240 305106
rect 592240 304982 593240 305050
rect 592240 304926 592310 304982
rect 592366 304926 592434 304982
rect 592490 304926 592558 304982
rect 592614 304926 592682 304982
rect 592738 304926 592806 304982
rect 592862 304926 592930 304982
rect 592986 304926 593054 304982
rect 593110 304926 593240 304982
rect 592240 281972 593240 304926
rect 633195 305786 633515 314284
rect 634790 307186 635110 314284
rect 634790 307130 634860 307186
rect 634916 307130 634984 307186
rect 635040 307130 635110 307186
rect 634790 307062 635110 307130
rect 634790 307006 634860 307062
rect 634916 307006 634984 307062
rect 635040 307006 635110 307062
rect 634790 306938 635110 307006
rect 634790 306882 634860 306938
rect 634916 306882 634984 306938
rect 635040 306882 635110 306938
rect 634790 306814 635110 306882
rect 634790 306758 634860 306814
rect 634916 306758 634984 306814
rect 635040 306758 635110 306814
rect 634790 306690 635110 306758
rect 634790 306634 634860 306690
rect 634916 306634 634984 306690
rect 635040 306634 635110 306690
rect 634790 306566 635110 306634
rect 634790 306510 634860 306566
rect 634916 306510 634984 306566
rect 635040 306510 635110 306566
rect 634790 306442 635110 306510
rect 634790 306386 634860 306442
rect 634916 306386 634984 306442
rect 635040 306386 635110 306442
rect 634790 306256 635110 306386
rect 633195 305730 633265 305786
rect 633321 305730 633389 305786
rect 633445 305730 633515 305786
rect 633195 305662 633515 305730
rect 633195 305606 633265 305662
rect 633321 305606 633389 305662
rect 633445 305606 633515 305662
rect 633195 305538 633515 305606
rect 633195 305482 633265 305538
rect 633321 305482 633389 305538
rect 633445 305482 633515 305538
rect 633195 305414 633515 305482
rect 633195 305358 633265 305414
rect 633321 305358 633389 305414
rect 633445 305358 633515 305414
rect 633195 305290 633515 305358
rect 633195 305234 633265 305290
rect 633321 305234 633389 305290
rect 633445 305234 633515 305290
rect 633195 305166 633515 305234
rect 633195 305110 633265 305166
rect 633321 305110 633389 305166
rect 633445 305110 633515 305166
rect 633195 305042 633515 305110
rect 633195 304986 633265 305042
rect 633321 304986 633389 305042
rect 633445 304986 633515 305042
rect 633195 304856 633515 304986
rect 636385 305786 636705 314284
rect 637980 307186 638300 314284
rect 637980 307130 638050 307186
rect 638106 307130 638174 307186
rect 638230 307130 638300 307186
rect 637980 307062 638300 307130
rect 637980 307006 638050 307062
rect 638106 307006 638174 307062
rect 638230 307006 638300 307062
rect 637980 306938 638300 307006
rect 637980 306882 638050 306938
rect 638106 306882 638174 306938
rect 638230 306882 638300 306938
rect 637980 306814 638300 306882
rect 637980 306758 638050 306814
rect 638106 306758 638174 306814
rect 638230 306758 638300 306814
rect 637980 306690 638300 306758
rect 637980 306634 638050 306690
rect 638106 306634 638174 306690
rect 638230 306634 638300 306690
rect 637980 306566 638300 306634
rect 637980 306510 638050 306566
rect 638106 306510 638174 306566
rect 638230 306510 638300 306566
rect 637980 306442 638300 306510
rect 637980 306386 638050 306442
rect 638106 306386 638174 306442
rect 638230 306386 638300 306442
rect 637980 306256 638300 306386
rect 636385 305730 636455 305786
rect 636511 305730 636579 305786
rect 636635 305730 636705 305786
rect 636385 305662 636705 305730
rect 636385 305606 636455 305662
rect 636511 305606 636579 305662
rect 636635 305606 636705 305662
rect 636385 305538 636705 305606
rect 636385 305482 636455 305538
rect 636511 305482 636579 305538
rect 636635 305482 636705 305538
rect 636385 305414 636705 305482
rect 636385 305358 636455 305414
rect 636511 305358 636579 305414
rect 636635 305358 636705 305414
rect 636385 305290 636705 305358
rect 636385 305234 636455 305290
rect 636511 305234 636579 305290
rect 636635 305234 636705 305290
rect 636385 305166 636705 305234
rect 636385 305110 636455 305166
rect 636511 305110 636579 305166
rect 636635 305110 636705 305166
rect 636385 305042 636705 305110
rect 636385 304986 636455 305042
rect 636511 304986 636579 305042
rect 636635 304986 636705 305042
rect 636385 304856 636705 304986
rect 639575 305786 639895 314284
rect 641170 307186 641490 314284
rect 641170 307130 641240 307186
rect 641296 307130 641364 307186
rect 641420 307130 641490 307186
rect 641170 307062 641490 307130
rect 641170 307006 641240 307062
rect 641296 307006 641364 307062
rect 641420 307006 641490 307062
rect 641170 306938 641490 307006
rect 641170 306882 641240 306938
rect 641296 306882 641364 306938
rect 641420 306882 641490 306938
rect 641170 306814 641490 306882
rect 641170 306758 641240 306814
rect 641296 306758 641364 306814
rect 641420 306758 641490 306814
rect 641170 306690 641490 306758
rect 641170 306634 641240 306690
rect 641296 306634 641364 306690
rect 641420 306634 641490 306690
rect 641170 306566 641490 306634
rect 641170 306510 641240 306566
rect 641296 306510 641364 306566
rect 641420 306510 641490 306566
rect 641170 306442 641490 306510
rect 641170 306386 641240 306442
rect 641296 306386 641364 306442
rect 641420 306386 641490 306442
rect 641170 306256 641490 306386
rect 639575 305730 639645 305786
rect 639701 305730 639769 305786
rect 639825 305730 639895 305786
rect 639575 305662 639895 305730
rect 639575 305606 639645 305662
rect 639701 305606 639769 305662
rect 639825 305606 639895 305662
rect 639575 305538 639895 305606
rect 639575 305482 639645 305538
rect 639701 305482 639769 305538
rect 639825 305482 639895 305538
rect 639575 305414 639895 305482
rect 639575 305358 639645 305414
rect 639701 305358 639769 305414
rect 639825 305358 639895 305414
rect 639575 305290 639895 305358
rect 639575 305234 639645 305290
rect 639701 305234 639769 305290
rect 639825 305234 639895 305290
rect 639575 305166 639895 305234
rect 639575 305110 639645 305166
rect 639701 305110 639769 305166
rect 639825 305110 639895 305166
rect 639575 305042 639895 305110
rect 639575 304986 639645 305042
rect 639701 304986 639769 305042
rect 639825 304986 639895 305042
rect 639575 304856 639895 304986
rect 642765 305786 643085 314284
rect 642765 305730 642835 305786
rect 642891 305730 642959 305786
rect 643015 305730 643085 305786
rect 642765 305662 643085 305730
rect 642765 305606 642835 305662
rect 642891 305606 642959 305662
rect 643015 305606 643085 305662
rect 642765 305538 643085 305606
rect 642765 305482 642835 305538
rect 642891 305482 642959 305538
rect 643015 305482 643085 305538
rect 642765 305414 643085 305482
rect 642765 305358 642835 305414
rect 642891 305358 642959 305414
rect 643015 305358 643085 305414
rect 642765 305290 643085 305358
rect 642765 305234 642835 305290
rect 642891 305234 642959 305290
rect 643015 305234 643085 305290
rect 642765 305166 643085 305234
rect 642765 305110 642835 305166
rect 642891 305110 642959 305166
rect 643015 305110 643085 305166
rect 642765 305042 643085 305110
rect 642765 304986 642835 305042
rect 642891 304986 642959 305042
rect 643015 304986 643085 305042
rect 642765 304856 643085 304986
rect 697922 313434 698922 320378
rect 697922 313378 698044 313434
rect 698100 313378 698344 313434
rect 698400 313378 698644 313434
rect 698700 313378 698922 313434
rect 697922 307186 698922 313378
rect 697922 307130 698052 307186
rect 698108 307130 698176 307186
rect 698232 307130 698300 307186
rect 698356 307130 698424 307186
rect 698480 307130 698548 307186
rect 698604 307130 698672 307186
rect 698728 307130 698796 307186
rect 698852 307130 698922 307186
rect 697922 307062 698922 307130
rect 697922 307006 698052 307062
rect 698108 307006 698176 307062
rect 698232 307006 698300 307062
rect 698356 307006 698424 307062
rect 698480 307006 698548 307062
rect 698604 307006 698672 307062
rect 698728 307006 698796 307062
rect 698852 307006 698922 307062
rect 697922 306938 698922 307006
rect 697922 306882 698052 306938
rect 698108 306882 698176 306938
rect 698232 306882 698300 306938
rect 698356 306882 698424 306938
rect 698480 306882 698548 306938
rect 698604 306882 698672 306938
rect 698728 306882 698796 306938
rect 698852 306882 698922 306938
rect 697922 306814 698922 306882
rect 697922 306758 698052 306814
rect 698108 306758 698176 306814
rect 698232 306758 698300 306814
rect 698356 306758 698424 306814
rect 698480 306758 698548 306814
rect 698604 306758 698672 306814
rect 698728 306758 698796 306814
rect 698852 306758 698922 306814
rect 697922 306690 698922 306758
rect 697922 306634 698052 306690
rect 698108 306634 698176 306690
rect 698232 306634 698300 306690
rect 698356 306634 698424 306690
rect 698480 306634 698548 306690
rect 698604 306634 698672 306690
rect 698728 306634 698796 306690
rect 698852 306634 698922 306690
rect 697922 306566 698922 306634
rect 697922 306510 698052 306566
rect 698108 306510 698176 306566
rect 698232 306510 698300 306566
rect 698356 306510 698424 306566
rect 698480 306510 698548 306566
rect 698604 306510 698672 306566
rect 698728 306510 698796 306566
rect 698852 306510 698922 306566
rect 697922 306442 698922 306510
rect 697922 306386 698052 306442
rect 698108 306386 698176 306442
rect 698232 306386 698300 306442
rect 698356 306386 698424 306442
rect 698480 306386 698548 306442
rect 698604 306386 698672 306442
rect 698728 306386 698796 306442
rect 698852 306386 698922 306442
rect 592240 281916 592370 281972
rect 592426 281916 592494 281972
rect 592550 281916 592618 281972
rect 592674 281916 592742 281972
rect 592798 281916 592866 281972
rect 592922 281916 592990 281972
rect 593046 281916 593114 281972
rect 593170 281916 593240 281972
rect 592240 281848 593240 281916
rect 592240 281792 592370 281848
rect 592426 281792 592494 281848
rect 592550 281792 592618 281848
rect 592674 281792 592742 281848
rect 592798 281792 592866 281848
rect 592922 281792 592990 281848
rect 593046 281792 593114 281848
rect 593170 281792 593240 281848
rect 592240 281724 593240 281792
rect 592240 281668 592370 281724
rect 592426 281668 592494 281724
rect 592550 281668 592618 281724
rect 592674 281668 592742 281724
rect 592798 281668 592866 281724
rect 592922 281668 592990 281724
rect 593046 281668 593114 281724
rect 593170 281668 593240 281724
rect 592240 281600 593240 281668
rect 592240 281544 592370 281600
rect 592426 281544 592494 281600
rect 592550 281544 592618 281600
rect 592674 281544 592742 281600
rect 592798 281544 592866 281600
rect 592922 281544 592990 281600
rect 593046 281544 593114 281600
rect 593170 281544 593240 281600
rect 592240 281476 593240 281544
rect 592240 281420 592370 281476
rect 592426 281420 592494 281476
rect 592550 281420 592618 281476
rect 592674 281420 592742 281476
rect 592798 281420 592866 281476
rect 592922 281420 592990 281476
rect 593046 281420 593114 281476
rect 593170 281420 593240 281476
rect 592240 281352 593240 281420
rect 592240 281296 592370 281352
rect 592426 281296 592494 281352
rect 592550 281296 592618 281352
rect 592674 281296 592742 281352
rect 592798 281296 592866 281352
rect 592922 281296 592990 281352
rect 593046 281296 593114 281352
rect 593170 281296 593240 281352
rect 592240 281228 593240 281296
rect 592240 281172 592370 281228
rect 592426 281172 592494 281228
rect 592550 281172 592618 281228
rect 592674 281172 592742 281228
rect 592798 281172 592866 281228
rect 592922 281172 592990 281228
rect 593046 281172 593114 281228
rect 593170 281172 593240 281228
rect 592240 268372 593240 281172
rect 592240 268316 592370 268372
rect 592426 268316 592494 268372
rect 592550 268316 592618 268372
rect 592674 268316 592742 268372
rect 592798 268316 592866 268372
rect 592922 268316 592990 268372
rect 593046 268316 593114 268372
rect 593170 268316 593240 268372
rect 592240 268248 593240 268316
rect 592240 268192 592370 268248
rect 592426 268192 592494 268248
rect 592550 268192 592618 268248
rect 592674 268192 592742 268248
rect 592798 268192 592866 268248
rect 592922 268192 592990 268248
rect 593046 268192 593114 268248
rect 593170 268192 593240 268248
rect 592240 242372 593240 268192
rect 592240 242316 592370 242372
rect 592426 242316 592494 242372
rect 592550 242316 592618 242372
rect 592674 242316 592742 242372
rect 592798 242316 592866 242372
rect 592922 242316 592990 242372
rect 593046 242316 593114 242372
rect 593170 242316 593240 242372
rect 592240 242248 593240 242316
rect 592240 242192 592370 242248
rect 592426 242192 592494 242248
rect 592550 242192 592618 242248
rect 592674 242192 592742 242248
rect 592798 242192 592866 242248
rect 592922 242192 592990 242248
rect 593046 242192 593114 242248
rect 593170 242192 593240 242248
rect 592240 216372 593240 242192
rect 592240 216316 592370 216372
rect 592426 216316 592494 216372
rect 592550 216316 592618 216372
rect 592674 216316 592742 216372
rect 592798 216316 592866 216372
rect 592922 216316 592990 216372
rect 593046 216316 593114 216372
rect 593170 216316 593240 216372
rect 592240 216248 593240 216316
rect 592240 216192 592370 216248
rect 592426 216192 592494 216248
rect 592550 216192 592618 216248
rect 592674 216192 592742 216248
rect 592798 216192 592866 216248
rect 592922 216192 592990 216248
rect 593046 216192 593114 216248
rect 593170 216192 593240 216248
rect 592240 190372 593240 216192
rect 592240 190316 592370 190372
rect 592426 190316 592494 190372
rect 592550 190316 592618 190372
rect 592674 190316 592742 190372
rect 592798 190316 592866 190372
rect 592922 190316 592990 190372
rect 593046 190316 593114 190372
rect 593170 190316 593240 190372
rect 592240 190248 593240 190316
rect 592240 190192 592370 190248
rect 592426 190192 592494 190248
rect 592550 190192 592618 190248
rect 592674 190192 592742 190248
rect 592798 190192 592866 190248
rect 592922 190192 592990 190248
rect 593046 190192 593114 190248
rect 593170 190192 593240 190248
rect 592240 164372 593240 190192
rect 592240 164316 592370 164372
rect 592426 164316 592494 164372
rect 592550 164316 592618 164372
rect 592674 164316 592742 164372
rect 592798 164316 592866 164372
rect 592922 164316 592990 164372
rect 593046 164316 593114 164372
rect 593170 164316 593240 164372
rect 592240 164248 593240 164316
rect 592240 164192 592370 164248
rect 592426 164192 592494 164248
rect 592550 164192 592618 164248
rect 592674 164192 592742 164248
rect 592798 164192 592866 164248
rect 592922 164192 592990 164248
rect 593046 164192 593114 164248
rect 593170 164192 593240 164248
rect 592240 138372 593240 164192
rect 592240 138316 592370 138372
rect 592426 138316 592494 138372
rect 592550 138316 592618 138372
rect 592674 138316 592742 138372
rect 592798 138316 592866 138372
rect 592922 138316 592990 138372
rect 593046 138316 593114 138372
rect 593170 138316 593240 138372
rect 592240 138248 593240 138316
rect 592240 138192 592370 138248
rect 592426 138192 592494 138248
rect 592550 138192 592618 138248
rect 592674 138192 592742 138248
rect 592798 138192 592866 138248
rect 592922 138192 592990 138248
rect 593046 138192 593114 138248
rect 593170 138192 593240 138248
rect 592240 121691 593240 138192
rect 592240 121635 592359 121691
rect 592415 121635 592659 121691
rect 592715 121635 592959 121691
rect 593015 121635 593240 121691
rect 592240 118583 593240 121635
rect 592240 118527 592359 118583
rect 592415 118527 592659 118583
rect 592715 118527 592959 118583
rect 593015 118527 593240 118583
rect 592240 115475 593240 118527
rect 592240 115419 592359 115475
rect 592415 115419 592659 115475
rect 592715 115419 592959 115475
rect 593015 115419 593240 115475
rect 592240 112372 593240 115419
rect 592240 112316 592370 112372
rect 592426 112316 592494 112372
rect 592550 112316 592618 112372
rect 592674 112316 592742 112372
rect 592798 112316 592866 112372
rect 592922 112316 592990 112372
rect 593046 112316 593114 112372
rect 593170 112316 593240 112372
rect 592240 112248 593240 112316
rect 592240 112192 592370 112248
rect 592426 112192 592494 112248
rect 592550 112192 592618 112248
rect 592674 112192 592742 112248
rect 592798 112192 592866 112248
rect 592922 112192 592990 112248
rect 593046 112192 593114 112248
rect 593170 112192 593240 112248
rect 592240 86372 593240 112192
rect 697922 290008 698922 306386
rect 697922 289952 698060 290008
rect 698116 289952 698360 290008
rect 698416 289952 698660 290008
rect 698716 289952 698922 290008
rect 697922 283925 698922 289952
rect 697922 283869 698044 283925
rect 698100 283869 698344 283925
rect 698400 283869 698644 283925
rect 698700 283869 698922 283925
rect 697922 277434 698922 283869
rect 697922 277378 698044 277434
rect 698100 277378 698344 277434
rect 698400 277378 698644 277434
rect 698700 277378 698922 277434
rect 697922 270434 698922 277378
rect 697922 270378 698044 270434
rect 698100 270378 698344 270434
rect 698400 270378 698644 270434
rect 698700 270378 698922 270434
rect 697922 263434 698922 270378
rect 697922 263378 698044 263434
rect 698100 263378 698344 263434
rect 698400 263378 698644 263434
rect 698700 263378 698922 263434
rect 697922 253289 698922 263378
rect 697922 253233 698044 253289
rect 698100 253233 698344 253289
rect 698400 253233 698644 253289
rect 698700 253233 698922 253289
rect 697922 247008 698922 253233
rect 697922 246952 698060 247008
rect 698116 246952 698360 247008
rect 698416 246952 698660 247008
rect 698716 246952 698922 247008
rect 697922 234434 698922 246952
rect 697922 234378 698044 234434
rect 698100 234378 698344 234434
rect 698400 234378 698644 234434
rect 698700 234378 698922 234434
rect 697922 227434 698922 234378
rect 697922 227378 698044 227434
rect 698100 227378 698344 227434
rect 698400 227378 698644 227434
rect 698700 227378 698922 227434
rect 697922 222653 698922 227378
rect 697922 222597 698044 222653
rect 698100 222597 698344 222653
rect 698400 222597 698644 222653
rect 698700 222597 698922 222653
rect 697922 220434 698922 222597
rect 697922 220378 698044 220434
rect 698100 220378 698344 220434
rect 698400 220378 698644 220434
rect 698700 220378 698922 220434
rect 697922 204008 698922 220378
rect 697922 203952 698060 204008
rect 698116 203952 698360 204008
rect 698416 203952 698660 204008
rect 698716 203952 698922 204008
rect 697922 192017 698922 203952
rect 697922 191961 698044 192017
rect 698100 191961 698344 192017
rect 698400 191961 698644 192017
rect 698700 191961 698922 192017
rect 697922 191434 698922 191961
rect 697922 191378 698044 191434
rect 698100 191378 698344 191434
rect 698400 191378 698644 191434
rect 698700 191378 698922 191434
rect 697922 184434 698922 191378
rect 697922 184378 698044 184434
rect 698100 184378 698344 184434
rect 698400 184378 698644 184434
rect 698700 184378 698922 184434
rect 697922 177434 698922 184378
rect 697922 177378 698044 177434
rect 698100 177378 698344 177434
rect 698400 177378 698644 177434
rect 698700 177378 698922 177434
rect 697922 161381 698922 177378
rect 697922 161325 698044 161381
rect 698100 161325 698344 161381
rect 698400 161325 698644 161381
rect 698700 161325 698922 161381
rect 697922 161008 698922 161325
rect 697922 160952 698060 161008
rect 698116 160952 698360 161008
rect 698416 160952 698660 161008
rect 698716 160952 698922 161008
rect 697922 148434 698922 160952
rect 697922 148378 698044 148434
rect 698100 148378 698344 148434
rect 698400 148378 698644 148434
rect 698700 148378 698922 148434
rect 697922 141434 698922 148378
rect 697922 141378 698044 141434
rect 698100 141378 698344 141434
rect 698400 141378 698644 141434
rect 698700 141378 698922 141434
rect 697922 134418 698922 141378
rect 697922 134362 698044 134418
rect 698100 134362 698344 134418
rect 698400 134362 698644 134418
rect 698700 134362 698922 134418
rect 697922 133003 698922 134362
rect 697922 132947 698044 133003
rect 698100 132947 698344 133003
rect 698400 132947 698644 133003
rect 698700 132947 698922 133003
rect 697922 118008 698922 132947
rect 697922 117952 698060 118008
rect 698116 117952 698360 118008
rect 698416 117952 698660 118008
rect 698716 117952 698922 118008
rect 697922 105434 698922 117952
rect 697922 105378 698044 105434
rect 698100 105378 698344 105434
rect 698400 105378 698644 105434
rect 698700 105378 698922 105434
rect 592240 86316 592370 86372
rect 592426 86316 592494 86372
rect 592550 86316 592618 86372
rect 592674 86316 592742 86372
rect 592798 86316 592866 86372
rect 592922 86316 592990 86372
rect 593046 86316 593114 86372
rect 593170 86316 593240 86372
rect 592240 86248 593240 86316
rect 592240 86192 592370 86248
rect 592426 86192 592494 86248
rect 592550 86192 592618 86248
rect 592674 86192 592742 86248
rect 592798 86192 592866 86248
rect 592922 86192 592990 86248
rect 593046 86192 593114 86248
rect 593170 86192 593240 86248
rect 554224 78552 554294 78608
rect 554350 78552 554418 78608
rect 554474 78552 554544 78608
rect 554224 78484 554544 78552
rect 554224 78428 554294 78484
rect 554350 78428 554418 78484
rect 554474 78428 554544 78484
rect 554224 78360 554544 78428
rect 554224 78304 554294 78360
rect 554350 78304 554418 78360
rect 554474 78304 554544 78360
rect 554224 78236 554544 78304
rect 554224 78180 554294 78236
rect 554350 78180 554418 78236
rect 554474 78180 554544 78236
rect 554224 78112 554544 78180
rect 554224 78056 554294 78112
rect 554350 78056 554418 78112
rect 554474 78056 554544 78112
rect 554224 77988 554544 78056
rect 554224 77932 554294 77988
rect 554350 77932 554418 77988
rect 554474 77932 554544 77988
rect 554224 77864 554544 77932
rect 554224 77808 554294 77864
rect 554350 77808 554418 77864
rect 554474 77808 554544 77864
rect 554224 77678 554544 77808
rect 592240 78608 593240 86192
rect 668002 99509 668802 99579
rect 668002 99453 668060 99509
rect 668116 99453 668184 99509
rect 668240 99453 668308 99509
rect 668364 99453 668432 99509
rect 668488 99453 668556 99509
rect 668612 99453 668680 99509
rect 668736 99453 668802 99509
rect 668002 99385 668802 99453
rect 668002 99329 668060 99385
rect 668116 99329 668184 99385
rect 668240 99329 668308 99385
rect 668364 99329 668432 99385
rect 668488 99329 668556 99385
rect 668612 99329 668680 99385
rect 668736 99329 668802 99385
rect 668002 99261 668802 99329
rect 668002 99205 668060 99261
rect 668116 99205 668184 99261
rect 668240 99205 668308 99261
rect 668364 99205 668432 99261
rect 668488 99205 668556 99261
rect 668612 99205 668680 99261
rect 668736 99205 668802 99261
rect 668002 99137 668802 99205
rect 668002 99081 668060 99137
rect 668116 99081 668184 99137
rect 668240 99081 668308 99137
rect 668364 99081 668432 99137
rect 668488 99081 668556 99137
rect 668612 99081 668680 99137
rect 668736 99081 668802 99137
rect 668002 99013 668802 99081
rect 668002 98957 668060 99013
rect 668116 98957 668184 99013
rect 668240 98957 668308 99013
rect 668364 98957 668432 99013
rect 668488 98957 668556 99013
rect 668612 98957 668680 99013
rect 668736 98957 668802 99013
rect 668002 98889 668802 98957
rect 668002 98833 668060 98889
rect 668116 98833 668184 98889
rect 668240 98833 668308 98889
rect 668364 98833 668432 98889
rect 668488 98833 668556 98889
rect 668612 98833 668680 98889
rect 668736 98833 668802 98889
rect 668002 98765 668802 98833
rect 668002 98709 668060 98765
rect 668116 98709 668184 98765
rect 668240 98709 668308 98765
rect 668364 98709 668432 98765
rect 668488 98709 668556 98765
rect 668612 98709 668680 98765
rect 668736 98709 668802 98765
rect 592240 78552 592370 78608
rect 592426 78552 592494 78608
rect 592550 78552 592618 78608
rect 592674 78552 592742 78608
rect 592798 78552 592866 78608
rect 592922 78552 592990 78608
rect 593046 78552 593114 78608
rect 593170 78552 593240 78608
rect 592240 78484 593240 78552
rect 592240 78428 592370 78484
rect 592426 78428 592494 78484
rect 592550 78428 592618 78484
rect 592674 78428 592742 78484
rect 592798 78428 592866 78484
rect 592922 78428 592990 78484
rect 593046 78428 593114 78484
rect 593170 78428 593240 78484
rect 592240 78360 593240 78428
rect 592240 78304 592370 78360
rect 592426 78304 592494 78360
rect 592550 78304 592618 78360
rect 592674 78304 592742 78360
rect 592798 78304 592866 78360
rect 592922 78304 592990 78360
rect 593046 78304 593114 78360
rect 593170 78304 593240 78360
rect 592240 78236 593240 78304
rect 592240 78180 592370 78236
rect 592426 78180 592494 78236
rect 592550 78180 592618 78236
rect 592674 78180 592742 78236
rect 592798 78180 592866 78236
rect 592922 78180 592990 78236
rect 593046 78180 593114 78236
rect 593170 78180 593240 78236
rect 592240 78112 593240 78180
rect 592240 78056 592370 78112
rect 592426 78056 592494 78112
rect 592550 78056 592618 78112
rect 592674 78056 592742 78112
rect 592798 78056 592866 78112
rect 592922 78056 592990 78112
rect 593046 78056 593114 78112
rect 593170 78056 593240 78112
rect 592240 77988 593240 78056
rect 592240 77932 592370 77988
rect 592426 77932 592494 77988
rect 592550 77932 592618 77988
rect 592674 77932 592742 77988
rect 592798 77932 592866 77988
rect 592922 77932 592990 77988
rect 593046 77932 593114 77988
rect 593170 77932 593240 77988
rect 592240 77864 593240 77932
rect 592240 77808 592370 77864
rect 592426 77808 592494 77864
rect 592550 77808 592618 77864
rect 592674 77808 592742 77864
rect 592798 77808 592866 77864
rect 592922 77808 592990 77864
rect 593046 77808 593114 77864
rect 593170 77808 593240 77864
rect 592240 77678 593240 77808
rect 602272 80008 604172 80078
rect 602272 79952 602330 80008
rect 602386 79952 602454 80008
rect 602510 79952 602578 80008
rect 602634 79952 602702 80008
rect 602758 79952 602826 80008
rect 602882 79952 602950 80008
rect 603006 79952 603074 80008
rect 603130 79952 603198 80008
rect 603254 79952 603322 80008
rect 603378 79952 603446 80008
rect 603502 79952 603570 80008
rect 603626 79952 603694 80008
rect 603750 79952 603818 80008
rect 603874 79952 603942 80008
rect 603998 79952 604066 80008
rect 604122 79952 604172 80008
rect 602272 79884 604172 79952
rect 602272 79828 602330 79884
rect 602386 79828 602454 79884
rect 602510 79828 602578 79884
rect 602634 79828 602702 79884
rect 602758 79828 602826 79884
rect 602882 79828 602950 79884
rect 603006 79828 603074 79884
rect 603130 79828 603198 79884
rect 603254 79828 603322 79884
rect 603378 79828 603446 79884
rect 603502 79828 603570 79884
rect 603626 79828 603694 79884
rect 603750 79828 603818 79884
rect 603874 79828 603942 79884
rect 603998 79828 604066 79884
rect 604122 79828 604172 79884
rect 602272 79760 604172 79828
rect 602272 79704 602330 79760
rect 602386 79704 602454 79760
rect 602510 79704 602578 79760
rect 602634 79704 602702 79760
rect 602758 79704 602826 79760
rect 602882 79704 602950 79760
rect 603006 79704 603074 79760
rect 603130 79704 603198 79760
rect 603254 79704 603322 79760
rect 603378 79704 603446 79760
rect 603502 79704 603570 79760
rect 603626 79704 603694 79760
rect 603750 79704 603818 79760
rect 603874 79704 603942 79760
rect 603998 79704 604066 79760
rect 604122 79704 604172 79760
rect 602272 79636 604172 79704
rect 602272 79580 602330 79636
rect 602386 79580 602454 79636
rect 602510 79580 602578 79636
rect 602634 79580 602702 79636
rect 602758 79580 602826 79636
rect 602882 79580 602950 79636
rect 603006 79580 603074 79636
rect 603130 79580 603198 79636
rect 603254 79580 603322 79636
rect 603378 79580 603446 79636
rect 603502 79580 603570 79636
rect 603626 79580 603694 79636
rect 603750 79580 603818 79636
rect 603874 79580 603942 79636
rect 603998 79580 604066 79636
rect 604122 79580 604172 79636
rect 602272 79512 604172 79580
rect 602272 79456 602330 79512
rect 602386 79456 602454 79512
rect 602510 79456 602578 79512
rect 602634 79456 602702 79512
rect 602758 79456 602826 79512
rect 602882 79456 602950 79512
rect 603006 79456 603074 79512
rect 603130 79456 603198 79512
rect 603254 79456 603322 79512
rect 603378 79456 603446 79512
rect 603502 79456 603570 79512
rect 603626 79456 603694 79512
rect 603750 79456 603818 79512
rect 603874 79456 603942 79512
rect 603998 79456 604066 79512
rect 604122 79456 604172 79512
rect 602272 79388 604172 79456
rect 602272 79332 602330 79388
rect 602386 79332 602454 79388
rect 602510 79332 602578 79388
rect 602634 79332 602702 79388
rect 602758 79332 602826 79388
rect 602882 79332 602950 79388
rect 603006 79332 603074 79388
rect 603130 79332 603198 79388
rect 603254 79332 603322 79388
rect 603378 79332 603446 79388
rect 603502 79332 603570 79388
rect 603626 79332 603694 79388
rect 603750 79332 603818 79388
rect 603874 79332 603942 79388
rect 603998 79332 604066 79388
rect 604122 79332 604172 79388
rect 602272 79264 604172 79332
rect 602272 79208 602330 79264
rect 602386 79208 602454 79264
rect 602510 79208 602578 79264
rect 602634 79208 602702 79264
rect 602758 79208 602826 79264
rect 602882 79208 602950 79264
rect 603006 79208 603074 79264
rect 603130 79208 603198 79264
rect 603254 79208 603322 79264
rect 603378 79208 603446 79264
rect 603502 79208 603570 79264
rect 603626 79208 603694 79264
rect 603750 79208 603818 79264
rect 603874 79208 603942 79264
rect 603998 79208 604066 79264
rect 604122 79208 604172 79264
rect 284828 70074 284866 70130
rect 284922 70074 284990 70130
rect 285046 70074 285114 70130
rect 285170 70074 285238 70130
rect 285294 70074 285362 70130
rect 285418 70074 285486 70130
rect 285542 70074 285610 70130
rect 285666 70074 285734 70130
rect 285790 70074 285858 70130
rect 285914 70074 285982 70130
rect 286038 70074 286106 70130
rect 286162 70074 286230 70130
rect 286286 70074 286354 70130
rect 286410 70074 286478 70130
rect 286534 70074 286602 70130
rect 286658 70074 286728 70130
rect 284828 70000 286728 70074
rect 602272 70130 604172 79208
rect 602272 70074 602342 70130
rect 602398 70074 602466 70130
rect 602522 70074 602590 70130
rect 602646 70074 602714 70130
rect 602770 70074 602838 70130
rect 602894 70074 602962 70130
rect 603018 70074 603086 70130
rect 603142 70074 603210 70130
rect 603266 70074 603334 70130
rect 603390 70074 603458 70130
rect 603514 70074 603582 70130
rect 603638 70074 603706 70130
rect 603762 70074 603830 70130
rect 603886 70074 603954 70130
rect 604010 70074 604078 70130
rect 604134 70074 604172 70130
rect 602272 70000 604172 70074
rect 604752 80008 606802 80078
rect 604752 79952 604810 80008
rect 604866 79952 604934 80008
rect 604990 79952 605058 80008
rect 605114 79952 605182 80008
rect 605238 79952 605306 80008
rect 605362 79952 605430 80008
rect 605486 79952 605554 80008
rect 605610 79952 605678 80008
rect 605734 79952 605802 80008
rect 605858 79952 605926 80008
rect 605982 79952 606050 80008
rect 606106 79952 606174 80008
rect 606230 79952 606298 80008
rect 606354 79952 606422 80008
rect 606478 79952 606546 80008
rect 606602 79952 606670 80008
rect 606726 79952 606802 80008
rect 604752 79884 606802 79952
rect 604752 79828 604810 79884
rect 604866 79828 604934 79884
rect 604990 79828 605058 79884
rect 605114 79828 605182 79884
rect 605238 79828 605306 79884
rect 605362 79828 605430 79884
rect 605486 79828 605554 79884
rect 605610 79828 605678 79884
rect 605734 79828 605802 79884
rect 605858 79828 605926 79884
rect 605982 79828 606050 79884
rect 606106 79828 606174 79884
rect 606230 79828 606298 79884
rect 606354 79828 606422 79884
rect 606478 79828 606546 79884
rect 606602 79828 606670 79884
rect 606726 79828 606802 79884
rect 604752 79760 606802 79828
rect 604752 79704 604810 79760
rect 604866 79704 604934 79760
rect 604990 79704 605058 79760
rect 605114 79704 605182 79760
rect 605238 79704 605306 79760
rect 605362 79704 605430 79760
rect 605486 79704 605554 79760
rect 605610 79704 605678 79760
rect 605734 79704 605802 79760
rect 605858 79704 605926 79760
rect 605982 79704 606050 79760
rect 606106 79704 606174 79760
rect 606230 79704 606298 79760
rect 606354 79704 606422 79760
rect 606478 79704 606546 79760
rect 606602 79704 606670 79760
rect 606726 79704 606802 79760
rect 604752 79636 606802 79704
rect 604752 79580 604810 79636
rect 604866 79580 604934 79636
rect 604990 79580 605058 79636
rect 605114 79580 605182 79636
rect 605238 79580 605306 79636
rect 605362 79580 605430 79636
rect 605486 79580 605554 79636
rect 605610 79580 605678 79636
rect 605734 79580 605802 79636
rect 605858 79580 605926 79636
rect 605982 79580 606050 79636
rect 606106 79580 606174 79636
rect 606230 79580 606298 79636
rect 606354 79580 606422 79636
rect 606478 79580 606546 79636
rect 606602 79580 606670 79636
rect 606726 79580 606802 79636
rect 604752 79512 606802 79580
rect 604752 79456 604810 79512
rect 604866 79456 604934 79512
rect 604990 79456 605058 79512
rect 605114 79456 605182 79512
rect 605238 79456 605306 79512
rect 605362 79456 605430 79512
rect 605486 79456 605554 79512
rect 605610 79456 605678 79512
rect 605734 79456 605802 79512
rect 605858 79456 605926 79512
rect 605982 79456 606050 79512
rect 606106 79456 606174 79512
rect 606230 79456 606298 79512
rect 606354 79456 606422 79512
rect 606478 79456 606546 79512
rect 606602 79456 606670 79512
rect 606726 79456 606802 79512
rect 604752 79388 606802 79456
rect 604752 79332 604810 79388
rect 604866 79332 604934 79388
rect 604990 79332 605058 79388
rect 605114 79332 605182 79388
rect 605238 79332 605306 79388
rect 605362 79332 605430 79388
rect 605486 79332 605554 79388
rect 605610 79332 605678 79388
rect 605734 79332 605802 79388
rect 605858 79332 605926 79388
rect 605982 79332 606050 79388
rect 606106 79332 606174 79388
rect 606230 79332 606298 79388
rect 606354 79332 606422 79388
rect 606478 79332 606546 79388
rect 606602 79332 606670 79388
rect 606726 79332 606802 79388
rect 604752 79264 606802 79332
rect 604752 79208 604810 79264
rect 604866 79208 604934 79264
rect 604990 79208 605058 79264
rect 605114 79208 605182 79264
rect 605238 79208 605306 79264
rect 605362 79208 605430 79264
rect 605486 79208 605554 79264
rect 605610 79208 605678 79264
rect 605734 79208 605802 79264
rect 605858 79208 605926 79264
rect 605982 79208 606050 79264
rect 606106 79208 606174 79264
rect 606230 79208 606298 79264
rect 606354 79208 606422 79264
rect 606478 79208 606546 79264
rect 606602 79208 606670 79264
rect 606726 79208 606802 79264
rect 604752 70130 606802 79208
rect 604752 70074 604822 70130
rect 604878 70074 604946 70130
rect 605002 70074 605070 70130
rect 605126 70074 605194 70130
rect 605250 70074 605318 70130
rect 605374 70074 605442 70130
rect 605498 70074 605566 70130
rect 605622 70074 605690 70130
rect 605746 70074 605814 70130
rect 605870 70074 605938 70130
rect 605994 70074 606062 70130
rect 606118 70074 606186 70130
rect 606242 70074 606310 70130
rect 606366 70074 606434 70130
rect 606490 70074 606558 70130
rect 606614 70074 606682 70130
rect 606738 70074 606802 70130
rect 604752 70000 606802 70074
rect 607122 80008 609172 80078
rect 607122 79952 607180 80008
rect 607236 79952 607304 80008
rect 607360 79952 607428 80008
rect 607484 79952 607552 80008
rect 607608 79952 607676 80008
rect 607732 79952 607800 80008
rect 607856 79952 607924 80008
rect 607980 79952 608048 80008
rect 608104 79952 608172 80008
rect 608228 79952 608296 80008
rect 608352 79952 608420 80008
rect 608476 79952 608544 80008
rect 608600 79952 608668 80008
rect 608724 79952 608792 80008
rect 608848 79952 608916 80008
rect 608972 79952 609040 80008
rect 609096 79952 609172 80008
rect 607122 79884 609172 79952
rect 607122 79828 607180 79884
rect 607236 79828 607304 79884
rect 607360 79828 607428 79884
rect 607484 79828 607552 79884
rect 607608 79828 607676 79884
rect 607732 79828 607800 79884
rect 607856 79828 607924 79884
rect 607980 79828 608048 79884
rect 608104 79828 608172 79884
rect 608228 79828 608296 79884
rect 608352 79828 608420 79884
rect 608476 79828 608544 79884
rect 608600 79828 608668 79884
rect 608724 79828 608792 79884
rect 608848 79828 608916 79884
rect 608972 79828 609040 79884
rect 609096 79828 609172 79884
rect 607122 79760 609172 79828
rect 607122 79704 607180 79760
rect 607236 79704 607304 79760
rect 607360 79704 607428 79760
rect 607484 79704 607552 79760
rect 607608 79704 607676 79760
rect 607732 79704 607800 79760
rect 607856 79704 607924 79760
rect 607980 79704 608048 79760
rect 608104 79704 608172 79760
rect 608228 79704 608296 79760
rect 608352 79704 608420 79760
rect 608476 79704 608544 79760
rect 608600 79704 608668 79760
rect 608724 79704 608792 79760
rect 608848 79704 608916 79760
rect 608972 79704 609040 79760
rect 609096 79704 609172 79760
rect 607122 79636 609172 79704
rect 607122 79580 607180 79636
rect 607236 79580 607304 79636
rect 607360 79580 607428 79636
rect 607484 79580 607552 79636
rect 607608 79580 607676 79636
rect 607732 79580 607800 79636
rect 607856 79580 607924 79636
rect 607980 79580 608048 79636
rect 608104 79580 608172 79636
rect 608228 79580 608296 79636
rect 608352 79580 608420 79636
rect 608476 79580 608544 79636
rect 608600 79580 608668 79636
rect 608724 79580 608792 79636
rect 608848 79580 608916 79636
rect 608972 79580 609040 79636
rect 609096 79580 609172 79636
rect 607122 79512 609172 79580
rect 607122 79456 607180 79512
rect 607236 79456 607304 79512
rect 607360 79456 607428 79512
rect 607484 79456 607552 79512
rect 607608 79456 607676 79512
rect 607732 79456 607800 79512
rect 607856 79456 607924 79512
rect 607980 79456 608048 79512
rect 608104 79456 608172 79512
rect 608228 79456 608296 79512
rect 608352 79456 608420 79512
rect 608476 79456 608544 79512
rect 608600 79456 608668 79512
rect 608724 79456 608792 79512
rect 608848 79456 608916 79512
rect 608972 79456 609040 79512
rect 609096 79456 609172 79512
rect 607122 79388 609172 79456
rect 607122 79332 607180 79388
rect 607236 79332 607304 79388
rect 607360 79332 607428 79388
rect 607484 79332 607552 79388
rect 607608 79332 607676 79388
rect 607732 79332 607800 79388
rect 607856 79332 607924 79388
rect 607980 79332 608048 79388
rect 608104 79332 608172 79388
rect 608228 79332 608296 79388
rect 608352 79332 608420 79388
rect 608476 79332 608544 79388
rect 608600 79332 608668 79388
rect 608724 79332 608792 79388
rect 608848 79332 608916 79388
rect 608972 79332 609040 79388
rect 609096 79332 609172 79388
rect 607122 79264 609172 79332
rect 607122 79208 607180 79264
rect 607236 79208 607304 79264
rect 607360 79208 607428 79264
rect 607484 79208 607552 79264
rect 607608 79208 607676 79264
rect 607732 79208 607800 79264
rect 607856 79208 607924 79264
rect 607980 79208 608048 79264
rect 608104 79208 608172 79264
rect 608228 79208 608296 79264
rect 608352 79208 608420 79264
rect 608476 79208 608544 79264
rect 608600 79208 608668 79264
rect 608724 79208 608792 79264
rect 608848 79208 608916 79264
rect 608972 79208 609040 79264
rect 609096 79208 609172 79264
rect 607122 70130 609172 79208
rect 607122 70074 607192 70130
rect 607248 70074 607316 70130
rect 607372 70074 607440 70130
rect 607496 70074 607564 70130
rect 607620 70074 607688 70130
rect 607744 70074 607812 70130
rect 607868 70074 607936 70130
rect 607992 70074 608060 70130
rect 608116 70074 608184 70130
rect 608240 70074 608308 70130
rect 608364 70074 608432 70130
rect 608488 70074 608556 70130
rect 608612 70074 608680 70130
rect 608736 70074 608804 70130
rect 608860 70074 608928 70130
rect 608984 70074 609052 70130
rect 609108 70074 609172 70130
rect 607122 70000 609172 70074
rect 609828 80008 611878 80078
rect 609828 79952 609886 80008
rect 609942 79952 610010 80008
rect 610066 79952 610134 80008
rect 610190 79952 610258 80008
rect 610314 79952 610382 80008
rect 610438 79952 610506 80008
rect 610562 79952 610630 80008
rect 610686 79952 610754 80008
rect 610810 79952 610878 80008
rect 610934 79952 611002 80008
rect 611058 79952 611126 80008
rect 611182 79952 611250 80008
rect 611306 79952 611374 80008
rect 611430 79952 611498 80008
rect 611554 79952 611622 80008
rect 611678 79952 611746 80008
rect 611802 79952 611878 80008
rect 609828 79884 611878 79952
rect 609828 79828 609886 79884
rect 609942 79828 610010 79884
rect 610066 79828 610134 79884
rect 610190 79828 610258 79884
rect 610314 79828 610382 79884
rect 610438 79828 610506 79884
rect 610562 79828 610630 79884
rect 610686 79828 610754 79884
rect 610810 79828 610878 79884
rect 610934 79828 611002 79884
rect 611058 79828 611126 79884
rect 611182 79828 611250 79884
rect 611306 79828 611374 79884
rect 611430 79828 611498 79884
rect 611554 79828 611622 79884
rect 611678 79828 611746 79884
rect 611802 79828 611878 79884
rect 609828 79760 611878 79828
rect 609828 79704 609886 79760
rect 609942 79704 610010 79760
rect 610066 79704 610134 79760
rect 610190 79704 610258 79760
rect 610314 79704 610382 79760
rect 610438 79704 610506 79760
rect 610562 79704 610630 79760
rect 610686 79704 610754 79760
rect 610810 79704 610878 79760
rect 610934 79704 611002 79760
rect 611058 79704 611126 79760
rect 611182 79704 611250 79760
rect 611306 79704 611374 79760
rect 611430 79704 611498 79760
rect 611554 79704 611622 79760
rect 611678 79704 611746 79760
rect 611802 79704 611878 79760
rect 609828 79636 611878 79704
rect 609828 79580 609886 79636
rect 609942 79580 610010 79636
rect 610066 79580 610134 79636
rect 610190 79580 610258 79636
rect 610314 79580 610382 79636
rect 610438 79580 610506 79636
rect 610562 79580 610630 79636
rect 610686 79580 610754 79636
rect 610810 79580 610878 79636
rect 610934 79580 611002 79636
rect 611058 79580 611126 79636
rect 611182 79580 611250 79636
rect 611306 79580 611374 79636
rect 611430 79580 611498 79636
rect 611554 79580 611622 79636
rect 611678 79580 611746 79636
rect 611802 79580 611878 79636
rect 609828 79512 611878 79580
rect 609828 79456 609886 79512
rect 609942 79456 610010 79512
rect 610066 79456 610134 79512
rect 610190 79456 610258 79512
rect 610314 79456 610382 79512
rect 610438 79456 610506 79512
rect 610562 79456 610630 79512
rect 610686 79456 610754 79512
rect 610810 79456 610878 79512
rect 610934 79456 611002 79512
rect 611058 79456 611126 79512
rect 611182 79456 611250 79512
rect 611306 79456 611374 79512
rect 611430 79456 611498 79512
rect 611554 79456 611622 79512
rect 611678 79456 611746 79512
rect 611802 79456 611878 79512
rect 609828 79388 611878 79456
rect 609828 79332 609886 79388
rect 609942 79332 610010 79388
rect 610066 79332 610134 79388
rect 610190 79332 610258 79388
rect 610314 79332 610382 79388
rect 610438 79332 610506 79388
rect 610562 79332 610630 79388
rect 610686 79332 610754 79388
rect 610810 79332 610878 79388
rect 610934 79332 611002 79388
rect 611058 79332 611126 79388
rect 611182 79332 611250 79388
rect 611306 79332 611374 79388
rect 611430 79332 611498 79388
rect 611554 79332 611622 79388
rect 611678 79332 611746 79388
rect 611802 79332 611878 79388
rect 609828 79264 611878 79332
rect 609828 79208 609886 79264
rect 609942 79208 610010 79264
rect 610066 79208 610134 79264
rect 610190 79208 610258 79264
rect 610314 79208 610382 79264
rect 610438 79208 610506 79264
rect 610562 79208 610630 79264
rect 610686 79208 610754 79264
rect 610810 79208 610878 79264
rect 610934 79208 611002 79264
rect 611058 79208 611126 79264
rect 611182 79208 611250 79264
rect 611306 79208 611374 79264
rect 611430 79208 611498 79264
rect 611554 79208 611622 79264
rect 611678 79208 611746 79264
rect 611802 79208 611878 79264
rect 609828 70130 611878 79208
rect 609828 70074 609892 70130
rect 609948 70074 610016 70130
rect 610072 70074 610140 70130
rect 610196 70074 610264 70130
rect 610320 70074 610388 70130
rect 610444 70074 610512 70130
rect 610568 70074 610636 70130
rect 610692 70074 610760 70130
rect 610816 70074 610884 70130
rect 610940 70074 611008 70130
rect 611064 70074 611132 70130
rect 611188 70074 611256 70130
rect 611312 70074 611380 70130
rect 611436 70074 611504 70130
rect 611560 70074 611628 70130
rect 611684 70074 611752 70130
rect 611808 70074 611878 70130
rect 609828 70000 611878 70074
rect 612198 80008 614248 80078
rect 612198 79952 612256 80008
rect 612312 79952 612380 80008
rect 612436 79952 612504 80008
rect 612560 79952 612628 80008
rect 612684 79952 612752 80008
rect 612808 79952 612876 80008
rect 612932 79952 613000 80008
rect 613056 79952 613124 80008
rect 613180 79952 613248 80008
rect 613304 79952 613372 80008
rect 613428 79952 613496 80008
rect 613552 79952 613620 80008
rect 613676 79952 613744 80008
rect 613800 79952 613868 80008
rect 613924 79952 613992 80008
rect 614048 79952 614116 80008
rect 614172 79952 614248 80008
rect 612198 79884 614248 79952
rect 612198 79828 612256 79884
rect 612312 79828 612380 79884
rect 612436 79828 612504 79884
rect 612560 79828 612628 79884
rect 612684 79828 612752 79884
rect 612808 79828 612876 79884
rect 612932 79828 613000 79884
rect 613056 79828 613124 79884
rect 613180 79828 613248 79884
rect 613304 79828 613372 79884
rect 613428 79828 613496 79884
rect 613552 79828 613620 79884
rect 613676 79828 613744 79884
rect 613800 79828 613868 79884
rect 613924 79828 613992 79884
rect 614048 79828 614116 79884
rect 614172 79828 614248 79884
rect 612198 79760 614248 79828
rect 612198 79704 612256 79760
rect 612312 79704 612380 79760
rect 612436 79704 612504 79760
rect 612560 79704 612628 79760
rect 612684 79704 612752 79760
rect 612808 79704 612876 79760
rect 612932 79704 613000 79760
rect 613056 79704 613124 79760
rect 613180 79704 613248 79760
rect 613304 79704 613372 79760
rect 613428 79704 613496 79760
rect 613552 79704 613620 79760
rect 613676 79704 613744 79760
rect 613800 79704 613868 79760
rect 613924 79704 613992 79760
rect 614048 79704 614116 79760
rect 614172 79704 614248 79760
rect 612198 79636 614248 79704
rect 612198 79580 612256 79636
rect 612312 79580 612380 79636
rect 612436 79580 612504 79636
rect 612560 79580 612628 79636
rect 612684 79580 612752 79636
rect 612808 79580 612876 79636
rect 612932 79580 613000 79636
rect 613056 79580 613124 79636
rect 613180 79580 613248 79636
rect 613304 79580 613372 79636
rect 613428 79580 613496 79636
rect 613552 79580 613620 79636
rect 613676 79580 613744 79636
rect 613800 79580 613868 79636
rect 613924 79580 613992 79636
rect 614048 79580 614116 79636
rect 614172 79580 614248 79636
rect 612198 79512 614248 79580
rect 612198 79456 612256 79512
rect 612312 79456 612380 79512
rect 612436 79456 612504 79512
rect 612560 79456 612628 79512
rect 612684 79456 612752 79512
rect 612808 79456 612876 79512
rect 612932 79456 613000 79512
rect 613056 79456 613124 79512
rect 613180 79456 613248 79512
rect 613304 79456 613372 79512
rect 613428 79456 613496 79512
rect 613552 79456 613620 79512
rect 613676 79456 613744 79512
rect 613800 79456 613868 79512
rect 613924 79456 613992 79512
rect 614048 79456 614116 79512
rect 614172 79456 614248 79512
rect 612198 79388 614248 79456
rect 612198 79332 612256 79388
rect 612312 79332 612380 79388
rect 612436 79332 612504 79388
rect 612560 79332 612628 79388
rect 612684 79332 612752 79388
rect 612808 79332 612876 79388
rect 612932 79332 613000 79388
rect 613056 79332 613124 79388
rect 613180 79332 613248 79388
rect 613304 79332 613372 79388
rect 613428 79332 613496 79388
rect 613552 79332 613620 79388
rect 613676 79332 613744 79388
rect 613800 79332 613868 79388
rect 613924 79332 613992 79388
rect 614048 79332 614116 79388
rect 614172 79332 614248 79388
rect 612198 79264 614248 79332
rect 612198 79208 612256 79264
rect 612312 79208 612380 79264
rect 612436 79208 612504 79264
rect 612560 79208 612628 79264
rect 612684 79208 612752 79264
rect 612808 79208 612876 79264
rect 612932 79208 613000 79264
rect 613056 79208 613124 79264
rect 613180 79208 613248 79264
rect 613304 79208 613372 79264
rect 613428 79208 613496 79264
rect 613552 79208 613620 79264
rect 613676 79208 613744 79264
rect 613800 79208 613868 79264
rect 613924 79208 613992 79264
rect 614048 79208 614116 79264
rect 614172 79208 614248 79264
rect 612198 70130 614248 79208
rect 612198 70074 612262 70130
rect 612318 70074 612386 70130
rect 612442 70074 612510 70130
rect 612566 70074 612634 70130
rect 612690 70074 612758 70130
rect 612814 70074 612882 70130
rect 612938 70074 613006 70130
rect 613062 70074 613130 70130
rect 613186 70074 613254 70130
rect 613310 70074 613378 70130
rect 613434 70074 613502 70130
rect 613558 70074 613626 70130
rect 613682 70074 613750 70130
rect 613806 70074 613874 70130
rect 613930 70074 613998 70130
rect 614054 70074 614122 70130
rect 614178 70074 614248 70130
rect 612198 70000 614248 70074
rect 614828 80008 616728 80078
rect 614828 79952 614860 80008
rect 614916 79952 614984 80008
rect 615040 79952 615108 80008
rect 615164 79952 615232 80008
rect 615288 79952 615356 80008
rect 615412 79952 615480 80008
rect 615536 79952 615604 80008
rect 615660 79952 615728 80008
rect 615784 79952 615852 80008
rect 615908 79952 615976 80008
rect 616032 79952 616100 80008
rect 616156 79952 616224 80008
rect 616280 79952 616348 80008
rect 616404 79952 616472 80008
rect 616528 79952 616596 80008
rect 616652 79952 616728 80008
rect 614828 79884 616728 79952
rect 614828 79828 614860 79884
rect 614916 79828 614984 79884
rect 615040 79828 615108 79884
rect 615164 79828 615232 79884
rect 615288 79828 615356 79884
rect 615412 79828 615480 79884
rect 615536 79828 615604 79884
rect 615660 79828 615728 79884
rect 615784 79828 615852 79884
rect 615908 79828 615976 79884
rect 616032 79828 616100 79884
rect 616156 79828 616224 79884
rect 616280 79828 616348 79884
rect 616404 79828 616472 79884
rect 616528 79828 616596 79884
rect 616652 79828 616728 79884
rect 614828 79760 616728 79828
rect 614828 79704 614860 79760
rect 614916 79704 614984 79760
rect 615040 79704 615108 79760
rect 615164 79704 615232 79760
rect 615288 79704 615356 79760
rect 615412 79704 615480 79760
rect 615536 79704 615604 79760
rect 615660 79704 615728 79760
rect 615784 79704 615852 79760
rect 615908 79704 615976 79760
rect 616032 79704 616100 79760
rect 616156 79704 616224 79760
rect 616280 79704 616348 79760
rect 616404 79704 616472 79760
rect 616528 79704 616596 79760
rect 616652 79704 616728 79760
rect 614828 79636 616728 79704
rect 614828 79580 614860 79636
rect 614916 79580 614984 79636
rect 615040 79580 615108 79636
rect 615164 79580 615232 79636
rect 615288 79580 615356 79636
rect 615412 79580 615480 79636
rect 615536 79580 615604 79636
rect 615660 79580 615728 79636
rect 615784 79580 615852 79636
rect 615908 79580 615976 79636
rect 616032 79580 616100 79636
rect 616156 79580 616224 79636
rect 616280 79580 616348 79636
rect 616404 79580 616472 79636
rect 616528 79580 616596 79636
rect 616652 79580 616728 79636
rect 614828 79512 616728 79580
rect 614828 79456 614860 79512
rect 614916 79456 614984 79512
rect 615040 79456 615108 79512
rect 615164 79456 615232 79512
rect 615288 79456 615356 79512
rect 615412 79456 615480 79512
rect 615536 79456 615604 79512
rect 615660 79456 615728 79512
rect 615784 79456 615852 79512
rect 615908 79456 615976 79512
rect 616032 79456 616100 79512
rect 616156 79456 616224 79512
rect 616280 79456 616348 79512
rect 616404 79456 616472 79512
rect 616528 79456 616596 79512
rect 616652 79456 616728 79512
rect 614828 79388 616728 79456
rect 614828 79332 614860 79388
rect 614916 79332 614984 79388
rect 615040 79332 615108 79388
rect 615164 79332 615232 79388
rect 615288 79332 615356 79388
rect 615412 79332 615480 79388
rect 615536 79332 615604 79388
rect 615660 79332 615728 79388
rect 615784 79332 615852 79388
rect 615908 79332 615976 79388
rect 616032 79332 616100 79388
rect 616156 79332 616224 79388
rect 616280 79332 616348 79388
rect 616404 79332 616472 79388
rect 616528 79332 616596 79388
rect 616652 79332 616728 79388
rect 614828 79264 616728 79332
rect 614828 79208 614860 79264
rect 614916 79208 614984 79264
rect 615040 79208 615108 79264
rect 615164 79208 615232 79264
rect 615288 79208 615356 79264
rect 615412 79208 615480 79264
rect 615536 79208 615604 79264
rect 615660 79208 615728 79264
rect 615784 79208 615852 79264
rect 615908 79208 615976 79264
rect 616032 79208 616100 79264
rect 616156 79208 616224 79264
rect 616280 79208 616348 79264
rect 616404 79208 616472 79264
rect 616528 79208 616596 79264
rect 616652 79208 616728 79264
rect 614828 70130 616728 79208
rect 624657 78608 624977 84750
rect 628627 80008 628947 84750
rect 628627 79952 628697 80008
rect 628753 79952 628821 80008
rect 628877 79952 628947 80008
rect 628627 79884 628947 79952
rect 628627 79828 628697 79884
rect 628753 79828 628821 79884
rect 628877 79828 628947 79884
rect 628627 79760 628947 79828
rect 628627 79704 628697 79760
rect 628753 79704 628821 79760
rect 628877 79704 628947 79760
rect 628627 79636 628947 79704
rect 628627 79580 628697 79636
rect 628753 79580 628821 79636
rect 628877 79580 628947 79636
rect 628627 79512 628947 79580
rect 628627 79456 628697 79512
rect 628753 79456 628821 79512
rect 628877 79456 628947 79512
rect 628627 79388 628947 79456
rect 628627 79332 628697 79388
rect 628753 79332 628821 79388
rect 628877 79332 628947 79388
rect 628627 79264 628947 79332
rect 628627 79208 628697 79264
rect 628753 79208 628821 79264
rect 628877 79208 628947 79264
rect 628627 79078 628947 79208
rect 624657 78552 624727 78608
rect 624783 78552 624851 78608
rect 624907 78552 624977 78608
rect 624657 78484 624977 78552
rect 624657 78428 624727 78484
rect 624783 78428 624851 78484
rect 624907 78428 624977 78484
rect 624657 78360 624977 78428
rect 624657 78304 624727 78360
rect 624783 78304 624851 78360
rect 624907 78304 624977 78360
rect 624657 78236 624977 78304
rect 624657 78180 624727 78236
rect 624783 78180 624851 78236
rect 624907 78180 624977 78236
rect 624657 78112 624977 78180
rect 624657 78056 624727 78112
rect 624783 78056 624851 78112
rect 624907 78056 624977 78112
rect 624657 77988 624977 78056
rect 624657 77932 624727 77988
rect 624783 77932 624851 77988
rect 624907 77932 624977 77988
rect 624657 77864 624977 77932
rect 624657 77808 624727 77864
rect 624783 77808 624851 77864
rect 624907 77808 624977 77864
rect 624657 77678 624977 77808
rect 632597 78608 632917 84750
rect 636567 80008 636887 84750
rect 636567 79952 636637 80008
rect 636693 79952 636761 80008
rect 636817 79952 636887 80008
rect 636567 79884 636887 79952
rect 636567 79828 636637 79884
rect 636693 79828 636761 79884
rect 636817 79828 636887 79884
rect 636567 79760 636887 79828
rect 636567 79704 636637 79760
rect 636693 79704 636761 79760
rect 636817 79704 636887 79760
rect 636567 79636 636887 79704
rect 636567 79580 636637 79636
rect 636693 79580 636761 79636
rect 636817 79580 636887 79636
rect 636567 79512 636887 79580
rect 636567 79456 636637 79512
rect 636693 79456 636761 79512
rect 636817 79456 636887 79512
rect 636567 79388 636887 79456
rect 636567 79332 636637 79388
rect 636693 79332 636761 79388
rect 636817 79332 636887 79388
rect 636567 79264 636887 79332
rect 636567 79208 636637 79264
rect 636693 79208 636761 79264
rect 636817 79208 636887 79264
rect 636567 79078 636887 79208
rect 632597 78552 632667 78608
rect 632723 78552 632791 78608
rect 632847 78552 632917 78608
rect 632597 78484 632917 78552
rect 632597 78428 632667 78484
rect 632723 78428 632791 78484
rect 632847 78428 632917 78484
rect 632597 78360 632917 78428
rect 632597 78304 632667 78360
rect 632723 78304 632791 78360
rect 632847 78304 632917 78360
rect 632597 78236 632917 78304
rect 632597 78180 632667 78236
rect 632723 78180 632791 78236
rect 632847 78180 632917 78236
rect 632597 78112 632917 78180
rect 632597 78056 632667 78112
rect 632723 78056 632791 78112
rect 632847 78056 632917 78112
rect 632597 77988 632917 78056
rect 632597 77932 632667 77988
rect 632723 77932 632791 77988
rect 632847 77932 632917 77988
rect 632597 77864 632917 77932
rect 632597 77808 632667 77864
rect 632723 77808 632791 77864
rect 632847 77808 632917 77864
rect 632597 77678 632917 77808
rect 640537 78608 640857 84750
rect 644507 80008 644827 84750
rect 644507 79952 644577 80008
rect 644633 79952 644701 80008
rect 644757 79952 644827 80008
rect 644507 79884 644827 79952
rect 644507 79828 644577 79884
rect 644633 79828 644701 79884
rect 644757 79828 644827 79884
rect 644507 79760 644827 79828
rect 644507 79704 644577 79760
rect 644633 79704 644701 79760
rect 644757 79704 644827 79760
rect 644507 79636 644827 79704
rect 644507 79580 644577 79636
rect 644633 79580 644701 79636
rect 644757 79580 644827 79636
rect 644507 79512 644827 79580
rect 644507 79456 644577 79512
rect 644633 79456 644701 79512
rect 644757 79456 644827 79512
rect 644507 79388 644827 79456
rect 644507 79332 644577 79388
rect 644633 79332 644701 79388
rect 644757 79332 644827 79388
rect 644507 79264 644827 79332
rect 644507 79208 644577 79264
rect 644633 79208 644701 79264
rect 644757 79208 644827 79264
rect 644507 79078 644827 79208
rect 640537 78552 640607 78608
rect 640663 78552 640731 78608
rect 640787 78552 640857 78608
rect 640537 78484 640857 78552
rect 640537 78428 640607 78484
rect 640663 78428 640731 78484
rect 640787 78428 640857 78484
rect 640537 78360 640857 78428
rect 640537 78304 640607 78360
rect 640663 78304 640731 78360
rect 640787 78304 640857 78360
rect 640537 78236 640857 78304
rect 640537 78180 640607 78236
rect 640663 78180 640731 78236
rect 640787 78180 640857 78236
rect 640537 78112 640857 78180
rect 640537 78056 640607 78112
rect 640663 78056 640731 78112
rect 640787 78056 640857 78112
rect 640537 77988 640857 78056
rect 640537 77932 640607 77988
rect 640663 77932 640731 77988
rect 640787 77932 640857 77988
rect 640537 77864 640857 77932
rect 640537 77808 640607 77864
rect 640663 77808 640731 77864
rect 640787 77808 640857 77864
rect 640537 77678 640857 77808
rect 648477 78608 648797 84750
rect 668002 78678 668802 98709
rect 670032 99509 670832 99579
rect 670032 99453 670090 99509
rect 670146 99453 670214 99509
rect 670270 99453 670338 99509
rect 670394 99453 670462 99509
rect 670518 99453 670586 99509
rect 670642 99453 670710 99509
rect 670766 99453 670832 99509
rect 670032 99385 670832 99453
rect 670032 99329 670090 99385
rect 670146 99329 670214 99385
rect 670270 99329 670338 99385
rect 670394 99329 670462 99385
rect 670518 99329 670586 99385
rect 670642 99329 670710 99385
rect 670766 99329 670832 99385
rect 670032 99261 670832 99329
rect 670032 99205 670090 99261
rect 670146 99205 670214 99261
rect 670270 99205 670338 99261
rect 670394 99205 670462 99261
rect 670518 99205 670586 99261
rect 670642 99205 670710 99261
rect 670766 99205 670832 99261
rect 670032 99137 670832 99205
rect 670032 99081 670090 99137
rect 670146 99081 670214 99137
rect 670270 99081 670338 99137
rect 670394 99081 670462 99137
rect 670518 99081 670586 99137
rect 670642 99081 670710 99137
rect 670766 99081 670832 99137
rect 670032 99013 670832 99081
rect 670032 98957 670090 99013
rect 670146 98957 670214 99013
rect 670270 98957 670338 99013
rect 670394 98957 670462 99013
rect 670518 98957 670586 99013
rect 670642 98957 670710 99013
rect 670766 98957 670832 99013
rect 670032 98889 670832 98957
rect 670032 98833 670090 98889
rect 670146 98833 670214 98889
rect 670270 98833 670338 98889
rect 670394 98833 670462 98889
rect 670518 98833 670586 98889
rect 670642 98833 670710 98889
rect 670766 98833 670832 98889
rect 670032 98765 670832 98833
rect 670032 98709 670090 98765
rect 670146 98709 670214 98765
rect 670270 98709 670338 98765
rect 670394 98709 670462 98765
rect 670518 98709 670586 98765
rect 670642 98709 670710 98765
rect 670766 98709 670832 98765
rect 670032 80008 670832 98709
rect 670032 79952 670090 80008
rect 670146 79952 670214 80008
rect 670270 79952 670338 80008
rect 670394 79952 670462 80008
rect 670518 79952 670586 80008
rect 670642 79952 670710 80008
rect 670766 79952 670832 80008
rect 670032 79884 670832 79952
rect 670032 79828 670090 79884
rect 670146 79828 670214 79884
rect 670270 79828 670338 79884
rect 670394 79828 670462 79884
rect 670518 79828 670586 79884
rect 670642 79828 670710 79884
rect 670766 79828 670832 79884
rect 670032 79760 670832 79828
rect 670032 79704 670090 79760
rect 670146 79704 670214 79760
rect 670270 79704 670338 79760
rect 670394 79704 670462 79760
rect 670518 79704 670586 79760
rect 670642 79704 670710 79760
rect 670766 79704 670832 79760
rect 670032 79636 670832 79704
rect 670032 79580 670090 79636
rect 670146 79580 670214 79636
rect 670270 79580 670338 79636
rect 670394 79580 670462 79636
rect 670518 79580 670586 79636
rect 670642 79580 670710 79636
rect 670766 79580 670832 79636
rect 670032 79512 670832 79580
rect 670032 79456 670090 79512
rect 670146 79456 670214 79512
rect 670270 79456 670338 79512
rect 670394 79456 670462 79512
rect 670518 79456 670586 79512
rect 670642 79456 670710 79512
rect 670766 79456 670832 79512
rect 670032 79388 670832 79456
rect 670032 79332 670090 79388
rect 670146 79332 670214 79388
rect 670270 79332 670338 79388
rect 670394 79332 670462 79388
rect 670518 79332 670586 79388
rect 670642 79332 670710 79388
rect 670766 79332 670832 79388
rect 670032 79264 670832 79332
rect 670032 79208 670090 79264
rect 670146 79208 670214 79264
rect 670270 79208 670338 79264
rect 670394 79208 670462 79264
rect 670518 79208 670586 79264
rect 670642 79208 670710 79264
rect 670766 79208 670832 79264
rect 670032 79078 670832 79208
rect 697922 98434 698922 105378
rect 697922 98378 698044 98434
rect 698100 98378 698344 98434
rect 698400 98378 698644 98434
rect 698700 98378 698922 98434
rect 697922 91434 698922 98378
rect 697922 91378 698044 91434
rect 698100 91378 698344 91434
rect 698400 91378 698644 91434
rect 698700 91378 698922 91434
rect 697922 80008 698922 91378
rect 697922 79952 698052 80008
rect 698108 79952 698176 80008
rect 698232 79952 698300 80008
rect 698356 79952 698424 80008
rect 698480 79952 698548 80008
rect 698604 79952 698672 80008
rect 698728 79952 698796 80008
rect 698852 79952 698922 80008
rect 697922 79884 698922 79952
rect 697922 79828 698052 79884
rect 698108 79828 698176 79884
rect 698232 79828 698300 79884
rect 698356 79828 698424 79884
rect 698480 79828 698548 79884
rect 698604 79828 698672 79884
rect 698728 79828 698796 79884
rect 698852 79828 698922 79884
rect 697922 79760 698922 79828
rect 697922 79704 698052 79760
rect 698108 79704 698176 79760
rect 698232 79704 698300 79760
rect 698356 79704 698424 79760
rect 698480 79704 698548 79760
rect 698604 79704 698672 79760
rect 698728 79704 698796 79760
rect 698852 79704 698922 79760
rect 697922 79636 698922 79704
rect 697922 79580 698052 79636
rect 698108 79580 698176 79636
rect 698232 79580 698300 79636
rect 698356 79580 698424 79636
rect 698480 79580 698548 79636
rect 698604 79580 698672 79636
rect 698728 79580 698796 79636
rect 698852 79580 698922 79636
rect 697922 79512 698922 79580
rect 697922 79456 698052 79512
rect 698108 79456 698176 79512
rect 698232 79456 698300 79512
rect 698356 79456 698424 79512
rect 698480 79456 698548 79512
rect 698604 79456 698672 79512
rect 698728 79456 698796 79512
rect 698852 79456 698922 79512
rect 697922 79388 698922 79456
rect 697922 79332 698052 79388
rect 698108 79332 698176 79388
rect 698232 79332 698300 79388
rect 698356 79332 698424 79388
rect 698480 79332 698548 79388
rect 698604 79332 698672 79388
rect 698728 79332 698796 79388
rect 698852 79332 698922 79388
rect 697922 79264 698922 79332
rect 697922 79208 698052 79264
rect 698108 79208 698176 79264
rect 698232 79208 698300 79264
rect 698356 79208 698424 79264
rect 698480 79208 698548 79264
rect 698604 79208 698672 79264
rect 698728 79208 698796 79264
rect 698852 79208 698922 79264
rect 648477 78552 648547 78608
rect 648603 78552 648671 78608
rect 648727 78552 648797 78608
rect 648477 78484 648797 78552
rect 648477 78428 648547 78484
rect 648603 78428 648671 78484
rect 648727 78428 648797 78484
rect 648477 78360 648797 78428
rect 648477 78304 648547 78360
rect 648603 78304 648671 78360
rect 648727 78304 648797 78360
rect 648477 78236 648797 78304
rect 648477 78180 648547 78236
rect 648603 78180 648671 78236
rect 648727 78180 648797 78236
rect 648477 78112 648797 78180
rect 648477 78056 648547 78112
rect 648603 78056 648671 78112
rect 648727 78056 648797 78112
rect 648477 77988 648797 78056
rect 648477 77932 648547 77988
rect 648603 77932 648671 77988
rect 648727 77932 648797 77988
rect 648477 77864 648797 77932
rect 648477 77808 648547 77864
rect 648603 77808 648671 77864
rect 648727 77808 648797 77864
rect 648477 77678 648797 77808
rect 657272 78608 659172 78678
rect 657272 78552 657330 78608
rect 657386 78552 657454 78608
rect 657510 78552 657578 78608
rect 657634 78552 657702 78608
rect 657758 78552 657826 78608
rect 657882 78552 657950 78608
rect 658006 78552 658074 78608
rect 658130 78552 658198 78608
rect 658254 78552 658322 78608
rect 658378 78552 658446 78608
rect 658502 78552 658570 78608
rect 658626 78552 658694 78608
rect 658750 78552 658818 78608
rect 658874 78552 658942 78608
rect 658998 78552 659066 78608
rect 659122 78552 659172 78608
rect 657272 78484 659172 78552
rect 657272 78428 657330 78484
rect 657386 78428 657454 78484
rect 657510 78428 657578 78484
rect 657634 78428 657702 78484
rect 657758 78428 657826 78484
rect 657882 78428 657950 78484
rect 658006 78428 658074 78484
rect 658130 78428 658198 78484
rect 658254 78428 658322 78484
rect 658378 78428 658446 78484
rect 658502 78428 658570 78484
rect 658626 78428 658694 78484
rect 658750 78428 658818 78484
rect 658874 78428 658942 78484
rect 658998 78428 659066 78484
rect 659122 78428 659172 78484
rect 657272 78360 659172 78428
rect 657272 78304 657330 78360
rect 657386 78304 657454 78360
rect 657510 78304 657578 78360
rect 657634 78304 657702 78360
rect 657758 78304 657826 78360
rect 657882 78304 657950 78360
rect 658006 78304 658074 78360
rect 658130 78304 658198 78360
rect 658254 78304 658322 78360
rect 658378 78304 658446 78360
rect 658502 78304 658570 78360
rect 658626 78304 658694 78360
rect 658750 78304 658818 78360
rect 658874 78304 658942 78360
rect 658998 78304 659066 78360
rect 659122 78304 659172 78360
rect 657272 78236 659172 78304
rect 657272 78180 657330 78236
rect 657386 78180 657454 78236
rect 657510 78180 657578 78236
rect 657634 78180 657702 78236
rect 657758 78180 657826 78236
rect 657882 78180 657950 78236
rect 658006 78180 658074 78236
rect 658130 78180 658198 78236
rect 658254 78180 658322 78236
rect 658378 78180 658446 78236
rect 658502 78180 658570 78236
rect 658626 78180 658694 78236
rect 658750 78180 658818 78236
rect 658874 78180 658942 78236
rect 658998 78180 659066 78236
rect 659122 78180 659172 78236
rect 657272 78112 659172 78180
rect 657272 78056 657330 78112
rect 657386 78056 657454 78112
rect 657510 78056 657578 78112
rect 657634 78056 657702 78112
rect 657758 78056 657826 78112
rect 657882 78056 657950 78112
rect 658006 78056 658074 78112
rect 658130 78056 658198 78112
rect 658254 78056 658322 78112
rect 658378 78056 658446 78112
rect 658502 78056 658570 78112
rect 658626 78056 658694 78112
rect 658750 78056 658818 78112
rect 658874 78056 658942 78112
rect 658998 78056 659066 78112
rect 659122 78056 659172 78112
rect 657272 77988 659172 78056
rect 657272 77932 657330 77988
rect 657386 77932 657454 77988
rect 657510 77932 657578 77988
rect 657634 77932 657702 77988
rect 657758 77932 657826 77988
rect 657882 77932 657950 77988
rect 658006 77932 658074 77988
rect 658130 77932 658198 77988
rect 658254 77932 658322 77988
rect 658378 77932 658446 77988
rect 658502 77932 658570 77988
rect 658626 77932 658694 77988
rect 658750 77932 658818 77988
rect 658874 77932 658942 77988
rect 658998 77932 659066 77988
rect 659122 77932 659172 77988
rect 657272 77864 659172 77932
rect 657272 77808 657330 77864
rect 657386 77808 657454 77864
rect 657510 77808 657578 77864
rect 657634 77808 657702 77864
rect 657758 77808 657826 77864
rect 657882 77808 657950 77864
rect 658006 77808 658074 77864
rect 658130 77808 658198 77864
rect 658254 77808 658322 77864
rect 658378 77808 658446 77864
rect 658502 77808 658570 77864
rect 658626 77808 658694 77864
rect 658750 77808 658818 77864
rect 658874 77808 658942 77864
rect 658998 77808 659066 77864
rect 659122 77808 659172 77864
rect 614828 70074 614866 70130
rect 614922 70074 614990 70130
rect 615046 70074 615114 70130
rect 615170 70074 615238 70130
rect 615294 70074 615362 70130
rect 615418 70074 615486 70130
rect 615542 70074 615610 70130
rect 615666 70074 615734 70130
rect 615790 70074 615858 70130
rect 615914 70074 615982 70130
rect 616038 70074 616106 70130
rect 616162 70074 616230 70130
rect 616286 70074 616354 70130
rect 616410 70074 616478 70130
rect 616534 70074 616602 70130
rect 616658 70074 616728 70130
rect 614828 70000 616728 70074
rect 657272 70130 659172 77808
rect 657272 70074 657342 70130
rect 657398 70074 657466 70130
rect 657522 70074 657590 70130
rect 657646 70074 657714 70130
rect 657770 70074 657838 70130
rect 657894 70074 657962 70130
rect 658018 70074 658086 70130
rect 658142 70074 658210 70130
rect 658266 70074 658334 70130
rect 658390 70074 658458 70130
rect 658514 70074 658582 70130
rect 658638 70074 658706 70130
rect 658762 70074 658830 70130
rect 658886 70074 658954 70130
rect 659010 70074 659078 70130
rect 659134 70074 659172 70130
rect 657272 70000 659172 70074
rect 659752 78608 661802 78678
rect 659752 78552 659810 78608
rect 659866 78552 659934 78608
rect 659990 78552 660058 78608
rect 660114 78552 660182 78608
rect 660238 78552 660306 78608
rect 660362 78552 660430 78608
rect 660486 78552 660554 78608
rect 660610 78552 660678 78608
rect 660734 78552 660802 78608
rect 660858 78552 660926 78608
rect 660982 78552 661050 78608
rect 661106 78552 661174 78608
rect 661230 78552 661298 78608
rect 661354 78552 661422 78608
rect 661478 78552 661546 78608
rect 661602 78552 661670 78608
rect 661726 78552 661802 78608
rect 659752 78484 661802 78552
rect 659752 78428 659810 78484
rect 659866 78428 659934 78484
rect 659990 78428 660058 78484
rect 660114 78428 660182 78484
rect 660238 78428 660306 78484
rect 660362 78428 660430 78484
rect 660486 78428 660554 78484
rect 660610 78428 660678 78484
rect 660734 78428 660802 78484
rect 660858 78428 660926 78484
rect 660982 78428 661050 78484
rect 661106 78428 661174 78484
rect 661230 78428 661298 78484
rect 661354 78428 661422 78484
rect 661478 78428 661546 78484
rect 661602 78428 661670 78484
rect 661726 78428 661802 78484
rect 659752 78360 661802 78428
rect 659752 78304 659810 78360
rect 659866 78304 659934 78360
rect 659990 78304 660058 78360
rect 660114 78304 660182 78360
rect 660238 78304 660306 78360
rect 660362 78304 660430 78360
rect 660486 78304 660554 78360
rect 660610 78304 660678 78360
rect 660734 78304 660802 78360
rect 660858 78304 660926 78360
rect 660982 78304 661050 78360
rect 661106 78304 661174 78360
rect 661230 78304 661298 78360
rect 661354 78304 661422 78360
rect 661478 78304 661546 78360
rect 661602 78304 661670 78360
rect 661726 78304 661802 78360
rect 659752 78236 661802 78304
rect 659752 78180 659810 78236
rect 659866 78180 659934 78236
rect 659990 78180 660058 78236
rect 660114 78180 660182 78236
rect 660238 78180 660306 78236
rect 660362 78180 660430 78236
rect 660486 78180 660554 78236
rect 660610 78180 660678 78236
rect 660734 78180 660802 78236
rect 660858 78180 660926 78236
rect 660982 78180 661050 78236
rect 661106 78180 661174 78236
rect 661230 78180 661298 78236
rect 661354 78180 661422 78236
rect 661478 78180 661546 78236
rect 661602 78180 661670 78236
rect 661726 78180 661802 78236
rect 659752 78112 661802 78180
rect 659752 78056 659810 78112
rect 659866 78056 659934 78112
rect 659990 78056 660058 78112
rect 660114 78056 660182 78112
rect 660238 78056 660306 78112
rect 660362 78056 660430 78112
rect 660486 78056 660554 78112
rect 660610 78056 660678 78112
rect 660734 78056 660802 78112
rect 660858 78056 660926 78112
rect 660982 78056 661050 78112
rect 661106 78056 661174 78112
rect 661230 78056 661298 78112
rect 661354 78056 661422 78112
rect 661478 78056 661546 78112
rect 661602 78056 661670 78112
rect 661726 78056 661802 78112
rect 659752 77988 661802 78056
rect 659752 77932 659810 77988
rect 659866 77932 659934 77988
rect 659990 77932 660058 77988
rect 660114 77932 660182 77988
rect 660238 77932 660306 77988
rect 660362 77932 660430 77988
rect 660486 77932 660554 77988
rect 660610 77932 660678 77988
rect 660734 77932 660802 77988
rect 660858 77932 660926 77988
rect 660982 77932 661050 77988
rect 661106 77932 661174 77988
rect 661230 77932 661298 77988
rect 661354 77932 661422 77988
rect 661478 77932 661546 77988
rect 661602 77932 661670 77988
rect 661726 77932 661802 77988
rect 659752 77864 661802 77932
rect 659752 77808 659810 77864
rect 659866 77808 659934 77864
rect 659990 77808 660058 77864
rect 660114 77808 660182 77864
rect 660238 77808 660306 77864
rect 660362 77808 660430 77864
rect 660486 77808 660554 77864
rect 660610 77808 660678 77864
rect 660734 77808 660802 77864
rect 660858 77808 660926 77864
rect 660982 77808 661050 77864
rect 661106 77808 661174 77864
rect 661230 77808 661298 77864
rect 661354 77808 661422 77864
rect 661478 77808 661546 77864
rect 661602 77808 661670 77864
rect 661726 77808 661802 77864
rect 659752 70130 661802 77808
rect 659752 70074 659822 70130
rect 659878 70074 659946 70130
rect 660002 70074 660070 70130
rect 660126 70074 660194 70130
rect 660250 70074 660318 70130
rect 660374 70074 660442 70130
rect 660498 70074 660566 70130
rect 660622 70074 660690 70130
rect 660746 70074 660814 70130
rect 660870 70074 660938 70130
rect 660994 70074 661062 70130
rect 661118 70074 661186 70130
rect 661242 70074 661310 70130
rect 661366 70074 661434 70130
rect 661490 70074 661558 70130
rect 661614 70074 661682 70130
rect 661738 70074 661802 70130
rect 659752 70000 661802 70074
rect 662122 78608 664172 78678
rect 662122 78552 662180 78608
rect 662236 78552 662304 78608
rect 662360 78552 662428 78608
rect 662484 78552 662552 78608
rect 662608 78552 662676 78608
rect 662732 78552 662800 78608
rect 662856 78552 662924 78608
rect 662980 78552 663048 78608
rect 663104 78552 663172 78608
rect 663228 78552 663296 78608
rect 663352 78552 663420 78608
rect 663476 78552 663544 78608
rect 663600 78552 663668 78608
rect 663724 78552 663792 78608
rect 663848 78552 663916 78608
rect 663972 78552 664040 78608
rect 664096 78552 664172 78608
rect 662122 78484 664172 78552
rect 662122 78428 662180 78484
rect 662236 78428 662304 78484
rect 662360 78428 662428 78484
rect 662484 78428 662552 78484
rect 662608 78428 662676 78484
rect 662732 78428 662800 78484
rect 662856 78428 662924 78484
rect 662980 78428 663048 78484
rect 663104 78428 663172 78484
rect 663228 78428 663296 78484
rect 663352 78428 663420 78484
rect 663476 78428 663544 78484
rect 663600 78428 663668 78484
rect 663724 78428 663792 78484
rect 663848 78428 663916 78484
rect 663972 78428 664040 78484
rect 664096 78428 664172 78484
rect 662122 78360 664172 78428
rect 662122 78304 662180 78360
rect 662236 78304 662304 78360
rect 662360 78304 662428 78360
rect 662484 78304 662552 78360
rect 662608 78304 662676 78360
rect 662732 78304 662800 78360
rect 662856 78304 662924 78360
rect 662980 78304 663048 78360
rect 663104 78304 663172 78360
rect 663228 78304 663296 78360
rect 663352 78304 663420 78360
rect 663476 78304 663544 78360
rect 663600 78304 663668 78360
rect 663724 78304 663792 78360
rect 663848 78304 663916 78360
rect 663972 78304 664040 78360
rect 664096 78304 664172 78360
rect 662122 78236 664172 78304
rect 662122 78180 662180 78236
rect 662236 78180 662304 78236
rect 662360 78180 662428 78236
rect 662484 78180 662552 78236
rect 662608 78180 662676 78236
rect 662732 78180 662800 78236
rect 662856 78180 662924 78236
rect 662980 78180 663048 78236
rect 663104 78180 663172 78236
rect 663228 78180 663296 78236
rect 663352 78180 663420 78236
rect 663476 78180 663544 78236
rect 663600 78180 663668 78236
rect 663724 78180 663792 78236
rect 663848 78180 663916 78236
rect 663972 78180 664040 78236
rect 664096 78180 664172 78236
rect 662122 78112 664172 78180
rect 662122 78056 662180 78112
rect 662236 78056 662304 78112
rect 662360 78056 662428 78112
rect 662484 78056 662552 78112
rect 662608 78056 662676 78112
rect 662732 78056 662800 78112
rect 662856 78056 662924 78112
rect 662980 78056 663048 78112
rect 663104 78056 663172 78112
rect 663228 78056 663296 78112
rect 663352 78056 663420 78112
rect 663476 78056 663544 78112
rect 663600 78056 663668 78112
rect 663724 78056 663792 78112
rect 663848 78056 663916 78112
rect 663972 78056 664040 78112
rect 664096 78056 664172 78112
rect 662122 77988 664172 78056
rect 662122 77932 662180 77988
rect 662236 77932 662304 77988
rect 662360 77932 662428 77988
rect 662484 77932 662552 77988
rect 662608 77932 662676 77988
rect 662732 77932 662800 77988
rect 662856 77932 662924 77988
rect 662980 77932 663048 77988
rect 663104 77932 663172 77988
rect 663228 77932 663296 77988
rect 663352 77932 663420 77988
rect 663476 77932 663544 77988
rect 663600 77932 663668 77988
rect 663724 77932 663792 77988
rect 663848 77932 663916 77988
rect 663972 77932 664040 77988
rect 664096 77932 664172 77988
rect 662122 77864 664172 77932
rect 662122 77808 662180 77864
rect 662236 77808 662304 77864
rect 662360 77808 662428 77864
rect 662484 77808 662552 77864
rect 662608 77808 662676 77864
rect 662732 77808 662800 77864
rect 662856 77808 662924 77864
rect 662980 77808 663048 77864
rect 663104 77808 663172 77864
rect 663228 77808 663296 77864
rect 663352 77808 663420 77864
rect 663476 77808 663544 77864
rect 663600 77808 663668 77864
rect 663724 77808 663792 77864
rect 663848 77808 663916 77864
rect 663972 77808 664040 77864
rect 664096 77808 664172 77864
rect 662122 70130 664172 77808
rect 662122 70074 662192 70130
rect 662248 70074 662316 70130
rect 662372 70074 662440 70130
rect 662496 70074 662564 70130
rect 662620 70074 662688 70130
rect 662744 70074 662812 70130
rect 662868 70074 662936 70130
rect 662992 70074 663060 70130
rect 663116 70074 663184 70130
rect 663240 70074 663308 70130
rect 663364 70074 663432 70130
rect 663488 70074 663556 70130
rect 663612 70074 663680 70130
rect 663736 70074 663804 70130
rect 663860 70074 663928 70130
rect 663984 70074 664052 70130
rect 664108 70074 664172 70130
rect 662122 70000 664172 70074
rect 664828 78608 666878 78678
rect 664828 78552 664886 78608
rect 664942 78552 665010 78608
rect 665066 78552 665134 78608
rect 665190 78552 665258 78608
rect 665314 78552 665382 78608
rect 665438 78552 665506 78608
rect 665562 78552 665630 78608
rect 665686 78552 665754 78608
rect 665810 78552 665878 78608
rect 665934 78552 666002 78608
rect 666058 78552 666126 78608
rect 666182 78552 666250 78608
rect 666306 78552 666374 78608
rect 666430 78552 666498 78608
rect 666554 78552 666622 78608
rect 666678 78552 666746 78608
rect 666802 78552 666878 78608
rect 664828 78484 666878 78552
rect 664828 78428 664886 78484
rect 664942 78428 665010 78484
rect 665066 78428 665134 78484
rect 665190 78428 665258 78484
rect 665314 78428 665382 78484
rect 665438 78428 665506 78484
rect 665562 78428 665630 78484
rect 665686 78428 665754 78484
rect 665810 78428 665878 78484
rect 665934 78428 666002 78484
rect 666058 78428 666126 78484
rect 666182 78428 666250 78484
rect 666306 78428 666374 78484
rect 666430 78428 666498 78484
rect 666554 78428 666622 78484
rect 666678 78428 666746 78484
rect 666802 78428 666878 78484
rect 664828 78360 666878 78428
rect 664828 78304 664886 78360
rect 664942 78304 665010 78360
rect 665066 78304 665134 78360
rect 665190 78304 665258 78360
rect 665314 78304 665382 78360
rect 665438 78304 665506 78360
rect 665562 78304 665630 78360
rect 665686 78304 665754 78360
rect 665810 78304 665878 78360
rect 665934 78304 666002 78360
rect 666058 78304 666126 78360
rect 666182 78304 666250 78360
rect 666306 78304 666374 78360
rect 666430 78304 666498 78360
rect 666554 78304 666622 78360
rect 666678 78304 666746 78360
rect 666802 78304 666878 78360
rect 664828 78236 666878 78304
rect 664828 78180 664886 78236
rect 664942 78180 665010 78236
rect 665066 78180 665134 78236
rect 665190 78180 665258 78236
rect 665314 78180 665382 78236
rect 665438 78180 665506 78236
rect 665562 78180 665630 78236
rect 665686 78180 665754 78236
rect 665810 78180 665878 78236
rect 665934 78180 666002 78236
rect 666058 78180 666126 78236
rect 666182 78180 666250 78236
rect 666306 78180 666374 78236
rect 666430 78180 666498 78236
rect 666554 78180 666622 78236
rect 666678 78180 666746 78236
rect 666802 78180 666878 78236
rect 664828 78112 666878 78180
rect 664828 78056 664886 78112
rect 664942 78056 665010 78112
rect 665066 78056 665134 78112
rect 665190 78056 665258 78112
rect 665314 78056 665382 78112
rect 665438 78056 665506 78112
rect 665562 78056 665630 78112
rect 665686 78056 665754 78112
rect 665810 78056 665878 78112
rect 665934 78056 666002 78112
rect 666058 78056 666126 78112
rect 666182 78056 666250 78112
rect 666306 78056 666374 78112
rect 666430 78056 666498 78112
rect 666554 78056 666622 78112
rect 666678 78056 666746 78112
rect 666802 78056 666878 78112
rect 664828 77988 666878 78056
rect 664828 77932 664886 77988
rect 664942 77932 665010 77988
rect 665066 77932 665134 77988
rect 665190 77932 665258 77988
rect 665314 77932 665382 77988
rect 665438 77932 665506 77988
rect 665562 77932 665630 77988
rect 665686 77932 665754 77988
rect 665810 77932 665878 77988
rect 665934 77932 666002 77988
rect 666058 77932 666126 77988
rect 666182 77932 666250 77988
rect 666306 77932 666374 77988
rect 666430 77932 666498 77988
rect 666554 77932 666622 77988
rect 666678 77932 666746 77988
rect 666802 77932 666878 77988
rect 664828 77864 666878 77932
rect 664828 77808 664886 77864
rect 664942 77808 665010 77864
rect 665066 77808 665134 77864
rect 665190 77808 665258 77864
rect 665314 77808 665382 77864
rect 665438 77808 665506 77864
rect 665562 77808 665630 77864
rect 665686 77808 665754 77864
rect 665810 77808 665878 77864
rect 665934 77808 666002 77864
rect 666058 77808 666126 77864
rect 666182 77808 666250 77864
rect 666306 77808 666374 77864
rect 666430 77808 666498 77864
rect 666554 77808 666622 77864
rect 666678 77808 666746 77864
rect 666802 77808 666878 77864
rect 664828 70130 666878 77808
rect 664828 70074 664892 70130
rect 664948 70074 665016 70130
rect 665072 70074 665140 70130
rect 665196 70074 665264 70130
rect 665320 70074 665388 70130
rect 665444 70074 665512 70130
rect 665568 70074 665636 70130
rect 665692 70074 665760 70130
rect 665816 70074 665884 70130
rect 665940 70074 666008 70130
rect 666064 70074 666132 70130
rect 666188 70074 666256 70130
rect 666312 70074 666380 70130
rect 666436 70074 666504 70130
rect 666560 70074 666628 70130
rect 666684 70074 666752 70130
rect 666808 70074 666878 70130
rect 664828 70000 666878 70074
rect 667198 78608 669248 78678
rect 667198 78552 667256 78608
rect 667312 78552 667380 78608
rect 667436 78552 667504 78608
rect 667560 78552 667628 78608
rect 667684 78552 667752 78608
rect 667808 78552 667876 78608
rect 667932 78552 668000 78608
rect 668056 78552 668124 78608
rect 668180 78552 668248 78608
rect 668304 78552 668372 78608
rect 668428 78552 668496 78608
rect 668552 78552 668620 78608
rect 668676 78552 668744 78608
rect 668800 78552 668868 78608
rect 668924 78552 668992 78608
rect 669048 78552 669116 78608
rect 669172 78552 669248 78608
rect 667198 78484 669248 78552
rect 667198 78428 667256 78484
rect 667312 78428 667380 78484
rect 667436 78428 667504 78484
rect 667560 78428 667628 78484
rect 667684 78428 667752 78484
rect 667808 78428 667876 78484
rect 667932 78428 668000 78484
rect 668056 78428 668124 78484
rect 668180 78428 668248 78484
rect 668304 78428 668372 78484
rect 668428 78428 668496 78484
rect 668552 78428 668620 78484
rect 668676 78428 668744 78484
rect 668800 78428 668868 78484
rect 668924 78428 668992 78484
rect 669048 78428 669116 78484
rect 669172 78428 669248 78484
rect 667198 78360 669248 78428
rect 667198 78304 667256 78360
rect 667312 78304 667380 78360
rect 667436 78304 667504 78360
rect 667560 78304 667628 78360
rect 667684 78304 667752 78360
rect 667808 78304 667876 78360
rect 667932 78304 668000 78360
rect 668056 78304 668124 78360
rect 668180 78304 668248 78360
rect 668304 78304 668372 78360
rect 668428 78304 668496 78360
rect 668552 78304 668620 78360
rect 668676 78304 668744 78360
rect 668800 78304 668868 78360
rect 668924 78304 668992 78360
rect 669048 78304 669116 78360
rect 669172 78304 669248 78360
rect 667198 78236 669248 78304
rect 667198 78180 667256 78236
rect 667312 78180 667380 78236
rect 667436 78180 667504 78236
rect 667560 78180 667628 78236
rect 667684 78180 667752 78236
rect 667808 78180 667876 78236
rect 667932 78180 668000 78236
rect 668056 78180 668124 78236
rect 668180 78180 668248 78236
rect 668304 78180 668372 78236
rect 668428 78180 668496 78236
rect 668552 78180 668620 78236
rect 668676 78180 668744 78236
rect 668800 78180 668868 78236
rect 668924 78180 668992 78236
rect 669048 78180 669116 78236
rect 669172 78180 669248 78236
rect 667198 78112 669248 78180
rect 667198 78056 667256 78112
rect 667312 78056 667380 78112
rect 667436 78056 667504 78112
rect 667560 78056 667628 78112
rect 667684 78056 667752 78112
rect 667808 78056 667876 78112
rect 667932 78056 668000 78112
rect 668056 78056 668124 78112
rect 668180 78056 668248 78112
rect 668304 78056 668372 78112
rect 668428 78056 668496 78112
rect 668552 78056 668620 78112
rect 668676 78056 668744 78112
rect 668800 78056 668868 78112
rect 668924 78056 668992 78112
rect 669048 78056 669116 78112
rect 669172 78056 669248 78112
rect 667198 77988 669248 78056
rect 667198 77932 667256 77988
rect 667312 77932 667380 77988
rect 667436 77932 667504 77988
rect 667560 77932 667628 77988
rect 667684 77932 667752 77988
rect 667808 77932 667876 77988
rect 667932 77932 668000 77988
rect 668056 77932 668124 77988
rect 668180 77932 668248 77988
rect 668304 77932 668372 77988
rect 668428 77932 668496 77988
rect 668552 77932 668620 77988
rect 668676 77932 668744 77988
rect 668800 77932 668868 77988
rect 668924 77932 668992 77988
rect 669048 77932 669116 77988
rect 669172 77932 669248 77988
rect 667198 77864 669248 77932
rect 667198 77808 667256 77864
rect 667312 77808 667380 77864
rect 667436 77808 667504 77864
rect 667560 77808 667628 77864
rect 667684 77808 667752 77864
rect 667808 77808 667876 77864
rect 667932 77808 668000 77864
rect 668056 77808 668124 77864
rect 668180 77808 668248 77864
rect 668304 77808 668372 77864
rect 668428 77808 668496 77864
rect 668552 77808 668620 77864
rect 668676 77808 668744 77864
rect 668800 77808 668868 77864
rect 668924 77808 668992 77864
rect 669048 77808 669116 77864
rect 669172 77808 669248 77864
rect 667198 70130 669248 77808
rect 667198 70074 667262 70130
rect 667318 70074 667386 70130
rect 667442 70074 667510 70130
rect 667566 70074 667634 70130
rect 667690 70074 667758 70130
rect 667814 70074 667882 70130
rect 667938 70074 668006 70130
rect 668062 70074 668130 70130
rect 668186 70074 668254 70130
rect 668310 70074 668378 70130
rect 668434 70074 668502 70130
rect 668558 70074 668626 70130
rect 668682 70074 668750 70130
rect 668806 70074 668874 70130
rect 668930 70074 668998 70130
rect 669054 70074 669122 70130
rect 669178 70074 669248 70130
rect 667198 70000 669248 70074
rect 669828 78608 671728 78678
rect 669828 78552 669860 78608
rect 669916 78552 669984 78608
rect 670040 78552 670108 78608
rect 670164 78552 670232 78608
rect 670288 78552 670356 78608
rect 670412 78552 670480 78608
rect 670536 78552 670604 78608
rect 670660 78552 670728 78608
rect 670784 78552 670852 78608
rect 670908 78552 670976 78608
rect 671032 78552 671100 78608
rect 671156 78552 671224 78608
rect 671280 78552 671348 78608
rect 671404 78552 671472 78608
rect 671528 78552 671596 78608
rect 671652 78552 671728 78608
rect 669828 78484 671728 78552
rect 669828 78428 669860 78484
rect 669916 78428 669984 78484
rect 670040 78428 670108 78484
rect 670164 78428 670232 78484
rect 670288 78428 670356 78484
rect 670412 78428 670480 78484
rect 670536 78428 670604 78484
rect 670660 78428 670728 78484
rect 670784 78428 670852 78484
rect 670908 78428 670976 78484
rect 671032 78428 671100 78484
rect 671156 78428 671224 78484
rect 671280 78428 671348 78484
rect 671404 78428 671472 78484
rect 671528 78428 671596 78484
rect 671652 78428 671728 78484
rect 669828 78360 671728 78428
rect 669828 78304 669860 78360
rect 669916 78304 669984 78360
rect 670040 78304 670108 78360
rect 670164 78304 670232 78360
rect 670288 78304 670356 78360
rect 670412 78304 670480 78360
rect 670536 78304 670604 78360
rect 670660 78304 670728 78360
rect 670784 78304 670852 78360
rect 670908 78304 670976 78360
rect 671032 78304 671100 78360
rect 671156 78304 671224 78360
rect 671280 78304 671348 78360
rect 671404 78304 671472 78360
rect 671528 78304 671596 78360
rect 671652 78304 671728 78360
rect 669828 78236 671728 78304
rect 669828 78180 669860 78236
rect 669916 78180 669984 78236
rect 670040 78180 670108 78236
rect 670164 78180 670232 78236
rect 670288 78180 670356 78236
rect 670412 78180 670480 78236
rect 670536 78180 670604 78236
rect 670660 78180 670728 78236
rect 670784 78180 670852 78236
rect 670908 78180 670976 78236
rect 671032 78180 671100 78236
rect 671156 78180 671224 78236
rect 671280 78180 671348 78236
rect 671404 78180 671472 78236
rect 671528 78180 671596 78236
rect 671652 78180 671728 78236
rect 669828 78112 671728 78180
rect 669828 78056 669860 78112
rect 669916 78056 669984 78112
rect 670040 78056 670108 78112
rect 670164 78056 670232 78112
rect 670288 78056 670356 78112
rect 670412 78056 670480 78112
rect 670536 78056 670604 78112
rect 670660 78056 670728 78112
rect 670784 78056 670852 78112
rect 670908 78056 670976 78112
rect 671032 78056 671100 78112
rect 671156 78056 671224 78112
rect 671280 78056 671348 78112
rect 671404 78056 671472 78112
rect 671528 78056 671596 78112
rect 671652 78056 671728 78112
rect 669828 77988 671728 78056
rect 669828 77932 669860 77988
rect 669916 77932 669984 77988
rect 670040 77932 670108 77988
rect 670164 77932 670232 77988
rect 670288 77932 670356 77988
rect 670412 77932 670480 77988
rect 670536 77932 670604 77988
rect 670660 77932 670728 77988
rect 670784 77932 670852 77988
rect 670908 77932 670976 77988
rect 671032 77932 671100 77988
rect 671156 77932 671224 77988
rect 671280 77932 671348 77988
rect 671404 77932 671472 77988
rect 671528 77932 671596 77988
rect 671652 77932 671728 77988
rect 669828 77864 671728 77932
rect 669828 77808 669860 77864
rect 669916 77808 669984 77864
rect 670040 77808 670108 77864
rect 670164 77808 670232 77864
rect 670288 77808 670356 77864
rect 670412 77808 670480 77864
rect 670536 77808 670604 77864
rect 670660 77808 670728 77864
rect 670784 77808 670852 77864
rect 670908 77808 670976 77864
rect 671032 77808 671100 77864
rect 671156 77808 671224 77864
rect 671280 77808 671348 77864
rect 671404 77808 671472 77864
rect 671528 77808 671596 77864
rect 671652 77808 671728 77864
rect 669828 70130 671728 77808
rect 697922 75008 698922 79208
rect 699322 925954 700322 941392
rect 699322 925898 699444 925954
rect 699500 925898 699744 925954
rect 699800 925898 700044 925954
rect 700100 925898 700322 925954
rect 699322 918954 700322 925898
rect 699322 918898 699444 918954
rect 699500 918898 699744 918954
rect 699800 918898 700044 918954
rect 700100 918898 700322 918954
rect 699322 914429 700322 918898
rect 699322 914373 699544 914429
rect 699600 914373 699844 914429
rect 699900 914373 700144 914429
rect 700200 914373 700322 914429
rect 699322 914229 700322 914373
rect 699322 914173 699544 914229
rect 699600 914173 699844 914229
rect 699900 914173 700144 914229
rect 700200 914173 700322 914229
rect 699322 911954 700322 914173
rect 699322 911898 699444 911954
rect 699500 911898 699744 911954
rect 699800 911898 700044 911954
rect 700100 911898 700322 911954
rect 699322 892423 700322 911898
rect 699322 892367 699497 892423
rect 699553 892367 699797 892423
rect 699853 892367 700097 892423
rect 700153 892367 700322 892423
rect 699322 883652 700322 892367
rect 699322 883596 699392 883652
rect 699448 883596 699516 883652
rect 699572 883596 699640 883652
rect 699696 883596 699764 883652
rect 699820 883596 699888 883652
rect 699944 883596 700012 883652
rect 700068 883596 700136 883652
rect 700192 883596 700322 883652
rect 699322 883528 700322 883596
rect 699322 883472 699392 883528
rect 699448 883472 699516 883528
rect 699572 883472 699640 883528
rect 699696 883472 699764 883528
rect 699820 883472 699888 883528
rect 699944 883472 700012 883528
rect 700068 883472 700136 883528
rect 700192 883472 700322 883528
rect 699322 883404 700322 883472
rect 699322 883348 699392 883404
rect 699448 883348 699516 883404
rect 699572 883348 699640 883404
rect 699696 883348 699764 883404
rect 699820 883348 699888 883404
rect 699944 883348 700012 883404
rect 700068 883348 700136 883404
rect 700192 883348 700322 883404
rect 699322 883280 700322 883348
rect 699322 883224 699392 883280
rect 699448 883224 699516 883280
rect 699572 883224 699640 883280
rect 699696 883224 699764 883280
rect 699820 883224 699888 883280
rect 699944 883224 700012 883280
rect 700068 883224 700136 883280
rect 700192 883224 700322 883280
rect 699322 883156 700322 883224
rect 699322 883100 699392 883156
rect 699448 883100 699516 883156
rect 699572 883100 699640 883156
rect 699696 883100 699764 883156
rect 699820 883100 699888 883156
rect 699944 883100 700012 883156
rect 700068 883100 700136 883156
rect 700192 883100 700322 883156
rect 699322 883032 700322 883100
rect 699322 882976 699392 883032
rect 699448 882976 699516 883032
rect 699572 882976 699640 883032
rect 699696 882976 699764 883032
rect 699820 882976 699888 883032
rect 699944 882976 700012 883032
rect 700068 882976 700136 883032
rect 700192 882976 700322 883032
rect 699322 882908 700322 882976
rect 699322 882852 699392 882908
rect 699448 882852 699516 882908
rect 699572 882852 699640 882908
rect 699696 882852 699764 882908
rect 699820 882852 699888 882908
rect 699944 882852 700012 882908
rect 700068 882852 700136 882908
rect 700192 882852 700322 882908
rect 699322 882784 700322 882852
rect 699322 882728 699392 882784
rect 699448 882728 699516 882784
rect 699572 882728 699640 882784
rect 699696 882728 699764 882784
rect 699820 882728 699888 882784
rect 699944 882728 700012 882784
rect 700068 882728 700136 882784
rect 700192 882728 700322 882784
rect 699322 882660 700322 882728
rect 699322 882604 699392 882660
rect 699448 882604 699516 882660
rect 699572 882604 699640 882660
rect 699696 882604 699764 882660
rect 699820 882604 699888 882660
rect 699944 882604 700012 882660
rect 700068 882604 700136 882660
rect 700192 882604 700322 882660
rect 699322 882536 700322 882604
rect 699322 882480 699392 882536
rect 699448 882480 699516 882536
rect 699572 882480 699640 882536
rect 699696 882480 699764 882536
rect 699820 882480 699888 882536
rect 699944 882480 700012 882536
rect 700068 882480 700136 882536
rect 700192 882480 700322 882536
rect 699322 882412 700322 882480
rect 699322 882356 699392 882412
rect 699448 882356 699516 882412
rect 699572 882356 699640 882412
rect 699696 882356 699764 882412
rect 699820 882356 699888 882412
rect 699944 882356 700012 882412
rect 700068 882356 700136 882412
rect 700192 882356 700322 882412
rect 699322 882288 700322 882356
rect 699322 882232 699392 882288
rect 699448 882232 699516 882288
rect 699572 882232 699640 882288
rect 699696 882232 699764 882288
rect 699820 882232 699888 882288
rect 699944 882232 700012 882288
rect 700068 882232 700136 882288
rect 700192 882232 700322 882288
rect 699322 882164 700322 882232
rect 699322 882108 699392 882164
rect 699448 882108 699516 882164
rect 699572 882108 699640 882164
rect 699696 882108 699764 882164
rect 699820 882108 699888 882164
rect 699944 882108 700012 882164
rect 700068 882108 700136 882164
rect 700192 882108 700322 882164
rect 699322 882040 700322 882108
rect 699322 881984 699392 882040
rect 699448 881984 699516 882040
rect 699572 881984 699640 882040
rect 699696 881984 699764 882040
rect 699820 881984 699888 882040
rect 699944 881984 700012 882040
rect 700068 881984 700136 882040
rect 700192 881984 700322 882040
rect 699322 881916 700322 881984
rect 699322 881860 699392 881916
rect 699448 881860 699516 881916
rect 699572 881860 699640 881916
rect 699696 881860 699764 881916
rect 699820 881860 699888 881916
rect 699944 881860 700012 881916
rect 700068 881860 700136 881916
rect 700192 881860 700322 881916
rect 699322 881172 700322 881860
rect 707800 883658 708000 883728
rect 707800 883602 707870 883658
rect 707926 883602 708000 883658
rect 707800 883534 708000 883602
rect 707800 883478 707870 883534
rect 707926 883478 708000 883534
rect 707800 883410 708000 883478
rect 707800 883354 707870 883410
rect 707926 883354 708000 883410
rect 707800 883286 708000 883354
rect 707800 883230 707870 883286
rect 707926 883230 708000 883286
rect 707800 883162 708000 883230
rect 707800 883106 707870 883162
rect 707926 883106 708000 883162
rect 707800 883038 708000 883106
rect 707800 882982 707870 883038
rect 707926 882982 708000 883038
rect 707800 882914 708000 882982
rect 707800 882858 707870 882914
rect 707926 882858 708000 882914
rect 707800 882790 708000 882858
rect 707800 882734 707870 882790
rect 707926 882734 708000 882790
rect 707800 882666 708000 882734
rect 707800 882610 707870 882666
rect 707926 882610 708000 882666
rect 707800 882542 708000 882610
rect 707800 882486 707870 882542
rect 707926 882486 708000 882542
rect 707800 882418 708000 882486
rect 707800 882362 707870 882418
rect 707926 882362 708000 882418
rect 707800 882294 708000 882362
rect 707800 882238 707870 882294
rect 707926 882238 708000 882294
rect 707800 882170 708000 882238
rect 707800 882114 707870 882170
rect 707926 882114 708000 882170
rect 707800 882046 708000 882114
rect 707800 881990 707870 882046
rect 707926 881990 708000 882046
rect 707800 881922 708000 881990
rect 707800 881866 707870 881922
rect 707926 881866 708000 881922
rect 707800 881828 708000 881866
rect 699322 881116 699392 881172
rect 699448 881116 699516 881172
rect 699572 881116 699640 881172
rect 699696 881116 699764 881172
rect 699820 881116 699888 881172
rect 699944 881116 700012 881172
rect 700068 881116 700136 881172
rect 700192 881116 700322 881172
rect 699322 881048 700322 881116
rect 699322 880992 699392 881048
rect 699448 880992 699516 881048
rect 699572 880992 699640 881048
rect 699696 880992 699764 881048
rect 699820 880992 699888 881048
rect 699944 880992 700012 881048
rect 700068 880992 700136 881048
rect 700192 880992 700322 881048
rect 699322 880924 700322 880992
rect 699322 880868 699392 880924
rect 699448 880868 699516 880924
rect 699572 880868 699640 880924
rect 699696 880868 699764 880924
rect 699820 880868 699888 880924
rect 699944 880868 700012 880924
rect 700068 880868 700136 880924
rect 700192 880868 700322 880924
rect 699322 880800 700322 880868
rect 699322 880744 699392 880800
rect 699448 880744 699516 880800
rect 699572 880744 699640 880800
rect 699696 880744 699764 880800
rect 699820 880744 699888 880800
rect 699944 880744 700012 880800
rect 700068 880744 700136 880800
rect 700192 880744 700322 880800
rect 699322 880676 700322 880744
rect 699322 880620 699392 880676
rect 699448 880620 699516 880676
rect 699572 880620 699640 880676
rect 699696 880620 699764 880676
rect 699820 880620 699888 880676
rect 699944 880620 700012 880676
rect 700068 880620 700136 880676
rect 700192 880620 700322 880676
rect 699322 880552 700322 880620
rect 699322 880496 699392 880552
rect 699448 880496 699516 880552
rect 699572 880496 699640 880552
rect 699696 880496 699764 880552
rect 699820 880496 699888 880552
rect 699944 880496 700012 880552
rect 700068 880496 700136 880552
rect 700192 880496 700322 880552
rect 699322 880428 700322 880496
rect 699322 880372 699392 880428
rect 699448 880372 699516 880428
rect 699572 880372 699640 880428
rect 699696 880372 699764 880428
rect 699820 880372 699888 880428
rect 699944 880372 700012 880428
rect 700068 880372 700136 880428
rect 700192 880372 700322 880428
rect 699322 880304 700322 880372
rect 699322 880248 699392 880304
rect 699448 880248 699516 880304
rect 699572 880248 699640 880304
rect 699696 880248 699764 880304
rect 699820 880248 699888 880304
rect 699944 880248 700012 880304
rect 700068 880248 700136 880304
rect 700192 880248 700322 880304
rect 699322 880180 700322 880248
rect 699322 880124 699392 880180
rect 699448 880124 699516 880180
rect 699572 880124 699640 880180
rect 699696 880124 699764 880180
rect 699820 880124 699888 880180
rect 699944 880124 700012 880180
rect 700068 880124 700136 880180
rect 700192 880124 700322 880180
rect 699322 880056 700322 880124
rect 699322 880000 699392 880056
rect 699448 880000 699516 880056
rect 699572 880000 699640 880056
rect 699696 880000 699764 880056
rect 699820 880000 699888 880056
rect 699944 880000 700012 880056
rect 700068 880000 700136 880056
rect 700192 880000 700322 880056
rect 699322 879932 700322 880000
rect 699322 879876 699392 879932
rect 699448 879876 699516 879932
rect 699572 879876 699640 879932
rect 699696 879876 699764 879932
rect 699820 879876 699888 879932
rect 699944 879876 700012 879932
rect 700068 879876 700136 879932
rect 700192 879876 700322 879932
rect 699322 879808 700322 879876
rect 699322 879752 699392 879808
rect 699448 879752 699516 879808
rect 699572 879752 699640 879808
rect 699696 879752 699764 879808
rect 699820 879752 699888 879808
rect 699944 879752 700012 879808
rect 700068 879752 700136 879808
rect 700192 879752 700322 879808
rect 699322 879684 700322 879752
rect 699322 879628 699392 879684
rect 699448 879628 699516 879684
rect 699572 879628 699640 879684
rect 699696 879628 699764 879684
rect 699820 879628 699888 879684
rect 699944 879628 700012 879684
rect 700068 879628 700136 879684
rect 700192 879628 700322 879684
rect 699322 879560 700322 879628
rect 699322 879504 699392 879560
rect 699448 879504 699516 879560
rect 699572 879504 699640 879560
rect 699696 879504 699764 879560
rect 699820 879504 699888 879560
rect 699944 879504 700012 879560
rect 700068 879504 700136 879560
rect 700192 879504 700322 879560
rect 699322 879436 700322 879504
rect 699322 879380 699392 879436
rect 699448 879380 699516 879436
rect 699572 879380 699640 879436
rect 699696 879380 699764 879436
rect 699820 879380 699888 879436
rect 699944 879380 700012 879436
rect 700068 879380 700136 879436
rect 700192 879380 700322 879436
rect 699322 879312 700322 879380
rect 699322 879256 699392 879312
rect 699448 879256 699516 879312
rect 699572 879256 699640 879312
rect 699696 879256 699764 879312
rect 699820 879256 699888 879312
rect 699944 879256 700012 879312
rect 700068 879256 700136 879312
rect 700192 879256 700322 879312
rect 699322 878802 700322 879256
rect 707800 881178 708000 881248
rect 707800 881122 707870 881178
rect 707926 881122 708000 881178
rect 707800 881054 708000 881122
rect 707800 880998 707870 881054
rect 707926 880998 708000 881054
rect 707800 880930 708000 880998
rect 707800 880874 707870 880930
rect 707926 880874 708000 880930
rect 707800 880806 708000 880874
rect 707800 880750 707870 880806
rect 707926 880750 708000 880806
rect 707800 880682 708000 880750
rect 707800 880626 707870 880682
rect 707926 880626 708000 880682
rect 707800 880558 708000 880626
rect 707800 880502 707870 880558
rect 707926 880502 708000 880558
rect 707800 880434 708000 880502
rect 707800 880378 707870 880434
rect 707926 880378 708000 880434
rect 707800 880310 708000 880378
rect 707800 880254 707870 880310
rect 707926 880254 708000 880310
rect 707800 880186 708000 880254
rect 707800 880130 707870 880186
rect 707926 880130 708000 880186
rect 707800 880062 708000 880130
rect 707800 880006 707870 880062
rect 707926 880006 708000 880062
rect 707800 879938 708000 880006
rect 707800 879882 707870 879938
rect 707926 879882 708000 879938
rect 707800 879814 708000 879882
rect 707800 879758 707870 879814
rect 707926 879758 708000 879814
rect 707800 879690 708000 879758
rect 707800 879634 707870 879690
rect 707926 879634 708000 879690
rect 707800 879566 708000 879634
rect 707800 879510 707870 879566
rect 707926 879510 708000 879566
rect 707800 879442 708000 879510
rect 707800 879386 707870 879442
rect 707926 879386 708000 879442
rect 707800 879318 708000 879386
rect 707800 879262 707870 879318
rect 707926 879262 708000 879318
rect 707800 879198 708000 879262
rect 699322 878746 699392 878802
rect 699448 878746 699516 878802
rect 699572 878746 699640 878802
rect 699696 878746 699764 878802
rect 699820 878746 699888 878802
rect 699944 878746 700012 878802
rect 700068 878746 700136 878802
rect 700192 878746 700322 878802
rect 699322 878678 700322 878746
rect 699322 878622 699392 878678
rect 699448 878622 699516 878678
rect 699572 878622 699640 878678
rect 699696 878622 699764 878678
rect 699820 878622 699888 878678
rect 699944 878622 700012 878678
rect 700068 878622 700136 878678
rect 700192 878622 700322 878678
rect 699322 878554 700322 878622
rect 699322 878498 699392 878554
rect 699448 878498 699516 878554
rect 699572 878498 699640 878554
rect 699696 878498 699764 878554
rect 699820 878498 699888 878554
rect 699944 878498 700012 878554
rect 700068 878498 700136 878554
rect 700192 878498 700322 878554
rect 699322 878430 700322 878498
rect 699322 878374 699392 878430
rect 699448 878374 699516 878430
rect 699572 878374 699640 878430
rect 699696 878374 699764 878430
rect 699820 878374 699888 878430
rect 699944 878374 700012 878430
rect 700068 878374 700136 878430
rect 700192 878374 700322 878430
rect 699322 878306 700322 878374
rect 699322 878250 699392 878306
rect 699448 878250 699516 878306
rect 699572 878250 699640 878306
rect 699696 878250 699764 878306
rect 699820 878250 699888 878306
rect 699944 878250 700012 878306
rect 700068 878250 700136 878306
rect 700192 878250 700322 878306
rect 699322 878182 700322 878250
rect 699322 878126 699392 878182
rect 699448 878126 699516 878182
rect 699572 878126 699640 878182
rect 699696 878126 699764 878182
rect 699820 878126 699888 878182
rect 699944 878126 700012 878182
rect 700068 878126 700136 878182
rect 700192 878126 700322 878182
rect 699322 878058 700322 878126
rect 699322 878002 699392 878058
rect 699448 878002 699516 878058
rect 699572 878002 699640 878058
rect 699696 878002 699764 878058
rect 699820 878002 699888 878058
rect 699944 878002 700012 878058
rect 700068 878002 700136 878058
rect 700192 878002 700322 878058
rect 699322 877934 700322 878002
rect 699322 877878 699392 877934
rect 699448 877878 699516 877934
rect 699572 877878 699640 877934
rect 699696 877878 699764 877934
rect 699820 877878 699888 877934
rect 699944 877878 700012 877934
rect 700068 877878 700136 877934
rect 700192 877878 700322 877934
rect 699322 877810 700322 877878
rect 699322 877754 699392 877810
rect 699448 877754 699516 877810
rect 699572 877754 699640 877810
rect 699696 877754 699764 877810
rect 699820 877754 699888 877810
rect 699944 877754 700012 877810
rect 700068 877754 700136 877810
rect 700192 877754 700322 877810
rect 699322 877686 700322 877754
rect 699322 877630 699392 877686
rect 699448 877630 699516 877686
rect 699572 877630 699640 877686
rect 699696 877630 699764 877686
rect 699820 877630 699888 877686
rect 699944 877630 700012 877686
rect 700068 877630 700136 877686
rect 700192 877630 700322 877686
rect 699322 877562 700322 877630
rect 699322 877506 699392 877562
rect 699448 877506 699516 877562
rect 699572 877506 699640 877562
rect 699696 877506 699764 877562
rect 699820 877506 699888 877562
rect 699944 877506 700012 877562
rect 700068 877506 700136 877562
rect 700192 877506 700322 877562
rect 699322 877438 700322 877506
rect 699322 877382 699392 877438
rect 699448 877382 699516 877438
rect 699572 877382 699640 877438
rect 699696 877382 699764 877438
rect 699820 877382 699888 877438
rect 699944 877382 700012 877438
rect 700068 877382 700136 877438
rect 700192 877382 700322 877438
rect 699322 877314 700322 877382
rect 699322 877258 699392 877314
rect 699448 877258 699516 877314
rect 699572 877258 699640 877314
rect 699696 877258 699764 877314
rect 699820 877258 699888 877314
rect 699944 877258 700012 877314
rect 700068 877258 700136 877314
rect 700192 877258 700322 877314
rect 699322 877190 700322 877258
rect 699322 877134 699392 877190
rect 699448 877134 699516 877190
rect 699572 877134 699640 877190
rect 699696 877134 699764 877190
rect 699820 877134 699888 877190
rect 699944 877134 700012 877190
rect 700068 877134 700136 877190
rect 700192 877134 700322 877190
rect 699322 877066 700322 877134
rect 699322 877010 699392 877066
rect 699448 877010 699516 877066
rect 699572 877010 699640 877066
rect 699696 877010 699764 877066
rect 699820 877010 699888 877066
rect 699944 877010 700012 877066
rect 700068 877010 700136 877066
rect 700192 877010 700322 877066
rect 699322 876942 700322 877010
rect 699322 876886 699392 876942
rect 699448 876886 699516 876942
rect 699572 876886 699640 876942
rect 699696 876886 699764 876942
rect 699820 876886 699888 876942
rect 699944 876886 700012 876942
rect 700068 876886 700136 876942
rect 700192 876886 700322 876942
rect 699322 876096 700322 876886
rect 707800 878808 708000 878878
rect 707800 878752 707870 878808
rect 707926 878752 708000 878808
rect 707800 878684 708000 878752
rect 707800 878628 707870 878684
rect 707926 878628 708000 878684
rect 707800 878560 708000 878628
rect 707800 878504 707870 878560
rect 707926 878504 708000 878560
rect 707800 878436 708000 878504
rect 707800 878380 707870 878436
rect 707926 878380 708000 878436
rect 707800 878312 708000 878380
rect 707800 878256 707870 878312
rect 707926 878256 708000 878312
rect 707800 878188 708000 878256
rect 707800 878132 707870 878188
rect 707926 878132 708000 878188
rect 707800 878064 708000 878132
rect 707800 878008 707870 878064
rect 707926 878008 708000 878064
rect 707800 877940 708000 878008
rect 707800 877884 707870 877940
rect 707926 877884 708000 877940
rect 707800 877816 708000 877884
rect 707800 877760 707870 877816
rect 707926 877760 708000 877816
rect 707800 877692 708000 877760
rect 707800 877636 707870 877692
rect 707926 877636 708000 877692
rect 707800 877568 708000 877636
rect 707800 877512 707870 877568
rect 707926 877512 708000 877568
rect 707800 877444 708000 877512
rect 707800 877388 707870 877444
rect 707926 877388 708000 877444
rect 707800 877320 708000 877388
rect 707800 877264 707870 877320
rect 707926 877264 708000 877320
rect 707800 877196 708000 877264
rect 707800 877140 707870 877196
rect 707926 877140 708000 877196
rect 707800 877072 708000 877140
rect 707800 877016 707870 877072
rect 707926 877016 708000 877072
rect 707800 876948 708000 877016
rect 707800 876892 707870 876948
rect 707926 876892 708000 876948
rect 707800 876828 708000 876892
rect 699322 876040 699392 876096
rect 699448 876040 699516 876096
rect 699572 876040 699640 876096
rect 699696 876040 699764 876096
rect 699820 876040 699888 876096
rect 699944 876040 700012 876096
rect 700068 876040 700136 876096
rect 700192 876040 700322 876096
rect 699322 875972 700322 876040
rect 699322 875916 699392 875972
rect 699448 875916 699516 875972
rect 699572 875916 699640 875972
rect 699696 875916 699764 875972
rect 699820 875916 699888 875972
rect 699944 875916 700012 875972
rect 700068 875916 700136 875972
rect 700192 875916 700322 875972
rect 699322 875848 700322 875916
rect 699322 875792 699392 875848
rect 699448 875792 699516 875848
rect 699572 875792 699640 875848
rect 699696 875792 699764 875848
rect 699820 875792 699888 875848
rect 699944 875792 700012 875848
rect 700068 875792 700136 875848
rect 700192 875792 700322 875848
rect 699322 875724 700322 875792
rect 699322 875668 699392 875724
rect 699448 875668 699516 875724
rect 699572 875668 699640 875724
rect 699696 875668 699764 875724
rect 699820 875668 699888 875724
rect 699944 875668 700012 875724
rect 700068 875668 700136 875724
rect 700192 875668 700322 875724
rect 699322 875600 700322 875668
rect 699322 875544 699392 875600
rect 699448 875544 699516 875600
rect 699572 875544 699640 875600
rect 699696 875544 699764 875600
rect 699820 875544 699888 875600
rect 699944 875544 700012 875600
rect 700068 875544 700136 875600
rect 700192 875544 700322 875600
rect 699322 875476 700322 875544
rect 699322 875420 699392 875476
rect 699448 875420 699516 875476
rect 699572 875420 699640 875476
rect 699696 875420 699764 875476
rect 699820 875420 699888 875476
rect 699944 875420 700012 875476
rect 700068 875420 700136 875476
rect 700192 875420 700322 875476
rect 699322 875352 700322 875420
rect 699322 875296 699392 875352
rect 699448 875296 699516 875352
rect 699572 875296 699640 875352
rect 699696 875296 699764 875352
rect 699820 875296 699888 875352
rect 699944 875296 700012 875352
rect 700068 875296 700136 875352
rect 700192 875296 700322 875352
rect 699322 875228 700322 875296
rect 699322 875172 699392 875228
rect 699448 875172 699516 875228
rect 699572 875172 699640 875228
rect 699696 875172 699764 875228
rect 699820 875172 699888 875228
rect 699944 875172 700012 875228
rect 700068 875172 700136 875228
rect 700192 875172 700322 875228
rect 699322 875104 700322 875172
rect 699322 875048 699392 875104
rect 699448 875048 699516 875104
rect 699572 875048 699640 875104
rect 699696 875048 699764 875104
rect 699820 875048 699888 875104
rect 699944 875048 700012 875104
rect 700068 875048 700136 875104
rect 700192 875048 700322 875104
rect 699322 874980 700322 875048
rect 699322 874924 699392 874980
rect 699448 874924 699516 874980
rect 699572 874924 699640 874980
rect 699696 874924 699764 874980
rect 699820 874924 699888 874980
rect 699944 874924 700012 874980
rect 700068 874924 700136 874980
rect 700192 874924 700322 874980
rect 699322 874856 700322 874924
rect 699322 874800 699392 874856
rect 699448 874800 699516 874856
rect 699572 874800 699640 874856
rect 699696 874800 699764 874856
rect 699820 874800 699888 874856
rect 699944 874800 700012 874856
rect 700068 874800 700136 874856
rect 700192 874800 700322 874856
rect 699322 874732 700322 874800
rect 699322 874676 699392 874732
rect 699448 874676 699516 874732
rect 699572 874676 699640 874732
rect 699696 874676 699764 874732
rect 699820 874676 699888 874732
rect 699944 874676 700012 874732
rect 700068 874676 700136 874732
rect 700192 874676 700322 874732
rect 699322 874608 700322 874676
rect 699322 874552 699392 874608
rect 699448 874552 699516 874608
rect 699572 874552 699640 874608
rect 699696 874552 699764 874608
rect 699820 874552 699888 874608
rect 699944 874552 700012 874608
rect 700068 874552 700136 874608
rect 700192 874552 700322 874608
rect 699322 874484 700322 874552
rect 699322 874428 699392 874484
rect 699448 874428 699516 874484
rect 699572 874428 699640 874484
rect 699696 874428 699764 874484
rect 699820 874428 699888 874484
rect 699944 874428 700012 874484
rect 700068 874428 700136 874484
rect 700192 874428 700322 874484
rect 699322 874360 700322 874428
rect 699322 874304 699392 874360
rect 699448 874304 699516 874360
rect 699572 874304 699640 874360
rect 699696 874304 699764 874360
rect 699820 874304 699888 874360
rect 699944 874304 700012 874360
rect 700068 874304 700136 874360
rect 700192 874304 700322 874360
rect 699322 874236 700322 874304
rect 699322 874180 699392 874236
rect 699448 874180 699516 874236
rect 699572 874180 699640 874236
rect 699696 874180 699764 874236
rect 699820 874180 699888 874236
rect 699944 874180 700012 874236
rect 700068 874180 700136 874236
rect 700192 874180 700322 874236
rect 699322 873726 700322 874180
rect 707800 876102 708000 876172
rect 707800 876046 707870 876102
rect 707926 876046 708000 876102
rect 707800 875978 708000 876046
rect 707800 875922 707870 875978
rect 707926 875922 708000 875978
rect 707800 875854 708000 875922
rect 707800 875798 707870 875854
rect 707926 875798 708000 875854
rect 707800 875730 708000 875798
rect 707800 875674 707870 875730
rect 707926 875674 708000 875730
rect 707800 875606 708000 875674
rect 707800 875550 707870 875606
rect 707926 875550 708000 875606
rect 707800 875482 708000 875550
rect 707800 875426 707870 875482
rect 707926 875426 708000 875482
rect 707800 875358 708000 875426
rect 707800 875302 707870 875358
rect 707926 875302 708000 875358
rect 707800 875234 708000 875302
rect 707800 875178 707870 875234
rect 707926 875178 708000 875234
rect 707800 875110 708000 875178
rect 707800 875054 707870 875110
rect 707926 875054 708000 875110
rect 707800 874986 708000 875054
rect 707800 874930 707870 874986
rect 707926 874930 708000 874986
rect 707800 874862 708000 874930
rect 707800 874806 707870 874862
rect 707926 874806 708000 874862
rect 707800 874738 708000 874806
rect 707800 874682 707870 874738
rect 707926 874682 708000 874738
rect 707800 874614 708000 874682
rect 707800 874558 707870 874614
rect 707926 874558 708000 874614
rect 707800 874490 708000 874558
rect 707800 874434 707870 874490
rect 707926 874434 708000 874490
rect 707800 874366 708000 874434
rect 707800 874310 707870 874366
rect 707926 874310 708000 874366
rect 707800 874242 708000 874310
rect 707800 874186 707870 874242
rect 707926 874186 708000 874242
rect 707800 874122 708000 874186
rect 699322 873670 699392 873726
rect 699448 873670 699516 873726
rect 699572 873670 699640 873726
rect 699696 873670 699764 873726
rect 699820 873670 699888 873726
rect 699944 873670 700012 873726
rect 700068 873670 700136 873726
rect 700192 873670 700322 873726
rect 699322 873602 700322 873670
rect 699322 873546 699392 873602
rect 699448 873546 699516 873602
rect 699572 873546 699640 873602
rect 699696 873546 699764 873602
rect 699820 873546 699888 873602
rect 699944 873546 700012 873602
rect 700068 873546 700136 873602
rect 700192 873546 700322 873602
rect 699322 873478 700322 873546
rect 699322 873422 699392 873478
rect 699448 873422 699516 873478
rect 699572 873422 699640 873478
rect 699696 873422 699764 873478
rect 699820 873422 699888 873478
rect 699944 873422 700012 873478
rect 700068 873422 700136 873478
rect 700192 873422 700322 873478
rect 699322 873354 700322 873422
rect 699322 873298 699392 873354
rect 699448 873298 699516 873354
rect 699572 873298 699640 873354
rect 699696 873298 699764 873354
rect 699820 873298 699888 873354
rect 699944 873298 700012 873354
rect 700068 873298 700136 873354
rect 700192 873298 700322 873354
rect 699322 873230 700322 873298
rect 699322 873174 699392 873230
rect 699448 873174 699516 873230
rect 699572 873174 699640 873230
rect 699696 873174 699764 873230
rect 699820 873174 699888 873230
rect 699944 873174 700012 873230
rect 700068 873174 700136 873230
rect 700192 873174 700322 873230
rect 699322 873106 700322 873174
rect 699322 873050 699392 873106
rect 699448 873050 699516 873106
rect 699572 873050 699640 873106
rect 699696 873050 699764 873106
rect 699820 873050 699888 873106
rect 699944 873050 700012 873106
rect 700068 873050 700136 873106
rect 700192 873050 700322 873106
rect 699322 872982 700322 873050
rect 699322 872926 699392 872982
rect 699448 872926 699516 872982
rect 699572 872926 699640 872982
rect 699696 872926 699764 872982
rect 699820 872926 699888 872982
rect 699944 872926 700012 872982
rect 700068 872926 700136 872982
rect 700192 872926 700322 872982
rect 699322 872858 700322 872926
rect 699322 872802 699392 872858
rect 699448 872802 699516 872858
rect 699572 872802 699640 872858
rect 699696 872802 699764 872858
rect 699820 872802 699888 872858
rect 699944 872802 700012 872858
rect 700068 872802 700136 872858
rect 700192 872802 700322 872858
rect 699322 872734 700322 872802
rect 699322 872678 699392 872734
rect 699448 872678 699516 872734
rect 699572 872678 699640 872734
rect 699696 872678 699764 872734
rect 699820 872678 699888 872734
rect 699944 872678 700012 872734
rect 700068 872678 700136 872734
rect 700192 872678 700322 872734
rect 699322 872610 700322 872678
rect 699322 872554 699392 872610
rect 699448 872554 699516 872610
rect 699572 872554 699640 872610
rect 699696 872554 699764 872610
rect 699820 872554 699888 872610
rect 699944 872554 700012 872610
rect 700068 872554 700136 872610
rect 700192 872554 700322 872610
rect 699322 872486 700322 872554
rect 699322 872430 699392 872486
rect 699448 872430 699516 872486
rect 699572 872430 699640 872486
rect 699696 872430 699764 872486
rect 699820 872430 699888 872486
rect 699944 872430 700012 872486
rect 700068 872430 700136 872486
rect 700192 872430 700322 872486
rect 699322 872362 700322 872430
rect 699322 872306 699392 872362
rect 699448 872306 699516 872362
rect 699572 872306 699640 872362
rect 699696 872306 699764 872362
rect 699820 872306 699888 872362
rect 699944 872306 700012 872362
rect 700068 872306 700136 872362
rect 700192 872306 700322 872362
rect 699322 872238 700322 872306
rect 699322 872182 699392 872238
rect 699448 872182 699516 872238
rect 699572 872182 699640 872238
rect 699696 872182 699764 872238
rect 699820 872182 699888 872238
rect 699944 872182 700012 872238
rect 700068 872182 700136 872238
rect 700192 872182 700322 872238
rect 699322 872114 700322 872182
rect 699322 872058 699392 872114
rect 699448 872058 699516 872114
rect 699572 872058 699640 872114
rect 699696 872058 699764 872114
rect 699820 872058 699888 872114
rect 699944 872058 700012 872114
rect 700068 872058 700136 872114
rect 700192 872058 700322 872114
rect 699322 871990 700322 872058
rect 699322 871934 699392 871990
rect 699448 871934 699516 871990
rect 699572 871934 699640 871990
rect 699696 871934 699764 871990
rect 699820 871934 699888 871990
rect 699944 871934 700012 871990
rect 700068 871934 700136 871990
rect 700192 871934 700322 871990
rect 699322 871866 700322 871934
rect 699322 871810 699392 871866
rect 699448 871810 699516 871866
rect 699572 871810 699640 871866
rect 699696 871810 699764 871866
rect 699820 871810 699888 871866
rect 699944 871810 700012 871866
rect 700068 871810 700136 871866
rect 700192 871810 700322 871866
rect 699322 871122 700322 871810
rect 707800 873732 708000 873802
rect 707800 873676 707870 873732
rect 707926 873676 708000 873732
rect 707800 873608 708000 873676
rect 707800 873552 707870 873608
rect 707926 873552 708000 873608
rect 707800 873484 708000 873552
rect 707800 873428 707870 873484
rect 707926 873428 708000 873484
rect 707800 873360 708000 873428
rect 707800 873304 707870 873360
rect 707926 873304 708000 873360
rect 707800 873236 708000 873304
rect 707800 873180 707870 873236
rect 707926 873180 708000 873236
rect 707800 873112 708000 873180
rect 707800 873056 707870 873112
rect 707926 873056 708000 873112
rect 707800 872988 708000 873056
rect 707800 872932 707870 872988
rect 707926 872932 708000 872988
rect 707800 872864 708000 872932
rect 707800 872808 707870 872864
rect 707926 872808 708000 872864
rect 707800 872740 708000 872808
rect 707800 872684 707870 872740
rect 707926 872684 708000 872740
rect 707800 872616 708000 872684
rect 707800 872560 707870 872616
rect 707926 872560 708000 872616
rect 707800 872492 708000 872560
rect 707800 872436 707870 872492
rect 707926 872436 708000 872492
rect 707800 872368 708000 872436
rect 707800 872312 707870 872368
rect 707926 872312 708000 872368
rect 707800 872244 708000 872312
rect 707800 872188 707870 872244
rect 707926 872188 708000 872244
rect 707800 872120 708000 872188
rect 707800 872064 707870 872120
rect 707926 872064 708000 872120
rect 707800 871996 708000 872064
rect 707800 871940 707870 871996
rect 707926 871940 708000 871996
rect 707800 871872 708000 871940
rect 707800 871816 707870 871872
rect 707926 871816 708000 871872
rect 707800 871752 708000 871816
rect 699322 871066 699392 871122
rect 699448 871066 699516 871122
rect 699572 871066 699640 871122
rect 699696 871066 699764 871122
rect 699820 871066 699888 871122
rect 699944 871066 700012 871122
rect 700068 871066 700136 871122
rect 700192 871066 700322 871122
rect 699322 870998 700322 871066
rect 699322 870942 699392 870998
rect 699448 870942 699516 870998
rect 699572 870942 699640 870998
rect 699696 870942 699764 870998
rect 699820 870942 699888 870998
rect 699944 870942 700012 870998
rect 700068 870942 700136 870998
rect 700192 870942 700322 870998
rect 699322 870874 700322 870942
rect 699322 870818 699392 870874
rect 699448 870818 699516 870874
rect 699572 870818 699640 870874
rect 699696 870818 699764 870874
rect 699820 870818 699888 870874
rect 699944 870818 700012 870874
rect 700068 870818 700136 870874
rect 700192 870818 700322 870874
rect 699322 870750 700322 870818
rect 699322 870694 699392 870750
rect 699448 870694 699516 870750
rect 699572 870694 699640 870750
rect 699696 870694 699764 870750
rect 699820 870694 699888 870750
rect 699944 870694 700012 870750
rect 700068 870694 700136 870750
rect 700192 870694 700322 870750
rect 699322 870626 700322 870694
rect 699322 870570 699392 870626
rect 699448 870570 699516 870626
rect 699572 870570 699640 870626
rect 699696 870570 699764 870626
rect 699820 870570 699888 870626
rect 699944 870570 700012 870626
rect 700068 870570 700136 870626
rect 700192 870570 700322 870626
rect 699322 870502 700322 870570
rect 699322 870446 699392 870502
rect 699448 870446 699516 870502
rect 699572 870446 699640 870502
rect 699696 870446 699764 870502
rect 699820 870446 699888 870502
rect 699944 870446 700012 870502
rect 700068 870446 700136 870502
rect 700192 870446 700322 870502
rect 699322 870378 700322 870446
rect 699322 870322 699392 870378
rect 699448 870322 699516 870378
rect 699572 870322 699640 870378
rect 699696 870322 699764 870378
rect 699820 870322 699888 870378
rect 699944 870322 700012 870378
rect 700068 870322 700136 870378
rect 700192 870322 700322 870378
rect 699322 870254 700322 870322
rect 699322 870198 699392 870254
rect 699448 870198 699516 870254
rect 699572 870198 699640 870254
rect 699696 870198 699764 870254
rect 699820 870198 699888 870254
rect 699944 870198 700012 870254
rect 700068 870198 700136 870254
rect 700192 870198 700322 870254
rect 699322 870130 700322 870198
rect 699322 870074 699392 870130
rect 699448 870074 699516 870130
rect 699572 870074 699640 870130
rect 699696 870074 699764 870130
rect 699820 870074 699888 870130
rect 699944 870074 700012 870130
rect 700068 870074 700136 870130
rect 700192 870074 700322 870130
rect 699322 870006 700322 870074
rect 699322 869950 699392 870006
rect 699448 869950 699516 870006
rect 699572 869950 699640 870006
rect 699696 869950 699764 870006
rect 699820 869950 699888 870006
rect 699944 869950 700012 870006
rect 700068 869950 700136 870006
rect 700192 869950 700322 870006
rect 699322 869882 700322 869950
rect 699322 869826 699392 869882
rect 699448 869826 699516 869882
rect 699572 869826 699640 869882
rect 699696 869826 699764 869882
rect 699820 869826 699888 869882
rect 699944 869826 700012 869882
rect 700068 869826 700136 869882
rect 700192 869826 700322 869882
rect 699322 869758 700322 869826
rect 699322 869702 699392 869758
rect 699448 869702 699516 869758
rect 699572 869702 699640 869758
rect 699696 869702 699764 869758
rect 699820 869702 699888 869758
rect 699944 869702 700012 869758
rect 700068 869702 700136 869758
rect 700192 869702 700322 869758
rect 699322 869634 700322 869702
rect 699322 869578 699392 869634
rect 699448 869578 699516 869634
rect 699572 869578 699640 869634
rect 699696 869578 699764 869634
rect 699820 869578 699888 869634
rect 699944 869578 700012 869634
rect 700068 869578 700136 869634
rect 700192 869578 700322 869634
rect 699322 869510 700322 869578
rect 699322 869454 699392 869510
rect 699448 869454 699516 869510
rect 699572 869454 699640 869510
rect 699696 869454 699764 869510
rect 699820 869454 699888 869510
rect 699944 869454 700012 869510
rect 700068 869454 700136 869510
rect 700192 869454 700322 869510
rect 699322 869386 700322 869454
rect 699322 869330 699392 869386
rect 699448 869330 699516 869386
rect 699572 869330 699640 869386
rect 699696 869330 699764 869386
rect 699820 869330 699888 869386
rect 699944 869330 700012 869386
rect 700068 869330 700136 869386
rect 700192 869330 700322 869386
rect 699322 842429 700322 869330
rect 707800 871134 708000 871172
rect 707800 871078 707870 871134
rect 707926 871078 708000 871134
rect 707800 871010 708000 871078
rect 707800 870954 707870 871010
rect 707926 870954 708000 871010
rect 707800 870886 708000 870954
rect 707800 870830 707870 870886
rect 707926 870830 708000 870886
rect 707800 870762 708000 870830
rect 707800 870706 707870 870762
rect 707926 870706 708000 870762
rect 707800 870638 708000 870706
rect 707800 870582 707870 870638
rect 707926 870582 708000 870638
rect 707800 870514 708000 870582
rect 707800 870458 707870 870514
rect 707926 870458 708000 870514
rect 707800 870390 708000 870458
rect 707800 870334 707870 870390
rect 707926 870334 708000 870390
rect 707800 870266 708000 870334
rect 707800 870210 707870 870266
rect 707926 870210 708000 870266
rect 707800 870142 708000 870210
rect 707800 870086 707870 870142
rect 707926 870086 708000 870142
rect 707800 870018 708000 870086
rect 707800 869962 707870 870018
rect 707926 869962 708000 870018
rect 707800 869894 708000 869962
rect 707800 869838 707870 869894
rect 707926 869838 708000 869894
rect 707800 869770 708000 869838
rect 707800 869714 707870 869770
rect 707926 869714 708000 869770
rect 707800 869646 708000 869714
rect 707800 869590 707870 869646
rect 707926 869590 708000 869646
rect 707800 869522 708000 869590
rect 707800 869466 707870 869522
rect 707926 869466 708000 869522
rect 707800 869398 708000 869466
rect 707800 869342 707870 869398
rect 707926 869342 708000 869398
rect 707800 869272 708000 869342
rect 699322 842373 699544 842429
rect 699600 842373 699844 842429
rect 699900 842373 700144 842429
rect 700200 842373 700322 842429
rect 699322 842229 700322 842373
rect 699322 842173 699544 842229
rect 699600 842173 699844 842229
rect 699900 842173 700144 842229
rect 700200 842173 700322 842229
rect 699322 839954 700322 842173
rect 699322 839898 699444 839954
rect 699500 839898 699744 839954
rect 699800 839898 700044 839954
rect 700100 839898 700322 839954
rect 699322 832954 700322 839898
rect 699322 832898 699444 832954
rect 699500 832898 699744 832954
rect 699800 832898 700044 832954
rect 700100 832898 700322 832954
rect 699322 825954 700322 832898
rect 699322 825898 699444 825954
rect 699500 825898 699744 825954
rect 699800 825898 700044 825954
rect 700100 825898 700322 825954
rect 699322 806423 700322 825898
rect 699322 806367 699497 806423
rect 699553 806367 699797 806423
rect 699853 806367 700097 806423
rect 700153 806367 700322 806423
rect 699322 797652 700322 806367
rect 699322 797596 699392 797652
rect 699448 797596 699516 797652
rect 699572 797596 699640 797652
rect 699696 797596 699764 797652
rect 699820 797596 699888 797652
rect 699944 797596 700012 797652
rect 700068 797596 700136 797652
rect 700192 797596 700322 797652
rect 699322 797528 700322 797596
rect 699322 797472 699392 797528
rect 699448 797472 699516 797528
rect 699572 797472 699640 797528
rect 699696 797472 699764 797528
rect 699820 797472 699888 797528
rect 699944 797472 700012 797528
rect 700068 797472 700136 797528
rect 700192 797472 700322 797528
rect 699322 797404 700322 797472
rect 699322 797348 699392 797404
rect 699448 797348 699516 797404
rect 699572 797348 699640 797404
rect 699696 797348 699764 797404
rect 699820 797348 699888 797404
rect 699944 797348 700012 797404
rect 700068 797348 700136 797404
rect 700192 797348 700322 797404
rect 699322 797280 700322 797348
rect 699322 797224 699392 797280
rect 699448 797224 699516 797280
rect 699572 797224 699640 797280
rect 699696 797224 699764 797280
rect 699820 797224 699888 797280
rect 699944 797224 700012 797280
rect 700068 797224 700136 797280
rect 700192 797224 700322 797280
rect 699322 797156 700322 797224
rect 699322 797100 699392 797156
rect 699448 797100 699516 797156
rect 699572 797100 699640 797156
rect 699696 797100 699764 797156
rect 699820 797100 699888 797156
rect 699944 797100 700012 797156
rect 700068 797100 700136 797156
rect 700192 797100 700322 797156
rect 699322 797032 700322 797100
rect 699322 796976 699392 797032
rect 699448 796976 699516 797032
rect 699572 796976 699640 797032
rect 699696 796976 699764 797032
rect 699820 796976 699888 797032
rect 699944 796976 700012 797032
rect 700068 796976 700136 797032
rect 700192 796976 700322 797032
rect 699322 796908 700322 796976
rect 699322 796852 699392 796908
rect 699448 796852 699516 796908
rect 699572 796852 699640 796908
rect 699696 796852 699764 796908
rect 699820 796852 699888 796908
rect 699944 796852 700012 796908
rect 700068 796852 700136 796908
rect 700192 796852 700322 796908
rect 699322 796784 700322 796852
rect 699322 796728 699392 796784
rect 699448 796728 699516 796784
rect 699572 796728 699640 796784
rect 699696 796728 699764 796784
rect 699820 796728 699888 796784
rect 699944 796728 700012 796784
rect 700068 796728 700136 796784
rect 700192 796728 700322 796784
rect 699322 796660 700322 796728
rect 699322 796604 699392 796660
rect 699448 796604 699516 796660
rect 699572 796604 699640 796660
rect 699696 796604 699764 796660
rect 699820 796604 699888 796660
rect 699944 796604 700012 796660
rect 700068 796604 700136 796660
rect 700192 796604 700322 796660
rect 699322 796536 700322 796604
rect 699322 796480 699392 796536
rect 699448 796480 699516 796536
rect 699572 796480 699640 796536
rect 699696 796480 699764 796536
rect 699820 796480 699888 796536
rect 699944 796480 700012 796536
rect 700068 796480 700136 796536
rect 700192 796480 700322 796536
rect 699322 796412 700322 796480
rect 699322 796356 699392 796412
rect 699448 796356 699516 796412
rect 699572 796356 699640 796412
rect 699696 796356 699764 796412
rect 699820 796356 699888 796412
rect 699944 796356 700012 796412
rect 700068 796356 700136 796412
rect 700192 796356 700322 796412
rect 699322 796288 700322 796356
rect 699322 796232 699392 796288
rect 699448 796232 699516 796288
rect 699572 796232 699640 796288
rect 699696 796232 699764 796288
rect 699820 796232 699888 796288
rect 699944 796232 700012 796288
rect 700068 796232 700136 796288
rect 700192 796232 700322 796288
rect 699322 796164 700322 796232
rect 699322 796108 699392 796164
rect 699448 796108 699516 796164
rect 699572 796108 699640 796164
rect 699696 796108 699764 796164
rect 699820 796108 699888 796164
rect 699944 796108 700012 796164
rect 700068 796108 700136 796164
rect 700192 796108 700322 796164
rect 699322 796040 700322 796108
rect 699322 795984 699392 796040
rect 699448 795984 699516 796040
rect 699572 795984 699640 796040
rect 699696 795984 699764 796040
rect 699820 795984 699888 796040
rect 699944 795984 700012 796040
rect 700068 795984 700136 796040
rect 700192 795984 700322 796040
rect 699322 795916 700322 795984
rect 699322 795860 699392 795916
rect 699448 795860 699516 795916
rect 699572 795860 699640 795916
rect 699696 795860 699764 795916
rect 699820 795860 699888 795916
rect 699944 795860 700012 795916
rect 700068 795860 700136 795916
rect 700192 795860 700322 795916
rect 699322 795172 700322 795860
rect 707800 797658 708000 797728
rect 707800 797602 707870 797658
rect 707926 797602 708000 797658
rect 707800 797534 708000 797602
rect 707800 797478 707870 797534
rect 707926 797478 708000 797534
rect 707800 797410 708000 797478
rect 707800 797354 707870 797410
rect 707926 797354 708000 797410
rect 707800 797286 708000 797354
rect 707800 797230 707870 797286
rect 707926 797230 708000 797286
rect 707800 797162 708000 797230
rect 707800 797106 707870 797162
rect 707926 797106 708000 797162
rect 707800 797038 708000 797106
rect 707800 796982 707870 797038
rect 707926 796982 708000 797038
rect 707800 796914 708000 796982
rect 707800 796858 707870 796914
rect 707926 796858 708000 796914
rect 707800 796790 708000 796858
rect 707800 796734 707870 796790
rect 707926 796734 708000 796790
rect 707800 796666 708000 796734
rect 707800 796610 707870 796666
rect 707926 796610 708000 796666
rect 707800 796542 708000 796610
rect 707800 796486 707870 796542
rect 707926 796486 708000 796542
rect 707800 796418 708000 796486
rect 707800 796362 707870 796418
rect 707926 796362 708000 796418
rect 707800 796294 708000 796362
rect 707800 796238 707870 796294
rect 707926 796238 708000 796294
rect 707800 796170 708000 796238
rect 707800 796114 707870 796170
rect 707926 796114 708000 796170
rect 707800 796046 708000 796114
rect 707800 795990 707870 796046
rect 707926 795990 708000 796046
rect 707800 795922 708000 795990
rect 707800 795866 707870 795922
rect 707926 795866 708000 795922
rect 707800 795828 708000 795866
rect 699322 795116 699392 795172
rect 699448 795116 699516 795172
rect 699572 795116 699640 795172
rect 699696 795116 699764 795172
rect 699820 795116 699888 795172
rect 699944 795116 700012 795172
rect 700068 795116 700136 795172
rect 700192 795116 700322 795172
rect 699322 795048 700322 795116
rect 699322 794992 699392 795048
rect 699448 794992 699516 795048
rect 699572 794992 699640 795048
rect 699696 794992 699764 795048
rect 699820 794992 699888 795048
rect 699944 794992 700012 795048
rect 700068 794992 700136 795048
rect 700192 794992 700322 795048
rect 699322 794924 700322 794992
rect 699322 794868 699392 794924
rect 699448 794868 699516 794924
rect 699572 794868 699640 794924
rect 699696 794868 699764 794924
rect 699820 794868 699888 794924
rect 699944 794868 700012 794924
rect 700068 794868 700136 794924
rect 700192 794868 700322 794924
rect 699322 794800 700322 794868
rect 699322 794744 699392 794800
rect 699448 794744 699516 794800
rect 699572 794744 699640 794800
rect 699696 794744 699764 794800
rect 699820 794744 699888 794800
rect 699944 794744 700012 794800
rect 700068 794744 700136 794800
rect 700192 794744 700322 794800
rect 699322 794676 700322 794744
rect 699322 794620 699392 794676
rect 699448 794620 699516 794676
rect 699572 794620 699640 794676
rect 699696 794620 699764 794676
rect 699820 794620 699888 794676
rect 699944 794620 700012 794676
rect 700068 794620 700136 794676
rect 700192 794620 700322 794676
rect 699322 794552 700322 794620
rect 699322 794496 699392 794552
rect 699448 794496 699516 794552
rect 699572 794496 699640 794552
rect 699696 794496 699764 794552
rect 699820 794496 699888 794552
rect 699944 794496 700012 794552
rect 700068 794496 700136 794552
rect 700192 794496 700322 794552
rect 699322 794428 700322 794496
rect 699322 794372 699392 794428
rect 699448 794372 699516 794428
rect 699572 794372 699640 794428
rect 699696 794372 699764 794428
rect 699820 794372 699888 794428
rect 699944 794372 700012 794428
rect 700068 794372 700136 794428
rect 700192 794372 700322 794428
rect 699322 794304 700322 794372
rect 699322 794248 699392 794304
rect 699448 794248 699516 794304
rect 699572 794248 699640 794304
rect 699696 794248 699764 794304
rect 699820 794248 699888 794304
rect 699944 794248 700012 794304
rect 700068 794248 700136 794304
rect 700192 794248 700322 794304
rect 699322 794180 700322 794248
rect 699322 794124 699392 794180
rect 699448 794124 699516 794180
rect 699572 794124 699640 794180
rect 699696 794124 699764 794180
rect 699820 794124 699888 794180
rect 699944 794124 700012 794180
rect 700068 794124 700136 794180
rect 700192 794124 700322 794180
rect 699322 794056 700322 794124
rect 699322 794000 699392 794056
rect 699448 794000 699516 794056
rect 699572 794000 699640 794056
rect 699696 794000 699764 794056
rect 699820 794000 699888 794056
rect 699944 794000 700012 794056
rect 700068 794000 700136 794056
rect 700192 794000 700322 794056
rect 699322 793932 700322 794000
rect 699322 793876 699392 793932
rect 699448 793876 699516 793932
rect 699572 793876 699640 793932
rect 699696 793876 699764 793932
rect 699820 793876 699888 793932
rect 699944 793876 700012 793932
rect 700068 793876 700136 793932
rect 700192 793876 700322 793932
rect 699322 793808 700322 793876
rect 699322 793752 699392 793808
rect 699448 793752 699516 793808
rect 699572 793752 699640 793808
rect 699696 793752 699764 793808
rect 699820 793752 699888 793808
rect 699944 793752 700012 793808
rect 700068 793752 700136 793808
rect 700192 793752 700322 793808
rect 699322 793684 700322 793752
rect 699322 793628 699392 793684
rect 699448 793628 699516 793684
rect 699572 793628 699640 793684
rect 699696 793628 699764 793684
rect 699820 793628 699888 793684
rect 699944 793628 700012 793684
rect 700068 793628 700136 793684
rect 700192 793628 700322 793684
rect 699322 793560 700322 793628
rect 699322 793504 699392 793560
rect 699448 793504 699516 793560
rect 699572 793504 699640 793560
rect 699696 793504 699764 793560
rect 699820 793504 699888 793560
rect 699944 793504 700012 793560
rect 700068 793504 700136 793560
rect 700192 793504 700322 793560
rect 699322 793436 700322 793504
rect 699322 793380 699392 793436
rect 699448 793380 699516 793436
rect 699572 793380 699640 793436
rect 699696 793380 699764 793436
rect 699820 793380 699888 793436
rect 699944 793380 700012 793436
rect 700068 793380 700136 793436
rect 700192 793380 700322 793436
rect 699322 793312 700322 793380
rect 699322 793256 699392 793312
rect 699448 793256 699516 793312
rect 699572 793256 699640 793312
rect 699696 793256 699764 793312
rect 699820 793256 699888 793312
rect 699944 793256 700012 793312
rect 700068 793256 700136 793312
rect 700192 793256 700322 793312
rect 699322 792802 700322 793256
rect 707800 795178 708000 795248
rect 707800 795122 707870 795178
rect 707926 795122 708000 795178
rect 707800 795054 708000 795122
rect 707800 794998 707870 795054
rect 707926 794998 708000 795054
rect 707800 794930 708000 794998
rect 707800 794874 707870 794930
rect 707926 794874 708000 794930
rect 707800 794806 708000 794874
rect 707800 794750 707870 794806
rect 707926 794750 708000 794806
rect 707800 794682 708000 794750
rect 707800 794626 707870 794682
rect 707926 794626 708000 794682
rect 707800 794558 708000 794626
rect 707800 794502 707870 794558
rect 707926 794502 708000 794558
rect 707800 794434 708000 794502
rect 707800 794378 707870 794434
rect 707926 794378 708000 794434
rect 707800 794310 708000 794378
rect 707800 794254 707870 794310
rect 707926 794254 708000 794310
rect 707800 794186 708000 794254
rect 707800 794130 707870 794186
rect 707926 794130 708000 794186
rect 707800 794062 708000 794130
rect 707800 794006 707870 794062
rect 707926 794006 708000 794062
rect 707800 793938 708000 794006
rect 707800 793882 707870 793938
rect 707926 793882 708000 793938
rect 707800 793814 708000 793882
rect 707800 793758 707870 793814
rect 707926 793758 708000 793814
rect 707800 793690 708000 793758
rect 707800 793634 707870 793690
rect 707926 793634 708000 793690
rect 707800 793566 708000 793634
rect 707800 793510 707870 793566
rect 707926 793510 708000 793566
rect 707800 793442 708000 793510
rect 707800 793386 707870 793442
rect 707926 793386 708000 793442
rect 707800 793318 708000 793386
rect 707800 793262 707870 793318
rect 707926 793262 708000 793318
rect 707800 793198 708000 793262
rect 699322 792746 699392 792802
rect 699448 792746 699516 792802
rect 699572 792746 699640 792802
rect 699696 792746 699764 792802
rect 699820 792746 699888 792802
rect 699944 792746 700012 792802
rect 700068 792746 700136 792802
rect 700192 792746 700322 792802
rect 699322 792678 700322 792746
rect 699322 792622 699392 792678
rect 699448 792622 699516 792678
rect 699572 792622 699640 792678
rect 699696 792622 699764 792678
rect 699820 792622 699888 792678
rect 699944 792622 700012 792678
rect 700068 792622 700136 792678
rect 700192 792622 700322 792678
rect 699322 792554 700322 792622
rect 699322 792498 699392 792554
rect 699448 792498 699516 792554
rect 699572 792498 699640 792554
rect 699696 792498 699764 792554
rect 699820 792498 699888 792554
rect 699944 792498 700012 792554
rect 700068 792498 700136 792554
rect 700192 792498 700322 792554
rect 699322 792430 700322 792498
rect 699322 792374 699392 792430
rect 699448 792374 699516 792430
rect 699572 792374 699640 792430
rect 699696 792374 699764 792430
rect 699820 792374 699888 792430
rect 699944 792374 700012 792430
rect 700068 792374 700136 792430
rect 700192 792374 700322 792430
rect 699322 792306 700322 792374
rect 699322 792250 699392 792306
rect 699448 792250 699516 792306
rect 699572 792250 699640 792306
rect 699696 792250 699764 792306
rect 699820 792250 699888 792306
rect 699944 792250 700012 792306
rect 700068 792250 700136 792306
rect 700192 792250 700322 792306
rect 699322 792182 700322 792250
rect 699322 792126 699392 792182
rect 699448 792126 699516 792182
rect 699572 792126 699640 792182
rect 699696 792126 699764 792182
rect 699820 792126 699888 792182
rect 699944 792126 700012 792182
rect 700068 792126 700136 792182
rect 700192 792126 700322 792182
rect 699322 792058 700322 792126
rect 699322 792002 699392 792058
rect 699448 792002 699516 792058
rect 699572 792002 699640 792058
rect 699696 792002 699764 792058
rect 699820 792002 699888 792058
rect 699944 792002 700012 792058
rect 700068 792002 700136 792058
rect 700192 792002 700322 792058
rect 699322 791934 700322 792002
rect 699322 791878 699392 791934
rect 699448 791878 699516 791934
rect 699572 791878 699640 791934
rect 699696 791878 699764 791934
rect 699820 791878 699888 791934
rect 699944 791878 700012 791934
rect 700068 791878 700136 791934
rect 700192 791878 700322 791934
rect 699322 791810 700322 791878
rect 699322 791754 699392 791810
rect 699448 791754 699516 791810
rect 699572 791754 699640 791810
rect 699696 791754 699764 791810
rect 699820 791754 699888 791810
rect 699944 791754 700012 791810
rect 700068 791754 700136 791810
rect 700192 791754 700322 791810
rect 699322 791686 700322 791754
rect 699322 791630 699392 791686
rect 699448 791630 699516 791686
rect 699572 791630 699640 791686
rect 699696 791630 699764 791686
rect 699820 791630 699888 791686
rect 699944 791630 700012 791686
rect 700068 791630 700136 791686
rect 700192 791630 700322 791686
rect 699322 791562 700322 791630
rect 699322 791506 699392 791562
rect 699448 791506 699516 791562
rect 699572 791506 699640 791562
rect 699696 791506 699764 791562
rect 699820 791506 699888 791562
rect 699944 791506 700012 791562
rect 700068 791506 700136 791562
rect 700192 791506 700322 791562
rect 699322 791438 700322 791506
rect 699322 791382 699392 791438
rect 699448 791382 699516 791438
rect 699572 791382 699640 791438
rect 699696 791382 699764 791438
rect 699820 791382 699888 791438
rect 699944 791382 700012 791438
rect 700068 791382 700136 791438
rect 700192 791382 700322 791438
rect 699322 791314 700322 791382
rect 699322 791258 699392 791314
rect 699448 791258 699516 791314
rect 699572 791258 699640 791314
rect 699696 791258 699764 791314
rect 699820 791258 699888 791314
rect 699944 791258 700012 791314
rect 700068 791258 700136 791314
rect 700192 791258 700322 791314
rect 699322 791190 700322 791258
rect 699322 791134 699392 791190
rect 699448 791134 699516 791190
rect 699572 791134 699640 791190
rect 699696 791134 699764 791190
rect 699820 791134 699888 791190
rect 699944 791134 700012 791190
rect 700068 791134 700136 791190
rect 700192 791134 700322 791190
rect 699322 791066 700322 791134
rect 699322 791010 699392 791066
rect 699448 791010 699516 791066
rect 699572 791010 699640 791066
rect 699696 791010 699764 791066
rect 699820 791010 699888 791066
rect 699944 791010 700012 791066
rect 700068 791010 700136 791066
rect 700192 791010 700322 791066
rect 699322 790942 700322 791010
rect 699322 790886 699392 790942
rect 699448 790886 699516 790942
rect 699572 790886 699640 790942
rect 699696 790886 699764 790942
rect 699820 790886 699888 790942
rect 699944 790886 700012 790942
rect 700068 790886 700136 790942
rect 700192 790886 700322 790942
rect 699322 790096 700322 790886
rect 707800 792808 708000 792878
rect 707800 792752 707870 792808
rect 707926 792752 708000 792808
rect 707800 792684 708000 792752
rect 707800 792628 707870 792684
rect 707926 792628 708000 792684
rect 707800 792560 708000 792628
rect 707800 792504 707870 792560
rect 707926 792504 708000 792560
rect 707800 792436 708000 792504
rect 707800 792380 707870 792436
rect 707926 792380 708000 792436
rect 707800 792312 708000 792380
rect 707800 792256 707870 792312
rect 707926 792256 708000 792312
rect 707800 792188 708000 792256
rect 707800 792132 707870 792188
rect 707926 792132 708000 792188
rect 707800 792064 708000 792132
rect 707800 792008 707870 792064
rect 707926 792008 708000 792064
rect 707800 791940 708000 792008
rect 707800 791884 707870 791940
rect 707926 791884 708000 791940
rect 707800 791816 708000 791884
rect 707800 791760 707870 791816
rect 707926 791760 708000 791816
rect 707800 791692 708000 791760
rect 707800 791636 707870 791692
rect 707926 791636 708000 791692
rect 707800 791568 708000 791636
rect 707800 791512 707870 791568
rect 707926 791512 708000 791568
rect 707800 791444 708000 791512
rect 707800 791388 707870 791444
rect 707926 791388 708000 791444
rect 707800 791320 708000 791388
rect 707800 791264 707870 791320
rect 707926 791264 708000 791320
rect 707800 791196 708000 791264
rect 707800 791140 707870 791196
rect 707926 791140 708000 791196
rect 707800 791072 708000 791140
rect 707800 791016 707870 791072
rect 707926 791016 708000 791072
rect 707800 790948 708000 791016
rect 707800 790892 707870 790948
rect 707926 790892 708000 790948
rect 707800 790828 708000 790892
rect 699322 790040 699392 790096
rect 699448 790040 699516 790096
rect 699572 790040 699640 790096
rect 699696 790040 699764 790096
rect 699820 790040 699888 790096
rect 699944 790040 700012 790096
rect 700068 790040 700136 790096
rect 700192 790040 700322 790096
rect 699322 789972 700322 790040
rect 699322 789916 699392 789972
rect 699448 789916 699516 789972
rect 699572 789916 699640 789972
rect 699696 789916 699764 789972
rect 699820 789916 699888 789972
rect 699944 789916 700012 789972
rect 700068 789916 700136 789972
rect 700192 789916 700322 789972
rect 699322 789848 700322 789916
rect 699322 789792 699392 789848
rect 699448 789792 699516 789848
rect 699572 789792 699640 789848
rect 699696 789792 699764 789848
rect 699820 789792 699888 789848
rect 699944 789792 700012 789848
rect 700068 789792 700136 789848
rect 700192 789792 700322 789848
rect 699322 789724 700322 789792
rect 699322 789668 699392 789724
rect 699448 789668 699516 789724
rect 699572 789668 699640 789724
rect 699696 789668 699764 789724
rect 699820 789668 699888 789724
rect 699944 789668 700012 789724
rect 700068 789668 700136 789724
rect 700192 789668 700322 789724
rect 699322 789600 700322 789668
rect 699322 789544 699392 789600
rect 699448 789544 699516 789600
rect 699572 789544 699640 789600
rect 699696 789544 699764 789600
rect 699820 789544 699888 789600
rect 699944 789544 700012 789600
rect 700068 789544 700136 789600
rect 700192 789544 700322 789600
rect 699322 789476 700322 789544
rect 699322 789420 699392 789476
rect 699448 789420 699516 789476
rect 699572 789420 699640 789476
rect 699696 789420 699764 789476
rect 699820 789420 699888 789476
rect 699944 789420 700012 789476
rect 700068 789420 700136 789476
rect 700192 789420 700322 789476
rect 699322 789352 700322 789420
rect 699322 789296 699392 789352
rect 699448 789296 699516 789352
rect 699572 789296 699640 789352
rect 699696 789296 699764 789352
rect 699820 789296 699888 789352
rect 699944 789296 700012 789352
rect 700068 789296 700136 789352
rect 700192 789296 700322 789352
rect 699322 789228 700322 789296
rect 699322 789172 699392 789228
rect 699448 789172 699516 789228
rect 699572 789172 699640 789228
rect 699696 789172 699764 789228
rect 699820 789172 699888 789228
rect 699944 789172 700012 789228
rect 700068 789172 700136 789228
rect 700192 789172 700322 789228
rect 699322 789104 700322 789172
rect 699322 789048 699392 789104
rect 699448 789048 699516 789104
rect 699572 789048 699640 789104
rect 699696 789048 699764 789104
rect 699820 789048 699888 789104
rect 699944 789048 700012 789104
rect 700068 789048 700136 789104
rect 700192 789048 700322 789104
rect 699322 788980 700322 789048
rect 699322 788924 699392 788980
rect 699448 788924 699516 788980
rect 699572 788924 699640 788980
rect 699696 788924 699764 788980
rect 699820 788924 699888 788980
rect 699944 788924 700012 788980
rect 700068 788924 700136 788980
rect 700192 788924 700322 788980
rect 699322 788856 700322 788924
rect 699322 788800 699392 788856
rect 699448 788800 699516 788856
rect 699572 788800 699640 788856
rect 699696 788800 699764 788856
rect 699820 788800 699888 788856
rect 699944 788800 700012 788856
rect 700068 788800 700136 788856
rect 700192 788800 700322 788856
rect 699322 788732 700322 788800
rect 699322 788676 699392 788732
rect 699448 788676 699516 788732
rect 699572 788676 699640 788732
rect 699696 788676 699764 788732
rect 699820 788676 699888 788732
rect 699944 788676 700012 788732
rect 700068 788676 700136 788732
rect 700192 788676 700322 788732
rect 699322 788608 700322 788676
rect 699322 788552 699392 788608
rect 699448 788552 699516 788608
rect 699572 788552 699640 788608
rect 699696 788552 699764 788608
rect 699820 788552 699888 788608
rect 699944 788552 700012 788608
rect 700068 788552 700136 788608
rect 700192 788552 700322 788608
rect 699322 788484 700322 788552
rect 699322 788428 699392 788484
rect 699448 788428 699516 788484
rect 699572 788428 699640 788484
rect 699696 788428 699764 788484
rect 699820 788428 699888 788484
rect 699944 788428 700012 788484
rect 700068 788428 700136 788484
rect 700192 788428 700322 788484
rect 699322 788360 700322 788428
rect 699322 788304 699392 788360
rect 699448 788304 699516 788360
rect 699572 788304 699640 788360
rect 699696 788304 699764 788360
rect 699820 788304 699888 788360
rect 699944 788304 700012 788360
rect 700068 788304 700136 788360
rect 700192 788304 700322 788360
rect 699322 788236 700322 788304
rect 699322 788180 699392 788236
rect 699448 788180 699516 788236
rect 699572 788180 699640 788236
rect 699696 788180 699764 788236
rect 699820 788180 699888 788236
rect 699944 788180 700012 788236
rect 700068 788180 700136 788236
rect 700192 788180 700322 788236
rect 699322 787726 700322 788180
rect 707800 790102 708000 790172
rect 707800 790046 707870 790102
rect 707926 790046 708000 790102
rect 707800 789978 708000 790046
rect 707800 789922 707870 789978
rect 707926 789922 708000 789978
rect 707800 789854 708000 789922
rect 707800 789798 707870 789854
rect 707926 789798 708000 789854
rect 707800 789730 708000 789798
rect 707800 789674 707870 789730
rect 707926 789674 708000 789730
rect 707800 789606 708000 789674
rect 707800 789550 707870 789606
rect 707926 789550 708000 789606
rect 707800 789482 708000 789550
rect 707800 789426 707870 789482
rect 707926 789426 708000 789482
rect 707800 789358 708000 789426
rect 707800 789302 707870 789358
rect 707926 789302 708000 789358
rect 707800 789234 708000 789302
rect 707800 789178 707870 789234
rect 707926 789178 708000 789234
rect 707800 789110 708000 789178
rect 707800 789054 707870 789110
rect 707926 789054 708000 789110
rect 707800 788986 708000 789054
rect 707800 788930 707870 788986
rect 707926 788930 708000 788986
rect 707800 788862 708000 788930
rect 707800 788806 707870 788862
rect 707926 788806 708000 788862
rect 707800 788738 708000 788806
rect 707800 788682 707870 788738
rect 707926 788682 708000 788738
rect 707800 788614 708000 788682
rect 707800 788558 707870 788614
rect 707926 788558 708000 788614
rect 707800 788490 708000 788558
rect 707800 788434 707870 788490
rect 707926 788434 708000 788490
rect 707800 788366 708000 788434
rect 707800 788310 707870 788366
rect 707926 788310 708000 788366
rect 707800 788242 708000 788310
rect 707800 788186 707870 788242
rect 707926 788186 708000 788242
rect 707800 788122 708000 788186
rect 699322 787670 699392 787726
rect 699448 787670 699516 787726
rect 699572 787670 699640 787726
rect 699696 787670 699764 787726
rect 699820 787670 699888 787726
rect 699944 787670 700012 787726
rect 700068 787670 700136 787726
rect 700192 787670 700322 787726
rect 699322 787602 700322 787670
rect 699322 787546 699392 787602
rect 699448 787546 699516 787602
rect 699572 787546 699640 787602
rect 699696 787546 699764 787602
rect 699820 787546 699888 787602
rect 699944 787546 700012 787602
rect 700068 787546 700136 787602
rect 700192 787546 700322 787602
rect 699322 787478 700322 787546
rect 699322 787422 699392 787478
rect 699448 787422 699516 787478
rect 699572 787422 699640 787478
rect 699696 787422 699764 787478
rect 699820 787422 699888 787478
rect 699944 787422 700012 787478
rect 700068 787422 700136 787478
rect 700192 787422 700322 787478
rect 699322 787354 700322 787422
rect 699322 787298 699392 787354
rect 699448 787298 699516 787354
rect 699572 787298 699640 787354
rect 699696 787298 699764 787354
rect 699820 787298 699888 787354
rect 699944 787298 700012 787354
rect 700068 787298 700136 787354
rect 700192 787298 700322 787354
rect 699322 787230 700322 787298
rect 699322 787174 699392 787230
rect 699448 787174 699516 787230
rect 699572 787174 699640 787230
rect 699696 787174 699764 787230
rect 699820 787174 699888 787230
rect 699944 787174 700012 787230
rect 700068 787174 700136 787230
rect 700192 787174 700322 787230
rect 699322 787106 700322 787174
rect 699322 787050 699392 787106
rect 699448 787050 699516 787106
rect 699572 787050 699640 787106
rect 699696 787050 699764 787106
rect 699820 787050 699888 787106
rect 699944 787050 700012 787106
rect 700068 787050 700136 787106
rect 700192 787050 700322 787106
rect 699322 786982 700322 787050
rect 699322 786926 699392 786982
rect 699448 786926 699516 786982
rect 699572 786926 699640 786982
rect 699696 786926 699764 786982
rect 699820 786926 699888 786982
rect 699944 786926 700012 786982
rect 700068 786926 700136 786982
rect 700192 786926 700322 786982
rect 699322 786858 700322 786926
rect 699322 786802 699392 786858
rect 699448 786802 699516 786858
rect 699572 786802 699640 786858
rect 699696 786802 699764 786858
rect 699820 786802 699888 786858
rect 699944 786802 700012 786858
rect 700068 786802 700136 786858
rect 700192 786802 700322 786858
rect 699322 786734 700322 786802
rect 699322 786678 699392 786734
rect 699448 786678 699516 786734
rect 699572 786678 699640 786734
rect 699696 786678 699764 786734
rect 699820 786678 699888 786734
rect 699944 786678 700012 786734
rect 700068 786678 700136 786734
rect 700192 786678 700322 786734
rect 699322 786610 700322 786678
rect 699322 786554 699392 786610
rect 699448 786554 699516 786610
rect 699572 786554 699640 786610
rect 699696 786554 699764 786610
rect 699820 786554 699888 786610
rect 699944 786554 700012 786610
rect 700068 786554 700136 786610
rect 700192 786554 700322 786610
rect 699322 786486 700322 786554
rect 699322 786430 699392 786486
rect 699448 786430 699516 786486
rect 699572 786430 699640 786486
rect 699696 786430 699764 786486
rect 699820 786430 699888 786486
rect 699944 786430 700012 786486
rect 700068 786430 700136 786486
rect 700192 786430 700322 786486
rect 699322 786362 700322 786430
rect 699322 786306 699392 786362
rect 699448 786306 699516 786362
rect 699572 786306 699640 786362
rect 699696 786306 699764 786362
rect 699820 786306 699888 786362
rect 699944 786306 700012 786362
rect 700068 786306 700136 786362
rect 700192 786306 700322 786362
rect 699322 786238 700322 786306
rect 699322 786182 699392 786238
rect 699448 786182 699516 786238
rect 699572 786182 699640 786238
rect 699696 786182 699764 786238
rect 699820 786182 699888 786238
rect 699944 786182 700012 786238
rect 700068 786182 700136 786238
rect 700192 786182 700322 786238
rect 699322 786114 700322 786182
rect 699322 786058 699392 786114
rect 699448 786058 699516 786114
rect 699572 786058 699640 786114
rect 699696 786058 699764 786114
rect 699820 786058 699888 786114
rect 699944 786058 700012 786114
rect 700068 786058 700136 786114
rect 700192 786058 700322 786114
rect 699322 785990 700322 786058
rect 699322 785934 699392 785990
rect 699448 785934 699516 785990
rect 699572 785934 699640 785990
rect 699696 785934 699764 785990
rect 699820 785934 699888 785990
rect 699944 785934 700012 785990
rect 700068 785934 700136 785990
rect 700192 785934 700322 785990
rect 699322 785866 700322 785934
rect 699322 785810 699392 785866
rect 699448 785810 699516 785866
rect 699572 785810 699640 785866
rect 699696 785810 699764 785866
rect 699820 785810 699888 785866
rect 699944 785810 700012 785866
rect 700068 785810 700136 785866
rect 700192 785810 700322 785866
rect 699322 785122 700322 785810
rect 707800 787732 708000 787802
rect 707800 787676 707870 787732
rect 707926 787676 708000 787732
rect 707800 787608 708000 787676
rect 707800 787552 707870 787608
rect 707926 787552 708000 787608
rect 707800 787484 708000 787552
rect 707800 787428 707870 787484
rect 707926 787428 708000 787484
rect 707800 787360 708000 787428
rect 707800 787304 707870 787360
rect 707926 787304 708000 787360
rect 707800 787236 708000 787304
rect 707800 787180 707870 787236
rect 707926 787180 708000 787236
rect 707800 787112 708000 787180
rect 707800 787056 707870 787112
rect 707926 787056 708000 787112
rect 707800 786988 708000 787056
rect 707800 786932 707870 786988
rect 707926 786932 708000 786988
rect 707800 786864 708000 786932
rect 707800 786808 707870 786864
rect 707926 786808 708000 786864
rect 707800 786740 708000 786808
rect 707800 786684 707870 786740
rect 707926 786684 708000 786740
rect 707800 786616 708000 786684
rect 707800 786560 707870 786616
rect 707926 786560 708000 786616
rect 707800 786492 708000 786560
rect 707800 786436 707870 786492
rect 707926 786436 708000 786492
rect 707800 786368 708000 786436
rect 707800 786312 707870 786368
rect 707926 786312 708000 786368
rect 707800 786244 708000 786312
rect 707800 786188 707870 786244
rect 707926 786188 708000 786244
rect 707800 786120 708000 786188
rect 707800 786064 707870 786120
rect 707926 786064 708000 786120
rect 707800 785996 708000 786064
rect 707800 785940 707870 785996
rect 707926 785940 708000 785996
rect 707800 785872 708000 785940
rect 707800 785816 707870 785872
rect 707926 785816 708000 785872
rect 707800 785752 708000 785816
rect 699322 785066 699392 785122
rect 699448 785066 699516 785122
rect 699572 785066 699640 785122
rect 699696 785066 699764 785122
rect 699820 785066 699888 785122
rect 699944 785066 700012 785122
rect 700068 785066 700136 785122
rect 700192 785066 700322 785122
rect 699322 784998 700322 785066
rect 699322 784942 699392 784998
rect 699448 784942 699516 784998
rect 699572 784942 699640 784998
rect 699696 784942 699764 784998
rect 699820 784942 699888 784998
rect 699944 784942 700012 784998
rect 700068 784942 700136 784998
rect 700192 784942 700322 784998
rect 699322 784874 700322 784942
rect 699322 784818 699392 784874
rect 699448 784818 699516 784874
rect 699572 784818 699640 784874
rect 699696 784818 699764 784874
rect 699820 784818 699888 784874
rect 699944 784818 700012 784874
rect 700068 784818 700136 784874
rect 700192 784818 700322 784874
rect 699322 784750 700322 784818
rect 699322 784694 699392 784750
rect 699448 784694 699516 784750
rect 699572 784694 699640 784750
rect 699696 784694 699764 784750
rect 699820 784694 699888 784750
rect 699944 784694 700012 784750
rect 700068 784694 700136 784750
rect 700192 784694 700322 784750
rect 699322 784626 700322 784694
rect 699322 784570 699392 784626
rect 699448 784570 699516 784626
rect 699572 784570 699640 784626
rect 699696 784570 699764 784626
rect 699820 784570 699888 784626
rect 699944 784570 700012 784626
rect 700068 784570 700136 784626
rect 700192 784570 700322 784626
rect 699322 784502 700322 784570
rect 699322 784446 699392 784502
rect 699448 784446 699516 784502
rect 699572 784446 699640 784502
rect 699696 784446 699764 784502
rect 699820 784446 699888 784502
rect 699944 784446 700012 784502
rect 700068 784446 700136 784502
rect 700192 784446 700322 784502
rect 699322 784378 700322 784446
rect 699322 784322 699392 784378
rect 699448 784322 699516 784378
rect 699572 784322 699640 784378
rect 699696 784322 699764 784378
rect 699820 784322 699888 784378
rect 699944 784322 700012 784378
rect 700068 784322 700136 784378
rect 700192 784322 700322 784378
rect 699322 784254 700322 784322
rect 699322 784198 699392 784254
rect 699448 784198 699516 784254
rect 699572 784198 699640 784254
rect 699696 784198 699764 784254
rect 699820 784198 699888 784254
rect 699944 784198 700012 784254
rect 700068 784198 700136 784254
rect 700192 784198 700322 784254
rect 699322 784130 700322 784198
rect 699322 784074 699392 784130
rect 699448 784074 699516 784130
rect 699572 784074 699640 784130
rect 699696 784074 699764 784130
rect 699820 784074 699888 784130
rect 699944 784074 700012 784130
rect 700068 784074 700136 784130
rect 700192 784074 700322 784130
rect 699322 784006 700322 784074
rect 699322 783950 699392 784006
rect 699448 783950 699516 784006
rect 699572 783950 699640 784006
rect 699696 783950 699764 784006
rect 699820 783950 699888 784006
rect 699944 783950 700012 784006
rect 700068 783950 700136 784006
rect 700192 783950 700322 784006
rect 699322 783882 700322 783950
rect 699322 783826 699392 783882
rect 699448 783826 699516 783882
rect 699572 783826 699640 783882
rect 699696 783826 699764 783882
rect 699820 783826 699888 783882
rect 699944 783826 700012 783882
rect 700068 783826 700136 783882
rect 700192 783826 700322 783882
rect 699322 783758 700322 783826
rect 699322 783702 699392 783758
rect 699448 783702 699516 783758
rect 699572 783702 699640 783758
rect 699696 783702 699764 783758
rect 699820 783702 699888 783758
rect 699944 783702 700012 783758
rect 700068 783702 700136 783758
rect 700192 783702 700322 783758
rect 699322 783634 700322 783702
rect 699322 783578 699392 783634
rect 699448 783578 699516 783634
rect 699572 783578 699640 783634
rect 699696 783578 699764 783634
rect 699820 783578 699888 783634
rect 699944 783578 700012 783634
rect 700068 783578 700136 783634
rect 700192 783578 700322 783634
rect 699322 783510 700322 783578
rect 699322 783454 699392 783510
rect 699448 783454 699516 783510
rect 699572 783454 699640 783510
rect 699696 783454 699764 783510
rect 699820 783454 699888 783510
rect 699944 783454 700012 783510
rect 700068 783454 700136 783510
rect 700192 783454 700322 783510
rect 699322 783386 700322 783454
rect 699322 783330 699392 783386
rect 699448 783330 699516 783386
rect 699572 783330 699640 783386
rect 699696 783330 699764 783386
rect 699820 783330 699888 783386
rect 699944 783330 700012 783386
rect 700068 783330 700136 783386
rect 700192 783330 700322 783386
rect 699322 770429 700322 783330
rect 707800 785134 708000 785172
rect 707800 785078 707870 785134
rect 707926 785078 708000 785134
rect 707800 785010 708000 785078
rect 707800 784954 707870 785010
rect 707926 784954 708000 785010
rect 707800 784886 708000 784954
rect 707800 784830 707870 784886
rect 707926 784830 708000 784886
rect 707800 784762 708000 784830
rect 707800 784706 707870 784762
rect 707926 784706 708000 784762
rect 707800 784638 708000 784706
rect 707800 784582 707870 784638
rect 707926 784582 708000 784638
rect 707800 784514 708000 784582
rect 707800 784458 707870 784514
rect 707926 784458 708000 784514
rect 707800 784390 708000 784458
rect 707800 784334 707870 784390
rect 707926 784334 708000 784390
rect 707800 784266 708000 784334
rect 707800 784210 707870 784266
rect 707926 784210 708000 784266
rect 707800 784142 708000 784210
rect 707800 784086 707870 784142
rect 707926 784086 708000 784142
rect 707800 784018 708000 784086
rect 707800 783962 707870 784018
rect 707926 783962 708000 784018
rect 707800 783894 708000 783962
rect 707800 783838 707870 783894
rect 707926 783838 708000 783894
rect 707800 783770 708000 783838
rect 707800 783714 707870 783770
rect 707926 783714 708000 783770
rect 707800 783646 708000 783714
rect 707800 783590 707870 783646
rect 707926 783590 708000 783646
rect 707800 783522 708000 783590
rect 707800 783466 707870 783522
rect 707926 783466 708000 783522
rect 707800 783398 708000 783466
rect 707800 783342 707870 783398
rect 707926 783342 708000 783398
rect 707800 783272 708000 783342
rect 699322 770373 699544 770429
rect 699600 770373 699844 770429
rect 699900 770373 700144 770429
rect 700200 770373 700322 770429
rect 699322 770229 700322 770373
rect 699322 770173 699544 770229
rect 699600 770173 699844 770229
rect 699900 770173 700144 770229
rect 700200 770173 700322 770229
rect 699322 753954 700322 770173
rect 699322 753898 699444 753954
rect 699500 753898 699744 753954
rect 699800 753898 700044 753954
rect 700100 753898 700322 753954
rect 699322 746954 700322 753898
rect 699322 746898 699444 746954
rect 699500 746898 699744 746954
rect 699800 746898 700044 746954
rect 700100 746898 700322 746954
rect 699322 739954 700322 746898
rect 699322 739898 699444 739954
rect 699500 739898 699744 739954
rect 699800 739898 700044 739954
rect 700100 739898 700322 739954
rect 699322 734429 700322 739898
rect 699322 734373 699544 734429
rect 699600 734373 699844 734429
rect 699900 734373 700144 734429
rect 700200 734373 700322 734429
rect 699322 734229 700322 734373
rect 699322 734173 699544 734229
rect 699600 734173 699844 734229
rect 699900 734173 700144 734229
rect 700200 734173 700322 734229
rect 699322 720423 700322 734173
rect 699322 720367 699497 720423
rect 699553 720367 699797 720423
rect 699853 720367 700097 720423
rect 700153 720367 700322 720423
rect 699322 710954 700322 720367
rect 699322 710898 699444 710954
rect 699500 710898 699744 710954
rect 699800 710898 700044 710954
rect 700100 710898 700322 710954
rect 699322 703954 700322 710898
rect 699322 703898 699444 703954
rect 699500 703898 699744 703954
rect 699800 703898 700044 703954
rect 700100 703898 700322 703954
rect 699322 698429 700322 703898
rect 699322 698373 699544 698429
rect 699600 698373 699844 698429
rect 699900 698373 700144 698429
rect 700200 698373 700322 698429
rect 699322 698229 700322 698373
rect 699322 698173 699544 698229
rect 699600 698173 699844 698229
rect 699900 698173 700144 698229
rect 700200 698173 700322 698229
rect 699322 696954 700322 698173
rect 699322 696898 699444 696954
rect 699500 696898 699744 696954
rect 699800 696898 700044 696954
rect 700100 696898 700322 696954
rect 699322 677423 700322 696898
rect 699322 677367 699497 677423
rect 699553 677367 699797 677423
rect 699853 677367 700097 677423
rect 700153 677367 700322 677423
rect 699322 667954 700322 677367
rect 699322 667898 699444 667954
rect 699500 667898 699744 667954
rect 699800 667898 700044 667954
rect 700100 667898 700322 667954
rect 699322 662429 700322 667898
rect 699322 662373 699544 662429
rect 699600 662373 699844 662429
rect 699900 662373 700144 662429
rect 700200 662373 700322 662429
rect 699322 662229 700322 662373
rect 699322 662173 699544 662229
rect 699600 662173 699844 662229
rect 699900 662173 700144 662229
rect 700200 662173 700322 662229
rect 699322 660954 700322 662173
rect 699322 660898 699444 660954
rect 699500 660898 699744 660954
rect 699800 660898 700044 660954
rect 700100 660898 700322 660954
rect 699322 653954 700322 660898
rect 699322 653898 699444 653954
rect 699500 653898 699744 653954
rect 699800 653898 700044 653954
rect 700100 653898 700322 653954
rect 699322 634423 700322 653898
rect 699322 634367 699497 634423
rect 699553 634367 699797 634423
rect 699853 634367 700097 634423
rect 700153 634367 700322 634423
rect 699322 626429 700322 634367
rect 699322 626373 699544 626429
rect 699600 626373 699844 626429
rect 699900 626373 700144 626429
rect 700200 626373 700322 626429
rect 699322 626229 700322 626373
rect 699322 626173 699544 626229
rect 699600 626173 699844 626229
rect 699900 626173 700144 626229
rect 700200 626173 700322 626229
rect 699322 624954 700322 626173
rect 699322 624898 699444 624954
rect 699500 624898 699744 624954
rect 699800 624898 700044 624954
rect 700100 624898 700322 624954
rect 699322 617954 700322 624898
rect 699322 617898 699444 617954
rect 699500 617898 699744 617954
rect 699800 617898 700044 617954
rect 700100 617898 700322 617954
rect 699322 610954 700322 617898
rect 699322 610898 699444 610954
rect 699500 610898 699744 610954
rect 699800 610898 700044 610954
rect 700100 610898 700322 610954
rect 699322 591423 700322 610898
rect 699322 591367 699497 591423
rect 699553 591367 699797 591423
rect 699853 591367 700097 591423
rect 700153 591367 700322 591423
rect 699322 590429 700322 591367
rect 699322 590373 699544 590429
rect 699600 590373 699844 590429
rect 699900 590373 700144 590429
rect 700200 590373 700322 590429
rect 699322 590229 700322 590373
rect 699322 590173 699544 590229
rect 699600 590173 699844 590229
rect 699900 590173 700144 590229
rect 700200 590173 700322 590229
rect 699322 581954 700322 590173
rect 699322 581898 699444 581954
rect 699500 581898 699744 581954
rect 699800 581898 700044 581954
rect 700100 581898 700322 581954
rect 699322 574954 700322 581898
rect 699322 574898 699444 574954
rect 699500 574898 699744 574954
rect 699800 574898 700044 574954
rect 700100 574898 700322 574954
rect 699322 567954 700322 574898
rect 699322 567898 699444 567954
rect 699500 567898 699744 567954
rect 699800 567898 700044 567954
rect 700100 567898 700322 567954
rect 699322 554429 700322 567898
rect 699322 554373 699544 554429
rect 699600 554373 699844 554429
rect 699900 554373 700144 554429
rect 700200 554373 700322 554429
rect 699322 554229 700322 554373
rect 699322 554173 699544 554229
rect 699600 554173 699844 554229
rect 699900 554173 700144 554229
rect 700200 554173 700322 554229
rect 699322 548423 700322 554173
rect 699322 548367 699497 548423
rect 699553 548367 699797 548423
rect 699853 548367 700097 548423
rect 700153 548367 700322 548423
rect 699322 538954 700322 548367
rect 699322 538898 699444 538954
rect 699500 538898 699744 538954
rect 699800 538898 700044 538954
rect 700100 538898 700322 538954
rect 699322 531954 700322 538898
rect 699322 531898 699444 531954
rect 699500 531898 699744 531954
rect 699800 531898 700044 531954
rect 700100 531898 700322 531954
rect 699322 524954 700322 531898
rect 699322 524898 699444 524954
rect 699500 524898 699744 524954
rect 699800 524898 700044 524954
rect 700100 524898 700322 524954
rect 699322 518429 700322 524898
rect 699322 518373 699544 518429
rect 699600 518373 699844 518429
rect 699900 518373 700144 518429
rect 700200 518373 700322 518429
rect 699322 518229 700322 518373
rect 699322 518173 699544 518229
rect 699600 518173 699844 518229
rect 699900 518173 700144 518229
rect 700200 518173 700322 518229
rect 699322 505423 700322 518173
rect 699322 505367 699497 505423
rect 699553 505367 699797 505423
rect 699853 505367 700097 505423
rect 700153 505367 700322 505423
rect 699322 496652 700322 505367
rect 699322 496596 699392 496652
rect 699448 496596 699516 496652
rect 699572 496596 699640 496652
rect 699696 496596 699764 496652
rect 699820 496596 699888 496652
rect 699944 496596 700012 496652
rect 700068 496596 700136 496652
rect 700192 496596 700322 496652
rect 699322 496528 700322 496596
rect 699322 496472 699392 496528
rect 699448 496472 699516 496528
rect 699572 496472 699640 496528
rect 699696 496472 699764 496528
rect 699820 496472 699888 496528
rect 699944 496472 700012 496528
rect 700068 496472 700136 496528
rect 700192 496472 700322 496528
rect 699322 496404 700322 496472
rect 699322 496348 699392 496404
rect 699448 496348 699516 496404
rect 699572 496348 699640 496404
rect 699696 496348 699764 496404
rect 699820 496348 699888 496404
rect 699944 496348 700012 496404
rect 700068 496348 700136 496404
rect 700192 496348 700322 496404
rect 699322 496280 700322 496348
rect 699322 496224 699392 496280
rect 699448 496224 699516 496280
rect 699572 496224 699640 496280
rect 699696 496224 699764 496280
rect 699820 496224 699888 496280
rect 699944 496224 700012 496280
rect 700068 496224 700136 496280
rect 700192 496224 700322 496280
rect 699322 496156 700322 496224
rect 699322 496100 699392 496156
rect 699448 496100 699516 496156
rect 699572 496100 699640 496156
rect 699696 496100 699764 496156
rect 699820 496100 699888 496156
rect 699944 496100 700012 496156
rect 700068 496100 700136 496156
rect 700192 496100 700322 496156
rect 699322 496032 700322 496100
rect 699322 495976 699392 496032
rect 699448 495976 699516 496032
rect 699572 495976 699640 496032
rect 699696 495976 699764 496032
rect 699820 495976 699888 496032
rect 699944 495976 700012 496032
rect 700068 495976 700136 496032
rect 700192 495976 700322 496032
rect 699322 495908 700322 495976
rect 699322 495852 699392 495908
rect 699448 495852 699516 495908
rect 699572 495852 699640 495908
rect 699696 495852 699764 495908
rect 699820 495852 699888 495908
rect 699944 495852 700012 495908
rect 700068 495852 700136 495908
rect 700192 495852 700322 495908
rect 699322 495784 700322 495852
rect 699322 495728 699392 495784
rect 699448 495728 699516 495784
rect 699572 495728 699640 495784
rect 699696 495728 699764 495784
rect 699820 495728 699888 495784
rect 699944 495728 700012 495784
rect 700068 495728 700136 495784
rect 700192 495728 700322 495784
rect 699322 495660 700322 495728
rect 699322 495604 699392 495660
rect 699448 495604 699516 495660
rect 699572 495604 699640 495660
rect 699696 495604 699764 495660
rect 699820 495604 699888 495660
rect 699944 495604 700012 495660
rect 700068 495604 700136 495660
rect 700192 495604 700322 495660
rect 699322 495536 700322 495604
rect 699322 495480 699392 495536
rect 699448 495480 699516 495536
rect 699572 495480 699640 495536
rect 699696 495480 699764 495536
rect 699820 495480 699888 495536
rect 699944 495480 700012 495536
rect 700068 495480 700136 495536
rect 700192 495480 700322 495536
rect 699322 495412 700322 495480
rect 699322 495356 699392 495412
rect 699448 495356 699516 495412
rect 699572 495356 699640 495412
rect 699696 495356 699764 495412
rect 699820 495356 699888 495412
rect 699944 495356 700012 495412
rect 700068 495356 700136 495412
rect 700192 495356 700322 495412
rect 699322 495288 700322 495356
rect 699322 495232 699392 495288
rect 699448 495232 699516 495288
rect 699572 495232 699640 495288
rect 699696 495232 699764 495288
rect 699820 495232 699888 495288
rect 699944 495232 700012 495288
rect 700068 495232 700136 495288
rect 700192 495232 700322 495288
rect 699322 495164 700322 495232
rect 699322 495108 699392 495164
rect 699448 495108 699516 495164
rect 699572 495108 699640 495164
rect 699696 495108 699764 495164
rect 699820 495108 699888 495164
rect 699944 495108 700012 495164
rect 700068 495108 700136 495164
rect 700192 495108 700322 495164
rect 699322 495040 700322 495108
rect 699322 494984 699392 495040
rect 699448 494984 699516 495040
rect 699572 494984 699640 495040
rect 699696 494984 699764 495040
rect 699820 494984 699888 495040
rect 699944 494984 700012 495040
rect 700068 494984 700136 495040
rect 700192 494984 700322 495040
rect 699322 494916 700322 494984
rect 699322 494860 699392 494916
rect 699448 494860 699516 494916
rect 699572 494860 699640 494916
rect 699696 494860 699764 494916
rect 699820 494860 699888 494916
rect 699944 494860 700012 494916
rect 700068 494860 700136 494916
rect 700192 494860 700322 494916
rect 699322 494172 700322 494860
rect 707800 496658 708000 496728
rect 707800 496602 707870 496658
rect 707926 496602 708000 496658
rect 707800 496534 708000 496602
rect 707800 496478 707870 496534
rect 707926 496478 708000 496534
rect 707800 496410 708000 496478
rect 707800 496354 707870 496410
rect 707926 496354 708000 496410
rect 707800 496286 708000 496354
rect 707800 496230 707870 496286
rect 707926 496230 708000 496286
rect 707800 496162 708000 496230
rect 707800 496106 707870 496162
rect 707926 496106 708000 496162
rect 707800 496038 708000 496106
rect 707800 495982 707870 496038
rect 707926 495982 708000 496038
rect 707800 495914 708000 495982
rect 707800 495858 707870 495914
rect 707926 495858 708000 495914
rect 707800 495790 708000 495858
rect 707800 495734 707870 495790
rect 707926 495734 708000 495790
rect 707800 495666 708000 495734
rect 707800 495610 707870 495666
rect 707926 495610 708000 495666
rect 707800 495542 708000 495610
rect 707800 495486 707870 495542
rect 707926 495486 708000 495542
rect 707800 495418 708000 495486
rect 707800 495362 707870 495418
rect 707926 495362 708000 495418
rect 707800 495294 708000 495362
rect 707800 495238 707870 495294
rect 707926 495238 708000 495294
rect 707800 495170 708000 495238
rect 707800 495114 707870 495170
rect 707926 495114 708000 495170
rect 707800 495046 708000 495114
rect 707800 494990 707870 495046
rect 707926 494990 708000 495046
rect 707800 494922 708000 494990
rect 707800 494866 707870 494922
rect 707926 494866 708000 494922
rect 707800 494828 708000 494866
rect 699322 494116 699392 494172
rect 699448 494116 699516 494172
rect 699572 494116 699640 494172
rect 699696 494116 699764 494172
rect 699820 494116 699888 494172
rect 699944 494116 700012 494172
rect 700068 494116 700136 494172
rect 700192 494116 700322 494172
rect 699322 494048 700322 494116
rect 699322 493992 699392 494048
rect 699448 493992 699516 494048
rect 699572 493992 699640 494048
rect 699696 493992 699764 494048
rect 699820 493992 699888 494048
rect 699944 493992 700012 494048
rect 700068 493992 700136 494048
rect 700192 493992 700322 494048
rect 699322 493924 700322 493992
rect 699322 493868 699392 493924
rect 699448 493868 699516 493924
rect 699572 493868 699640 493924
rect 699696 493868 699764 493924
rect 699820 493868 699888 493924
rect 699944 493868 700012 493924
rect 700068 493868 700136 493924
rect 700192 493868 700322 493924
rect 699322 493800 700322 493868
rect 699322 493744 699392 493800
rect 699448 493744 699516 493800
rect 699572 493744 699640 493800
rect 699696 493744 699764 493800
rect 699820 493744 699888 493800
rect 699944 493744 700012 493800
rect 700068 493744 700136 493800
rect 700192 493744 700322 493800
rect 699322 493676 700322 493744
rect 699322 493620 699392 493676
rect 699448 493620 699516 493676
rect 699572 493620 699640 493676
rect 699696 493620 699764 493676
rect 699820 493620 699888 493676
rect 699944 493620 700012 493676
rect 700068 493620 700136 493676
rect 700192 493620 700322 493676
rect 699322 493552 700322 493620
rect 699322 493496 699392 493552
rect 699448 493496 699516 493552
rect 699572 493496 699640 493552
rect 699696 493496 699764 493552
rect 699820 493496 699888 493552
rect 699944 493496 700012 493552
rect 700068 493496 700136 493552
rect 700192 493496 700322 493552
rect 699322 493428 700322 493496
rect 699322 493372 699392 493428
rect 699448 493372 699516 493428
rect 699572 493372 699640 493428
rect 699696 493372 699764 493428
rect 699820 493372 699888 493428
rect 699944 493372 700012 493428
rect 700068 493372 700136 493428
rect 700192 493372 700322 493428
rect 699322 493304 700322 493372
rect 699322 493248 699392 493304
rect 699448 493248 699516 493304
rect 699572 493248 699640 493304
rect 699696 493248 699764 493304
rect 699820 493248 699888 493304
rect 699944 493248 700012 493304
rect 700068 493248 700136 493304
rect 700192 493248 700322 493304
rect 699322 493180 700322 493248
rect 699322 493124 699392 493180
rect 699448 493124 699516 493180
rect 699572 493124 699640 493180
rect 699696 493124 699764 493180
rect 699820 493124 699888 493180
rect 699944 493124 700012 493180
rect 700068 493124 700136 493180
rect 700192 493124 700322 493180
rect 699322 493056 700322 493124
rect 699322 493000 699392 493056
rect 699448 493000 699516 493056
rect 699572 493000 699640 493056
rect 699696 493000 699764 493056
rect 699820 493000 699888 493056
rect 699944 493000 700012 493056
rect 700068 493000 700136 493056
rect 700192 493000 700322 493056
rect 699322 492932 700322 493000
rect 699322 492876 699392 492932
rect 699448 492876 699516 492932
rect 699572 492876 699640 492932
rect 699696 492876 699764 492932
rect 699820 492876 699888 492932
rect 699944 492876 700012 492932
rect 700068 492876 700136 492932
rect 700192 492876 700322 492932
rect 699322 492808 700322 492876
rect 699322 492752 699392 492808
rect 699448 492752 699516 492808
rect 699572 492752 699640 492808
rect 699696 492752 699764 492808
rect 699820 492752 699888 492808
rect 699944 492752 700012 492808
rect 700068 492752 700136 492808
rect 700192 492752 700322 492808
rect 699322 492684 700322 492752
rect 699322 492628 699392 492684
rect 699448 492628 699516 492684
rect 699572 492628 699640 492684
rect 699696 492628 699764 492684
rect 699820 492628 699888 492684
rect 699944 492628 700012 492684
rect 700068 492628 700136 492684
rect 700192 492628 700322 492684
rect 699322 492560 700322 492628
rect 699322 492504 699392 492560
rect 699448 492504 699516 492560
rect 699572 492504 699640 492560
rect 699696 492504 699764 492560
rect 699820 492504 699888 492560
rect 699944 492504 700012 492560
rect 700068 492504 700136 492560
rect 700192 492504 700322 492560
rect 699322 492436 700322 492504
rect 699322 492380 699392 492436
rect 699448 492380 699516 492436
rect 699572 492380 699640 492436
rect 699696 492380 699764 492436
rect 699820 492380 699888 492436
rect 699944 492380 700012 492436
rect 700068 492380 700136 492436
rect 700192 492380 700322 492436
rect 699322 492312 700322 492380
rect 699322 492256 699392 492312
rect 699448 492256 699516 492312
rect 699572 492256 699640 492312
rect 699696 492256 699764 492312
rect 699820 492256 699888 492312
rect 699944 492256 700012 492312
rect 700068 492256 700136 492312
rect 700192 492256 700322 492312
rect 699322 491802 700322 492256
rect 707800 494178 708000 494248
rect 707800 494122 707870 494178
rect 707926 494122 708000 494178
rect 707800 494054 708000 494122
rect 707800 493998 707870 494054
rect 707926 493998 708000 494054
rect 707800 493930 708000 493998
rect 707800 493874 707870 493930
rect 707926 493874 708000 493930
rect 707800 493806 708000 493874
rect 707800 493750 707870 493806
rect 707926 493750 708000 493806
rect 707800 493682 708000 493750
rect 707800 493626 707870 493682
rect 707926 493626 708000 493682
rect 707800 493558 708000 493626
rect 707800 493502 707870 493558
rect 707926 493502 708000 493558
rect 707800 493434 708000 493502
rect 707800 493378 707870 493434
rect 707926 493378 708000 493434
rect 707800 493310 708000 493378
rect 707800 493254 707870 493310
rect 707926 493254 708000 493310
rect 707800 493186 708000 493254
rect 707800 493130 707870 493186
rect 707926 493130 708000 493186
rect 707800 493062 708000 493130
rect 707800 493006 707870 493062
rect 707926 493006 708000 493062
rect 707800 492938 708000 493006
rect 707800 492882 707870 492938
rect 707926 492882 708000 492938
rect 707800 492814 708000 492882
rect 707800 492758 707870 492814
rect 707926 492758 708000 492814
rect 707800 492690 708000 492758
rect 707800 492634 707870 492690
rect 707926 492634 708000 492690
rect 707800 492566 708000 492634
rect 707800 492510 707870 492566
rect 707926 492510 708000 492566
rect 707800 492442 708000 492510
rect 707800 492386 707870 492442
rect 707926 492386 708000 492442
rect 707800 492318 708000 492386
rect 707800 492262 707870 492318
rect 707926 492262 708000 492318
rect 707800 492198 708000 492262
rect 699322 491746 699392 491802
rect 699448 491746 699516 491802
rect 699572 491746 699640 491802
rect 699696 491746 699764 491802
rect 699820 491746 699888 491802
rect 699944 491746 700012 491802
rect 700068 491746 700136 491802
rect 700192 491746 700322 491802
rect 699322 491678 700322 491746
rect 699322 491622 699392 491678
rect 699448 491622 699516 491678
rect 699572 491622 699640 491678
rect 699696 491622 699764 491678
rect 699820 491622 699888 491678
rect 699944 491622 700012 491678
rect 700068 491622 700136 491678
rect 700192 491622 700322 491678
rect 699322 491554 700322 491622
rect 699322 491498 699392 491554
rect 699448 491498 699516 491554
rect 699572 491498 699640 491554
rect 699696 491498 699764 491554
rect 699820 491498 699888 491554
rect 699944 491498 700012 491554
rect 700068 491498 700136 491554
rect 700192 491498 700322 491554
rect 699322 491430 700322 491498
rect 699322 491374 699392 491430
rect 699448 491374 699516 491430
rect 699572 491374 699640 491430
rect 699696 491374 699764 491430
rect 699820 491374 699888 491430
rect 699944 491374 700012 491430
rect 700068 491374 700136 491430
rect 700192 491374 700322 491430
rect 699322 491306 700322 491374
rect 699322 491250 699392 491306
rect 699448 491250 699516 491306
rect 699572 491250 699640 491306
rect 699696 491250 699764 491306
rect 699820 491250 699888 491306
rect 699944 491250 700012 491306
rect 700068 491250 700136 491306
rect 700192 491250 700322 491306
rect 699322 491182 700322 491250
rect 699322 491126 699392 491182
rect 699448 491126 699516 491182
rect 699572 491126 699640 491182
rect 699696 491126 699764 491182
rect 699820 491126 699888 491182
rect 699944 491126 700012 491182
rect 700068 491126 700136 491182
rect 700192 491126 700322 491182
rect 699322 491058 700322 491126
rect 699322 491002 699392 491058
rect 699448 491002 699516 491058
rect 699572 491002 699640 491058
rect 699696 491002 699764 491058
rect 699820 491002 699888 491058
rect 699944 491002 700012 491058
rect 700068 491002 700136 491058
rect 700192 491002 700322 491058
rect 699322 490934 700322 491002
rect 699322 490878 699392 490934
rect 699448 490878 699516 490934
rect 699572 490878 699640 490934
rect 699696 490878 699764 490934
rect 699820 490878 699888 490934
rect 699944 490878 700012 490934
rect 700068 490878 700136 490934
rect 700192 490878 700322 490934
rect 699322 490810 700322 490878
rect 699322 490754 699392 490810
rect 699448 490754 699516 490810
rect 699572 490754 699640 490810
rect 699696 490754 699764 490810
rect 699820 490754 699888 490810
rect 699944 490754 700012 490810
rect 700068 490754 700136 490810
rect 700192 490754 700322 490810
rect 699322 490686 700322 490754
rect 699322 490630 699392 490686
rect 699448 490630 699516 490686
rect 699572 490630 699640 490686
rect 699696 490630 699764 490686
rect 699820 490630 699888 490686
rect 699944 490630 700012 490686
rect 700068 490630 700136 490686
rect 700192 490630 700322 490686
rect 699322 490562 700322 490630
rect 699322 490506 699392 490562
rect 699448 490506 699516 490562
rect 699572 490506 699640 490562
rect 699696 490506 699764 490562
rect 699820 490506 699888 490562
rect 699944 490506 700012 490562
rect 700068 490506 700136 490562
rect 700192 490506 700322 490562
rect 699322 490438 700322 490506
rect 699322 490382 699392 490438
rect 699448 490382 699516 490438
rect 699572 490382 699640 490438
rect 699696 490382 699764 490438
rect 699820 490382 699888 490438
rect 699944 490382 700012 490438
rect 700068 490382 700136 490438
rect 700192 490382 700322 490438
rect 699322 490314 700322 490382
rect 699322 490258 699392 490314
rect 699448 490258 699516 490314
rect 699572 490258 699640 490314
rect 699696 490258 699764 490314
rect 699820 490258 699888 490314
rect 699944 490258 700012 490314
rect 700068 490258 700136 490314
rect 700192 490258 700322 490314
rect 699322 490190 700322 490258
rect 699322 490134 699392 490190
rect 699448 490134 699516 490190
rect 699572 490134 699640 490190
rect 699696 490134 699764 490190
rect 699820 490134 699888 490190
rect 699944 490134 700012 490190
rect 700068 490134 700136 490190
rect 700192 490134 700322 490190
rect 699322 490066 700322 490134
rect 699322 490010 699392 490066
rect 699448 490010 699516 490066
rect 699572 490010 699640 490066
rect 699696 490010 699764 490066
rect 699820 490010 699888 490066
rect 699944 490010 700012 490066
rect 700068 490010 700136 490066
rect 700192 490010 700322 490066
rect 699322 489942 700322 490010
rect 699322 489886 699392 489942
rect 699448 489886 699516 489942
rect 699572 489886 699640 489942
rect 699696 489886 699764 489942
rect 699820 489886 699888 489942
rect 699944 489886 700012 489942
rect 700068 489886 700136 489942
rect 700192 489886 700322 489942
rect 699322 489096 700322 489886
rect 707800 491808 708000 491878
rect 707800 491752 707870 491808
rect 707926 491752 708000 491808
rect 707800 491684 708000 491752
rect 707800 491628 707870 491684
rect 707926 491628 708000 491684
rect 707800 491560 708000 491628
rect 707800 491504 707870 491560
rect 707926 491504 708000 491560
rect 707800 491436 708000 491504
rect 707800 491380 707870 491436
rect 707926 491380 708000 491436
rect 707800 491312 708000 491380
rect 707800 491256 707870 491312
rect 707926 491256 708000 491312
rect 707800 491188 708000 491256
rect 707800 491132 707870 491188
rect 707926 491132 708000 491188
rect 707800 491064 708000 491132
rect 707800 491008 707870 491064
rect 707926 491008 708000 491064
rect 707800 490940 708000 491008
rect 707800 490884 707870 490940
rect 707926 490884 708000 490940
rect 707800 490816 708000 490884
rect 707800 490760 707870 490816
rect 707926 490760 708000 490816
rect 707800 490692 708000 490760
rect 707800 490636 707870 490692
rect 707926 490636 708000 490692
rect 707800 490568 708000 490636
rect 707800 490512 707870 490568
rect 707926 490512 708000 490568
rect 707800 490444 708000 490512
rect 707800 490388 707870 490444
rect 707926 490388 708000 490444
rect 707800 490320 708000 490388
rect 707800 490264 707870 490320
rect 707926 490264 708000 490320
rect 707800 490196 708000 490264
rect 707800 490140 707870 490196
rect 707926 490140 708000 490196
rect 707800 490072 708000 490140
rect 707800 490016 707870 490072
rect 707926 490016 708000 490072
rect 707800 489948 708000 490016
rect 707800 489892 707870 489948
rect 707926 489892 708000 489948
rect 707800 489828 708000 489892
rect 699322 489040 699392 489096
rect 699448 489040 699516 489096
rect 699572 489040 699640 489096
rect 699696 489040 699764 489096
rect 699820 489040 699888 489096
rect 699944 489040 700012 489096
rect 700068 489040 700136 489096
rect 700192 489040 700322 489096
rect 699322 488972 700322 489040
rect 699322 488916 699392 488972
rect 699448 488916 699516 488972
rect 699572 488916 699640 488972
rect 699696 488916 699764 488972
rect 699820 488916 699888 488972
rect 699944 488916 700012 488972
rect 700068 488916 700136 488972
rect 700192 488916 700322 488972
rect 699322 488848 700322 488916
rect 699322 488792 699392 488848
rect 699448 488792 699516 488848
rect 699572 488792 699640 488848
rect 699696 488792 699764 488848
rect 699820 488792 699888 488848
rect 699944 488792 700012 488848
rect 700068 488792 700136 488848
rect 700192 488792 700322 488848
rect 699322 488724 700322 488792
rect 699322 488668 699392 488724
rect 699448 488668 699516 488724
rect 699572 488668 699640 488724
rect 699696 488668 699764 488724
rect 699820 488668 699888 488724
rect 699944 488668 700012 488724
rect 700068 488668 700136 488724
rect 700192 488668 700322 488724
rect 699322 488600 700322 488668
rect 699322 488544 699392 488600
rect 699448 488544 699516 488600
rect 699572 488544 699640 488600
rect 699696 488544 699764 488600
rect 699820 488544 699888 488600
rect 699944 488544 700012 488600
rect 700068 488544 700136 488600
rect 700192 488544 700322 488600
rect 699322 488476 700322 488544
rect 699322 488420 699392 488476
rect 699448 488420 699516 488476
rect 699572 488420 699640 488476
rect 699696 488420 699764 488476
rect 699820 488420 699888 488476
rect 699944 488420 700012 488476
rect 700068 488420 700136 488476
rect 700192 488420 700322 488476
rect 699322 488352 700322 488420
rect 699322 488296 699392 488352
rect 699448 488296 699516 488352
rect 699572 488296 699640 488352
rect 699696 488296 699764 488352
rect 699820 488296 699888 488352
rect 699944 488296 700012 488352
rect 700068 488296 700136 488352
rect 700192 488296 700322 488352
rect 699322 488228 700322 488296
rect 699322 488172 699392 488228
rect 699448 488172 699516 488228
rect 699572 488172 699640 488228
rect 699696 488172 699764 488228
rect 699820 488172 699888 488228
rect 699944 488172 700012 488228
rect 700068 488172 700136 488228
rect 700192 488172 700322 488228
rect 699322 488104 700322 488172
rect 699322 488048 699392 488104
rect 699448 488048 699516 488104
rect 699572 488048 699640 488104
rect 699696 488048 699764 488104
rect 699820 488048 699888 488104
rect 699944 488048 700012 488104
rect 700068 488048 700136 488104
rect 700192 488048 700322 488104
rect 699322 487980 700322 488048
rect 699322 487924 699392 487980
rect 699448 487924 699516 487980
rect 699572 487924 699640 487980
rect 699696 487924 699764 487980
rect 699820 487924 699888 487980
rect 699944 487924 700012 487980
rect 700068 487924 700136 487980
rect 700192 487924 700322 487980
rect 699322 487856 700322 487924
rect 699322 487800 699392 487856
rect 699448 487800 699516 487856
rect 699572 487800 699640 487856
rect 699696 487800 699764 487856
rect 699820 487800 699888 487856
rect 699944 487800 700012 487856
rect 700068 487800 700136 487856
rect 700192 487800 700322 487856
rect 699322 487732 700322 487800
rect 699322 487676 699392 487732
rect 699448 487676 699516 487732
rect 699572 487676 699640 487732
rect 699696 487676 699764 487732
rect 699820 487676 699888 487732
rect 699944 487676 700012 487732
rect 700068 487676 700136 487732
rect 700192 487676 700322 487732
rect 699322 487608 700322 487676
rect 699322 487552 699392 487608
rect 699448 487552 699516 487608
rect 699572 487552 699640 487608
rect 699696 487552 699764 487608
rect 699820 487552 699888 487608
rect 699944 487552 700012 487608
rect 700068 487552 700136 487608
rect 700192 487552 700322 487608
rect 699322 487484 700322 487552
rect 699322 487428 699392 487484
rect 699448 487428 699516 487484
rect 699572 487428 699640 487484
rect 699696 487428 699764 487484
rect 699820 487428 699888 487484
rect 699944 487428 700012 487484
rect 700068 487428 700136 487484
rect 700192 487428 700322 487484
rect 699322 487360 700322 487428
rect 699322 487304 699392 487360
rect 699448 487304 699516 487360
rect 699572 487304 699640 487360
rect 699696 487304 699764 487360
rect 699820 487304 699888 487360
rect 699944 487304 700012 487360
rect 700068 487304 700136 487360
rect 700192 487304 700322 487360
rect 699322 487236 700322 487304
rect 699322 487180 699392 487236
rect 699448 487180 699516 487236
rect 699572 487180 699640 487236
rect 699696 487180 699764 487236
rect 699820 487180 699888 487236
rect 699944 487180 700012 487236
rect 700068 487180 700136 487236
rect 700192 487180 700322 487236
rect 699322 486726 700322 487180
rect 707800 489102 708000 489172
rect 707800 489046 707870 489102
rect 707926 489046 708000 489102
rect 707800 488978 708000 489046
rect 707800 488922 707870 488978
rect 707926 488922 708000 488978
rect 707800 488854 708000 488922
rect 707800 488798 707870 488854
rect 707926 488798 708000 488854
rect 707800 488730 708000 488798
rect 707800 488674 707870 488730
rect 707926 488674 708000 488730
rect 707800 488606 708000 488674
rect 707800 488550 707870 488606
rect 707926 488550 708000 488606
rect 707800 488482 708000 488550
rect 707800 488426 707870 488482
rect 707926 488426 708000 488482
rect 707800 488358 708000 488426
rect 707800 488302 707870 488358
rect 707926 488302 708000 488358
rect 707800 488234 708000 488302
rect 707800 488178 707870 488234
rect 707926 488178 708000 488234
rect 707800 488110 708000 488178
rect 707800 488054 707870 488110
rect 707926 488054 708000 488110
rect 707800 487986 708000 488054
rect 707800 487930 707870 487986
rect 707926 487930 708000 487986
rect 707800 487862 708000 487930
rect 707800 487806 707870 487862
rect 707926 487806 708000 487862
rect 707800 487738 708000 487806
rect 707800 487682 707870 487738
rect 707926 487682 708000 487738
rect 707800 487614 708000 487682
rect 707800 487558 707870 487614
rect 707926 487558 708000 487614
rect 707800 487490 708000 487558
rect 707800 487434 707870 487490
rect 707926 487434 708000 487490
rect 707800 487366 708000 487434
rect 707800 487310 707870 487366
rect 707926 487310 708000 487366
rect 707800 487242 708000 487310
rect 707800 487186 707870 487242
rect 707926 487186 708000 487242
rect 707800 487122 708000 487186
rect 699322 486670 699392 486726
rect 699448 486670 699516 486726
rect 699572 486670 699640 486726
rect 699696 486670 699764 486726
rect 699820 486670 699888 486726
rect 699944 486670 700012 486726
rect 700068 486670 700136 486726
rect 700192 486670 700322 486726
rect 699322 486602 700322 486670
rect 699322 486546 699392 486602
rect 699448 486546 699516 486602
rect 699572 486546 699640 486602
rect 699696 486546 699764 486602
rect 699820 486546 699888 486602
rect 699944 486546 700012 486602
rect 700068 486546 700136 486602
rect 700192 486546 700322 486602
rect 699322 486478 700322 486546
rect 699322 486422 699392 486478
rect 699448 486422 699516 486478
rect 699572 486422 699640 486478
rect 699696 486422 699764 486478
rect 699820 486422 699888 486478
rect 699944 486422 700012 486478
rect 700068 486422 700136 486478
rect 700192 486422 700322 486478
rect 699322 486354 700322 486422
rect 699322 486298 699392 486354
rect 699448 486298 699516 486354
rect 699572 486298 699640 486354
rect 699696 486298 699764 486354
rect 699820 486298 699888 486354
rect 699944 486298 700012 486354
rect 700068 486298 700136 486354
rect 700192 486298 700322 486354
rect 699322 486230 700322 486298
rect 699322 486174 699392 486230
rect 699448 486174 699516 486230
rect 699572 486174 699640 486230
rect 699696 486174 699764 486230
rect 699820 486174 699888 486230
rect 699944 486174 700012 486230
rect 700068 486174 700136 486230
rect 700192 486174 700322 486230
rect 699322 486106 700322 486174
rect 699322 486050 699392 486106
rect 699448 486050 699516 486106
rect 699572 486050 699640 486106
rect 699696 486050 699764 486106
rect 699820 486050 699888 486106
rect 699944 486050 700012 486106
rect 700068 486050 700136 486106
rect 700192 486050 700322 486106
rect 699322 485982 700322 486050
rect 699322 485926 699392 485982
rect 699448 485926 699516 485982
rect 699572 485926 699640 485982
rect 699696 485926 699764 485982
rect 699820 485926 699888 485982
rect 699944 485926 700012 485982
rect 700068 485926 700136 485982
rect 700192 485926 700322 485982
rect 699322 485858 700322 485926
rect 699322 485802 699392 485858
rect 699448 485802 699516 485858
rect 699572 485802 699640 485858
rect 699696 485802 699764 485858
rect 699820 485802 699888 485858
rect 699944 485802 700012 485858
rect 700068 485802 700136 485858
rect 700192 485802 700322 485858
rect 699322 485734 700322 485802
rect 699322 485678 699392 485734
rect 699448 485678 699516 485734
rect 699572 485678 699640 485734
rect 699696 485678 699764 485734
rect 699820 485678 699888 485734
rect 699944 485678 700012 485734
rect 700068 485678 700136 485734
rect 700192 485678 700322 485734
rect 699322 485610 700322 485678
rect 699322 485554 699392 485610
rect 699448 485554 699516 485610
rect 699572 485554 699640 485610
rect 699696 485554 699764 485610
rect 699820 485554 699888 485610
rect 699944 485554 700012 485610
rect 700068 485554 700136 485610
rect 700192 485554 700322 485610
rect 699322 485486 700322 485554
rect 699322 485430 699392 485486
rect 699448 485430 699516 485486
rect 699572 485430 699640 485486
rect 699696 485430 699764 485486
rect 699820 485430 699888 485486
rect 699944 485430 700012 485486
rect 700068 485430 700136 485486
rect 700192 485430 700322 485486
rect 699322 485362 700322 485430
rect 699322 485306 699392 485362
rect 699448 485306 699516 485362
rect 699572 485306 699640 485362
rect 699696 485306 699764 485362
rect 699820 485306 699888 485362
rect 699944 485306 700012 485362
rect 700068 485306 700136 485362
rect 700192 485306 700322 485362
rect 699322 485238 700322 485306
rect 699322 485182 699392 485238
rect 699448 485182 699516 485238
rect 699572 485182 699640 485238
rect 699696 485182 699764 485238
rect 699820 485182 699888 485238
rect 699944 485182 700012 485238
rect 700068 485182 700136 485238
rect 700192 485182 700322 485238
rect 699322 485114 700322 485182
rect 699322 485058 699392 485114
rect 699448 485058 699516 485114
rect 699572 485058 699640 485114
rect 699696 485058 699764 485114
rect 699820 485058 699888 485114
rect 699944 485058 700012 485114
rect 700068 485058 700136 485114
rect 700192 485058 700322 485114
rect 699322 484990 700322 485058
rect 699322 484934 699392 484990
rect 699448 484934 699516 484990
rect 699572 484934 699640 484990
rect 699696 484934 699764 484990
rect 699820 484934 699888 484990
rect 699944 484934 700012 484990
rect 700068 484934 700136 484990
rect 700192 484934 700322 484990
rect 699322 484866 700322 484934
rect 699322 484810 699392 484866
rect 699448 484810 699516 484866
rect 699572 484810 699640 484866
rect 699696 484810 699764 484866
rect 699820 484810 699888 484866
rect 699944 484810 700012 484866
rect 700068 484810 700136 484866
rect 700192 484810 700322 484866
rect 699322 484122 700322 484810
rect 707800 486732 708000 486802
rect 707800 486676 707870 486732
rect 707926 486676 708000 486732
rect 707800 486608 708000 486676
rect 707800 486552 707870 486608
rect 707926 486552 708000 486608
rect 707800 486484 708000 486552
rect 707800 486428 707870 486484
rect 707926 486428 708000 486484
rect 707800 486360 708000 486428
rect 707800 486304 707870 486360
rect 707926 486304 708000 486360
rect 707800 486236 708000 486304
rect 707800 486180 707870 486236
rect 707926 486180 708000 486236
rect 707800 486112 708000 486180
rect 707800 486056 707870 486112
rect 707926 486056 708000 486112
rect 707800 485988 708000 486056
rect 707800 485932 707870 485988
rect 707926 485932 708000 485988
rect 707800 485864 708000 485932
rect 707800 485808 707870 485864
rect 707926 485808 708000 485864
rect 707800 485740 708000 485808
rect 707800 485684 707870 485740
rect 707926 485684 708000 485740
rect 707800 485616 708000 485684
rect 707800 485560 707870 485616
rect 707926 485560 708000 485616
rect 707800 485492 708000 485560
rect 707800 485436 707870 485492
rect 707926 485436 708000 485492
rect 707800 485368 708000 485436
rect 707800 485312 707870 485368
rect 707926 485312 708000 485368
rect 707800 485244 708000 485312
rect 707800 485188 707870 485244
rect 707926 485188 708000 485244
rect 707800 485120 708000 485188
rect 707800 485064 707870 485120
rect 707926 485064 708000 485120
rect 707800 484996 708000 485064
rect 707800 484940 707870 484996
rect 707926 484940 708000 484996
rect 707800 484872 708000 484940
rect 707800 484816 707870 484872
rect 707926 484816 708000 484872
rect 707800 484752 708000 484816
rect 699322 484066 699392 484122
rect 699448 484066 699516 484122
rect 699572 484066 699640 484122
rect 699696 484066 699764 484122
rect 699820 484066 699888 484122
rect 699944 484066 700012 484122
rect 700068 484066 700136 484122
rect 700192 484066 700322 484122
rect 699322 483998 700322 484066
rect 699322 483942 699392 483998
rect 699448 483942 699516 483998
rect 699572 483942 699640 483998
rect 699696 483942 699764 483998
rect 699820 483942 699888 483998
rect 699944 483942 700012 483998
rect 700068 483942 700136 483998
rect 700192 483942 700322 483998
rect 699322 483874 700322 483942
rect 699322 483818 699392 483874
rect 699448 483818 699516 483874
rect 699572 483818 699640 483874
rect 699696 483818 699764 483874
rect 699820 483818 699888 483874
rect 699944 483818 700012 483874
rect 700068 483818 700136 483874
rect 700192 483818 700322 483874
rect 699322 483750 700322 483818
rect 699322 483694 699392 483750
rect 699448 483694 699516 483750
rect 699572 483694 699640 483750
rect 699696 483694 699764 483750
rect 699820 483694 699888 483750
rect 699944 483694 700012 483750
rect 700068 483694 700136 483750
rect 700192 483694 700322 483750
rect 699322 483626 700322 483694
rect 699322 483570 699392 483626
rect 699448 483570 699516 483626
rect 699572 483570 699640 483626
rect 699696 483570 699764 483626
rect 699820 483570 699888 483626
rect 699944 483570 700012 483626
rect 700068 483570 700136 483626
rect 700192 483570 700322 483626
rect 699322 483502 700322 483570
rect 699322 483446 699392 483502
rect 699448 483446 699516 483502
rect 699572 483446 699640 483502
rect 699696 483446 699764 483502
rect 699820 483446 699888 483502
rect 699944 483446 700012 483502
rect 700068 483446 700136 483502
rect 700192 483446 700322 483502
rect 699322 483378 700322 483446
rect 699322 483322 699392 483378
rect 699448 483322 699516 483378
rect 699572 483322 699640 483378
rect 699696 483322 699764 483378
rect 699820 483322 699888 483378
rect 699944 483322 700012 483378
rect 700068 483322 700136 483378
rect 700192 483322 700322 483378
rect 699322 483254 700322 483322
rect 699322 483198 699392 483254
rect 699448 483198 699516 483254
rect 699572 483198 699640 483254
rect 699696 483198 699764 483254
rect 699820 483198 699888 483254
rect 699944 483198 700012 483254
rect 700068 483198 700136 483254
rect 700192 483198 700322 483254
rect 699322 483130 700322 483198
rect 699322 483074 699392 483130
rect 699448 483074 699516 483130
rect 699572 483074 699640 483130
rect 699696 483074 699764 483130
rect 699820 483074 699888 483130
rect 699944 483074 700012 483130
rect 700068 483074 700136 483130
rect 700192 483074 700322 483130
rect 699322 483006 700322 483074
rect 699322 482950 699392 483006
rect 699448 482950 699516 483006
rect 699572 482950 699640 483006
rect 699696 482950 699764 483006
rect 699820 482950 699888 483006
rect 699944 482950 700012 483006
rect 700068 482950 700136 483006
rect 700192 482950 700322 483006
rect 699322 482882 700322 482950
rect 699322 482826 699392 482882
rect 699448 482826 699516 482882
rect 699572 482826 699640 482882
rect 699696 482826 699764 482882
rect 699820 482826 699888 482882
rect 699944 482826 700012 482882
rect 700068 482826 700136 482882
rect 700192 482826 700322 482882
rect 699322 482758 700322 482826
rect 699322 482702 699392 482758
rect 699448 482702 699516 482758
rect 699572 482702 699640 482758
rect 699696 482702 699764 482758
rect 699820 482702 699888 482758
rect 699944 482702 700012 482758
rect 700068 482702 700136 482758
rect 700192 482702 700322 482758
rect 699322 482634 700322 482702
rect 699322 482578 699392 482634
rect 699448 482578 699516 482634
rect 699572 482578 699640 482634
rect 699696 482578 699764 482634
rect 699820 482578 699888 482634
rect 699944 482578 700012 482634
rect 700068 482578 700136 482634
rect 700192 482578 700322 482634
rect 699322 482510 700322 482578
rect 699322 482454 699392 482510
rect 699448 482454 699516 482510
rect 699572 482454 699640 482510
rect 699696 482454 699764 482510
rect 699820 482454 699888 482510
rect 699944 482454 700012 482510
rect 700068 482454 700136 482510
rect 700192 482454 700322 482510
rect 699322 482386 700322 482454
rect 699322 482330 699392 482386
rect 699448 482330 699516 482386
rect 699572 482330 699640 482386
rect 699696 482330 699764 482386
rect 699820 482330 699888 482386
rect 699944 482330 700012 482386
rect 700068 482330 700136 482386
rect 700192 482330 700322 482386
rect 699322 374429 700322 482330
rect 707800 484134 708000 484172
rect 707800 484078 707870 484134
rect 707926 484078 708000 484134
rect 707800 484010 708000 484078
rect 707800 483954 707870 484010
rect 707926 483954 708000 484010
rect 707800 483886 708000 483954
rect 707800 483830 707870 483886
rect 707926 483830 708000 483886
rect 707800 483762 708000 483830
rect 707800 483706 707870 483762
rect 707926 483706 708000 483762
rect 707800 483638 708000 483706
rect 707800 483582 707870 483638
rect 707926 483582 708000 483638
rect 707800 483514 708000 483582
rect 707800 483458 707870 483514
rect 707926 483458 708000 483514
rect 707800 483390 708000 483458
rect 707800 483334 707870 483390
rect 707926 483334 708000 483390
rect 707800 483266 708000 483334
rect 707800 483210 707870 483266
rect 707926 483210 708000 483266
rect 707800 483142 708000 483210
rect 707800 483086 707870 483142
rect 707926 483086 708000 483142
rect 707800 483018 708000 483086
rect 707800 482962 707870 483018
rect 707926 482962 708000 483018
rect 707800 482894 708000 482962
rect 707800 482838 707870 482894
rect 707926 482838 708000 482894
rect 707800 482770 708000 482838
rect 707800 482714 707870 482770
rect 707926 482714 708000 482770
rect 707800 482646 708000 482714
rect 707800 482590 707870 482646
rect 707926 482590 708000 482646
rect 707800 482522 708000 482590
rect 707800 482466 707870 482522
rect 707926 482466 708000 482522
rect 707800 482398 708000 482466
rect 707800 482342 707870 482398
rect 707926 482342 708000 482398
rect 707800 482272 708000 482342
rect 707801 453658 708001 453728
rect 707801 453602 707870 453658
rect 707926 453602 708001 453658
rect 707801 453534 708001 453602
rect 707801 453478 707870 453534
rect 707926 453478 708001 453534
rect 707801 453410 708001 453478
rect 707801 453354 707870 453410
rect 707926 453354 708001 453410
rect 707801 453286 708001 453354
rect 707801 453230 707870 453286
rect 707926 453230 708001 453286
rect 707801 453162 708001 453230
rect 707801 453106 707870 453162
rect 707926 453106 708001 453162
rect 707801 453038 708001 453106
rect 707801 452982 707870 453038
rect 707926 452982 708001 453038
rect 707801 452914 708001 452982
rect 707801 452858 707870 452914
rect 707926 452858 708001 452914
rect 707801 452790 708001 452858
rect 707801 452734 707870 452790
rect 707926 452734 708001 452790
rect 707801 452666 708001 452734
rect 707801 452610 707870 452666
rect 707926 452610 708001 452666
rect 707801 452542 708001 452610
rect 707801 452486 707870 452542
rect 707926 452486 708001 452542
rect 707801 452418 708001 452486
rect 707801 452362 707870 452418
rect 707926 452362 708001 452418
rect 707801 452294 708001 452362
rect 707801 452238 707870 452294
rect 707926 452238 708001 452294
rect 707801 452170 708001 452238
rect 707801 452114 707870 452170
rect 707926 452114 708001 452170
rect 707801 452046 708001 452114
rect 707801 451990 707870 452046
rect 707926 451990 708001 452046
rect 707801 451922 708001 451990
rect 707801 451866 707870 451922
rect 707926 451866 708001 451922
rect 707801 451828 708001 451866
rect 707801 451178 708001 451248
rect 707801 451122 707870 451178
rect 707926 451122 708001 451178
rect 707801 451054 708001 451122
rect 707801 450998 707870 451054
rect 707926 450998 708001 451054
rect 707801 450930 708001 450998
rect 707801 450874 707870 450930
rect 707926 450874 708001 450930
rect 707801 450806 708001 450874
rect 707801 450750 707870 450806
rect 707926 450750 708001 450806
rect 707801 450682 708001 450750
rect 707801 450626 707870 450682
rect 707926 450626 708001 450682
rect 707801 450558 708001 450626
rect 707801 450502 707870 450558
rect 707926 450502 708001 450558
rect 707801 450434 708001 450502
rect 707801 450378 707870 450434
rect 707926 450378 708001 450434
rect 707801 450310 708001 450378
rect 707801 450254 707870 450310
rect 707926 450254 708001 450310
rect 707801 450186 708001 450254
rect 707801 450130 707870 450186
rect 707926 450130 708001 450186
rect 707801 450062 708001 450130
rect 707801 450006 707870 450062
rect 707926 450006 708001 450062
rect 707801 449938 708001 450006
rect 707801 449882 707870 449938
rect 707926 449882 708001 449938
rect 707801 449814 708001 449882
rect 707801 449758 707870 449814
rect 707926 449758 708001 449814
rect 707801 449690 708001 449758
rect 707801 449634 707870 449690
rect 707926 449634 708001 449690
rect 707801 449566 708001 449634
rect 707801 449510 707870 449566
rect 707926 449510 708001 449566
rect 707801 449442 708001 449510
rect 707801 449386 707870 449442
rect 707926 449386 708001 449442
rect 707801 449318 708001 449386
rect 707801 449262 707870 449318
rect 707926 449262 708001 449318
rect 707801 449198 708001 449262
rect 707801 448808 708001 448878
rect 707801 448752 707870 448808
rect 707926 448752 708001 448808
rect 707801 448684 708001 448752
rect 707801 448628 707870 448684
rect 707926 448628 708001 448684
rect 707801 448560 708001 448628
rect 707801 448504 707870 448560
rect 707926 448504 708001 448560
rect 707801 448436 708001 448504
rect 707801 448380 707870 448436
rect 707926 448380 708001 448436
rect 707801 448312 708001 448380
rect 707801 448256 707870 448312
rect 707926 448256 708001 448312
rect 707801 448188 708001 448256
rect 707801 448132 707870 448188
rect 707926 448132 708001 448188
rect 707801 448064 708001 448132
rect 707801 448008 707870 448064
rect 707926 448008 708001 448064
rect 707801 447940 708001 448008
rect 707801 447884 707870 447940
rect 707926 447884 708001 447940
rect 707801 447816 708001 447884
rect 707801 447760 707870 447816
rect 707926 447760 708001 447816
rect 707801 447692 708001 447760
rect 707801 447636 707870 447692
rect 707926 447636 708001 447692
rect 707801 447568 708001 447636
rect 707801 447512 707870 447568
rect 707926 447512 708001 447568
rect 707801 447444 708001 447512
rect 707801 447388 707870 447444
rect 707926 447388 708001 447444
rect 707801 447320 708001 447388
rect 707801 447264 707870 447320
rect 707926 447264 708001 447320
rect 707801 447196 708001 447264
rect 707801 447140 707870 447196
rect 707926 447140 708001 447196
rect 707801 447072 708001 447140
rect 707801 447016 707870 447072
rect 707926 447016 708001 447072
rect 707801 446948 708001 447016
rect 707801 446892 707870 446948
rect 707926 446892 708001 446948
rect 707801 446828 708001 446892
rect 707801 446102 708001 446172
rect 707801 446046 707870 446102
rect 707926 446046 708001 446102
rect 707801 445978 708001 446046
rect 707801 445922 707870 445978
rect 707926 445922 708001 445978
rect 707801 445854 708001 445922
rect 707801 445798 707870 445854
rect 707926 445798 708001 445854
rect 707801 445730 708001 445798
rect 707801 445674 707870 445730
rect 707926 445674 708001 445730
rect 707801 445606 708001 445674
rect 707801 445550 707870 445606
rect 707926 445550 708001 445606
rect 707801 445482 708001 445550
rect 707801 445426 707870 445482
rect 707926 445426 708001 445482
rect 707801 445358 708001 445426
rect 707801 445302 707870 445358
rect 707926 445302 708001 445358
rect 707801 445234 708001 445302
rect 707801 445178 707870 445234
rect 707926 445178 708001 445234
rect 707801 445110 708001 445178
rect 707801 445054 707870 445110
rect 707926 445054 708001 445110
rect 707801 444986 708001 445054
rect 707801 444930 707870 444986
rect 707926 444930 708001 444986
rect 707801 444862 708001 444930
rect 707801 444806 707870 444862
rect 707926 444806 708001 444862
rect 707801 444738 708001 444806
rect 707801 444682 707870 444738
rect 707926 444682 708001 444738
rect 707801 444614 708001 444682
rect 707801 444558 707870 444614
rect 707926 444558 708001 444614
rect 707801 444490 708001 444558
rect 707801 444434 707870 444490
rect 707926 444434 708001 444490
rect 707801 444366 708001 444434
rect 707801 444310 707870 444366
rect 707926 444310 708001 444366
rect 707801 444242 708001 444310
rect 707801 444186 707870 444242
rect 707926 444186 708001 444242
rect 707801 444122 708001 444186
rect 707801 443732 708001 443802
rect 707801 443676 707870 443732
rect 707926 443676 708001 443732
rect 707801 443608 708001 443676
rect 707801 443552 707870 443608
rect 707926 443552 708001 443608
rect 707801 443484 708001 443552
rect 707801 443428 707870 443484
rect 707926 443428 708001 443484
rect 707801 443360 708001 443428
rect 707801 443304 707870 443360
rect 707926 443304 708001 443360
rect 707801 443236 708001 443304
rect 707801 443180 707870 443236
rect 707926 443180 708001 443236
rect 707801 443112 708001 443180
rect 707801 443056 707870 443112
rect 707926 443056 708001 443112
rect 707801 442988 708001 443056
rect 707801 442932 707870 442988
rect 707926 442932 708001 442988
rect 707801 442864 708001 442932
rect 707801 442808 707870 442864
rect 707926 442808 708001 442864
rect 707801 442740 708001 442808
rect 707801 442684 707870 442740
rect 707926 442684 708001 442740
rect 707801 442616 708001 442684
rect 707801 442560 707870 442616
rect 707926 442560 708001 442616
rect 707801 442492 708001 442560
rect 707801 442436 707870 442492
rect 707926 442436 708001 442492
rect 707801 442368 708001 442436
rect 707801 442312 707870 442368
rect 707926 442312 708001 442368
rect 707801 442244 708001 442312
rect 707801 442188 707870 442244
rect 707926 442188 708001 442244
rect 707801 442120 708001 442188
rect 707801 442064 707870 442120
rect 707926 442064 708001 442120
rect 707801 441996 708001 442064
rect 707801 441940 707870 441996
rect 707926 441940 708001 441996
rect 707801 441872 708001 441940
rect 707801 441816 707870 441872
rect 707926 441816 708001 441872
rect 707801 441752 708001 441816
rect 707801 441134 708001 441172
rect 707801 441078 707870 441134
rect 707926 441078 708001 441134
rect 707801 441010 708001 441078
rect 707801 440954 707870 441010
rect 707926 440954 708001 441010
rect 707801 440886 708001 440954
rect 707801 440830 707870 440886
rect 707926 440830 708001 440886
rect 707801 440762 708001 440830
rect 707801 440706 707870 440762
rect 707926 440706 708001 440762
rect 707801 440638 708001 440706
rect 707801 440582 707870 440638
rect 707926 440582 708001 440638
rect 707801 440514 708001 440582
rect 707801 440458 707870 440514
rect 707926 440458 708001 440514
rect 707801 440390 708001 440458
rect 707801 440334 707870 440390
rect 707926 440334 708001 440390
rect 707801 440266 708001 440334
rect 707801 440210 707870 440266
rect 707926 440210 708001 440266
rect 707801 440142 708001 440210
rect 707801 440086 707870 440142
rect 707926 440086 708001 440142
rect 707801 440018 708001 440086
rect 707801 439962 707870 440018
rect 707926 439962 708001 440018
rect 707801 439894 708001 439962
rect 707801 439838 707870 439894
rect 707926 439838 708001 439894
rect 707801 439770 708001 439838
rect 707801 439714 707870 439770
rect 707926 439714 708001 439770
rect 707801 439646 708001 439714
rect 707801 439590 707870 439646
rect 707926 439590 708001 439646
rect 707801 439522 708001 439590
rect 707801 439466 707870 439522
rect 707926 439466 708001 439522
rect 707801 439398 708001 439466
rect 707801 439342 707870 439398
rect 707926 439342 708001 439398
rect 707801 439272 708001 439342
rect 707800 410658 708000 410728
rect 707800 410602 707870 410658
rect 707926 410602 708000 410658
rect 707800 410534 708000 410602
rect 707800 410478 707870 410534
rect 707926 410478 708000 410534
rect 707800 410410 708000 410478
rect 707800 410354 707870 410410
rect 707926 410354 708000 410410
rect 707800 410286 708000 410354
rect 707800 410230 707870 410286
rect 707926 410230 708000 410286
rect 707800 410162 708000 410230
rect 707800 410106 707870 410162
rect 707926 410106 708000 410162
rect 707800 410038 708000 410106
rect 707800 409982 707870 410038
rect 707926 409982 708000 410038
rect 707800 409914 708000 409982
rect 707800 409858 707870 409914
rect 707926 409858 708000 409914
rect 707800 409790 708000 409858
rect 707800 409734 707870 409790
rect 707926 409734 708000 409790
rect 707800 409666 708000 409734
rect 707800 409610 707870 409666
rect 707926 409610 708000 409666
rect 707800 409542 708000 409610
rect 707800 409486 707870 409542
rect 707926 409486 708000 409542
rect 707800 409418 708000 409486
rect 707800 409362 707870 409418
rect 707926 409362 708000 409418
rect 707800 409294 708000 409362
rect 707800 409238 707870 409294
rect 707926 409238 708000 409294
rect 707800 409170 708000 409238
rect 707800 409114 707870 409170
rect 707926 409114 708000 409170
rect 707800 409046 708000 409114
rect 707800 408990 707870 409046
rect 707926 408990 708000 409046
rect 707800 408922 708000 408990
rect 707800 408866 707870 408922
rect 707926 408866 708000 408922
rect 707800 408828 708000 408866
rect 707800 408178 708000 408248
rect 707800 408122 707870 408178
rect 707926 408122 708000 408178
rect 707800 408054 708000 408122
rect 707800 407998 707870 408054
rect 707926 407998 708000 408054
rect 707800 407930 708000 407998
rect 707800 407874 707870 407930
rect 707926 407874 708000 407930
rect 707800 407806 708000 407874
rect 707800 407750 707870 407806
rect 707926 407750 708000 407806
rect 707800 407682 708000 407750
rect 707800 407626 707870 407682
rect 707926 407626 708000 407682
rect 707800 407558 708000 407626
rect 707800 407502 707870 407558
rect 707926 407502 708000 407558
rect 707800 407434 708000 407502
rect 707800 407378 707870 407434
rect 707926 407378 708000 407434
rect 707800 407310 708000 407378
rect 707800 407254 707870 407310
rect 707926 407254 708000 407310
rect 707800 407186 708000 407254
rect 707800 407130 707870 407186
rect 707926 407130 708000 407186
rect 707800 407062 708000 407130
rect 707800 407006 707870 407062
rect 707926 407006 708000 407062
rect 707800 406938 708000 407006
rect 707800 406882 707870 406938
rect 707926 406882 708000 406938
rect 707800 406814 708000 406882
rect 707800 406758 707870 406814
rect 707926 406758 708000 406814
rect 707800 406690 708000 406758
rect 707800 406634 707870 406690
rect 707926 406634 708000 406690
rect 707800 406566 708000 406634
rect 707800 406510 707870 406566
rect 707926 406510 708000 406566
rect 707800 406442 708000 406510
rect 707800 406386 707870 406442
rect 707926 406386 708000 406442
rect 707800 406318 708000 406386
rect 707800 406262 707870 406318
rect 707926 406262 708000 406318
rect 707800 406198 708000 406262
rect 707800 405808 708000 405878
rect 707800 405752 707870 405808
rect 707926 405752 708000 405808
rect 707800 405684 708000 405752
rect 707800 405628 707870 405684
rect 707926 405628 708000 405684
rect 707800 405560 708000 405628
rect 707800 405504 707870 405560
rect 707926 405504 708000 405560
rect 707800 405436 708000 405504
rect 707800 405380 707870 405436
rect 707926 405380 708000 405436
rect 707800 405312 708000 405380
rect 707800 405256 707870 405312
rect 707926 405256 708000 405312
rect 707800 405188 708000 405256
rect 707800 405132 707870 405188
rect 707926 405132 708000 405188
rect 707800 405064 708000 405132
rect 707800 405008 707870 405064
rect 707926 405008 708000 405064
rect 707800 404940 708000 405008
rect 707800 404884 707870 404940
rect 707926 404884 708000 404940
rect 707800 404816 708000 404884
rect 707800 404760 707870 404816
rect 707926 404760 708000 404816
rect 707800 404692 708000 404760
rect 707800 404636 707870 404692
rect 707926 404636 708000 404692
rect 707800 404568 708000 404636
rect 707800 404512 707870 404568
rect 707926 404512 708000 404568
rect 707800 404444 708000 404512
rect 707800 404388 707870 404444
rect 707926 404388 708000 404444
rect 707800 404320 708000 404388
rect 707800 404264 707870 404320
rect 707926 404264 708000 404320
rect 707800 404196 708000 404264
rect 707800 404140 707870 404196
rect 707926 404140 708000 404196
rect 707800 404072 708000 404140
rect 707800 404016 707870 404072
rect 707926 404016 708000 404072
rect 707800 403948 708000 404016
rect 707800 403892 707870 403948
rect 707926 403892 708000 403948
rect 707800 403828 708000 403892
rect 707800 403102 708000 403172
rect 707800 403046 707870 403102
rect 707926 403046 708000 403102
rect 707800 402978 708000 403046
rect 707800 402922 707870 402978
rect 707926 402922 708000 402978
rect 707800 402854 708000 402922
rect 707800 402798 707870 402854
rect 707926 402798 708000 402854
rect 707800 402730 708000 402798
rect 707800 402674 707870 402730
rect 707926 402674 708000 402730
rect 707800 402606 708000 402674
rect 707800 402550 707870 402606
rect 707926 402550 708000 402606
rect 707800 402482 708000 402550
rect 707800 402426 707870 402482
rect 707926 402426 708000 402482
rect 707800 402358 708000 402426
rect 707800 402302 707870 402358
rect 707926 402302 708000 402358
rect 707800 402234 708000 402302
rect 707800 402178 707870 402234
rect 707926 402178 708000 402234
rect 707800 402110 708000 402178
rect 707800 402054 707870 402110
rect 707926 402054 708000 402110
rect 707800 401986 708000 402054
rect 707800 401930 707870 401986
rect 707926 401930 708000 401986
rect 707800 401862 708000 401930
rect 707800 401806 707870 401862
rect 707926 401806 708000 401862
rect 707800 401738 708000 401806
rect 707800 401682 707870 401738
rect 707926 401682 708000 401738
rect 707800 401614 708000 401682
rect 707800 401558 707870 401614
rect 707926 401558 708000 401614
rect 707800 401490 708000 401558
rect 707800 401434 707870 401490
rect 707926 401434 708000 401490
rect 707800 401366 708000 401434
rect 707800 401310 707870 401366
rect 707926 401310 708000 401366
rect 707800 401242 708000 401310
rect 707800 401186 707870 401242
rect 707926 401186 708000 401242
rect 707800 401122 708000 401186
rect 707800 400732 708000 400802
rect 707800 400676 707870 400732
rect 707926 400676 708000 400732
rect 707800 400608 708000 400676
rect 707800 400552 707870 400608
rect 707926 400552 708000 400608
rect 707800 400484 708000 400552
rect 707800 400428 707870 400484
rect 707926 400428 708000 400484
rect 707800 400360 708000 400428
rect 707800 400304 707870 400360
rect 707926 400304 708000 400360
rect 707800 400236 708000 400304
rect 707800 400180 707870 400236
rect 707926 400180 708000 400236
rect 707800 400112 708000 400180
rect 707800 400056 707870 400112
rect 707926 400056 708000 400112
rect 707800 399988 708000 400056
rect 707800 399932 707870 399988
rect 707926 399932 708000 399988
rect 707800 399864 708000 399932
rect 707800 399808 707870 399864
rect 707926 399808 708000 399864
rect 707800 399740 708000 399808
rect 707800 399684 707870 399740
rect 707926 399684 708000 399740
rect 707800 399616 708000 399684
rect 707800 399560 707870 399616
rect 707926 399560 708000 399616
rect 707800 399492 708000 399560
rect 707800 399436 707870 399492
rect 707926 399436 708000 399492
rect 707800 399368 708000 399436
rect 707800 399312 707870 399368
rect 707926 399312 708000 399368
rect 707800 399244 708000 399312
rect 707800 399188 707870 399244
rect 707926 399188 708000 399244
rect 707800 399120 708000 399188
rect 707800 399064 707870 399120
rect 707926 399064 708000 399120
rect 707800 398996 708000 399064
rect 707800 398940 707870 398996
rect 707926 398940 708000 398996
rect 707800 398872 708000 398940
rect 707800 398816 707870 398872
rect 707926 398816 708000 398872
rect 707800 398752 708000 398816
rect 707800 398134 708000 398172
rect 707800 398078 707870 398134
rect 707926 398078 708000 398134
rect 707800 398010 708000 398078
rect 707800 397954 707870 398010
rect 707926 397954 708000 398010
rect 707800 397886 708000 397954
rect 707800 397830 707870 397886
rect 707926 397830 708000 397886
rect 707800 397762 708000 397830
rect 707800 397706 707870 397762
rect 707926 397706 708000 397762
rect 707800 397638 708000 397706
rect 707800 397582 707870 397638
rect 707926 397582 708000 397638
rect 707800 397514 708000 397582
rect 707800 397458 707870 397514
rect 707926 397458 708000 397514
rect 707800 397390 708000 397458
rect 707800 397334 707870 397390
rect 707926 397334 708000 397390
rect 707800 397266 708000 397334
rect 707800 397210 707870 397266
rect 707926 397210 708000 397266
rect 707800 397142 708000 397210
rect 707800 397086 707870 397142
rect 707926 397086 708000 397142
rect 707800 397018 708000 397086
rect 707800 396962 707870 397018
rect 707926 396962 708000 397018
rect 707800 396894 708000 396962
rect 707800 396838 707870 396894
rect 707926 396838 708000 396894
rect 707800 396770 708000 396838
rect 707800 396714 707870 396770
rect 707926 396714 708000 396770
rect 707800 396646 708000 396714
rect 707800 396590 707870 396646
rect 707926 396590 708000 396646
rect 707800 396522 708000 396590
rect 707800 396466 707870 396522
rect 707926 396466 708000 396522
rect 707800 396398 708000 396466
rect 707800 396342 707870 396398
rect 707926 396342 708000 396398
rect 707800 396272 708000 396342
rect 699322 374373 699544 374429
rect 699600 374373 699844 374429
rect 699900 374373 700144 374429
rect 700200 374373 700322 374429
rect 699322 374229 700322 374373
rect 699322 374173 699544 374229
rect 699600 374173 699844 374229
rect 699900 374173 700144 374229
rect 700200 374173 700322 374229
rect 699322 366954 700322 374173
rect 699322 366898 699444 366954
rect 699500 366898 699744 366954
rect 699800 366898 700044 366954
rect 700100 366898 700322 366954
rect 699322 359954 700322 366898
rect 699322 359898 699444 359954
rect 699500 359898 699744 359954
rect 699800 359898 700044 359954
rect 700100 359898 700322 359954
rect 699322 352954 700322 359898
rect 699322 352898 699444 352954
rect 699500 352898 699744 352954
rect 699800 352898 700044 352954
rect 700100 352898 700322 352954
rect 699322 338429 700322 352898
rect 699322 338373 699544 338429
rect 699600 338373 699844 338429
rect 699900 338373 700144 338429
rect 700200 338373 700322 338429
rect 699322 338229 700322 338373
rect 699322 338173 699544 338229
rect 699600 338173 699844 338229
rect 699900 338173 700144 338229
rect 700200 338173 700322 338229
rect 699322 333423 700322 338173
rect 699322 333367 699497 333423
rect 699553 333367 699797 333423
rect 699853 333367 700097 333423
rect 700153 333367 700322 333423
rect 699322 329640 700322 333367
rect 699322 329584 699452 329640
rect 699508 329584 699576 329640
rect 699632 329584 699700 329640
rect 699756 329584 699824 329640
rect 699880 329584 699948 329640
rect 700004 329584 700072 329640
rect 700128 329584 700196 329640
rect 700252 329584 700322 329640
rect 699322 329516 700322 329584
rect 699322 329460 699452 329516
rect 699508 329460 699576 329516
rect 699632 329460 699700 329516
rect 699756 329460 699824 329516
rect 699880 329460 699948 329516
rect 700004 329460 700072 329516
rect 700128 329460 700196 329516
rect 700252 329460 700322 329516
rect 699322 329392 700322 329460
rect 699322 329336 699452 329392
rect 699508 329336 699576 329392
rect 699632 329336 699700 329392
rect 699756 329336 699824 329392
rect 699880 329336 699948 329392
rect 700004 329336 700072 329392
rect 700128 329336 700196 329392
rect 700252 329336 700322 329392
rect 699322 329268 700322 329336
rect 699322 329212 699452 329268
rect 699508 329212 699576 329268
rect 699632 329212 699700 329268
rect 699756 329212 699824 329268
rect 699880 329212 699948 329268
rect 700004 329212 700072 329268
rect 700128 329212 700196 329268
rect 700252 329212 700322 329268
rect 699322 329144 700322 329212
rect 699322 329088 699452 329144
rect 699508 329088 699576 329144
rect 699632 329088 699700 329144
rect 699756 329088 699824 329144
rect 699880 329088 699948 329144
rect 700004 329088 700072 329144
rect 700128 329088 700196 329144
rect 700252 329088 700322 329144
rect 699322 329020 700322 329088
rect 699322 328964 699452 329020
rect 699508 328964 699576 329020
rect 699632 328964 699700 329020
rect 699756 328964 699824 329020
rect 699880 328964 699948 329020
rect 700004 328964 700072 329020
rect 700128 328964 700196 329020
rect 700252 328964 700322 329020
rect 699322 328896 700322 328964
rect 699322 328840 699452 328896
rect 699508 328840 699576 328896
rect 699632 328840 699700 328896
rect 699756 328840 699824 328896
rect 699880 328840 699948 328896
rect 700004 328840 700072 328896
rect 700128 328840 700196 328896
rect 700252 328840 700322 328896
rect 699322 323954 700322 328840
rect 699322 323898 699444 323954
rect 699500 323898 699744 323954
rect 699800 323898 700044 323954
rect 700100 323898 700322 323954
rect 699322 316954 700322 323898
rect 699322 316898 699444 316954
rect 699500 316898 699744 316954
rect 699800 316898 700044 316954
rect 700100 316898 700322 316954
rect 699322 309954 700322 316898
rect 699322 309898 699444 309954
rect 699500 309898 699744 309954
rect 699800 309898 700044 309954
rect 700100 309898 700322 309954
rect 699322 305786 700322 309898
rect 699322 305730 699452 305786
rect 699508 305730 699576 305786
rect 699632 305730 699700 305786
rect 699756 305730 699824 305786
rect 699880 305730 699948 305786
rect 700004 305730 700072 305786
rect 700128 305730 700196 305786
rect 700252 305730 700322 305786
rect 699322 305662 700322 305730
rect 699322 305606 699452 305662
rect 699508 305606 699576 305662
rect 699632 305606 699700 305662
rect 699756 305606 699824 305662
rect 699880 305606 699948 305662
rect 700004 305606 700072 305662
rect 700128 305606 700196 305662
rect 700252 305606 700322 305662
rect 699322 305538 700322 305606
rect 699322 305482 699452 305538
rect 699508 305482 699576 305538
rect 699632 305482 699700 305538
rect 699756 305482 699824 305538
rect 699880 305482 699948 305538
rect 700004 305482 700072 305538
rect 700128 305482 700196 305538
rect 700252 305482 700322 305538
rect 699322 305414 700322 305482
rect 699322 305358 699452 305414
rect 699508 305358 699576 305414
rect 699632 305358 699700 305414
rect 699756 305358 699824 305414
rect 699880 305358 699948 305414
rect 700004 305358 700072 305414
rect 700128 305358 700196 305414
rect 700252 305358 700322 305414
rect 699322 305290 700322 305358
rect 699322 305234 699452 305290
rect 699508 305234 699576 305290
rect 699632 305234 699700 305290
rect 699756 305234 699824 305290
rect 699880 305234 699948 305290
rect 700004 305234 700072 305290
rect 700128 305234 700196 305290
rect 700252 305234 700322 305290
rect 699322 305166 700322 305234
rect 699322 305110 699452 305166
rect 699508 305110 699576 305166
rect 699632 305110 699700 305166
rect 699756 305110 699824 305166
rect 699880 305110 699948 305166
rect 700004 305110 700072 305166
rect 700128 305110 700196 305166
rect 700252 305110 700322 305166
rect 699322 305042 700322 305110
rect 699322 304986 699452 305042
rect 699508 304986 699576 305042
rect 699632 304986 699700 305042
rect 699756 304986 699824 305042
rect 699880 304986 699948 305042
rect 700004 304986 700072 305042
rect 700128 304986 700196 305042
rect 700252 304986 700322 305042
rect 699322 290423 700322 304986
rect 699322 290367 699497 290423
rect 699553 290367 699797 290423
rect 699853 290367 700097 290423
rect 700153 290367 700322 290423
rect 699322 280954 700322 290367
rect 699322 280898 699444 280954
rect 699500 280898 699744 280954
rect 699800 280898 700044 280954
rect 700100 280898 700322 280954
rect 699322 273954 700322 280898
rect 699322 273898 699444 273954
rect 699500 273898 699744 273954
rect 699800 273898 700044 273954
rect 700100 273898 700322 273954
rect 699322 268607 700322 273898
rect 699322 268551 699444 268607
rect 699500 268551 699744 268607
rect 699800 268551 700044 268607
rect 700100 268551 700322 268607
rect 699322 266954 700322 268551
rect 699322 266898 699444 266954
rect 699500 266898 699744 266954
rect 699800 266898 700044 266954
rect 700100 266898 700322 266954
rect 699322 247423 700322 266898
rect 699322 247367 699497 247423
rect 699553 247367 699797 247423
rect 699853 247367 700097 247423
rect 700153 247367 700322 247423
rect 699322 237971 700322 247367
rect 699322 237915 699444 237971
rect 699500 237915 699744 237971
rect 699800 237915 700044 237971
rect 700100 237915 700322 237971
rect 699322 230954 700322 237915
rect 699322 230898 699444 230954
rect 699500 230898 699744 230954
rect 699800 230898 700044 230954
rect 700100 230898 700322 230954
rect 699322 223954 700322 230898
rect 699322 223898 699444 223954
rect 699500 223898 699744 223954
rect 699800 223898 700044 223954
rect 700100 223898 700322 223954
rect 699322 207335 700322 223898
rect 699322 207279 699444 207335
rect 699500 207279 699744 207335
rect 699800 207279 700044 207335
rect 700100 207279 700322 207335
rect 699322 204423 700322 207279
rect 699322 204367 699497 204423
rect 699553 204367 699797 204423
rect 699853 204367 700097 204423
rect 700153 204367 700322 204423
rect 699322 194954 700322 204367
rect 699322 194898 699444 194954
rect 699500 194898 699744 194954
rect 699800 194898 700044 194954
rect 700100 194898 700322 194954
rect 699322 187954 700322 194898
rect 699322 187898 699444 187954
rect 699500 187898 699744 187954
rect 699800 187898 700044 187954
rect 700100 187898 700322 187954
rect 699322 180954 700322 187898
rect 699322 180898 699444 180954
rect 699500 180898 699744 180954
rect 699800 180898 700044 180954
rect 700100 180898 700322 180954
rect 699322 176699 700322 180898
rect 699322 176643 699444 176699
rect 699500 176643 699744 176699
rect 699800 176643 700044 176699
rect 700100 176643 700322 176699
rect 699322 161423 700322 176643
rect 699322 161367 699497 161423
rect 699553 161367 699797 161423
rect 699853 161367 700097 161423
rect 700153 161367 700322 161423
rect 699322 151954 700322 161367
rect 699322 151898 699444 151954
rect 699500 151898 699744 151954
rect 699800 151898 700044 151954
rect 700100 151898 700322 151954
rect 699322 146063 700322 151898
rect 699322 146007 699444 146063
rect 699500 146007 699744 146063
rect 699800 146007 700044 146063
rect 700100 146007 700322 146063
rect 699322 144954 700322 146007
rect 699322 144898 699444 144954
rect 699500 144898 699744 144954
rect 699800 144898 700044 144954
rect 700100 144898 700322 144954
rect 699322 137954 700322 144898
rect 699322 137898 699444 137954
rect 699500 137898 699744 137954
rect 699800 137898 700044 137954
rect 700100 137898 700322 137954
rect 699322 133803 700322 137898
rect 699322 133747 699444 133803
rect 699500 133747 699744 133803
rect 699800 133747 700044 133803
rect 700100 133747 700322 133803
rect 699322 118423 700322 133747
rect 699322 118367 699497 118423
rect 699553 118367 699797 118423
rect 699853 118367 700097 118423
rect 700153 118367 700322 118423
rect 699322 108954 700322 118367
rect 699322 108898 699444 108954
rect 699500 108898 699744 108954
rect 699800 108898 700044 108954
rect 700100 108898 700322 108954
rect 699322 101954 700322 108898
rect 699322 101898 699444 101954
rect 699500 101898 699744 101954
rect 699800 101898 700044 101954
rect 700100 101898 700322 101954
rect 699322 94954 700322 101898
rect 699322 94898 699444 94954
rect 699500 94898 699744 94954
rect 699800 94898 700044 94954
rect 700100 94898 700322 94954
rect 699322 78608 700322 94898
rect 699322 78552 699452 78608
rect 699508 78552 699576 78608
rect 699632 78552 699700 78608
rect 699756 78552 699824 78608
rect 699880 78552 699948 78608
rect 700004 78552 700072 78608
rect 700128 78552 700196 78608
rect 700252 78552 700322 78608
rect 699322 78484 700322 78552
rect 699322 78428 699452 78484
rect 699508 78428 699576 78484
rect 699632 78428 699700 78484
rect 699756 78428 699824 78484
rect 699880 78428 699948 78484
rect 700004 78428 700072 78484
rect 700128 78428 700196 78484
rect 700252 78428 700322 78484
rect 699322 78360 700322 78428
rect 699322 78304 699452 78360
rect 699508 78304 699576 78360
rect 699632 78304 699700 78360
rect 699756 78304 699824 78360
rect 699880 78304 699948 78360
rect 700004 78304 700072 78360
rect 700128 78304 700196 78360
rect 700252 78304 700322 78360
rect 699322 78236 700322 78304
rect 699322 78180 699452 78236
rect 699508 78180 699576 78236
rect 699632 78180 699700 78236
rect 699756 78180 699824 78236
rect 699880 78180 699948 78236
rect 700004 78180 700072 78236
rect 700128 78180 700196 78236
rect 700252 78180 700322 78236
rect 699322 78112 700322 78180
rect 699322 78056 699452 78112
rect 699508 78056 699576 78112
rect 699632 78056 699700 78112
rect 699756 78056 699824 78112
rect 699880 78056 699948 78112
rect 700004 78056 700072 78112
rect 700128 78056 700196 78112
rect 700252 78056 700322 78112
rect 699322 77988 700322 78056
rect 699322 77932 699452 77988
rect 699508 77932 699576 77988
rect 699632 77932 699700 77988
rect 699756 77932 699824 77988
rect 699880 77932 699948 77988
rect 700004 77932 700072 77988
rect 700128 77932 700196 77988
rect 700252 77932 700322 77988
rect 699322 77864 700322 77932
rect 699322 77808 699452 77864
rect 699508 77808 699576 77864
rect 699632 77808 699700 77864
rect 699756 77808 699824 77864
rect 699880 77808 699948 77864
rect 700004 77808 700072 77864
rect 700128 77808 700196 77864
rect 700252 77808 700322 77864
rect 699322 75423 700322 77808
rect 699322 75367 699497 75423
rect 699553 75367 699797 75423
rect 699853 75367 700097 75423
rect 700153 75367 700322 75423
rect 699322 75290 700322 75367
rect 697922 74952 698060 75008
rect 698116 74952 698360 75008
rect 698416 74952 698660 75008
rect 698716 74952 698922 75008
rect 697922 74890 698922 74952
rect 669828 70074 669866 70130
rect 669922 70074 669990 70130
rect 670046 70074 670114 70130
rect 670170 70074 670238 70130
rect 670294 70074 670362 70130
rect 670418 70074 670486 70130
rect 670542 70074 670610 70130
rect 670666 70074 670734 70130
rect 670790 70074 670858 70130
rect 670914 70074 670982 70130
rect 671038 70074 671106 70130
rect 671162 70074 671230 70130
rect 671286 70074 671354 70130
rect 671410 70074 671478 70130
rect 671534 70074 671602 70130
rect 671658 70074 671728 70130
rect 669828 70000 671728 70074
<< via4 >>
rect 79284 945992 79340 946048
rect 79584 945992 79640 946048
rect 79884 945992 79940 946048
rect 77847 945577 77903 945633
rect 78147 945577 78203 945633
rect 78447 945577 78503 945633
rect 77748 942196 77804 942252
rect 77872 942196 77928 942252
rect 77996 942196 78052 942252
rect 78120 942196 78176 942252
rect 78244 942196 78300 942252
rect 78368 942196 78424 942252
rect 78492 942196 78548 942252
rect 77748 942072 77804 942128
rect 77872 942072 77928 942128
rect 77996 942072 78052 942128
rect 78120 942072 78176 942128
rect 78244 942072 78300 942128
rect 78368 942072 78424 942128
rect 78492 942072 78548 942128
rect 77748 941948 77804 942004
rect 77872 941948 77928 942004
rect 77996 941948 78052 942004
rect 78120 941948 78176 942004
rect 78244 941948 78300 942004
rect 78368 941948 78424 942004
rect 78492 941948 78548 942004
rect 77748 941824 77804 941880
rect 77872 941824 77928 941880
rect 77996 941824 78052 941880
rect 78120 941824 78176 941880
rect 78244 941824 78300 941880
rect 78368 941824 78424 941880
rect 78492 941824 78548 941880
rect 77748 941700 77804 941756
rect 77872 941700 77928 941756
rect 77996 941700 78052 941756
rect 78120 941700 78176 941756
rect 78244 941700 78300 941756
rect 78368 941700 78424 941756
rect 78492 941700 78548 941756
rect 77748 941576 77804 941632
rect 77872 941576 77928 941632
rect 77996 941576 78052 941632
rect 78120 941576 78176 941632
rect 78244 941576 78300 941632
rect 78368 941576 78424 941632
rect 78492 941576 78548 941632
rect 77748 941452 77804 941508
rect 77872 941452 77928 941508
rect 77996 941452 78052 941508
rect 78120 941452 78176 941508
rect 78244 941452 78300 941508
rect 78368 941452 78424 941508
rect 78492 941452 78548 941508
rect 77900 926046 77956 926102
rect 78200 926046 78256 926102
rect 78500 926046 78556 926102
rect 77900 919046 77956 919102
rect 78200 919046 78256 919102
rect 78500 919046 78556 919102
rect 77800 914373 77856 914429
rect 78100 914373 78156 914429
rect 78400 914373 78456 914429
rect 77800 914173 77856 914229
rect 78100 914173 78156 914229
rect 78400 914173 78456 914229
rect 77900 912046 77956 912102
rect 78200 912046 78256 912102
rect 78500 912046 78556 912102
rect 70074 884602 70130 884658
rect 70074 884478 70130 884534
rect 70074 884354 70130 884410
rect 70074 884230 70130 884286
rect 70074 884106 70130 884162
rect 70074 883982 70130 884038
rect 70074 883858 70130 883914
rect 70074 883734 70130 883790
rect 70074 883610 70130 883666
rect 70074 883486 70130 883542
rect 70074 883362 70130 883418
rect 70074 883238 70130 883294
rect 70074 883114 70130 883170
rect 70074 882990 70130 883046
rect 70074 882866 70130 882922
rect 77808 884614 77864 884670
rect 77932 884614 77988 884670
rect 78056 884614 78112 884670
rect 78180 884614 78236 884670
rect 78304 884614 78360 884670
rect 78428 884614 78484 884670
rect 78552 884614 78608 884670
rect 77808 884490 77864 884546
rect 77932 884490 77988 884546
rect 78056 884490 78112 884546
rect 78180 884490 78236 884546
rect 78304 884490 78360 884546
rect 78428 884490 78484 884546
rect 78552 884490 78608 884546
rect 77808 884366 77864 884422
rect 77932 884366 77988 884422
rect 78056 884366 78112 884422
rect 78180 884366 78236 884422
rect 78304 884366 78360 884422
rect 78428 884366 78484 884422
rect 78552 884366 78608 884422
rect 77808 884242 77864 884298
rect 77932 884242 77988 884298
rect 78056 884242 78112 884298
rect 78180 884242 78236 884298
rect 78304 884242 78360 884298
rect 78428 884242 78484 884298
rect 78552 884242 78608 884298
rect 77808 884118 77864 884174
rect 77932 884118 77988 884174
rect 78056 884118 78112 884174
rect 78180 884118 78236 884174
rect 78304 884118 78360 884174
rect 78428 884118 78484 884174
rect 78552 884118 78608 884174
rect 77808 883994 77864 884050
rect 77932 883994 77988 884050
rect 78056 883994 78112 884050
rect 78180 883994 78236 884050
rect 78304 883994 78360 884050
rect 78428 883994 78484 884050
rect 78552 883994 78608 884050
rect 77808 883870 77864 883926
rect 77932 883870 77988 883926
rect 78056 883870 78112 883926
rect 78180 883870 78236 883926
rect 78304 883870 78360 883926
rect 78428 883870 78484 883926
rect 78552 883870 78608 883926
rect 77808 883746 77864 883802
rect 77932 883746 77988 883802
rect 78056 883746 78112 883802
rect 78180 883746 78236 883802
rect 78304 883746 78360 883802
rect 78428 883746 78484 883802
rect 78552 883746 78608 883802
rect 77808 883622 77864 883678
rect 77932 883622 77988 883678
rect 78056 883622 78112 883678
rect 78180 883622 78236 883678
rect 78304 883622 78360 883678
rect 78428 883622 78484 883678
rect 78552 883622 78608 883678
rect 77808 883498 77864 883554
rect 77932 883498 77988 883554
rect 78056 883498 78112 883554
rect 78180 883498 78236 883554
rect 78304 883498 78360 883554
rect 78428 883498 78484 883554
rect 78552 883498 78608 883554
rect 77808 883374 77864 883430
rect 77932 883374 77988 883430
rect 78056 883374 78112 883430
rect 78180 883374 78236 883430
rect 78304 883374 78360 883430
rect 78428 883374 78484 883430
rect 78552 883374 78608 883430
rect 77808 883250 77864 883306
rect 77932 883250 77988 883306
rect 78056 883250 78112 883306
rect 78180 883250 78236 883306
rect 78304 883250 78360 883306
rect 78428 883250 78484 883306
rect 78552 883250 78608 883306
rect 77808 883126 77864 883182
rect 77932 883126 77988 883182
rect 78056 883126 78112 883182
rect 78180 883126 78236 883182
rect 78304 883126 78360 883182
rect 78428 883126 78484 883182
rect 78552 883126 78608 883182
rect 77808 883002 77864 883058
rect 77932 883002 77988 883058
rect 78056 883002 78112 883058
rect 78180 883002 78236 883058
rect 78304 883002 78360 883058
rect 78428 883002 78484 883058
rect 78552 883002 78608 883058
rect 77808 882878 77864 882934
rect 77932 882878 77988 882934
rect 78056 882878 78112 882934
rect 78180 882878 78236 882934
rect 78304 882878 78360 882934
rect 78428 882878 78484 882934
rect 78552 882878 78608 882934
rect 70074 882128 70130 882184
rect 70074 882004 70130 882060
rect 70074 881880 70130 881936
rect 70074 881756 70130 881812
rect 70074 881632 70130 881688
rect 70074 881508 70130 881564
rect 70074 881384 70130 881440
rect 70074 881260 70130 881316
rect 70074 881136 70130 881192
rect 70074 881012 70130 881068
rect 70074 880888 70130 880944
rect 70074 880764 70130 880820
rect 70074 880640 70130 880696
rect 70074 880516 70130 880572
rect 70074 880392 70130 880448
rect 70074 880268 70130 880324
rect 77808 882134 77864 882190
rect 77932 882134 77988 882190
rect 78056 882134 78112 882190
rect 78180 882134 78236 882190
rect 78304 882134 78360 882190
rect 78428 882134 78484 882190
rect 78552 882134 78608 882190
rect 77808 882010 77864 882066
rect 77932 882010 77988 882066
rect 78056 882010 78112 882066
rect 78180 882010 78236 882066
rect 78304 882010 78360 882066
rect 78428 882010 78484 882066
rect 78552 882010 78608 882066
rect 77808 881886 77864 881942
rect 77932 881886 77988 881942
rect 78056 881886 78112 881942
rect 78180 881886 78236 881942
rect 78304 881886 78360 881942
rect 78428 881886 78484 881942
rect 78552 881886 78608 881942
rect 77808 881762 77864 881818
rect 77932 881762 77988 881818
rect 78056 881762 78112 881818
rect 78180 881762 78236 881818
rect 78304 881762 78360 881818
rect 78428 881762 78484 881818
rect 78552 881762 78608 881818
rect 77808 881638 77864 881694
rect 77932 881638 77988 881694
rect 78056 881638 78112 881694
rect 78180 881638 78236 881694
rect 78304 881638 78360 881694
rect 78428 881638 78484 881694
rect 78552 881638 78608 881694
rect 77808 881514 77864 881570
rect 77932 881514 77988 881570
rect 78056 881514 78112 881570
rect 78180 881514 78236 881570
rect 78304 881514 78360 881570
rect 78428 881514 78484 881570
rect 78552 881514 78608 881570
rect 77808 881390 77864 881446
rect 77932 881390 77988 881446
rect 78056 881390 78112 881446
rect 78180 881390 78236 881446
rect 78304 881390 78360 881446
rect 78428 881390 78484 881446
rect 78552 881390 78608 881446
rect 77808 881266 77864 881322
rect 77932 881266 77988 881322
rect 78056 881266 78112 881322
rect 78180 881266 78236 881322
rect 78304 881266 78360 881322
rect 78428 881266 78484 881322
rect 78552 881266 78608 881322
rect 77808 881142 77864 881198
rect 77932 881142 77988 881198
rect 78056 881142 78112 881198
rect 78180 881142 78236 881198
rect 78304 881142 78360 881198
rect 78428 881142 78484 881198
rect 78552 881142 78608 881198
rect 77808 881018 77864 881074
rect 77932 881018 77988 881074
rect 78056 881018 78112 881074
rect 78180 881018 78236 881074
rect 78304 881018 78360 881074
rect 78428 881018 78484 881074
rect 78552 881018 78608 881074
rect 77808 880894 77864 880950
rect 77932 880894 77988 880950
rect 78056 880894 78112 880950
rect 78180 880894 78236 880950
rect 78304 880894 78360 880950
rect 78428 880894 78484 880950
rect 78552 880894 78608 880950
rect 77808 880770 77864 880826
rect 77932 880770 77988 880826
rect 78056 880770 78112 880826
rect 78180 880770 78236 880826
rect 78304 880770 78360 880826
rect 78428 880770 78484 880826
rect 78552 880770 78608 880826
rect 77808 880646 77864 880702
rect 77932 880646 77988 880702
rect 78056 880646 78112 880702
rect 78180 880646 78236 880702
rect 78304 880646 78360 880702
rect 78428 880646 78484 880702
rect 78552 880646 78608 880702
rect 77808 880522 77864 880578
rect 77932 880522 77988 880578
rect 78056 880522 78112 880578
rect 78180 880522 78236 880578
rect 78304 880522 78360 880578
rect 78428 880522 78484 880578
rect 78552 880522 78608 880578
rect 77808 880398 77864 880454
rect 77932 880398 77988 880454
rect 78056 880398 78112 880454
rect 78180 880398 78236 880454
rect 78304 880398 78360 880454
rect 78428 880398 78484 880454
rect 78552 880398 78608 880454
rect 77808 880274 77864 880330
rect 77932 880274 77988 880330
rect 78056 880274 78112 880330
rect 78180 880274 78236 880330
rect 78304 880274 78360 880330
rect 78428 880274 78484 880330
rect 78552 880274 78608 880330
rect 70074 879758 70130 879814
rect 70074 879634 70130 879690
rect 70074 879510 70130 879566
rect 70074 879386 70130 879442
rect 70074 879262 70130 879318
rect 70074 879138 70130 879194
rect 70074 879014 70130 879070
rect 70074 878890 70130 878946
rect 70074 878766 70130 878822
rect 70074 878642 70130 878698
rect 70074 878518 70130 878574
rect 70074 878394 70130 878450
rect 70074 878270 70130 878326
rect 70074 878146 70130 878202
rect 70074 878022 70130 878078
rect 70074 877898 70130 877954
rect 77808 879764 77864 879820
rect 77932 879764 77988 879820
rect 78056 879764 78112 879820
rect 78180 879764 78236 879820
rect 78304 879764 78360 879820
rect 78428 879764 78484 879820
rect 78552 879764 78608 879820
rect 77808 879640 77864 879696
rect 77932 879640 77988 879696
rect 78056 879640 78112 879696
rect 78180 879640 78236 879696
rect 78304 879640 78360 879696
rect 78428 879640 78484 879696
rect 78552 879640 78608 879696
rect 77808 879516 77864 879572
rect 77932 879516 77988 879572
rect 78056 879516 78112 879572
rect 78180 879516 78236 879572
rect 78304 879516 78360 879572
rect 78428 879516 78484 879572
rect 78552 879516 78608 879572
rect 77808 879392 77864 879448
rect 77932 879392 77988 879448
rect 78056 879392 78112 879448
rect 78180 879392 78236 879448
rect 78304 879392 78360 879448
rect 78428 879392 78484 879448
rect 78552 879392 78608 879448
rect 77808 879268 77864 879324
rect 77932 879268 77988 879324
rect 78056 879268 78112 879324
rect 78180 879268 78236 879324
rect 78304 879268 78360 879324
rect 78428 879268 78484 879324
rect 78552 879268 78608 879324
rect 77808 879144 77864 879200
rect 77932 879144 77988 879200
rect 78056 879144 78112 879200
rect 78180 879144 78236 879200
rect 78304 879144 78360 879200
rect 78428 879144 78484 879200
rect 78552 879144 78608 879200
rect 77808 879020 77864 879076
rect 77932 879020 77988 879076
rect 78056 879020 78112 879076
rect 78180 879020 78236 879076
rect 78304 879020 78360 879076
rect 78428 879020 78484 879076
rect 78552 879020 78608 879076
rect 77808 878896 77864 878952
rect 77932 878896 77988 878952
rect 78056 878896 78112 878952
rect 78180 878896 78236 878952
rect 78304 878896 78360 878952
rect 78428 878896 78484 878952
rect 78552 878896 78608 878952
rect 77808 878772 77864 878828
rect 77932 878772 77988 878828
rect 78056 878772 78112 878828
rect 78180 878772 78236 878828
rect 78304 878772 78360 878828
rect 78428 878772 78484 878828
rect 78552 878772 78608 878828
rect 77808 878648 77864 878704
rect 77932 878648 77988 878704
rect 78056 878648 78112 878704
rect 78180 878648 78236 878704
rect 78304 878648 78360 878704
rect 78428 878648 78484 878704
rect 78552 878648 78608 878704
rect 77808 878524 77864 878580
rect 77932 878524 77988 878580
rect 78056 878524 78112 878580
rect 78180 878524 78236 878580
rect 78304 878524 78360 878580
rect 78428 878524 78484 878580
rect 78552 878524 78608 878580
rect 77808 878400 77864 878456
rect 77932 878400 77988 878456
rect 78056 878400 78112 878456
rect 78180 878400 78236 878456
rect 78304 878400 78360 878456
rect 78428 878400 78484 878456
rect 78552 878400 78608 878456
rect 77808 878276 77864 878332
rect 77932 878276 77988 878332
rect 78056 878276 78112 878332
rect 78180 878276 78236 878332
rect 78304 878276 78360 878332
rect 78428 878276 78484 878332
rect 78552 878276 78608 878332
rect 77808 878152 77864 878208
rect 77932 878152 77988 878208
rect 78056 878152 78112 878208
rect 78180 878152 78236 878208
rect 78304 878152 78360 878208
rect 78428 878152 78484 878208
rect 78552 878152 78608 878208
rect 77808 878028 77864 878084
rect 77932 878028 77988 878084
rect 78056 878028 78112 878084
rect 78180 878028 78236 878084
rect 78304 878028 78360 878084
rect 78428 878028 78484 878084
rect 78552 878028 78608 878084
rect 77808 877904 77864 877960
rect 77932 877904 77988 877960
rect 78056 877904 78112 877960
rect 78180 877904 78236 877960
rect 78304 877904 78360 877960
rect 78428 877904 78484 877960
rect 78552 877904 78608 877960
rect 70074 877052 70130 877108
rect 70074 876928 70130 876984
rect 70074 876804 70130 876860
rect 70074 876680 70130 876736
rect 70074 876556 70130 876612
rect 70074 876432 70130 876488
rect 70074 876308 70130 876364
rect 70074 876184 70130 876240
rect 70074 876060 70130 876116
rect 70074 875936 70130 875992
rect 70074 875812 70130 875868
rect 70074 875688 70130 875744
rect 70074 875564 70130 875620
rect 70074 875440 70130 875496
rect 70074 875316 70130 875372
rect 70074 875192 70130 875248
rect 77808 877058 77864 877114
rect 77932 877058 77988 877114
rect 78056 877058 78112 877114
rect 78180 877058 78236 877114
rect 78304 877058 78360 877114
rect 78428 877058 78484 877114
rect 78552 877058 78608 877114
rect 77808 876934 77864 876990
rect 77932 876934 77988 876990
rect 78056 876934 78112 876990
rect 78180 876934 78236 876990
rect 78304 876934 78360 876990
rect 78428 876934 78484 876990
rect 78552 876934 78608 876990
rect 77808 876810 77864 876866
rect 77932 876810 77988 876866
rect 78056 876810 78112 876866
rect 78180 876810 78236 876866
rect 78304 876810 78360 876866
rect 78428 876810 78484 876866
rect 78552 876810 78608 876866
rect 77808 876686 77864 876742
rect 77932 876686 77988 876742
rect 78056 876686 78112 876742
rect 78180 876686 78236 876742
rect 78304 876686 78360 876742
rect 78428 876686 78484 876742
rect 78552 876686 78608 876742
rect 77808 876562 77864 876618
rect 77932 876562 77988 876618
rect 78056 876562 78112 876618
rect 78180 876562 78236 876618
rect 78304 876562 78360 876618
rect 78428 876562 78484 876618
rect 78552 876562 78608 876618
rect 77808 876438 77864 876494
rect 77932 876438 77988 876494
rect 78056 876438 78112 876494
rect 78180 876438 78236 876494
rect 78304 876438 78360 876494
rect 78428 876438 78484 876494
rect 78552 876438 78608 876494
rect 77808 876314 77864 876370
rect 77932 876314 77988 876370
rect 78056 876314 78112 876370
rect 78180 876314 78236 876370
rect 78304 876314 78360 876370
rect 78428 876314 78484 876370
rect 78552 876314 78608 876370
rect 77808 876190 77864 876246
rect 77932 876190 77988 876246
rect 78056 876190 78112 876246
rect 78180 876190 78236 876246
rect 78304 876190 78360 876246
rect 78428 876190 78484 876246
rect 78552 876190 78608 876246
rect 77808 876066 77864 876122
rect 77932 876066 77988 876122
rect 78056 876066 78112 876122
rect 78180 876066 78236 876122
rect 78304 876066 78360 876122
rect 78428 876066 78484 876122
rect 78552 876066 78608 876122
rect 77808 875942 77864 875998
rect 77932 875942 77988 875998
rect 78056 875942 78112 875998
rect 78180 875942 78236 875998
rect 78304 875942 78360 875998
rect 78428 875942 78484 875998
rect 78552 875942 78608 875998
rect 77808 875818 77864 875874
rect 77932 875818 77988 875874
rect 78056 875818 78112 875874
rect 78180 875818 78236 875874
rect 78304 875818 78360 875874
rect 78428 875818 78484 875874
rect 78552 875818 78608 875874
rect 77808 875694 77864 875750
rect 77932 875694 77988 875750
rect 78056 875694 78112 875750
rect 78180 875694 78236 875750
rect 78304 875694 78360 875750
rect 78428 875694 78484 875750
rect 78552 875694 78608 875750
rect 77808 875570 77864 875626
rect 77932 875570 77988 875626
rect 78056 875570 78112 875626
rect 78180 875570 78236 875626
rect 78304 875570 78360 875626
rect 78428 875570 78484 875626
rect 78552 875570 78608 875626
rect 77808 875446 77864 875502
rect 77932 875446 77988 875502
rect 78056 875446 78112 875502
rect 78180 875446 78236 875502
rect 78304 875446 78360 875502
rect 78428 875446 78484 875502
rect 78552 875446 78608 875502
rect 77808 875322 77864 875378
rect 77932 875322 77988 875378
rect 78056 875322 78112 875378
rect 78180 875322 78236 875378
rect 78304 875322 78360 875378
rect 78428 875322 78484 875378
rect 78552 875322 78608 875378
rect 77808 875198 77864 875254
rect 77932 875198 77988 875254
rect 78056 875198 78112 875254
rect 78180 875198 78236 875254
rect 78304 875198 78360 875254
rect 78428 875198 78484 875254
rect 78552 875198 78608 875254
rect 70074 874682 70130 874738
rect 70074 874558 70130 874614
rect 70074 874434 70130 874490
rect 70074 874310 70130 874366
rect 70074 874186 70130 874242
rect 70074 874062 70130 874118
rect 70074 873938 70130 873994
rect 70074 873814 70130 873870
rect 70074 873690 70130 873746
rect 70074 873566 70130 873622
rect 70074 873442 70130 873498
rect 70074 873318 70130 873374
rect 70074 873194 70130 873250
rect 70074 873070 70130 873126
rect 70074 872946 70130 873002
rect 70074 872822 70130 872878
rect 77808 874688 77864 874744
rect 77932 874688 77988 874744
rect 78056 874688 78112 874744
rect 78180 874688 78236 874744
rect 78304 874688 78360 874744
rect 78428 874688 78484 874744
rect 78552 874688 78608 874744
rect 77808 874564 77864 874620
rect 77932 874564 77988 874620
rect 78056 874564 78112 874620
rect 78180 874564 78236 874620
rect 78304 874564 78360 874620
rect 78428 874564 78484 874620
rect 78552 874564 78608 874620
rect 77808 874440 77864 874496
rect 77932 874440 77988 874496
rect 78056 874440 78112 874496
rect 78180 874440 78236 874496
rect 78304 874440 78360 874496
rect 78428 874440 78484 874496
rect 78552 874440 78608 874496
rect 77808 874316 77864 874372
rect 77932 874316 77988 874372
rect 78056 874316 78112 874372
rect 78180 874316 78236 874372
rect 78304 874316 78360 874372
rect 78428 874316 78484 874372
rect 78552 874316 78608 874372
rect 77808 874192 77864 874248
rect 77932 874192 77988 874248
rect 78056 874192 78112 874248
rect 78180 874192 78236 874248
rect 78304 874192 78360 874248
rect 78428 874192 78484 874248
rect 78552 874192 78608 874248
rect 77808 874068 77864 874124
rect 77932 874068 77988 874124
rect 78056 874068 78112 874124
rect 78180 874068 78236 874124
rect 78304 874068 78360 874124
rect 78428 874068 78484 874124
rect 78552 874068 78608 874124
rect 77808 873944 77864 874000
rect 77932 873944 77988 874000
rect 78056 873944 78112 874000
rect 78180 873944 78236 874000
rect 78304 873944 78360 874000
rect 78428 873944 78484 874000
rect 78552 873944 78608 874000
rect 77808 873820 77864 873876
rect 77932 873820 77988 873876
rect 78056 873820 78112 873876
rect 78180 873820 78236 873876
rect 78304 873820 78360 873876
rect 78428 873820 78484 873876
rect 78552 873820 78608 873876
rect 77808 873696 77864 873752
rect 77932 873696 77988 873752
rect 78056 873696 78112 873752
rect 78180 873696 78236 873752
rect 78304 873696 78360 873752
rect 78428 873696 78484 873752
rect 78552 873696 78608 873752
rect 77808 873572 77864 873628
rect 77932 873572 77988 873628
rect 78056 873572 78112 873628
rect 78180 873572 78236 873628
rect 78304 873572 78360 873628
rect 78428 873572 78484 873628
rect 78552 873572 78608 873628
rect 77808 873448 77864 873504
rect 77932 873448 77988 873504
rect 78056 873448 78112 873504
rect 78180 873448 78236 873504
rect 78304 873448 78360 873504
rect 78428 873448 78484 873504
rect 78552 873448 78608 873504
rect 77808 873324 77864 873380
rect 77932 873324 77988 873380
rect 78056 873324 78112 873380
rect 78180 873324 78236 873380
rect 78304 873324 78360 873380
rect 78428 873324 78484 873380
rect 78552 873324 78608 873380
rect 77808 873200 77864 873256
rect 77932 873200 77988 873256
rect 78056 873200 78112 873256
rect 78180 873200 78236 873256
rect 78304 873200 78360 873256
rect 78428 873200 78484 873256
rect 78552 873200 78608 873256
rect 77808 873076 77864 873132
rect 77932 873076 77988 873132
rect 78056 873076 78112 873132
rect 78180 873076 78236 873132
rect 78304 873076 78360 873132
rect 78428 873076 78484 873132
rect 78552 873076 78608 873132
rect 77808 872952 77864 873008
rect 77932 872952 77988 873008
rect 78056 872952 78112 873008
rect 78180 872952 78236 873008
rect 78304 872952 78360 873008
rect 78428 872952 78484 873008
rect 78552 872952 78608 873008
rect 77808 872828 77864 872884
rect 77932 872828 77988 872884
rect 78056 872828 78112 872884
rect 78180 872828 78236 872884
rect 78304 872828 78360 872884
rect 78428 872828 78484 872884
rect 78552 872828 78608 872884
rect 70074 872078 70130 872134
rect 70074 871954 70130 872010
rect 70074 871830 70130 871886
rect 70074 871706 70130 871762
rect 70074 871582 70130 871638
rect 70074 871458 70130 871514
rect 70074 871334 70130 871390
rect 70074 871210 70130 871266
rect 70074 871086 70130 871142
rect 70074 870962 70130 871018
rect 70074 870838 70130 870894
rect 70074 870714 70130 870770
rect 70074 870590 70130 870646
rect 70074 870466 70130 870522
rect 70074 870342 70130 870398
rect 77808 872084 77864 872140
rect 77932 872084 77988 872140
rect 78056 872084 78112 872140
rect 78180 872084 78236 872140
rect 78304 872084 78360 872140
rect 78428 872084 78484 872140
rect 78552 872084 78608 872140
rect 77808 871960 77864 872016
rect 77932 871960 77988 872016
rect 78056 871960 78112 872016
rect 78180 871960 78236 872016
rect 78304 871960 78360 872016
rect 78428 871960 78484 872016
rect 78552 871960 78608 872016
rect 77808 871836 77864 871892
rect 77932 871836 77988 871892
rect 78056 871836 78112 871892
rect 78180 871836 78236 871892
rect 78304 871836 78360 871892
rect 78428 871836 78484 871892
rect 78552 871836 78608 871892
rect 77808 871712 77864 871768
rect 77932 871712 77988 871768
rect 78056 871712 78112 871768
rect 78180 871712 78236 871768
rect 78304 871712 78360 871768
rect 78428 871712 78484 871768
rect 78552 871712 78608 871768
rect 77808 871588 77864 871644
rect 77932 871588 77988 871644
rect 78056 871588 78112 871644
rect 78180 871588 78236 871644
rect 78304 871588 78360 871644
rect 78428 871588 78484 871644
rect 78552 871588 78608 871644
rect 77808 871464 77864 871520
rect 77932 871464 77988 871520
rect 78056 871464 78112 871520
rect 78180 871464 78236 871520
rect 78304 871464 78360 871520
rect 78428 871464 78484 871520
rect 78552 871464 78608 871520
rect 77808 871340 77864 871396
rect 77932 871340 77988 871396
rect 78056 871340 78112 871396
rect 78180 871340 78236 871396
rect 78304 871340 78360 871396
rect 78428 871340 78484 871396
rect 78552 871340 78608 871396
rect 77808 871216 77864 871272
rect 77932 871216 77988 871272
rect 78056 871216 78112 871272
rect 78180 871216 78236 871272
rect 78304 871216 78360 871272
rect 78428 871216 78484 871272
rect 78552 871216 78608 871272
rect 77808 871092 77864 871148
rect 77932 871092 77988 871148
rect 78056 871092 78112 871148
rect 78180 871092 78236 871148
rect 78304 871092 78360 871148
rect 78428 871092 78484 871148
rect 78552 871092 78608 871148
rect 77808 870968 77864 871024
rect 77932 870968 77988 871024
rect 78056 870968 78112 871024
rect 78180 870968 78236 871024
rect 78304 870968 78360 871024
rect 78428 870968 78484 871024
rect 78552 870968 78608 871024
rect 77808 870844 77864 870900
rect 77932 870844 77988 870900
rect 78056 870844 78112 870900
rect 78180 870844 78236 870900
rect 78304 870844 78360 870900
rect 78428 870844 78484 870900
rect 78552 870844 78608 870900
rect 77808 870720 77864 870776
rect 77932 870720 77988 870776
rect 78056 870720 78112 870776
rect 78180 870720 78236 870776
rect 78304 870720 78360 870776
rect 78428 870720 78484 870776
rect 78552 870720 78608 870776
rect 77808 870596 77864 870652
rect 77932 870596 77988 870652
rect 78056 870596 78112 870652
rect 78180 870596 78236 870652
rect 78304 870596 78360 870652
rect 78428 870596 78484 870652
rect 78552 870596 78608 870652
rect 77808 870472 77864 870528
rect 77932 870472 77988 870528
rect 78056 870472 78112 870528
rect 78180 870472 78236 870528
rect 78304 870472 78360 870528
rect 78428 870472 78484 870528
rect 78552 870472 78608 870528
rect 77808 870348 77864 870404
rect 77932 870348 77988 870404
rect 78056 870348 78112 870404
rect 78180 870348 78236 870404
rect 78304 870348 78360 870404
rect 78428 870348 78484 870404
rect 78552 870348 78608 870404
rect 70074 843602 70130 843658
rect 70074 843478 70130 843534
rect 70074 843354 70130 843410
rect 70074 843230 70130 843286
rect 70074 843106 70130 843162
rect 70074 842982 70130 843038
rect 70074 842858 70130 842914
rect 70074 842734 70130 842790
rect 70074 842610 70130 842666
rect 70074 842486 70130 842542
rect 70074 842362 70130 842418
rect 70074 842238 70130 842294
rect 70074 842114 70130 842170
rect 70074 841990 70130 842046
rect 70074 841866 70130 841922
rect 77808 843614 77864 843670
rect 77932 843614 77988 843670
rect 78056 843614 78112 843670
rect 78180 843614 78236 843670
rect 78304 843614 78360 843670
rect 78428 843614 78484 843670
rect 78552 843614 78608 843670
rect 77808 843490 77864 843546
rect 77932 843490 77988 843546
rect 78056 843490 78112 843546
rect 78180 843490 78236 843546
rect 78304 843490 78360 843546
rect 78428 843490 78484 843546
rect 78552 843490 78608 843546
rect 77808 843366 77864 843422
rect 77932 843366 77988 843422
rect 78056 843366 78112 843422
rect 78180 843366 78236 843422
rect 78304 843366 78360 843422
rect 78428 843366 78484 843422
rect 78552 843366 78608 843422
rect 77808 843242 77864 843298
rect 77932 843242 77988 843298
rect 78056 843242 78112 843298
rect 78180 843242 78236 843298
rect 78304 843242 78360 843298
rect 78428 843242 78484 843298
rect 78552 843242 78608 843298
rect 77808 843118 77864 843174
rect 77932 843118 77988 843174
rect 78056 843118 78112 843174
rect 78180 843118 78236 843174
rect 78304 843118 78360 843174
rect 78428 843118 78484 843174
rect 78552 843118 78608 843174
rect 77808 842994 77864 843050
rect 77932 842994 77988 843050
rect 78056 842994 78112 843050
rect 78180 842994 78236 843050
rect 78304 842994 78360 843050
rect 78428 842994 78484 843050
rect 78552 842994 78608 843050
rect 77808 842870 77864 842926
rect 77932 842870 77988 842926
rect 78056 842870 78112 842926
rect 78180 842870 78236 842926
rect 78304 842870 78360 842926
rect 78428 842870 78484 842926
rect 78552 842870 78608 842926
rect 77808 842746 77864 842802
rect 77932 842746 77988 842802
rect 78056 842746 78112 842802
rect 78180 842746 78236 842802
rect 78304 842746 78360 842802
rect 78428 842746 78484 842802
rect 78552 842746 78608 842802
rect 77808 842622 77864 842678
rect 77932 842622 77988 842678
rect 78056 842622 78112 842678
rect 78180 842622 78236 842678
rect 78304 842622 78360 842678
rect 78428 842622 78484 842678
rect 78552 842622 78608 842678
rect 77808 842498 77864 842554
rect 77932 842498 77988 842554
rect 78056 842498 78112 842554
rect 78180 842498 78236 842554
rect 78304 842498 78360 842554
rect 78428 842498 78484 842554
rect 78552 842498 78608 842554
rect 77808 842374 77864 842430
rect 77932 842374 77988 842430
rect 78056 842374 78112 842430
rect 78180 842374 78236 842430
rect 78304 842374 78360 842430
rect 78428 842374 78484 842430
rect 78552 842374 78608 842430
rect 77808 842250 77864 842306
rect 77932 842250 77988 842306
rect 78056 842250 78112 842306
rect 78180 842250 78236 842306
rect 78304 842250 78360 842306
rect 78428 842250 78484 842306
rect 78552 842250 78608 842306
rect 77808 842126 77864 842182
rect 77932 842126 77988 842182
rect 78056 842126 78112 842182
rect 78180 842126 78236 842182
rect 78304 842126 78360 842182
rect 78428 842126 78484 842182
rect 78552 842126 78608 842182
rect 77808 842002 77864 842058
rect 77932 842002 77988 842058
rect 78056 842002 78112 842058
rect 78180 842002 78236 842058
rect 78304 842002 78360 842058
rect 78428 842002 78484 842058
rect 78552 842002 78608 842058
rect 77808 841878 77864 841934
rect 77932 841878 77988 841934
rect 78056 841878 78112 841934
rect 78180 841878 78236 841934
rect 78304 841878 78360 841934
rect 78428 841878 78484 841934
rect 78552 841878 78608 841934
rect 70074 841128 70130 841184
rect 70074 841004 70130 841060
rect 70074 840880 70130 840936
rect 70074 840756 70130 840812
rect 70074 840632 70130 840688
rect 70074 840508 70130 840564
rect 70074 840384 70130 840440
rect 70074 840260 70130 840316
rect 70074 840136 70130 840192
rect 70074 840012 70130 840068
rect 70074 839888 70130 839944
rect 70074 839764 70130 839820
rect 70074 839640 70130 839696
rect 70074 839516 70130 839572
rect 70074 839392 70130 839448
rect 70074 839268 70130 839324
rect 77808 841134 77864 841190
rect 77932 841134 77988 841190
rect 78056 841134 78112 841190
rect 78180 841134 78236 841190
rect 78304 841134 78360 841190
rect 78428 841134 78484 841190
rect 78552 841134 78608 841190
rect 77808 841010 77864 841066
rect 77932 841010 77988 841066
rect 78056 841010 78112 841066
rect 78180 841010 78236 841066
rect 78304 841010 78360 841066
rect 78428 841010 78484 841066
rect 78552 841010 78608 841066
rect 77808 840886 77864 840942
rect 77932 840886 77988 840942
rect 78056 840886 78112 840942
rect 78180 840886 78236 840942
rect 78304 840886 78360 840942
rect 78428 840886 78484 840942
rect 78552 840886 78608 840942
rect 77808 840762 77864 840818
rect 77932 840762 77988 840818
rect 78056 840762 78112 840818
rect 78180 840762 78236 840818
rect 78304 840762 78360 840818
rect 78428 840762 78484 840818
rect 78552 840762 78608 840818
rect 77808 840638 77864 840694
rect 77932 840638 77988 840694
rect 78056 840638 78112 840694
rect 78180 840638 78236 840694
rect 78304 840638 78360 840694
rect 78428 840638 78484 840694
rect 78552 840638 78608 840694
rect 77808 840514 77864 840570
rect 77932 840514 77988 840570
rect 78056 840514 78112 840570
rect 78180 840514 78236 840570
rect 78304 840514 78360 840570
rect 78428 840514 78484 840570
rect 78552 840514 78608 840570
rect 77808 840390 77864 840446
rect 77932 840390 77988 840446
rect 78056 840390 78112 840446
rect 78180 840390 78236 840446
rect 78304 840390 78360 840446
rect 78428 840390 78484 840446
rect 78552 840390 78608 840446
rect 77808 840266 77864 840322
rect 77932 840266 77988 840322
rect 78056 840266 78112 840322
rect 78180 840266 78236 840322
rect 78304 840266 78360 840322
rect 78428 840266 78484 840322
rect 78552 840266 78608 840322
rect 77808 840142 77864 840198
rect 77932 840142 77988 840198
rect 78056 840142 78112 840198
rect 78180 840142 78236 840198
rect 78304 840142 78360 840198
rect 78428 840142 78484 840198
rect 78552 840142 78608 840198
rect 77808 840018 77864 840074
rect 77932 840018 77988 840074
rect 78056 840018 78112 840074
rect 78180 840018 78236 840074
rect 78304 840018 78360 840074
rect 78428 840018 78484 840074
rect 78552 840018 78608 840074
rect 77808 839894 77864 839950
rect 77932 839894 77988 839950
rect 78056 839894 78112 839950
rect 78180 839894 78236 839950
rect 78304 839894 78360 839950
rect 78428 839894 78484 839950
rect 78552 839894 78608 839950
rect 77808 839770 77864 839826
rect 77932 839770 77988 839826
rect 78056 839770 78112 839826
rect 78180 839770 78236 839826
rect 78304 839770 78360 839826
rect 78428 839770 78484 839826
rect 78552 839770 78608 839826
rect 77808 839646 77864 839702
rect 77932 839646 77988 839702
rect 78056 839646 78112 839702
rect 78180 839646 78236 839702
rect 78304 839646 78360 839702
rect 78428 839646 78484 839702
rect 78552 839646 78608 839702
rect 77808 839522 77864 839578
rect 77932 839522 77988 839578
rect 78056 839522 78112 839578
rect 78180 839522 78236 839578
rect 78304 839522 78360 839578
rect 78428 839522 78484 839578
rect 78552 839522 78608 839578
rect 77808 839398 77864 839454
rect 77932 839398 77988 839454
rect 78056 839398 78112 839454
rect 78180 839398 78236 839454
rect 78304 839398 78360 839454
rect 78428 839398 78484 839454
rect 78552 839398 78608 839454
rect 77808 839274 77864 839330
rect 77932 839274 77988 839330
rect 78056 839274 78112 839330
rect 78180 839274 78236 839330
rect 78304 839274 78360 839330
rect 78428 839274 78484 839330
rect 78552 839274 78608 839330
rect 70074 838758 70130 838814
rect 70074 838634 70130 838690
rect 70074 838510 70130 838566
rect 70074 838386 70130 838442
rect 70074 838262 70130 838318
rect 70074 838138 70130 838194
rect 70074 838014 70130 838070
rect 70074 837890 70130 837946
rect 70074 837766 70130 837822
rect 70074 837642 70130 837698
rect 70074 837518 70130 837574
rect 70074 837394 70130 837450
rect 70074 837270 70130 837326
rect 70074 837146 70130 837202
rect 70074 837022 70130 837078
rect 70074 836898 70130 836954
rect 77808 838764 77864 838820
rect 77932 838764 77988 838820
rect 78056 838764 78112 838820
rect 78180 838764 78236 838820
rect 78304 838764 78360 838820
rect 78428 838764 78484 838820
rect 78552 838764 78608 838820
rect 77808 838640 77864 838696
rect 77932 838640 77988 838696
rect 78056 838640 78112 838696
rect 78180 838640 78236 838696
rect 78304 838640 78360 838696
rect 78428 838640 78484 838696
rect 78552 838640 78608 838696
rect 77808 838516 77864 838572
rect 77932 838516 77988 838572
rect 78056 838516 78112 838572
rect 78180 838516 78236 838572
rect 78304 838516 78360 838572
rect 78428 838516 78484 838572
rect 78552 838516 78608 838572
rect 77808 838392 77864 838448
rect 77932 838392 77988 838448
rect 78056 838392 78112 838448
rect 78180 838392 78236 838448
rect 78304 838392 78360 838448
rect 78428 838392 78484 838448
rect 78552 838392 78608 838448
rect 77808 838268 77864 838324
rect 77932 838268 77988 838324
rect 78056 838268 78112 838324
rect 78180 838268 78236 838324
rect 78304 838268 78360 838324
rect 78428 838268 78484 838324
rect 78552 838268 78608 838324
rect 77808 838144 77864 838200
rect 77932 838144 77988 838200
rect 78056 838144 78112 838200
rect 78180 838144 78236 838200
rect 78304 838144 78360 838200
rect 78428 838144 78484 838200
rect 78552 838144 78608 838200
rect 77808 838020 77864 838076
rect 77932 838020 77988 838076
rect 78056 838020 78112 838076
rect 78180 838020 78236 838076
rect 78304 838020 78360 838076
rect 78428 838020 78484 838076
rect 78552 838020 78608 838076
rect 77808 837896 77864 837952
rect 77932 837896 77988 837952
rect 78056 837896 78112 837952
rect 78180 837896 78236 837952
rect 78304 837896 78360 837952
rect 78428 837896 78484 837952
rect 78552 837896 78608 837952
rect 77808 837772 77864 837828
rect 77932 837772 77988 837828
rect 78056 837772 78112 837828
rect 78180 837772 78236 837828
rect 78304 837772 78360 837828
rect 78428 837772 78484 837828
rect 78552 837772 78608 837828
rect 77808 837648 77864 837704
rect 77932 837648 77988 837704
rect 78056 837648 78112 837704
rect 78180 837648 78236 837704
rect 78304 837648 78360 837704
rect 78428 837648 78484 837704
rect 78552 837648 78608 837704
rect 77808 837524 77864 837580
rect 77932 837524 77988 837580
rect 78056 837524 78112 837580
rect 78180 837524 78236 837580
rect 78304 837524 78360 837580
rect 78428 837524 78484 837580
rect 78552 837524 78608 837580
rect 77808 837400 77864 837456
rect 77932 837400 77988 837456
rect 78056 837400 78112 837456
rect 78180 837400 78236 837456
rect 78304 837400 78360 837456
rect 78428 837400 78484 837456
rect 78552 837400 78608 837456
rect 77808 837276 77864 837332
rect 77932 837276 77988 837332
rect 78056 837276 78112 837332
rect 78180 837276 78236 837332
rect 78304 837276 78360 837332
rect 78428 837276 78484 837332
rect 78552 837276 78608 837332
rect 77808 837152 77864 837208
rect 77932 837152 77988 837208
rect 78056 837152 78112 837208
rect 78180 837152 78236 837208
rect 78304 837152 78360 837208
rect 78428 837152 78484 837208
rect 78552 837152 78608 837208
rect 77808 837028 77864 837084
rect 77932 837028 77988 837084
rect 78056 837028 78112 837084
rect 78180 837028 78236 837084
rect 78304 837028 78360 837084
rect 78428 837028 78484 837084
rect 78552 837028 78608 837084
rect 77808 836904 77864 836960
rect 77932 836904 77988 836960
rect 78056 836904 78112 836960
rect 78180 836904 78236 836960
rect 78304 836904 78360 836960
rect 78428 836904 78484 836960
rect 78552 836904 78608 836960
rect 70074 836052 70130 836108
rect 70074 835928 70130 835984
rect 70074 835804 70130 835860
rect 70074 835680 70130 835736
rect 70074 835556 70130 835612
rect 70074 835432 70130 835488
rect 70074 835308 70130 835364
rect 70074 835184 70130 835240
rect 70074 835060 70130 835116
rect 70074 834936 70130 834992
rect 70074 834812 70130 834868
rect 70074 834688 70130 834744
rect 70074 834564 70130 834620
rect 70074 834440 70130 834496
rect 70074 834316 70130 834372
rect 70074 834192 70130 834248
rect 77808 836058 77864 836114
rect 77932 836058 77988 836114
rect 78056 836058 78112 836114
rect 78180 836058 78236 836114
rect 78304 836058 78360 836114
rect 78428 836058 78484 836114
rect 78552 836058 78608 836114
rect 77808 835934 77864 835990
rect 77932 835934 77988 835990
rect 78056 835934 78112 835990
rect 78180 835934 78236 835990
rect 78304 835934 78360 835990
rect 78428 835934 78484 835990
rect 78552 835934 78608 835990
rect 77808 835810 77864 835866
rect 77932 835810 77988 835866
rect 78056 835810 78112 835866
rect 78180 835810 78236 835866
rect 78304 835810 78360 835866
rect 78428 835810 78484 835866
rect 78552 835810 78608 835866
rect 77808 835686 77864 835742
rect 77932 835686 77988 835742
rect 78056 835686 78112 835742
rect 78180 835686 78236 835742
rect 78304 835686 78360 835742
rect 78428 835686 78484 835742
rect 78552 835686 78608 835742
rect 77808 835562 77864 835618
rect 77932 835562 77988 835618
rect 78056 835562 78112 835618
rect 78180 835562 78236 835618
rect 78304 835562 78360 835618
rect 78428 835562 78484 835618
rect 78552 835562 78608 835618
rect 77808 835438 77864 835494
rect 77932 835438 77988 835494
rect 78056 835438 78112 835494
rect 78180 835438 78236 835494
rect 78304 835438 78360 835494
rect 78428 835438 78484 835494
rect 78552 835438 78608 835494
rect 77808 835314 77864 835370
rect 77932 835314 77988 835370
rect 78056 835314 78112 835370
rect 78180 835314 78236 835370
rect 78304 835314 78360 835370
rect 78428 835314 78484 835370
rect 78552 835314 78608 835370
rect 77808 835190 77864 835246
rect 77932 835190 77988 835246
rect 78056 835190 78112 835246
rect 78180 835190 78236 835246
rect 78304 835190 78360 835246
rect 78428 835190 78484 835246
rect 78552 835190 78608 835246
rect 77808 835066 77864 835122
rect 77932 835066 77988 835122
rect 78056 835066 78112 835122
rect 78180 835066 78236 835122
rect 78304 835066 78360 835122
rect 78428 835066 78484 835122
rect 78552 835066 78608 835122
rect 77808 834942 77864 834998
rect 77932 834942 77988 834998
rect 78056 834942 78112 834998
rect 78180 834942 78236 834998
rect 78304 834942 78360 834998
rect 78428 834942 78484 834998
rect 78552 834942 78608 834998
rect 77808 834818 77864 834874
rect 77932 834818 77988 834874
rect 78056 834818 78112 834874
rect 78180 834818 78236 834874
rect 78304 834818 78360 834874
rect 78428 834818 78484 834874
rect 78552 834818 78608 834874
rect 77808 834694 77864 834750
rect 77932 834694 77988 834750
rect 78056 834694 78112 834750
rect 78180 834694 78236 834750
rect 78304 834694 78360 834750
rect 78428 834694 78484 834750
rect 78552 834694 78608 834750
rect 77808 834570 77864 834626
rect 77932 834570 77988 834626
rect 78056 834570 78112 834626
rect 78180 834570 78236 834626
rect 78304 834570 78360 834626
rect 78428 834570 78484 834626
rect 78552 834570 78608 834626
rect 77808 834446 77864 834502
rect 77932 834446 77988 834502
rect 78056 834446 78112 834502
rect 78180 834446 78236 834502
rect 78304 834446 78360 834502
rect 78428 834446 78484 834502
rect 78552 834446 78608 834502
rect 77808 834322 77864 834378
rect 77932 834322 77988 834378
rect 78056 834322 78112 834378
rect 78180 834322 78236 834378
rect 78304 834322 78360 834378
rect 78428 834322 78484 834378
rect 78552 834322 78608 834378
rect 77808 834198 77864 834254
rect 77932 834198 77988 834254
rect 78056 834198 78112 834254
rect 78180 834198 78236 834254
rect 78304 834198 78360 834254
rect 78428 834198 78484 834254
rect 78552 834198 78608 834254
rect 70074 833682 70130 833738
rect 70074 833558 70130 833614
rect 70074 833434 70130 833490
rect 70074 833310 70130 833366
rect 70074 833186 70130 833242
rect 70074 833062 70130 833118
rect 70074 832938 70130 832994
rect 70074 832814 70130 832870
rect 70074 832690 70130 832746
rect 70074 832566 70130 832622
rect 70074 832442 70130 832498
rect 70074 832318 70130 832374
rect 70074 832194 70130 832250
rect 70074 832070 70130 832126
rect 70074 831946 70130 832002
rect 70074 831822 70130 831878
rect 77808 833688 77864 833744
rect 77932 833688 77988 833744
rect 78056 833688 78112 833744
rect 78180 833688 78236 833744
rect 78304 833688 78360 833744
rect 78428 833688 78484 833744
rect 78552 833688 78608 833744
rect 77808 833564 77864 833620
rect 77932 833564 77988 833620
rect 78056 833564 78112 833620
rect 78180 833564 78236 833620
rect 78304 833564 78360 833620
rect 78428 833564 78484 833620
rect 78552 833564 78608 833620
rect 77808 833440 77864 833496
rect 77932 833440 77988 833496
rect 78056 833440 78112 833496
rect 78180 833440 78236 833496
rect 78304 833440 78360 833496
rect 78428 833440 78484 833496
rect 78552 833440 78608 833496
rect 77808 833316 77864 833372
rect 77932 833316 77988 833372
rect 78056 833316 78112 833372
rect 78180 833316 78236 833372
rect 78304 833316 78360 833372
rect 78428 833316 78484 833372
rect 78552 833316 78608 833372
rect 77808 833192 77864 833248
rect 77932 833192 77988 833248
rect 78056 833192 78112 833248
rect 78180 833192 78236 833248
rect 78304 833192 78360 833248
rect 78428 833192 78484 833248
rect 78552 833192 78608 833248
rect 77808 833068 77864 833124
rect 77932 833068 77988 833124
rect 78056 833068 78112 833124
rect 78180 833068 78236 833124
rect 78304 833068 78360 833124
rect 78428 833068 78484 833124
rect 78552 833068 78608 833124
rect 77808 832944 77864 833000
rect 77932 832944 77988 833000
rect 78056 832944 78112 833000
rect 78180 832944 78236 833000
rect 78304 832944 78360 833000
rect 78428 832944 78484 833000
rect 78552 832944 78608 833000
rect 77808 832820 77864 832876
rect 77932 832820 77988 832876
rect 78056 832820 78112 832876
rect 78180 832820 78236 832876
rect 78304 832820 78360 832876
rect 78428 832820 78484 832876
rect 78552 832820 78608 832876
rect 77808 832696 77864 832752
rect 77932 832696 77988 832752
rect 78056 832696 78112 832752
rect 78180 832696 78236 832752
rect 78304 832696 78360 832752
rect 78428 832696 78484 832752
rect 78552 832696 78608 832752
rect 77808 832572 77864 832628
rect 77932 832572 77988 832628
rect 78056 832572 78112 832628
rect 78180 832572 78236 832628
rect 78304 832572 78360 832628
rect 78428 832572 78484 832628
rect 78552 832572 78608 832628
rect 77808 832448 77864 832504
rect 77932 832448 77988 832504
rect 78056 832448 78112 832504
rect 78180 832448 78236 832504
rect 78304 832448 78360 832504
rect 78428 832448 78484 832504
rect 78552 832448 78608 832504
rect 77808 832324 77864 832380
rect 77932 832324 77988 832380
rect 78056 832324 78112 832380
rect 78180 832324 78236 832380
rect 78304 832324 78360 832380
rect 78428 832324 78484 832380
rect 78552 832324 78608 832380
rect 77808 832200 77864 832256
rect 77932 832200 77988 832256
rect 78056 832200 78112 832256
rect 78180 832200 78236 832256
rect 78304 832200 78360 832256
rect 78428 832200 78484 832256
rect 78552 832200 78608 832256
rect 77808 832076 77864 832132
rect 77932 832076 77988 832132
rect 78056 832076 78112 832132
rect 78180 832076 78236 832132
rect 78304 832076 78360 832132
rect 78428 832076 78484 832132
rect 78552 832076 78608 832132
rect 77808 831952 77864 832008
rect 77932 831952 77988 832008
rect 78056 831952 78112 832008
rect 78180 831952 78236 832008
rect 78304 831952 78360 832008
rect 78428 831952 78484 832008
rect 78552 831952 78608 832008
rect 77808 831828 77864 831884
rect 77932 831828 77988 831884
rect 78056 831828 78112 831884
rect 78180 831828 78236 831884
rect 78304 831828 78360 831884
rect 78428 831828 78484 831884
rect 78552 831828 78608 831884
rect 70074 831078 70130 831134
rect 70074 830954 70130 831010
rect 70074 830830 70130 830886
rect 70074 830706 70130 830762
rect 70074 830582 70130 830638
rect 70074 830458 70130 830514
rect 70074 830334 70130 830390
rect 70074 830210 70130 830266
rect 70074 830086 70130 830142
rect 70074 829962 70130 830018
rect 70074 829838 70130 829894
rect 70074 829714 70130 829770
rect 70074 829590 70130 829646
rect 70074 829466 70130 829522
rect 70074 829342 70130 829398
rect 77808 831084 77864 831140
rect 77932 831084 77988 831140
rect 78056 831084 78112 831140
rect 78180 831084 78236 831140
rect 78304 831084 78360 831140
rect 78428 831084 78484 831140
rect 78552 831084 78608 831140
rect 77808 830960 77864 831016
rect 77932 830960 77988 831016
rect 78056 830960 78112 831016
rect 78180 830960 78236 831016
rect 78304 830960 78360 831016
rect 78428 830960 78484 831016
rect 78552 830960 78608 831016
rect 77808 830836 77864 830892
rect 77932 830836 77988 830892
rect 78056 830836 78112 830892
rect 78180 830836 78236 830892
rect 78304 830836 78360 830892
rect 78428 830836 78484 830892
rect 78552 830836 78608 830892
rect 77808 830712 77864 830768
rect 77932 830712 77988 830768
rect 78056 830712 78112 830768
rect 78180 830712 78236 830768
rect 78304 830712 78360 830768
rect 78428 830712 78484 830768
rect 78552 830712 78608 830768
rect 77808 830588 77864 830644
rect 77932 830588 77988 830644
rect 78056 830588 78112 830644
rect 78180 830588 78236 830644
rect 78304 830588 78360 830644
rect 78428 830588 78484 830644
rect 78552 830588 78608 830644
rect 77808 830464 77864 830520
rect 77932 830464 77988 830520
rect 78056 830464 78112 830520
rect 78180 830464 78236 830520
rect 78304 830464 78360 830520
rect 78428 830464 78484 830520
rect 78552 830464 78608 830520
rect 77808 830340 77864 830396
rect 77932 830340 77988 830396
rect 78056 830340 78112 830396
rect 78180 830340 78236 830396
rect 78304 830340 78360 830396
rect 78428 830340 78484 830396
rect 78552 830340 78608 830396
rect 77808 830216 77864 830272
rect 77932 830216 77988 830272
rect 78056 830216 78112 830272
rect 78180 830216 78236 830272
rect 78304 830216 78360 830272
rect 78428 830216 78484 830272
rect 78552 830216 78608 830272
rect 77808 830092 77864 830148
rect 77932 830092 77988 830148
rect 78056 830092 78112 830148
rect 78180 830092 78236 830148
rect 78304 830092 78360 830148
rect 78428 830092 78484 830148
rect 78552 830092 78608 830148
rect 77808 829968 77864 830024
rect 77932 829968 77988 830024
rect 78056 829968 78112 830024
rect 78180 829968 78236 830024
rect 78304 829968 78360 830024
rect 78428 829968 78484 830024
rect 78552 829968 78608 830024
rect 77808 829844 77864 829900
rect 77932 829844 77988 829900
rect 78056 829844 78112 829900
rect 78180 829844 78236 829900
rect 78304 829844 78360 829900
rect 78428 829844 78484 829900
rect 78552 829844 78608 829900
rect 77808 829720 77864 829776
rect 77932 829720 77988 829776
rect 78056 829720 78112 829776
rect 78180 829720 78236 829776
rect 78304 829720 78360 829776
rect 78428 829720 78484 829776
rect 78552 829720 78608 829776
rect 77808 829596 77864 829652
rect 77932 829596 77988 829652
rect 78056 829596 78112 829652
rect 78180 829596 78236 829652
rect 78304 829596 78360 829652
rect 78428 829596 78484 829652
rect 78552 829596 78608 829652
rect 77808 829472 77864 829528
rect 77932 829472 77988 829528
rect 78056 829472 78112 829528
rect 78180 829472 78236 829528
rect 78304 829472 78360 829528
rect 78428 829472 78484 829528
rect 78552 829472 78608 829528
rect 77808 829348 77864 829404
rect 77932 829348 77988 829404
rect 78056 829348 78112 829404
rect 78180 829348 78236 829404
rect 78304 829348 78360 829404
rect 78428 829348 78484 829404
rect 78552 829348 78608 829404
rect 77800 806373 77856 806429
rect 78100 806373 78156 806429
rect 78400 806373 78456 806429
rect 77800 806173 77856 806229
rect 78100 806173 78156 806229
rect 78400 806173 78456 806229
rect 70074 802602 70130 802658
rect 70074 802478 70130 802534
rect 70074 802354 70130 802410
rect 70074 802230 70130 802286
rect 70074 802106 70130 802162
rect 70074 801982 70130 802038
rect 70074 801858 70130 801914
rect 70074 801734 70130 801790
rect 70074 801610 70130 801666
rect 70074 801486 70130 801542
rect 70074 801362 70130 801418
rect 70074 801238 70130 801294
rect 70074 801114 70130 801170
rect 70074 800990 70130 801046
rect 70074 800866 70130 800922
rect 70074 800128 70130 800184
rect 70074 800004 70130 800060
rect 70074 799880 70130 799936
rect 70074 799756 70130 799812
rect 70074 799632 70130 799688
rect 70074 799508 70130 799564
rect 70074 799384 70130 799440
rect 70074 799260 70130 799316
rect 70074 799136 70130 799192
rect 70074 799012 70130 799068
rect 70074 798888 70130 798944
rect 70074 798764 70130 798820
rect 70074 798640 70130 798696
rect 70074 798516 70130 798572
rect 70074 798392 70130 798448
rect 70074 798268 70130 798324
rect 70074 797758 70130 797814
rect 70074 797634 70130 797690
rect 70074 797510 70130 797566
rect 70074 797386 70130 797442
rect 70074 797262 70130 797318
rect 70074 797138 70130 797194
rect 70074 797014 70130 797070
rect 70074 796890 70130 796946
rect 70074 796766 70130 796822
rect 70074 796642 70130 796698
rect 70074 796518 70130 796574
rect 70074 796394 70130 796450
rect 70074 796270 70130 796326
rect 70074 796146 70130 796202
rect 70074 796022 70130 796078
rect 70074 795898 70130 795954
rect 70074 795052 70130 795108
rect 70074 794928 70130 794984
rect 70074 794804 70130 794860
rect 70074 794680 70130 794736
rect 70074 794556 70130 794612
rect 70074 794432 70130 794488
rect 70074 794308 70130 794364
rect 70074 794184 70130 794240
rect 70074 794060 70130 794116
rect 70074 793936 70130 793992
rect 70074 793812 70130 793868
rect 70074 793688 70130 793744
rect 70074 793564 70130 793620
rect 70074 793440 70130 793496
rect 70074 793316 70130 793372
rect 70074 793192 70130 793248
rect 70074 792682 70130 792738
rect 70074 792558 70130 792614
rect 70074 792434 70130 792490
rect 70074 792310 70130 792366
rect 70074 792186 70130 792242
rect 70074 792062 70130 792118
rect 70074 791938 70130 791994
rect 70074 791814 70130 791870
rect 70074 791690 70130 791746
rect 70074 791566 70130 791622
rect 70074 791442 70130 791498
rect 70074 791318 70130 791374
rect 70074 791194 70130 791250
rect 70074 791070 70130 791126
rect 70074 790946 70130 791002
rect 70074 790822 70130 790878
rect 70074 790078 70130 790134
rect 70074 789954 70130 790010
rect 70074 789830 70130 789886
rect 70074 789706 70130 789762
rect 70074 789582 70130 789638
rect 70074 789458 70130 789514
rect 70074 789334 70130 789390
rect 70074 789210 70130 789266
rect 70074 789086 70130 789142
rect 70074 788962 70130 789018
rect 70074 788838 70130 788894
rect 70074 788714 70130 788770
rect 70074 788590 70130 788646
rect 70074 788466 70130 788522
rect 70074 788342 70130 788398
rect 77847 781577 77903 781633
rect 78147 781577 78203 781633
rect 78447 781577 78503 781633
rect 77800 770373 77856 770429
rect 78100 770373 78156 770429
rect 78400 770373 78456 770429
rect 77800 770173 77856 770229
rect 78100 770173 78156 770229
rect 78400 770173 78456 770229
rect 77900 762046 77956 762102
rect 78200 762046 78256 762102
rect 78500 762046 78556 762102
rect 77900 755046 77956 755102
rect 78200 755046 78256 755102
rect 78500 755046 78556 755102
rect 77900 748046 77956 748102
rect 78200 748046 78256 748102
rect 78500 748046 78556 748102
rect 77847 740577 77903 740633
rect 78147 740577 78203 740633
rect 78447 740577 78503 740633
rect 77800 734373 77856 734429
rect 78100 734373 78156 734429
rect 78400 734373 78456 734429
rect 77800 734173 77856 734229
rect 78100 734173 78156 734229
rect 78400 734173 78456 734229
rect 77900 721046 77956 721102
rect 78200 721046 78256 721102
rect 78500 721046 78556 721102
rect 77900 714046 77956 714102
rect 78200 714046 78256 714102
rect 78500 714046 78556 714102
rect 77900 707046 77956 707102
rect 78200 707046 78256 707102
rect 78500 707046 78556 707102
rect 77847 699577 77903 699633
rect 78147 699577 78203 699633
rect 78447 699577 78503 699633
rect 77800 698373 77856 698429
rect 78100 698373 78156 698429
rect 78400 698373 78456 698429
rect 77800 698173 77856 698229
rect 78100 698173 78156 698229
rect 78400 698173 78456 698229
rect 77900 680046 77956 680102
rect 78200 680046 78256 680102
rect 78500 680046 78556 680102
rect 77900 673046 77956 673102
rect 78200 673046 78256 673102
rect 78500 673046 78556 673102
rect 77900 666046 77956 666102
rect 78200 666046 78256 666102
rect 78500 666046 78556 666102
rect 77800 662373 77856 662429
rect 78100 662373 78156 662429
rect 78400 662373 78456 662429
rect 77800 662173 77856 662229
rect 78100 662173 78156 662229
rect 78400 662173 78456 662229
rect 77847 658577 77903 658633
rect 78147 658577 78203 658633
rect 78447 658577 78503 658633
rect 77900 639046 77956 639102
rect 78200 639046 78256 639102
rect 78500 639046 78556 639102
rect 77900 632046 77956 632102
rect 78200 632046 78256 632102
rect 78500 632046 78556 632102
rect 77800 626373 77856 626429
rect 78100 626373 78156 626429
rect 78400 626373 78456 626429
rect 77800 626173 77856 626229
rect 78100 626173 78156 626229
rect 78400 626173 78456 626229
rect 77900 625046 77956 625102
rect 78200 625046 78256 625102
rect 78500 625046 78556 625102
rect 77847 617577 77903 617633
rect 78147 617577 78203 617633
rect 78447 617577 78503 617633
rect 77900 598046 77956 598102
rect 78200 598046 78256 598102
rect 78500 598046 78556 598102
rect 77900 591046 77956 591102
rect 78200 591046 78256 591102
rect 78500 591046 78556 591102
rect 77800 590373 77856 590429
rect 78100 590373 78156 590429
rect 78400 590373 78456 590429
rect 77800 590173 77856 590229
rect 78100 590173 78156 590229
rect 78400 590173 78456 590229
rect 77900 584046 77956 584102
rect 78200 584046 78256 584102
rect 78500 584046 78556 584102
rect 77847 576577 77903 576633
rect 78147 576577 78203 576633
rect 78447 576577 78503 576633
rect 77900 557046 77956 557102
rect 78200 557046 78256 557102
rect 78500 557046 78556 557102
rect 77800 554373 77856 554429
rect 78100 554373 78156 554429
rect 78400 554373 78456 554429
rect 77800 554173 77856 554229
rect 78100 554173 78156 554229
rect 78400 554173 78456 554229
rect 77900 550046 77956 550102
rect 78200 550046 78256 550102
rect 78500 550046 78556 550102
rect 77900 543046 77956 543102
rect 78200 543046 78256 543102
rect 78500 543046 78556 543102
rect 77847 535577 77903 535633
rect 78147 535577 78203 535633
rect 78447 535577 78503 535633
rect 77800 518373 77856 518429
rect 78100 518373 78156 518429
rect 78400 518373 78456 518429
rect 77800 518173 77856 518229
rect 78100 518173 78156 518229
rect 78400 518173 78456 518229
rect 77900 516046 77956 516102
rect 78200 516046 78256 516102
rect 78500 516046 78556 516102
rect 77900 509046 77956 509102
rect 78200 509046 78256 509102
rect 78500 509046 78556 509102
rect 77900 502046 77956 502102
rect 78200 502046 78256 502102
rect 78500 502046 78556 502102
rect 77800 482373 77856 482429
rect 78100 482373 78156 482429
rect 78400 482373 78456 482429
rect 77800 482173 77856 482229
rect 78100 482173 78156 482229
rect 78400 482173 78456 482229
rect 70074 474602 70130 474658
rect 70074 474478 70130 474534
rect 70074 474354 70130 474410
rect 70074 474230 70130 474286
rect 70074 474106 70130 474162
rect 70074 473982 70130 474038
rect 70074 473858 70130 473914
rect 70074 473734 70130 473790
rect 70074 473610 70130 473666
rect 70074 473486 70130 473542
rect 70074 473362 70130 473418
rect 70074 473238 70130 473294
rect 70074 473114 70130 473170
rect 70074 472990 70130 473046
rect 70074 472866 70130 472922
rect 77808 474614 77864 474670
rect 77932 474614 77988 474670
rect 78056 474614 78112 474670
rect 78180 474614 78236 474670
rect 78304 474614 78360 474670
rect 78428 474614 78484 474670
rect 78552 474614 78608 474670
rect 77808 474490 77864 474546
rect 77932 474490 77988 474546
rect 78056 474490 78112 474546
rect 78180 474490 78236 474546
rect 78304 474490 78360 474546
rect 78428 474490 78484 474546
rect 78552 474490 78608 474546
rect 77808 474366 77864 474422
rect 77932 474366 77988 474422
rect 78056 474366 78112 474422
rect 78180 474366 78236 474422
rect 78304 474366 78360 474422
rect 78428 474366 78484 474422
rect 78552 474366 78608 474422
rect 77808 474242 77864 474298
rect 77932 474242 77988 474298
rect 78056 474242 78112 474298
rect 78180 474242 78236 474298
rect 78304 474242 78360 474298
rect 78428 474242 78484 474298
rect 78552 474242 78608 474298
rect 77808 474118 77864 474174
rect 77932 474118 77988 474174
rect 78056 474118 78112 474174
rect 78180 474118 78236 474174
rect 78304 474118 78360 474174
rect 78428 474118 78484 474174
rect 78552 474118 78608 474174
rect 77808 473994 77864 474050
rect 77932 473994 77988 474050
rect 78056 473994 78112 474050
rect 78180 473994 78236 474050
rect 78304 473994 78360 474050
rect 78428 473994 78484 474050
rect 78552 473994 78608 474050
rect 77808 473870 77864 473926
rect 77932 473870 77988 473926
rect 78056 473870 78112 473926
rect 78180 473870 78236 473926
rect 78304 473870 78360 473926
rect 78428 473870 78484 473926
rect 78552 473870 78608 473926
rect 77808 473746 77864 473802
rect 77932 473746 77988 473802
rect 78056 473746 78112 473802
rect 78180 473746 78236 473802
rect 78304 473746 78360 473802
rect 78428 473746 78484 473802
rect 78552 473746 78608 473802
rect 77808 473622 77864 473678
rect 77932 473622 77988 473678
rect 78056 473622 78112 473678
rect 78180 473622 78236 473678
rect 78304 473622 78360 473678
rect 78428 473622 78484 473678
rect 78552 473622 78608 473678
rect 77808 473498 77864 473554
rect 77932 473498 77988 473554
rect 78056 473498 78112 473554
rect 78180 473498 78236 473554
rect 78304 473498 78360 473554
rect 78428 473498 78484 473554
rect 78552 473498 78608 473554
rect 77808 473374 77864 473430
rect 77932 473374 77988 473430
rect 78056 473374 78112 473430
rect 78180 473374 78236 473430
rect 78304 473374 78360 473430
rect 78428 473374 78484 473430
rect 78552 473374 78608 473430
rect 77808 473250 77864 473306
rect 77932 473250 77988 473306
rect 78056 473250 78112 473306
rect 78180 473250 78236 473306
rect 78304 473250 78360 473306
rect 78428 473250 78484 473306
rect 78552 473250 78608 473306
rect 77808 473126 77864 473182
rect 77932 473126 77988 473182
rect 78056 473126 78112 473182
rect 78180 473126 78236 473182
rect 78304 473126 78360 473182
rect 78428 473126 78484 473182
rect 78552 473126 78608 473182
rect 77808 473002 77864 473058
rect 77932 473002 77988 473058
rect 78056 473002 78112 473058
rect 78180 473002 78236 473058
rect 78304 473002 78360 473058
rect 78428 473002 78484 473058
rect 78552 473002 78608 473058
rect 77808 472878 77864 472934
rect 77932 472878 77988 472934
rect 78056 472878 78112 472934
rect 78180 472878 78236 472934
rect 78304 472878 78360 472934
rect 78428 472878 78484 472934
rect 78552 472878 78608 472934
rect 70074 472128 70130 472184
rect 70074 472004 70130 472060
rect 70074 471880 70130 471936
rect 70074 471756 70130 471812
rect 70074 471632 70130 471688
rect 70074 471508 70130 471564
rect 70074 471384 70130 471440
rect 70074 471260 70130 471316
rect 70074 471136 70130 471192
rect 70074 471012 70130 471068
rect 70074 470888 70130 470944
rect 70074 470764 70130 470820
rect 70074 470640 70130 470696
rect 70074 470516 70130 470572
rect 70074 470392 70130 470448
rect 70074 470268 70130 470324
rect 77808 472134 77864 472190
rect 77932 472134 77988 472190
rect 78056 472134 78112 472190
rect 78180 472134 78236 472190
rect 78304 472134 78360 472190
rect 78428 472134 78484 472190
rect 78552 472134 78608 472190
rect 77808 472010 77864 472066
rect 77932 472010 77988 472066
rect 78056 472010 78112 472066
rect 78180 472010 78236 472066
rect 78304 472010 78360 472066
rect 78428 472010 78484 472066
rect 78552 472010 78608 472066
rect 77808 471886 77864 471942
rect 77932 471886 77988 471942
rect 78056 471886 78112 471942
rect 78180 471886 78236 471942
rect 78304 471886 78360 471942
rect 78428 471886 78484 471942
rect 78552 471886 78608 471942
rect 77808 471762 77864 471818
rect 77932 471762 77988 471818
rect 78056 471762 78112 471818
rect 78180 471762 78236 471818
rect 78304 471762 78360 471818
rect 78428 471762 78484 471818
rect 78552 471762 78608 471818
rect 77808 471638 77864 471694
rect 77932 471638 77988 471694
rect 78056 471638 78112 471694
rect 78180 471638 78236 471694
rect 78304 471638 78360 471694
rect 78428 471638 78484 471694
rect 78552 471638 78608 471694
rect 77808 471514 77864 471570
rect 77932 471514 77988 471570
rect 78056 471514 78112 471570
rect 78180 471514 78236 471570
rect 78304 471514 78360 471570
rect 78428 471514 78484 471570
rect 78552 471514 78608 471570
rect 77808 471390 77864 471446
rect 77932 471390 77988 471446
rect 78056 471390 78112 471446
rect 78180 471390 78236 471446
rect 78304 471390 78360 471446
rect 78428 471390 78484 471446
rect 78552 471390 78608 471446
rect 77808 471266 77864 471322
rect 77932 471266 77988 471322
rect 78056 471266 78112 471322
rect 78180 471266 78236 471322
rect 78304 471266 78360 471322
rect 78428 471266 78484 471322
rect 78552 471266 78608 471322
rect 77808 471142 77864 471198
rect 77932 471142 77988 471198
rect 78056 471142 78112 471198
rect 78180 471142 78236 471198
rect 78304 471142 78360 471198
rect 78428 471142 78484 471198
rect 78552 471142 78608 471198
rect 77808 471018 77864 471074
rect 77932 471018 77988 471074
rect 78056 471018 78112 471074
rect 78180 471018 78236 471074
rect 78304 471018 78360 471074
rect 78428 471018 78484 471074
rect 78552 471018 78608 471074
rect 77808 470894 77864 470950
rect 77932 470894 77988 470950
rect 78056 470894 78112 470950
rect 78180 470894 78236 470950
rect 78304 470894 78360 470950
rect 78428 470894 78484 470950
rect 78552 470894 78608 470950
rect 77808 470770 77864 470826
rect 77932 470770 77988 470826
rect 78056 470770 78112 470826
rect 78180 470770 78236 470826
rect 78304 470770 78360 470826
rect 78428 470770 78484 470826
rect 78552 470770 78608 470826
rect 77808 470646 77864 470702
rect 77932 470646 77988 470702
rect 78056 470646 78112 470702
rect 78180 470646 78236 470702
rect 78304 470646 78360 470702
rect 78428 470646 78484 470702
rect 78552 470646 78608 470702
rect 77808 470522 77864 470578
rect 77932 470522 77988 470578
rect 78056 470522 78112 470578
rect 78180 470522 78236 470578
rect 78304 470522 78360 470578
rect 78428 470522 78484 470578
rect 78552 470522 78608 470578
rect 77808 470398 77864 470454
rect 77932 470398 77988 470454
rect 78056 470398 78112 470454
rect 78180 470398 78236 470454
rect 78304 470398 78360 470454
rect 78428 470398 78484 470454
rect 78552 470398 78608 470454
rect 77808 470274 77864 470330
rect 77932 470274 77988 470330
rect 78056 470274 78112 470330
rect 78180 470274 78236 470330
rect 78304 470274 78360 470330
rect 78428 470274 78484 470330
rect 78552 470274 78608 470330
rect 70074 469758 70130 469814
rect 70074 469634 70130 469690
rect 70074 469510 70130 469566
rect 70074 469386 70130 469442
rect 70074 469262 70130 469318
rect 70074 469138 70130 469194
rect 70074 469014 70130 469070
rect 70074 468890 70130 468946
rect 70074 468766 70130 468822
rect 70074 468642 70130 468698
rect 70074 468518 70130 468574
rect 70074 468394 70130 468450
rect 70074 468270 70130 468326
rect 70074 468146 70130 468202
rect 70074 468022 70130 468078
rect 70074 467898 70130 467954
rect 77808 469764 77864 469820
rect 77932 469764 77988 469820
rect 78056 469764 78112 469820
rect 78180 469764 78236 469820
rect 78304 469764 78360 469820
rect 78428 469764 78484 469820
rect 78552 469764 78608 469820
rect 77808 469640 77864 469696
rect 77932 469640 77988 469696
rect 78056 469640 78112 469696
rect 78180 469640 78236 469696
rect 78304 469640 78360 469696
rect 78428 469640 78484 469696
rect 78552 469640 78608 469696
rect 77808 469516 77864 469572
rect 77932 469516 77988 469572
rect 78056 469516 78112 469572
rect 78180 469516 78236 469572
rect 78304 469516 78360 469572
rect 78428 469516 78484 469572
rect 78552 469516 78608 469572
rect 77808 469392 77864 469448
rect 77932 469392 77988 469448
rect 78056 469392 78112 469448
rect 78180 469392 78236 469448
rect 78304 469392 78360 469448
rect 78428 469392 78484 469448
rect 78552 469392 78608 469448
rect 77808 469268 77864 469324
rect 77932 469268 77988 469324
rect 78056 469268 78112 469324
rect 78180 469268 78236 469324
rect 78304 469268 78360 469324
rect 78428 469268 78484 469324
rect 78552 469268 78608 469324
rect 77808 469144 77864 469200
rect 77932 469144 77988 469200
rect 78056 469144 78112 469200
rect 78180 469144 78236 469200
rect 78304 469144 78360 469200
rect 78428 469144 78484 469200
rect 78552 469144 78608 469200
rect 77808 469020 77864 469076
rect 77932 469020 77988 469076
rect 78056 469020 78112 469076
rect 78180 469020 78236 469076
rect 78304 469020 78360 469076
rect 78428 469020 78484 469076
rect 78552 469020 78608 469076
rect 77808 468896 77864 468952
rect 77932 468896 77988 468952
rect 78056 468896 78112 468952
rect 78180 468896 78236 468952
rect 78304 468896 78360 468952
rect 78428 468896 78484 468952
rect 78552 468896 78608 468952
rect 77808 468772 77864 468828
rect 77932 468772 77988 468828
rect 78056 468772 78112 468828
rect 78180 468772 78236 468828
rect 78304 468772 78360 468828
rect 78428 468772 78484 468828
rect 78552 468772 78608 468828
rect 77808 468648 77864 468704
rect 77932 468648 77988 468704
rect 78056 468648 78112 468704
rect 78180 468648 78236 468704
rect 78304 468648 78360 468704
rect 78428 468648 78484 468704
rect 78552 468648 78608 468704
rect 77808 468524 77864 468580
rect 77932 468524 77988 468580
rect 78056 468524 78112 468580
rect 78180 468524 78236 468580
rect 78304 468524 78360 468580
rect 78428 468524 78484 468580
rect 78552 468524 78608 468580
rect 77808 468400 77864 468456
rect 77932 468400 77988 468456
rect 78056 468400 78112 468456
rect 78180 468400 78236 468456
rect 78304 468400 78360 468456
rect 78428 468400 78484 468456
rect 78552 468400 78608 468456
rect 77808 468276 77864 468332
rect 77932 468276 77988 468332
rect 78056 468276 78112 468332
rect 78180 468276 78236 468332
rect 78304 468276 78360 468332
rect 78428 468276 78484 468332
rect 78552 468276 78608 468332
rect 77808 468152 77864 468208
rect 77932 468152 77988 468208
rect 78056 468152 78112 468208
rect 78180 468152 78236 468208
rect 78304 468152 78360 468208
rect 78428 468152 78484 468208
rect 78552 468152 78608 468208
rect 77808 468028 77864 468084
rect 77932 468028 77988 468084
rect 78056 468028 78112 468084
rect 78180 468028 78236 468084
rect 78304 468028 78360 468084
rect 78428 468028 78484 468084
rect 78552 468028 78608 468084
rect 77808 467904 77864 467960
rect 77932 467904 77988 467960
rect 78056 467904 78112 467960
rect 78180 467904 78236 467960
rect 78304 467904 78360 467960
rect 78428 467904 78484 467960
rect 78552 467904 78608 467960
rect 70074 467052 70130 467108
rect 70074 466928 70130 466984
rect 70074 466804 70130 466860
rect 70074 466680 70130 466736
rect 70074 466556 70130 466612
rect 70074 466432 70130 466488
rect 70074 466308 70130 466364
rect 70074 466184 70130 466240
rect 70074 466060 70130 466116
rect 70074 465936 70130 465992
rect 70074 465812 70130 465868
rect 70074 465688 70130 465744
rect 70074 465564 70130 465620
rect 70074 465440 70130 465496
rect 70074 465316 70130 465372
rect 70074 465192 70130 465248
rect 77808 467058 77864 467114
rect 77932 467058 77988 467114
rect 78056 467058 78112 467114
rect 78180 467058 78236 467114
rect 78304 467058 78360 467114
rect 78428 467058 78484 467114
rect 78552 467058 78608 467114
rect 77808 466934 77864 466990
rect 77932 466934 77988 466990
rect 78056 466934 78112 466990
rect 78180 466934 78236 466990
rect 78304 466934 78360 466990
rect 78428 466934 78484 466990
rect 78552 466934 78608 466990
rect 77808 466810 77864 466866
rect 77932 466810 77988 466866
rect 78056 466810 78112 466866
rect 78180 466810 78236 466866
rect 78304 466810 78360 466866
rect 78428 466810 78484 466866
rect 78552 466810 78608 466866
rect 77808 466686 77864 466742
rect 77932 466686 77988 466742
rect 78056 466686 78112 466742
rect 78180 466686 78236 466742
rect 78304 466686 78360 466742
rect 78428 466686 78484 466742
rect 78552 466686 78608 466742
rect 77808 466562 77864 466618
rect 77932 466562 77988 466618
rect 78056 466562 78112 466618
rect 78180 466562 78236 466618
rect 78304 466562 78360 466618
rect 78428 466562 78484 466618
rect 78552 466562 78608 466618
rect 77808 466438 77864 466494
rect 77932 466438 77988 466494
rect 78056 466438 78112 466494
rect 78180 466438 78236 466494
rect 78304 466438 78360 466494
rect 78428 466438 78484 466494
rect 78552 466438 78608 466494
rect 77808 466314 77864 466370
rect 77932 466314 77988 466370
rect 78056 466314 78112 466370
rect 78180 466314 78236 466370
rect 78304 466314 78360 466370
rect 78428 466314 78484 466370
rect 78552 466314 78608 466370
rect 77808 466190 77864 466246
rect 77932 466190 77988 466246
rect 78056 466190 78112 466246
rect 78180 466190 78236 466246
rect 78304 466190 78360 466246
rect 78428 466190 78484 466246
rect 78552 466190 78608 466246
rect 77808 466066 77864 466122
rect 77932 466066 77988 466122
rect 78056 466066 78112 466122
rect 78180 466066 78236 466122
rect 78304 466066 78360 466122
rect 78428 466066 78484 466122
rect 78552 466066 78608 466122
rect 77808 465942 77864 465998
rect 77932 465942 77988 465998
rect 78056 465942 78112 465998
rect 78180 465942 78236 465998
rect 78304 465942 78360 465998
rect 78428 465942 78484 465998
rect 78552 465942 78608 465998
rect 77808 465818 77864 465874
rect 77932 465818 77988 465874
rect 78056 465818 78112 465874
rect 78180 465818 78236 465874
rect 78304 465818 78360 465874
rect 78428 465818 78484 465874
rect 78552 465818 78608 465874
rect 77808 465694 77864 465750
rect 77932 465694 77988 465750
rect 78056 465694 78112 465750
rect 78180 465694 78236 465750
rect 78304 465694 78360 465750
rect 78428 465694 78484 465750
rect 78552 465694 78608 465750
rect 77808 465570 77864 465626
rect 77932 465570 77988 465626
rect 78056 465570 78112 465626
rect 78180 465570 78236 465626
rect 78304 465570 78360 465626
rect 78428 465570 78484 465626
rect 78552 465570 78608 465626
rect 77808 465446 77864 465502
rect 77932 465446 77988 465502
rect 78056 465446 78112 465502
rect 78180 465446 78236 465502
rect 78304 465446 78360 465502
rect 78428 465446 78484 465502
rect 78552 465446 78608 465502
rect 77808 465322 77864 465378
rect 77932 465322 77988 465378
rect 78056 465322 78112 465378
rect 78180 465322 78236 465378
rect 78304 465322 78360 465378
rect 78428 465322 78484 465378
rect 78552 465322 78608 465378
rect 77808 465198 77864 465254
rect 77932 465198 77988 465254
rect 78056 465198 78112 465254
rect 78180 465198 78236 465254
rect 78304 465198 78360 465254
rect 78428 465198 78484 465254
rect 78552 465198 78608 465254
rect 70074 464682 70130 464738
rect 70074 464558 70130 464614
rect 70074 464434 70130 464490
rect 70074 464310 70130 464366
rect 70074 464186 70130 464242
rect 70074 464062 70130 464118
rect 70074 463938 70130 463994
rect 70074 463814 70130 463870
rect 70074 463690 70130 463746
rect 70074 463566 70130 463622
rect 70074 463442 70130 463498
rect 70074 463318 70130 463374
rect 70074 463194 70130 463250
rect 70074 463070 70130 463126
rect 70074 462946 70130 463002
rect 70074 462822 70130 462878
rect 77808 464688 77864 464744
rect 77932 464688 77988 464744
rect 78056 464688 78112 464744
rect 78180 464688 78236 464744
rect 78304 464688 78360 464744
rect 78428 464688 78484 464744
rect 78552 464688 78608 464744
rect 77808 464564 77864 464620
rect 77932 464564 77988 464620
rect 78056 464564 78112 464620
rect 78180 464564 78236 464620
rect 78304 464564 78360 464620
rect 78428 464564 78484 464620
rect 78552 464564 78608 464620
rect 77808 464440 77864 464496
rect 77932 464440 77988 464496
rect 78056 464440 78112 464496
rect 78180 464440 78236 464496
rect 78304 464440 78360 464496
rect 78428 464440 78484 464496
rect 78552 464440 78608 464496
rect 77808 464316 77864 464372
rect 77932 464316 77988 464372
rect 78056 464316 78112 464372
rect 78180 464316 78236 464372
rect 78304 464316 78360 464372
rect 78428 464316 78484 464372
rect 78552 464316 78608 464372
rect 77808 464192 77864 464248
rect 77932 464192 77988 464248
rect 78056 464192 78112 464248
rect 78180 464192 78236 464248
rect 78304 464192 78360 464248
rect 78428 464192 78484 464248
rect 78552 464192 78608 464248
rect 77808 464068 77864 464124
rect 77932 464068 77988 464124
rect 78056 464068 78112 464124
rect 78180 464068 78236 464124
rect 78304 464068 78360 464124
rect 78428 464068 78484 464124
rect 78552 464068 78608 464124
rect 77808 463944 77864 464000
rect 77932 463944 77988 464000
rect 78056 463944 78112 464000
rect 78180 463944 78236 464000
rect 78304 463944 78360 464000
rect 78428 463944 78484 464000
rect 78552 463944 78608 464000
rect 77808 463820 77864 463876
rect 77932 463820 77988 463876
rect 78056 463820 78112 463876
rect 78180 463820 78236 463876
rect 78304 463820 78360 463876
rect 78428 463820 78484 463876
rect 78552 463820 78608 463876
rect 77808 463696 77864 463752
rect 77932 463696 77988 463752
rect 78056 463696 78112 463752
rect 78180 463696 78236 463752
rect 78304 463696 78360 463752
rect 78428 463696 78484 463752
rect 78552 463696 78608 463752
rect 77808 463572 77864 463628
rect 77932 463572 77988 463628
rect 78056 463572 78112 463628
rect 78180 463572 78236 463628
rect 78304 463572 78360 463628
rect 78428 463572 78484 463628
rect 78552 463572 78608 463628
rect 77808 463448 77864 463504
rect 77932 463448 77988 463504
rect 78056 463448 78112 463504
rect 78180 463448 78236 463504
rect 78304 463448 78360 463504
rect 78428 463448 78484 463504
rect 78552 463448 78608 463504
rect 77808 463324 77864 463380
rect 77932 463324 77988 463380
rect 78056 463324 78112 463380
rect 78180 463324 78236 463380
rect 78304 463324 78360 463380
rect 78428 463324 78484 463380
rect 78552 463324 78608 463380
rect 77808 463200 77864 463256
rect 77932 463200 77988 463256
rect 78056 463200 78112 463256
rect 78180 463200 78236 463256
rect 78304 463200 78360 463256
rect 78428 463200 78484 463256
rect 78552 463200 78608 463256
rect 77808 463076 77864 463132
rect 77932 463076 77988 463132
rect 78056 463076 78112 463132
rect 78180 463076 78236 463132
rect 78304 463076 78360 463132
rect 78428 463076 78484 463132
rect 78552 463076 78608 463132
rect 77808 462952 77864 463008
rect 77932 462952 77988 463008
rect 78056 462952 78112 463008
rect 78180 462952 78236 463008
rect 78304 462952 78360 463008
rect 78428 462952 78484 463008
rect 78552 462952 78608 463008
rect 77808 462828 77864 462884
rect 77932 462828 77988 462884
rect 78056 462828 78112 462884
rect 78180 462828 78236 462884
rect 78304 462828 78360 462884
rect 78428 462828 78484 462884
rect 78552 462828 78608 462884
rect 70074 462078 70130 462134
rect 70074 461954 70130 462010
rect 70074 461830 70130 461886
rect 70074 461706 70130 461762
rect 70074 461582 70130 461638
rect 70074 461458 70130 461514
rect 70074 461334 70130 461390
rect 70074 461210 70130 461266
rect 70074 461086 70130 461142
rect 70074 460962 70130 461018
rect 70074 460838 70130 460894
rect 70074 460714 70130 460770
rect 70074 460590 70130 460646
rect 70074 460466 70130 460522
rect 70074 460342 70130 460398
rect 77808 462084 77864 462140
rect 77932 462084 77988 462140
rect 78056 462084 78112 462140
rect 78180 462084 78236 462140
rect 78304 462084 78360 462140
rect 78428 462084 78484 462140
rect 78552 462084 78608 462140
rect 77808 461960 77864 462016
rect 77932 461960 77988 462016
rect 78056 461960 78112 462016
rect 78180 461960 78236 462016
rect 78304 461960 78360 462016
rect 78428 461960 78484 462016
rect 78552 461960 78608 462016
rect 77808 461836 77864 461892
rect 77932 461836 77988 461892
rect 78056 461836 78112 461892
rect 78180 461836 78236 461892
rect 78304 461836 78360 461892
rect 78428 461836 78484 461892
rect 78552 461836 78608 461892
rect 77808 461712 77864 461768
rect 77932 461712 77988 461768
rect 78056 461712 78112 461768
rect 78180 461712 78236 461768
rect 78304 461712 78360 461768
rect 78428 461712 78484 461768
rect 78552 461712 78608 461768
rect 77808 461588 77864 461644
rect 77932 461588 77988 461644
rect 78056 461588 78112 461644
rect 78180 461588 78236 461644
rect 78304 461588 78360 461644
rect 78428 461588 78484 461644
rect 78552 461588 78608 461644
rect 77808 461464 77864 461520
rect 77932 461464 77988 461520
rect 78056 461464 78112 461520
rect 78180 461464 78236 461520
rect 78304 461464 78360 461520
rect 78428 461464 78484 461520
rect 78552 461464 78608 461520
rect 77808 461340 77864 461396
rect 77932 461340 77988 461396
rect 78056 461340 78112 461396
rect 78180 461340 78236 461396
rect 78304 461340 78360 461396
rect 78428 461340 78484 461396
rect 78552 461340 78608 461396
rect 77808 461216 77864 461272
rect 77932 461216 77988 461272
rect 78056 461216 78112 461272
rect 78180 461216 78236 461272
rect 78304 461216 78360 461272
rect 78428 461216 78484 461272
rect 78552 461216 78608 461272
rect 77808 461092 77864 461148
rect 77932 461092 77988 461148
rect 78056 461092 78112 461148
rect 78180 461092 78236 461148
rect 78304 461092 78360 461148
rect 78428 461092 78484 461148
rect 78552 461092 78608 461148
rect 77808 460968 77864 461024
rect 77932 460968 77988 461024
rect 78056 460968 78112 461024
rect 78180 460968 78236 461024
rect 78304 460968 78360 461024
rect 78428 460968 78484 461024
rect 78552 460968 78608 461024
rect 77808 460844 77864 460900
rect 77932 460844 77988 460900
rect 78056 460844 78112 460900
rect 78180 460844 78236 460900
rect 78304 460844 78360 460900
rect 78428 460844 78484 460900
rect 78552 460844 78608 460900
rect 77808 460720 77864 460776
rect 77932 460720 77988 460776
rect 78056 460720 78112 460776
rect 78180 460720 78236 460776
rect 78304 460720 78360 460776
rect 78428 460720 78484 460776
rect 78552 460720 78608 460776
rect 77808 460596 77864 460652
rect 77932 460596 77988 460652
rect 78056 460596 78112 460652
rect 78180 460596 78236 460652
rect 78304 460596 78360 460652
rect 78428 460596 78484 460652
rect 78552 460596 78608 460652
rect 77808 460472 77864 460528
rect 77932 460472 77988 460528
rect 78056 460472 78112 460528
rect 78180 460472 78236 460528
rect 78304 460472 78360 460528
rect 78428 460472 78484 460528
rect 78552 460472 78608 460528
rect 77808 460348 77864 460404
rect 77932 460348 77988 460404
rect 78056 460348 78112 460404
rect 78180 460348 78236 460404
rect 78304 460348 78360 460404
rect 78428 460348 78484 460404
rect 78552 460348 78608 460404
rect 77800 446373 77856 446429
rect 78100 446373 78156 446429
rect 78400 446373 78456 446429
rect 77800 446173 77856 446229
rect 78100 446173 78156 446229
rect 78400 446173 78456 446229
rect 70074 433602 70130 433658
rect 70074 433478 70130 433534
rect 70074 433354 70130 433410
rect 70074 433230 70130 433286
rect 70074 433106 70130 433162
rect 70074 432982 70130 433038
rect 70074 432858 70130 432914
rect 70074 432734 70130 432790
rect 70074 432610 70130 432666
rect 70074 432486 70130 432542
rect 70074 432362 70130 432418
rect 70074 432238 70130 432294
rect 70074 432114 70130 432170
rect 70074 431990 70130 432046
rect 70074 431866 70130 431922
rect 70074 431128 70130 431184
rect 70074 431004 70130 431060
rect 70074 430880 70130 430936
rect 70074 430756 70130 430812
rect 70074 430632 70130 430688
rect 70074 430508 70130 430564
rect 70074 430384 70130 430440
rect 70074 430260 70130 430316
rect 70074 430136 70130 430192
rect 70074 430012 70130 430068
rect 70074 429888 70130 429944
rect 70074 429764 70130 429820
rect 70074 429640 70130 429696
rect 70074 429516 70130 429572
rect 70074 429392 70130 429448
rect 70074 429268 70130 429324
rect 70074 428758 70130 428814
rect 70074 428634 70130 428690
rect 70074 428510 70130 428566
rect 70074 428386 70130 428442
rect 70074 428262 70130 428318
rect 70074 428138 70130 428194
rect 70074 428014 70130 428070
rect 70074 427890 70130 427946
rect 70074 427766 70130 427822
rect 70074 427642 70130 427698
rect 70074 427518 70130 427574
rect 70074 427394 70130 427450
rect 70074 427270 70130 427326
rect 70074 427146 70130 427202
rect 70074 427022 70130 427078
rect 70074 426898 70130 426954
rect 70074 426052 70130 426108
rect 70074 425928 70130 425984
rect 70074 425804 70130 425860
rect 70074 425680 70130 425736
rect 70074 425556 70130 425612
rect 70074 425432 70130 425488
rect 70074 425308 70130 425364
rect 70074 425184 70130 425240
rect 70074 425060 70130 425116
rect 70074 424936 70130 424992
rect 70074 424812 70130 424868
rect 70074 424688 70130 424744
rect 70074 424564 70130 424620
rect 70074 424440 70130 424496
rect 70074 424316 70130 424372
rect 70074 424192 70130 424248
rect 70074 423682 70130 423738
rect 70074 423558 70130 423614
rect 70074 423434 70130 423490
rect 70074 423310 70130 423366
rect 70074 423186 70130 423242
rect 70074 423062 70130 423118
rect 70074 422938 70130 422994
rect 70074 422814 70130 422870
rect 70074 422690 70130 422746
rect 70074 422566 70130 422622
rect 70074 422442 70130 422498
rect 70074 422318 70130 422374
rect 70074 422194 70130 422250
rect 70074 422070 70130 422126
rect 70074 421946 70130 422002
rect 70074 421822 70130 421878
rect 70074 421078 70130 421134
rect 70074 420954 70130 421010
rect 70074 420830 70130 420886
rect 70074 420706 70130 420762
rect 70074 420582 70130 420638
rect 70074 420458 70130 420514
rect 70074 420334 70130 420390
rect 70074 420210 70130 420266
rect 70074 420086 70130 420142
rect 70074 419962 70130 420018
rect 70074 419838 70130 419894
rect 70074 419714 70130 419770
rect 70074 419590 70130 419646
rect 70074 419466 70130 419522
rect 70074 419342 70130 419398
rect 77847 412577 77903 412633
rect 78147 412577 78203 412633
rect 78447 412577 78503 412633
rect 77800 410373 77856 410429
rect 78100 410373 78156 410429
rect 78400 410373 78456 410429
rect 77800 410173 77856 410229
rect 78100 410173 78156 410229
rect 78400 410173 78456 410229
rect 77900 393046 77956 393102
rect 78200 393046 78256 393102
rect 78500 393046 78556 393102
rect 77900 386046 77956 386102
rect 78200 386046 78256 386102
rect 78500 386046 78556 386102
rect 77900 379046 77956 379102
rect 78200 379046 78256 379102
rect 78500 379046 78556 379102
rect 77800 374373 77856 374429
rect 78100 374373 78156 374429
rect 78400 374373 78456 374429
rect 77800 374173 77856 374229
rect 78100 374173 78156 374229
rect 78400 374173 78456 374229
rect 77847 371577 77903 371633
rect 78147 371577 78203 371633
rect 78447 371577 78503 371633
rect 77900 352046 77956 352102
rect 78200 352046 78256 352102
rect 78500 352046 78556 352102
rect 77900 345046 77956 345102
rect 78200 345046 78256 345102
rect 78500 345046 78556 345102
rect 77800 338373 77856 338429
rect 78100 338373 78156 338429
rect 78400 338373 78456 338429
rect 77800 338173 77856 338229
rect 78100 338173 78156 338229
rect 78400 338173 78456 338229
rect 77900 338046 77956 338102
rect 78200 338046 78256 338102
rect 78500 338046 78556 338102
rect 77847 330577 77903 330633
rect 78147 330577 78203 330633
rect 78447 330577 78503 330633
rect 77808 329584 77864 329640
rect 77932 329584 77988 329640
rect 78056 329584 78112 329640
rect 78180 329584 78236 329640
rect 78304 329584 78360 329640
rect 78428 329584 78484 329640
rect 78552 329584 78608 329640
rect 77808 329460 77864 329516
rect 77932 329460 77988 329516
rect 78056 329460 78112 329516
rect 78180 329460 78236 329516
rect 78304 329460 78360 329516
rect 78428 329460 78484 329516
rect 78552 329460 78608 329516
rect 77808 329336 77864 329392
rect 77932 329336 77988 329392
rect 78056 329336 78112 329392
rect 78180 329336 78236 329392
rect 78304 329336 78360 329392
rect 78428 329336 78484 329392
rect 78552 329336 78608 329392
rect 77808 329212 77864 329268
rect 77932 329212 77988 329268
rect 78056 329212 78112 329268
rect 78180 329212 78236 329268
rect 78304 329212 78360 329268
rect 78428 329212 78484 329268
rect 78552 329212 78608 329268
rect 77808 329088 77864 329144
rect 77932 329088 77988 329144
rect 78056 329088 78112 329144
rect 78180 329088 78236 329144
rect 78304 329088 78360 329144
rect 78428 329088 78484 329144
rect 78552 329088 78608 329144
rect 77808 328964 77864 329020
rect 77932 328964 77988 329020
rect 78056 328964 78112 329020
rect 78180 328964 78236 329020
rect 78304 328964 78360 329020
rect 78428 328964 78484 329020
rect 78552 328964 78608 329020
rect 77808 328840 77864 328896
rect 77932 328840 77988 328896
rect 78056 328840 78112 328896
rect 78180 328840 78236 328896
rect 78304 328840 78360 328896
rect 78428 328840 78484 328896
rect 78552 328840 78608 328896
rect 77900 311046 77956 311102
rect 78200 311046 78256 311102
rect 78500 311046 78556 311102
rect 77808 305730 77864 305786
rect 77932 305730 77988 305786
rect 78056 305730 78112 305786
rect 78180 305730 78236 305786
rect 78304 305730 78360 305786
rect 78428 305730 78484 305786
rect 78552 305730 78608 305786
rect 77808 305606 77864 305662
rect 77932 305606 77988 305662
rect 78056 305606 78112 305662
rect 78180 305606 78236 305662
rect 78304 305606 78360 305662
rect 78428 305606 78484 305662
rect 78552 305606 78608 305662
rect 77808 305482 77864 305538
rect 77932 305482 77988 305538
rect 78056 305482 78112 305538
rect 78180 305482 78236 305538
rect 78304 305482 78360 305538
rect 78428 305482 78484 305538
rect 78552 305482 78608 305538
rect 77808 305358 77864 305414
rect 77932 305358 77988 305414
rect 78056 305358 78112 305414
rect 78180 305358 78236 305414
rect 78304 305358 78360 305414
rect 78428 305358 78484 305414
rect 78552 305358 78608 305414
rect 77808 305234 77864 305290
rect 77932 305234 77988 305290
rect 78056 305234 78112 305290
rect 78180 305234 78236 305290
rect 78304 305234 78360 305290
rect 78428 305234 78484 305290
rect 78552 305234 78608 305290
rect 77808 305110 77864 305166
rect 77932 305110 77988 305166
rect 78056 305110 78112 305166
rect 78180 305110 78236 305166
rect 78304 305110 78360 305166
rect 78428 305110 78484 305166
rect 78552 305110 78608 305166
rect 77808 304986 77864 305042
rect 77932 304986 77988 305042
rect 78056 304986 78112 305042
rect 78180 304986 78236 305042
rect 78304 304986 78360 305042
rect 78428 304986 78484 305042
rect 78552 304986 78608 305042
rect 77800 304066 77856 304122
rect 78100 304066 78156 304122
rect 78400 304066 78456 304122
rect 77900 297046 77956 297102
rect 78200 297046 78256 297102
rect 78500 297046 78556 297102
rect 77847 289577 77903 289633
rect 78147 289577 78203 289633
rect 78447 289577 78503 289633
rect 77808 281916 77864 281972
rect 77932 281916 77988 281972
rect 78056 281916 78112 281972
rect 78180 281916 78236 281972
rect 78304 281916 78360 281972
rect 78428 281916 78484 281972
rect 78552 281916 78608 281972
rect 77808 281792 77864 281848
rect 77932 281792 77988 281848
rect 78056 281792 78112 281848
rect 78180 281792 78236 281848
rect 78304 281792 78360 281848
rect 78428 281792 78484 281848
rect 78552 281792 78608 281848
rect 77808 281668 77864 281724
rect 77932 281668 77988 281724
rect 78056 281668 78112 281724
rect 78180 281668 78236 281724
rect 78304 281668 78360 281724
rect 78428 281668 78484 281724
rect 78552 281668 78608 281724
rect 77808 281544 77864 281600
rect 77932 281544 77988 281600
rect 78056 281544 78112 281600
rect 78180 281544 78236 281600
rect 78304 281544 78360 281600
rect 78428 281544 78484 281600
rect 78552 281544 78608 281600
rect 77808 281420 77864 281476
rect 77932 281420 77988 281476
rect 78056 281420 78112 281476
rect 78180 281420 78236 281476
rect 78304 281420 78360 281476
rect 78428 281420 78484 281476
rect 78552 281420 78608 281476
rect 77808 281296 77864 281352
rect 77932 281296 77988 281352
rect 78056 281296 78112 281352
rect 78180 281296 78236 281352
rect 78304 281296 78360 281352
rect 78428 281296 78484 281352
rect 78552 281296 78608 281352
rect 77808 281172 77864 281228
rect 77932 281172 77988 281228
rect 78056 281172 78112 281228
rect 78180 281172 78236 281228
rect 78304 281172 78360 281228
rect 78428 281172 78484 281228
rect 78552 281172 78608 281228
rect 77900 270046 77956 270102
rect 78200 270046 78256 270102
rect 78500 270046 78556 270102
rect 77748 268316 77804 268372
rect 77872 268316 77928 268372
rect 77996 268316 78052 268372
rect 78120 268316 78176 268372
rect 78244 268316 78300 268372
rect 78368 268316 78424 268372
rect 78492 268316 78548 268372
rect 77748 268192 77804 268248
rect 77872 268192 77928 268248
rect 77996 268192 78052 268248
rect 78120 268192 78176 268248
rect 78244 268192 78300 268248
rect 78368 268192 78424 268248
rect 78492 268192 78548 268248
rect 77900 263046 77956 263102
rect 78200 263046 78256 263102
rect 78500 263046 78556 263102
rect 77900 256046 77956 256102
rect 78200 256046 78256 256102
rect 78500 256046 78556 256102
rect 77847 248577 77903 248633
rect 78147 248577 78203 248633
rect 78447 248577 78503 248633
rect 77748 242316 77804 242372
rect 77872 242316 77928 242372
rect 77996 242316 78052 242372
rect 78120 242316 78176 242372
rect 78244 242316 78300 242372
rect 78368 242316 78424 242372
rect 78492 242316 78548 242372
rect 77748 242192 77804 242248
rect 77872 242192 77928 242248
rect 77996 242192 78052 242248
rect 78120 242192 78176 242248
rect 78244 242192 78300 242248
rect 78368 242192 78424 242248
rect 78492 242192 78548 242248
rect 77900 229046 77956 229102
rect 78200 229046 78256 229102
rect 78500 229046 78556 229102
rect 77900 222046 77956 222102
rect 78200 222046 78256 222102
rect 78500 222046 78556 222102
rect 77748 216316 77804 216372
rect 77872 216316 77928 216372
rect 77996 216316 78052 216372
rect 78120 216316 78176 216372
rect 78244 216316 78300 216372
rect 78368 216316 78424 216372
rect 78492 216316 78548 216372
rect 77748 216192 77804 216248
rect 77872 216192 77928 216248
rect 77996 216192 78052 216248
rect 78120 216192 78176 216248
rect 78244 216192 78300 216248
rect 78368 216192 78424 216248
rect 78492 216192 78548 216248
rect 77900 215046 77956 215102
rect 78200 215046 78256 215102
rect 78500 215046 78556 215102
rect 77847 207577 77903 207633
rect 78147 207577 78203 207633
rect 78447 207577 78503 207633
rect 77748 190316 77804 190372
rect 77872 190316 77928 190372
rect 77996 190316 78052 190372
rect 78120 190316 78176 190372
rect 78244 190316 78300 190372
rect 78368 190316 78424 190372
rect 78492 190316 78548 190372
rect 77748 190192 77804 190248
rect 77872 190192 77928 190248
rect 77996 190192 78052 190248
rect 78120 190192 78176 190248
rect 78244 190192 78300 190248
rect 78368 190192 78424 190248
rect 78492 190192 78548 190248
rect 77900 188046 77956 188102
rect 78200 188046 78256 188102
rect 78500 188046 78556 188102
rect 77900 181046 77956 181102
rect 78200 181046 78256 181102
rect 78500 181046 78556 181102
rect 77900 174046 77956 174102
rect 78200 174046 78256 174102
rect 78500 174046 78556 174102
rect 77748 164316 77804 164372
rect 77872 164316 77928 164372
rect 77996 164316 78052 164372
rect 78120 164316 78176 164372
rect 78244 164316 78300 164372
rect 78368 164316 78424 164372
rect 78492 164316 78548 164372
rect 77748 164192 77804 164248
rect 77872 164192 77928 164248
rect 77996 164192 78052 164248
rect 78120 164192 78176 164248
rect 78244 164192 78300 164248
rect 78368 164192 78424 164248
rect 78492 164192 78548 164248
rect 70074 146602 70130 146658
rect 70074 146478 70130 146534
rect 70074 146354 70130 146410
rect 70074 146230 70130 146286
rect 70074 146106 70130 146162
rect 70074 145982 70130 146038
rect 70074 145858 70130 145914
rect 70074 145734 70130 145790
rect 70074 145610 70130 145666
rect 70074 145486 70130 145542
rect 70074 145362 70130 145418
rect 70074 145238 70130 145294
rect 70074 145114 70130 145170
rect 70074 144990 70130 145046
rect 70074 144866 70130 144922
rect 77808 146614 77864 146670
rect 77932 146614 77988 146670
rect 78056 146614 78112 146670
rect 78180 146614 78236 146670
rect 78304 146614 78360 146670
rect 78428 146614 78484 146670
rect 78552 146614 78608 146670
rect 77808 146490 77864 146546
rect 77932 146490 77988 146546
rect 78056 146490 78112 146546
rect 78180 146490 78236 146546
rect 78304 146490 78360 146546
rect 78428 146490 78484 146546
rect 78552 146490 78608 146546
rect 77808 146366 77864 146422
rect 77932 146366 77988 146422
rect 78056 146366 78112 146422
rect 78180 146366 78236 146422
rect 78304 146366 78360 146422
rect 78428 146366 78484 146422
rect 78552 146366 78608 146422
rect 77808 146242 77864 146298
rect 77932 146242 77988 146298
rect 78056 146242 78112 146298
rect 78180 146242 78236 146298
rect 78304 146242 78360 146298
rect 78428 146242 78484 146298
rect 78552 146242 78608 146298
rect 77808 146118 77864 146174
rect 77932 146118 77988 146174
rect 78056 146118 78112 146174
rect 78180 146118 78236 146174
rect 78304 146118 78360 146174
rect 78428 146118 78484 146174
rect 78552 146118 78608 146174
rect 77808 145994 77864 146050
rect 77932 145994 77988 146050
rect 78056 145994 78112 146050
rect 78180 145994 78236 146050
rect 78304 145994 78360 146050
rect 78428 145994 78484 146050
rect 78552 145994 78608 146050
rect 77808 145870 77864 145926
rect 77932 145870 77988 145926
rect 78056 145870 78112 145926
rect 78180 145870 78236 145926
rect 78304 145870 78360 145926
rect 78428 145870 78484 145926
rect 78552 145870 78608 145926
rect 77808 145746 77864 145802
rect 77932 145746 77988 145802
rect 78056 145746 78112 145802
rect 78180 145746 78236 145802
rect 78304 145746 78360 145802
rect 78428 145746 78484 145802
rect 78552 145746 78608 145802
rect 77808 145622 77864 145678
rect 77932 145622 77988 145678
rect 78056 145622 78112 145678
rect 78180 145622 78236 145678
rect 78304 145622 78360 145678
rect 78428 145622 78484 145678
rect 78552 145622 78608 145678
rect 77808 145498 77864 145554
rect 77932 145498 77988 145554
rect 78056 145498 78112 145554
rect 78180 145498 78236 145554
rect 78304 145498 78360 145554
rect 78428 145498 78484 145554
rect 78552 145498 78608 145554
rect 77808 145374 77864 145430
rect 77932 145374 77988 145430
rect 78056 145374 78112 145430
rect 78180 145374 78236 145430
rect 78304 145374 78360 145430
rect 78428 145374 78484 145430
rect 78552 145374 78608 145430
rect 77808 145250 77864 145306
rect 77932 145250 77988 145306
rect 78056 145250 78112 145306
rect 78180 145250 78236 145306
rect 78304 145250 78360 145306
rect 78428 145250 78484 145306
rect 78552 145250 78608 145306
rect 77808 145126 77864 145182
rect 77932 145126 77988 145182
rect 78056 145126 78112 145182
rect 78180 145126 78236 145182
rect 78304 145126 78360 145182
rect 78428 145126 78484 145182
rect 78552 145126 78608 145182
rect 77808 145002 77864 145058
rect 77932 145002 77988 145058
rect 78056 145002 78112 145058
rect 78180 145002 78236 145058
rect 78304 145002 78360 145058
rect 78428 145002 78484 145058
rect 78552 145002 78608 145058
rect 77808 144878 77864 144934
rect 77932 144878 77988 144934
rect 78056 144878 78112 144934
rect 78180 144878 78236 144934
rect 78304 144878 78360 144934
rect 78428 144878 78484 144934
rect 78552 144878 78608 144934
rect 70074 144128 70130 144184
rect 70074 144004 70130 144060
rect 70074 143880 70130 143936
rect 70074 143756 70130 143812
rect 70074 143632 70130 143688
rect 70074 143508 70130 143564
rect 70074 143384 70130 143440
rect 70074 143260 70130 143316
rect 70074 143136 70130 143192
rect 70074 143012 70130 143068
rect 70074 142888 70130 142944
rect 70074 142764 70130 142820
rect 70074 142640 70130 142696
rect 70074 142516 70130 142572
rect 70074 142392 70130 142448
rect 70074 142268 70130 142324
rect 77808 144134 77864 144190
rect 77932 144134 77988 144190
rect 78056 144134 78112 144190
rect 78180 144134 78236 144190
rect 78304 144134 78360 144190
rect 78428 144134 78484 144190
rect 78552 144134 78608 144190
rect 77808 144010 77864 144066
rect 77932 144010 77988 144066
rect 78056 144010 78112 144066
rect 78180 144010 78236 144066
rect 78304 144010 78360 144066
rect 78428 144010 78484 144066
rect 78552 144010 78608 144066
rect 77808 143886 77864 143942
rect 77932 143886 77988 143942
rect 78056 143886 78112 143942
rect 78180 143886 78236 143942
rect 78304 143886 78360 143942
rect 78428 143886 78484 143942
rect 78552 143886 78608 143942
rect 77808 143762 77864 143818
rect 77932 143762 77988 143818
rect 78056 143762 78112 143818
rect 78180 143762 78236 143818
rect 78304 143762 78360 143818
rect 78428 143762 78484 143818
rect 78552 143762 78608 143818
rect 77808 143638 77864 143694
rect 77932 143638 77988 143694
rect 78056 143638 78112 143694
rect 78180 143638 78236 143694
rect 78304 143638 78360 143694
rect 78428 143638 78484 143694
rect 78552 143638 78608 143694
rect 77808 143514 77864 143570
rect 77932 143514 77988 143570
rect 78056 143514 78112 143570
rect 78180 143514 78236 143570
rect 78304 143514 78360 143570
rect 78428 143514 78484 143570
rect 78552 143514 78608 143570
rect 77808 143390 77864 143446
rect 77932 143390 77988 143446
rect 78056 143390 78112 143446
rect 78180 143390 78236 143446
rect 78304 143390 78360 143446
rect 78428 143390 78484 143446
rect 78552 143390 78608 143446
rect 77808 143266 77864 143322
rect 77932 143266 77988 143322
rect 78056 143266 78112 143322
rect 78180 143266 78236 143322
rect 78304 143266 78360 143322
rect 78428 143266 78484 143322
rect 78552 143266 78608 143322
rect 77808 143142 77864 143198
rect 77932 143142 77988 143198
rect 78056 143142 78112 143198
rect 78180 143142 78236 143198
rect 78304 143142 78360 143198
rect 78428 143142 78484 143198
rect 78552 143142 78608 143198
rect 77808 143018 77864 143074
rect 77932 143018 77988 143074
rect 78056 143018 78112 143074
rect 78180 143018 78236 143074
rect 78304 143018 78360 143074
rect 78428 143018 78484 143074
rect 78552 143018 78608 143074
rect 77808 142894 77864 142950
rect 77932 142894 77988 142950
rect 78056 142894 78112 142950
rect 78180 142894 78236 142950
rect 78304 142894 78360 142950
rect 78428 142894 78484 142950
rect 78552 142894 78608 142950
rect 77808 142770 77864 142826
rect 77932 142770 77988 142826
rect 78056 142770 78112 142826
rect 78180 142770 78236 142826
rect 78304 142770 78360 142826
rect 78428 142770 78484 142826
rect 78552 142770 78608 142826
rect 77808 142646 77864 142702
rect 77932 142646 77988 142702
rect 78056 142646 78112 142702
rect 78180 142646 78236 142702
rect 78304 142646 78360 142702
rect 78428 142646 78484 142702
rect 78552 142646 78608 142702
rect 77808 142522 77864 142578
rect 77932 142522 77988 142578
rect 78056 142522 78112 142578
rect 78180 142522 78236 142578
rect 78304 142522 78360 142578
rect 78428 142522 78484 142578
rect 78552 142522 78608 142578
rect 77808 142398 77864 142454
rect 77932 142398 77988 142454
rect 78056 142398 78112 142454
rect 78180 142398 78236 142454
rect 78304 142398 78360 142454
rect 78428 142398 78484 142454
rect 78552 142398 78608 142454
rect 77808 142274 77864 142330
rect 77932 142274 77988 142330
rect 78056 142274 78112 142330
rect 78180 142274 78236 142330
rect 78304 142274 78360 142330
rect 78428 142274 78484 142330
rect 78552 142274 78608 142330
rect 70074 141758 70130 141814
rect 70074 141634 70130 141690
rect 70074 141510 70130 141566
rect 70074 141386 70130 141442
rect 70074 141262 70130 141318
rect 70074 141138 70130 141194
rect 70074 141014 70130 141070
rect 70074 140890 70130 140946
rect 70074 140766 70130 140822
rect 70074 140642 70130 140698
rect 70074 140518 70130 140574
rect 70074 140394 70130 140450
rect 70074 140270 70130 140326
rect 70074 140146 70130 140202
rect 70074 140022 70130 140078
rect 70074 139898 70130 139954
rect 77808 141764 77864 141820
rect 77932 141764 77988 141820
rect 78056 141764 78112 141820
rect 78180 141764 78236 141820
rect 78304 141764 78360 141820
rect 78428 141764 78484 141820
rect 78552 141764 78608 141820
rect 77808 141640 77864 141696
rect 77932 141640 77988 141696
rect 78056 141640 78112 141696
rect 78180 141640 78236 141696
rect 78304 141640 78360 141696
rect 78428 141640 78484 141696
rect 78552 141640 78608 141696
rect 77808 141516 77864 141572
rect 77932 141516 77988 141572
rect 78056 141516 78112 141572
rect 78180 141516 78236 141572
rect 78304 141516 78360 141572
rect 78428 141516 78484 141572
rect 78552 141516 78608 141572
rect 77808 141392 77864 141448
rect 77932 141392 77988 141448
rect 78056 141392 78112 141448
rect 78180 141392 78236 141448
rect 78304 141392 78360 141448
rect 78428 141392 78484 141448
rect 78552 141392 78608 141448
rect 77808 141268 77864 141324
rect 77932 141268 77988 141324
rect 78056 141268 78112 141324
rect 78180 141268 78236 141324
rect 78304 141268 78360 141324
rect 78428 141268 78484 141324
rect 78552 141268 78608 141324
rect 77808 141144 77864 141200
rect 77932 141144 77988 141200
rect 78056 141144 78112 141200
rect 78180 141144 78236 141200
rect 78304 141144 78360 141200
rect 78428 141144 78484 141200
rect 78552 141144 78608 141200
rect 77808 141020 77864 141076
rect 77932 141020 77988 141076
rect 78056 141020 78112 141076
rect 78180 141020 78236 141076
rect 78304 141020 78360 141076
rect 78428 141020 78484 141076
rect 78552 141020 78608 141076
rect 77808 140896 77864 140952
rect 77932 140896 77988 140952
rect 78056 140896 78112 140952
rect 78180 140896 78236 140952
rect 78304 140896 78360 140952
rect 78428 140896 78484 140952
rect 78552 140896 78608 140952
rect 77808 140772 77864 140828
rect 77932 140772 77988 140828
rect 78056 140772 78112 140828
rect 78180 140772 78236 140828
rect 78304 140772 78360 140828
rect 78428 140772 78484 140828
rect 78552 140772 78608 140828
rect 77808 140648 77864 140704
rect 77932 140648 77988 140704
rect 78056 140648 78112 140704
rect 78180 140648 78236 140704
rect 78304 140648 78360 140704
rect 78428 140648 78484 140704
rect 78552 140648 78608 140704
rect 77808 140524 77864 140580
rect 77932 140524 77988 140580
rect 78056 140524 78112 140580
rect 78180 140524 78236 140580
rect 78304 140524 78360 140580
rect 78428 140524 78484 140580
rect 78552 140524 78608 140580
rect 77808 140400 77864 140456
rect 77932 140400 77988 140456
rect 78056 140400 78112 140456
rect 78180 140400 78236 140456
rect 78304 140400 78360 140456
rect 78428 140400 78484 140456
rect 78552 140400 78608 140456
rect 77808 140276 77864 140332
rect 77932 140276 77988 140332
rect 78056 140276 78112 140332
rect 78180 140276 78236 140332
rect 78304 140276 78360 140332
rect 78428 140276 78484 140332
rect 78552 140276 78608 140332
rect 77808 140152 77864 140208
rect 77932 140152 77988 140208
rect 78056 140152 78112 140208
rect 78180 140152 78236 140208
rect 78304 140152 78360 140208
rect 78428 140152 78484 140208
rect 78552 140152 78608 140208
rect 77808 140028 77864 140084
rect 77932 140028 77988 140084
rect 78056 140028 78112 140084
rect 78180 140028 78236 140084
rect 78304 140028 78360 140084
rect 78428 140028 78484 140084
rect 78552 140028 78608 140084
rect 77808 139904 77864 139960
rect 77932 139904 77988 139960
rect 78056 139904 78112 139960
rect 78180 139904 78236 139960
rect 78304 139904 78360 139960
rect 78428 139904 78484 139960
rect 78552 139904 78608 139960
rect 70074 139052 70130 139108
rect 70074 138928 70130 138984
rect 70074 138804 70130 138860
rect 70074 138680 70130 138736
rect 70074 138556 70130 138612
rect 70074 138432 70130 138488
rect 70074 138308 70130 138364
rect 70074 138184 70130 138240
rect 70074 138060 70130 138116
rect 70074 137936 70130 137992
rect 70074 137812 70130 137868
rect 70074 137688 70130 137744
rect 70074 137564 70130 137620
rect 70074 137440 70130 137496
rect 70074 137316 70130 137372
rect 70074 137192 70130 137248
rect 77808 139058 77864 139114
rect 77932 139058 77988 139114
rect 78056 139058 78112 139114
rect 78180 139058 78236 139114
rect 78304 139058 78360 139114
rect 78428 139058 78484 139114
rect 78552 139058 78608 139114
rect 77808 138934 77864 138990
rect 77932 138934 77988 138990
rect 78056 138934 78112 138990
rect 78180 138934 78236 138990
rect 78304 138934 78360 138990
rect 78428 138934 78484 138990
rect 78552 138934 78608 138990
rect 77808 138810 77864 138866
rect 77932 138810 77988 138866
rect 78056 138810 78112 138866
rect 78180 138810 78236 138866
rect 78304 138810 78360 138866
rect 78428 138810 78484 138866
rect 78552 138810 78608 138866
rect 77808 138686 77864 138742
rect 77932 138686 77988 138742
rect 78056 138686 78112 138742
rect 78180 138686 78236 138742
rect 78304 138686 78360 138742
rect 78428 138686 78484 138742
rect 78552 138686 78608 138742
rect 77808 138562 77864 138618
rect 77932 138562 77988 138618
rect 78056 138562 78112 138618
rect 78180 138562 78236 138618
rect 78304 138562 78360 138618
rect 78428 138562 78484 138618
rect 78552 138562 78608 138618
rect 77808 138438 77864 138494
rect 77932 138438 77988 138494
rect 78056 138438 78112 138494
rect 78180 138438 78236 138494
rect 78304 138438 78360 138494
rect 78428 138438 78484 138494
rect 78552 138438 78608 138494
rect 77808 138314 77864 138370
rect 77932 138314 77988 138370
rect 78056 138314 78112 138370
rect 78180 138314 78236 138370
rect 78304 138314 78360 138370
rect 78428 138314 78484 138370
rect 78552 138314 78608 138370
rect 77808 138190 77864 138246
rect 77932 138190 77988 138246
rect 78056 138190 78112 138246
rect 78180 138190 78236 138246
rect 78304 138190 78360 138246
rect 78428 138190 78484 138246
rect 78552 138190 78608 138246
rect 77808 138066 77864 138122
rect 77932 138066 77988 138122
rect 78056 138066 78112 138122
rect 78180 138066 78236 138122
rect 78304 138066 78360 138122
rect 78428 138066 78484 138122
rect 78552 138066 78608 138122
rect 77808 137942 77864 137998
rect 77932 137942 77988 137998
rect 78056 137942 78112 137998
rect 78180 137942 78236 137998
rect 78304 137942 78360 137998
rect 78428 137942 78484 137998
rect 78552 137942 78608 137998
rect 77808 137818 77864 137874
rect 77932 137818 77988 137874
rect 78056 137818 78112 137874
rect 78180 137818 78236 137874
rect 78304 137818 78360 137874
rect 78428 137818 78484 137874
rect 78552 137818 78608 137874
rect 77808 137694 77864 137750
rect 77932 137694 77988 137750
rect 78056 137694 78112 137750
rect 78180 137694 78236 137750
rect 78304 137694 78360 137750
rect 78428 137694 78484 137750
rect 78552 137694 78608 137750
rect 77808 137570 77864 137626
rect 77932 137570 77988 137626
rect 78056 137570 78112 137626
rect 78180 137570 78236 137626
rect 78304 137570 78360 137626
rect 78428 137570 78484 137626
rect 78552 137570 78608 137626
rect 77808 137446 77864 137502
rect 77932 137446 77988 137502
rect 78056 137446 78112 137502
rect 78180 137446 78236 137502
rect 78304 137446 78360 137502
rect 78428 137446 78484 137502
rect 78552 137446 78608 137502
rect 77808 137322 77864 137378
rect 77932 137322 77988 137378
rect 78056 137322 78112 137378
rect 78180 137322 78236 137378
rect 78304 137322 78360 137378
rect 78428 137322 78484 137378
rect 78552 137322 78608 137378
rect 77808 137198 77864 137254
rect 77932 137198 77988 137254
rect 78056 137198 78112 137254
rect 78180 137198 78236 137254
rect 78304 137198 78360 137254
rect 78428 137198 78484 137254
rect 78552 137198 78608 137254
rect 70074 136682 70130 136738
rect 70074 136558 70130 136614
rect 70074 136434 70130 136490
rect 70074 136310 70130 136366
rect 70074 136186 70130 136242
rect 70074 136062 70130 136118
rect 70074 135938 70130 135994
rect 70074 135814 70130 135870
rect 70074 135690 70130 135746
rect 70074 135566 70130 135622
rect 70074 135442 70130 135498
rect 70074 135318 70130 135374
rect 70074 135194 70130 135250
rect 70074 135070 70130 135126
rect 70074 134946 70130 135002
rect 70074 134822 70130 134878
rect 77808 136688 77864 136744
rect 77932 136688 77988 136744
rect 78056 136688 78112 136744
rect 78180 136688 78236 136744
rect 78304 136688 78360 136744
rect 78428 136688 78484 136744
rect 78552 136688 78608 136744
rect 77808 136564 77864 136620
rect 77932 136564 77988 136620
rect 78056 136564 78112 136620
rect 78180 136564 78236 136620
rect 78304 136564 78360 136620
rect 78428 136564 78484 136620
rect 78552 136564 78608 136620
rect 77808 136440 77864 136496
rect 77932 136440 77988 136496
rect 78056 136440 78112 136496
rect 78180 136440 78236 136496
rect 78304 136440 78360 136496
rect 78428 136440 78484 136496
rect 78552 136440 78608 136496
rect 77808 136316 77864 136372
rect 77932 136316 77988 136372
rect 78056 136316 78112 136372
rect 78180 136316 78236 136372
rect 78304 136316 78360 136372
rect 78428 136316 78484 136372
rect 78552 136316 78608 136372
rect 77808 136192 77864 136248
rect 77932 136192 77988 136248
rect 78056 136192 78112 136248
rect 78180 136192 78236 136248
rect 78304 136192 78360 136248
rect 78428 136192 78484 136248
rect 78552 136192 78608 136248
rect 77808 136068 77864 136124
rect 77932 136068 77988 136124
rect 78056 136068 78112 136124
rect 78180 136068 78236 136124
rect 78304 136068 78360 136124
rect 78428 136068 78484 136124
rect 78552 136068 78608 136124
rect 77808 135944 77864 136000
rect 77932 135944 77988 136000
rect 78056 135944 78112 136000
rect 78180 135944 78236 136000
rect 78304 135944 78360 136000
rect 78428 135944 78484 136000
rect 78552 135944 78608 136000
rect 77808 135820 77864 135876
rect 77932 135820 77988 135876
rect 78056 135820 78112 135876
rect 78180 135820 78236 135876
rect 78304 135820 78360 135876
rect 78428 135820 78484 135876
rect 78552 135820 78608 135876
rect 77808 135696 77864 135752
rect 77932 135696 77988 135752
rect 78056 135696 78112 135752
rect 78180 135696 78236 135752
rect 78304 135696 78360 135752
rect 78428 135696 78484 135752
rect 78552 135696 78608 135752
rect 77808 135572 77864 135628
rect 77932 135572 77988 135628
rect 78056 135572 78112 135628
rect 78180 135572 78236 135628
rect 78304 135572 78360 135628
rect 78428 135572 78484 135628
rect 78552 135572 78608 135628
rect 77808 135448 77864 135504
rect 77932 135448 77988 135504
rect 78056 135448 78112 135504
rect 78180 135448 78236 135504
rect 78304 135448 78360 135504
rect 78428 135448 78484 135504
rect 78552 135448 78608 135504
rect 77808 135324 77864 135380
rect 77932 135324 77988 135380
rect 78056 135324 78112 135380
rect 78180 135324 78236 135380
rect 78304 135324 78360 135380
rect 78428 135324 78484 135380
rect 78552 135324 78608 135380
rect 77808 135200 77864 135256
rect 77932 135200 77988 135256
rect 78056 135200 78112 135256
rect 78180 135200 78236 135256
rect 78304 135200 78360 135256
rect 78428 135200 78484 135256
rect 78552 135200 78608 135256
rect 77808 135076 77864 135132
rect 77932 135076 77988 135132
rect 78056 135076 78112 135132
rect 78180 135076 78236 135132
rect 78304 135076 78360 135132
rect 78428 135076 78484 135132
rect 78552 135076 78608 135132
rect 77808 134952 77864 135008
rect 77932 134952 77988 135008
rect 78056 134952 78112 135008
rect 78180 134952 78236 135008
rect 78304 134952 78360 135008
rect 78428 134952 78484 135008
rect 78552 134952 78608 135008
rect 77808 134828 77864 134884
rect 77932 134828 77988 134884
rect 78056 134828 78112 134884
rect 78180 134828 78236 134884
rect 78304 134828 78360 134884
rect 78428 134828 78484 134884
rect 78552 134828 78608 134884
rect 70074 134078 70130 134134
rect 70074 133954 70130 134010
rect 70074 133830 70130 133886
rect 70074 133706 70130 133762
rect 70074 133582 70130 133638
rect 70074 133458 70130 133514
rect 70074 133334 70130 133390
rect 70074 133210 70130 133266
rect 70074 133086 70130 133142
rect 70074 132962 70130 133018
rect 70074 132838 70130 132894
rect 70074 132714 70130 132770
rect 70074 132590 70130 132646
rect 70074 132466 70130 132522
rect 70074 132342 70130 132398
rect 77808 134084 77864 134140
rect 77932 134084 77988 134140
rect 78056 134084 78112 134140
rect 78180 134084 78236 134140
rect 78304 134084 78360 134140
rect 78428 134084 78484 134140
rect 78552 134084 78608 134140
rect 77808 133960 77864 134016
rect 77932 133960 77988 134016
rect 78056 133960 78112 134016
rect 78180 133960 78236 134016
rect 78304 133960 78360 134016
rect 78428 133960 78484 134016
rect 78552 133960 78608 134016
rect 77808 133836 77864 133892
rect 77932 133836 77988 133892
rect 78056 133836 78112 133892
rect 78180 133836 78236 133892
rect 78304 133836 78360 133892
rect 78428 133836 78484 133892
rect 78552 133836 78608 133892
rect 77808 133712 77864 133768
rect 77932 133712 77988 133768
rect 78056 133712 78112 133768
rect 78180 133712 78236 133768
rect 78304 133712 78360 133768
rect 78428 133712 78484 133768
rect 78552 133712 78608 133768
rect 77808 133588 77864 133644
rect 77932 133588 77988 133644
rect 78056 133588 78112 133644
rect 78180 133588 78236 133644
rect 78304 133588 78360 133644
rect 78428 133588 78484 133644
rect 78552 133588 78608 133644
rect 77808 133464 77864 133520
rect 77932 133464 77988 133520
rect 78056 133464 78112 133520
rect 78180 133464 78236 133520
rect 78304 133464 78360 133520
rect 78428 133464 78484 133520
rect 78552 133464 78608 133520
rect 77808 133340 77864 133396
rect 77932 133340 77988 133396
rect 78056 133340 78112 133396
rect 78180 133340 78236 133396
rect 78304 133340 78360 133396
rect 78428 133340 78484 133396
rect 78552 133340 78608 133396
rect 77808 133216 77864 133272
rect 77932 133216 77988 133272
rect 78056 133216 78112 133272
rect 78180 133216 78236 133272
rect 78304 133216 78360 133272
rect 78428 133216 78484 133272
rect 78552 133216 78608 133272
rect 77808 133092 77864 133148
rect 77932 133092 77988 133148
rect 78056 133092 78112 133148
rect 78180 133092 78236 133148
rect 78304 133092 78360 133148
rect 78428 133092 78484 133148
rect 78552 133092 78608 133148
rect 77808 132968 77864 133024
rect 77932 132968 77988 133024
rect 78056 132968 78112 133024
rect 78180 132968 78236 133024
rect 78304 132968 78360 133024
rect 78428 132968 78484 133024
rect 78552 132968 78608 133024
rect 77808 132844 77864 132900
rect 77932 132844 77988 132900
rect 78056 132844 78112 132900
rect 78180 132844 78236 132900
rect 78304 132844 78360 132900
rect 78428 132844 78484 132900
rect 78552 132844 78608 132900
rect 77808 132720 77864 132776
rect 77932 132720 77988 132776
rect 78056 132720 78112 132776
rect 78180 132720 78236 132776
rect 78304 132720 78360 132776
rect 78428 132720 78484 132776
rect 78552 132720 78608 132776
rect 77808 132596 77864 132652
rect 77932 132596 77988 132652
rect 78056 132596 78112 132652
rect 78180 132596 78236 132652
rect 78304 132596 78360 132652
rect 78428 132596 78484 132652
rect 78552 132596 78608 132652
rect 77808 132472 77864 132528
rect 77932 132472 77988 132528
rect 78056 132472 78112 132528
rect 78180 132472 78236 132528
rect 78304 132472 78360 132528
rect 78428 132472 78484 132528
rect 78552 132472 78608 132528
rect 77808 132348 77864 132404
rect 77932 132348 77988 132404
rect 78056 132348 78112 132404
rect 78180 132348 78236 132404
rect 78304 132348 78360 132404
rect 78428 132348 78484 132404
rect 78552 132348 78608 132404
rect 77748 112316 77804 112372
rect 77872 112316 77928 112372
rect 77996 112316 78052 112372
rect 78120 112316 78176 112372
rect 78244 112316 78300 112372
rect 78368 112316 78424 112372
rect 78492 112316 78548 112372
rect 77748 112192 77804 112248
rect 77872 112192 77928 112248
rect 77996 112192 78052 112248
rect 78120 112192 78176 112248
rect 78244 112192 78300 112248
rect 78368 112192 78424 112248
rect 78492 112192 78548 112248
rect 70074 105602 70130 105658
rect 70074 105478 70130 105534
rect 70074 105354 70130 105410
rect 70074 105230 70130 105286
rect 70074 105106 70130 105162
rect 70074 104982 70130 105038
rect 70074 104858 70130 104914
rect 70074 104734 70130 104790
rect 70074 104610 70130 104666
rect 70074 104486 70130 104542
rect 70074 104362 70130 104418
rect 70074 104238 70130 104294
rect 70074 104114 70130 104170
rect 70074 103990 70130 104046
rect 70074 103866 70130 103922
rect 77808 105614 77864 105670
rect 77932 105614 77988 105670
rect 78056 105614 78112 105670
rect 78180 105614 78236 105670
rect 78304 105614 78360 105670
rect 78428 105614 78484 105670
rect 78552 105614 78608 105670
rect 77808 105490 77864 105546
rect 77932 105490 77988 105546
rect 78056 105490 78112 105546
rect 78180 105490 78236 105546
rect 78304 105490 78360 105546
rect 78428 105490 78484 105546
rect 78552 105490 78608 105546
rect 77808 105366 77864 105422
rect 77932 105366 77988 105422
rect 78056 105366 78112 105422
rect 78180 105366 78236 105422
rect 78304 105366 78360 105422
rect 78428 105366 78484 105422
rect 78552 105366 78608 105422
rect 77808 105242 77864 105298
rect 77932 105242 77988 105298
rect 78056 105242 78112 105298
rect 78180 105242 78236 105298
rect 78304 105242 78360 105298
rect 78428 105242 78484 105298
rect 78552 105242 78608 105298
rect 77808 105118 77864 105174
rect 77932 105118 77988 105174
rect 78056 105118 78112 105174
rect 78180 105118 78236 105174
rect 78304 105118 78360 105174
rect 78428 105118 78484 105174
rect 78552 105118 78608 105174
rect 77808 104994 77864 105050
rect 77932 104994 77988 105050
rect 78056 104994 78112 105050
rect 78180 104994 78236 105050
rect 78304 104994 78360 105050
rect 78428 104994 78484 105050
rect 78552 104994 78608 105050
rect 77808 104870 77864 104926
rect 77932 104870 77988 104926
rect 78056 104870 78112 104926
rect 78180 104870 78236 104926
rect 78304 104870 78360 104926
rect 78428 104870 78484 104926
rect 78552 104870 78608 104926
rect 77808 104746 77864 104802
rect 77932 104746 77988 104802
rect 78056 104746 78112 104802
rect 78180 104746 78236 104802
rect 78304 104746 78360 104802
rect 78428 104746 78484 104802
rect 78552 104746 78608 104802
rect 77808 104622 77864 104678
rect 77932 104622 77988 104678
rect 78056 104622 78112 104678
rect 78180 104622 78236 104678
rect 78304 104622 78360 104678
rect 78428 104622 78484 104678
rect 78552 104622 78608 104678
rect 77808 104498 77864 104554
rect 77932 104498 77988 104554
rect 78056 104498 78112 104554
rect 78180 104498 78236 104554
rect 78304 104498 78360 104554
rect 78428 104498 78484 104554
rect 78552 104498 78608 104554
rect 77808 104374 77864 104430
rect 77932 104374 77988 104430
rect 78056 104374 78112 104430
rect 78180 104374 78236 104430
rect 78304 104374 78360 104430
rect 78428 104374 78484 104430
rect 78552 104374 78608 104430
rect 77808 104250 77864 104306
rect 77932 104250 77988 104306
rect 78056 104250 78112 104306
rect 78180 104250 78236 104306
rect 78304 104250 78360 104306
rect 78428 104250 78484 104306
rect 78552 104250 78608 104306
rect 77808 104126 77864 104182
rect 77932 104126 77988 104182
rect 78056 104126 78112 104182
rect 78180 104126 78236 104182
rect 78304 104126 78360 104182
rect 78428 104126 78484 104182
rect 78552 104126 78608 104182
rect 77808 104002 77864 104058
rect 77932 104002 77988 104058
rect 78056 104002 78112 104058
rect 78180 104002 78236 104058
rect 78304 104002 78360 104058
rect 78428 104002 78484 104058
rect 78552 104002 78608 104058
rect 77808 103878 77864 103934
rect 77932 103878 77988 103934
rect 78056 103878 78112 103934
rect 78180 103878 78236 103934
rect 78304 103878 78360 103934
rect 78428 103878 78484 103934
rect 78552 103878 78608 103934
rect 70074 103128 70130 103184
rect 70074 103004 70130 103060
rect 70074 102880 70130 102936
rect 70074 102756 70130 102812
rect 70074 102632 70130 102688
rect 70074 102508 70130 102564
rect 70074 102384 70130 102440
rect 70074 102260 70130 102316
rect 70074 102136 70130 102192
rect 70074 102012 70130 102068
rect 70074 101888 70130 101944
rect 70074 101764 70130 101820
rect 70074 101640 70130 101696
rect 70074 101516 70130 101572
rect 70074 101392 70130 101448
rect 70074 101268 70130 101324
rect 77808 103134 77864 103190
rect 77932 103134 77988 103190
rect 78056 103134 78112 103190
rect 78180 103134 78236 103190
rect 78304 103134 78360 103190
rect 78428 103134 78484 103190
rect 78552 103134 78608 103190
rect 77808 103010 77864 103066
rect 77932 103010 77988 103066
rect 78056 103010 78112 103066
rect 78180 103010 78236 103066
rect 78304 103010 78360 103066
rect 78428 103010 78484 103066
rect 78552 103010 78608 103066
rect 77808 102886 77864 102942
rect 77932 102886 77988 102942
rect 78056 102886 78112 102942
rect 78180 102886 78236 102942
rect 78304 102886 78360 102942
rect 78428 102886 78484 102942
rect 78552 102886 78608 102942
rect 77808 102762 77864 102818
rect 77932 102762 77988 102818
rect 78056 102762 78112 102818
rect 78180 102762 78236 102818
rect 78304 102762 78360 102818
rect 78428 102762 78484 102818
rect 78552 102762 78608 102818
rect 77808 102638 77864 102694
rect 77932 102638 77988 102694
rect 78056 102638 78112 102694
rect 78180 102638 78236 102694
rect 78304 102638 78360 102694
rect 78428 102638 78484 102694
rect 78552 102638 78608 102694
rect 77808 102514 77864 102570
rect 77932 102514 77988 102570
rect 78056 102514 78112 102570
rect 78180 102514 78236 102570
rect 78304 102514 78360 102570
rect 78428 102514 78484 102570
rect 78552 102514 78608 102570
rect 77808 102390 77864 102446
rect 77932 102390 77988 102446
rect 78056 102390 78112 102446
rect 78180 102390 78236 102446
rect 78304 102390 78360 102446
rect 78428 102390 78484 102446
rect 78552 102390 78608 102446
rect 77808 102266 77864 102322
rect 77932 102266 77988 102322
rect 78056 102266 78112 102322
rect 78180 102266 78236 102322
rect 78304 102266 78360 102322
rect 78428 102266 78484 102322
rect 78552 102266 78608 102322
rect 77808 102142 77864 102198
rect 77932 102142 77988 102198
rect 78056 102142 78112 102198
rect 78180 102142 78236 102198
rect 78304 102142 78360 102198
rect 78428 102142 78484 102198
rect 78552 102142 78608 102198
rect 77808 102018 77864 102074
rect 77932 102018 77988 102074
rect 78056 102018 78112 102074
rect 78180 102018 78236 102074
rect 78304 102018 78360 102074
rect 78428 102018 78484 102074
rect 78552 102018 78608 102074
rect 77808 101894 77864 101950
rect 77932 101894 77988 101950
rect 78056 101894 78112 101950
rect 78180 101894 78236 101950
rect 78304 101894 78360 101950
rect 78428 101894 78484 101950
rect 78552 101894 78608 101950
rect 77808 101770 77864 101826
rect 77932 101770 77988 101826
rect 78056 101770 78112 101826
rect 78180 101770 78236 101826
rect 78304 101770 78360 101826
rect 78428 101770 78484 101826
rect 78552 101770 78608 101826
rect 77808 101646 77864 101702
rect 77932 101646 77988 101702
rect 78056 101646 78112 101702
rect 78180 101646 78236 101702
rect 78304 101646 78360 101702
rect 78428 101646 78484 101702
rect 78552 101646 78608 101702
rect 77808 101522 77864 101578
rect 77932 101522 77988 101578
rect 78056 101522 78112 101578
rect 78180 101522 78236 101578
rect 78304 101522 78360 101578
rect 78428 101522 78484 101578
rect 78552 101522 78608 101578
rect 77808 101398 77864 101454
rect 77932 101398 77988 101454
rect 78056 101398 78112 101454
rect 78180 101398 78236 101454
rect 78304 101398 78360 101454
rect 78428 101398 78484 101454
rect 78552 101398 78608 101454
rect 77808 101274 77864 101330
rect 77932 101274 77988 101330
rect 78056 101274 78112 101330
rect 78180 101274 78236 101330
rect 78304 101274 78360 101330
rect 78428 101274 78484 101330
rect 78552 101274 78608 101330
rect 70074 100758 70130 100814
rect 70074 100634 70130 100690
rect 70074 100510 70130 100566
rect 70074 100386 70130 100442
rect 70074 100262 70130 100318
rect 70074 100138 70130 100194
rect 70074 100014 70130 100070
rect 70074 99890 70130 99946
rect 70074 99766 70130 99822
rect 70074 99642 70130 99698
rect 70074 99518 70130 99574
rect 70074 99394 70130 99450
rect 70074 99270 70130 99326
rect 70074 99146 70130 99202
rect 70074 99022 70130 99078
rect 70074 98898 70130 98954
rect 77808 100764 77864 100820
rect 77932 100764 77988 100820
rect 78056 100764 78112 100820
rect 78180 100764 78236 100820
rect 78304 100764 78360 100820
rect 78428 100764 78484 100820
rect 78552 100764 78608 100820
rect 77808 100640 77864 100696
rect 77932 100640 77988 100696
rect 78056 100640 78112 100696
rect 78180 100640 78236 100696
rect 78304 100640 78360 100696
rect 78428 100640 78484 100696
rect 78552 100640 78608 100696
rect 77808 100516 77864 100572
rect 77932 100516 77988 100572
rect 78056 100516 78112 100572
rect 78180 100516 78236 100572
rect 78304 100516 78360 100572
rect 78428 100516 78484 100572
rect 78552 100516 78608 100572
rect 77808 100392 77864 100448
rect 77932 100392 77988 100448
rect 78056 100392 78112 100448
rect 78180 100392 78236 100448
rect 78304 100392 78360 100448
rect 78428 100392 78484 100448
rect 78552 100392 78608 100448
rect 77808 100268 77864 100324
rect 77932 100268 77988 100324
rect 78056 100268 78112 100324
rect 78180 100268 78236 100324
rect 78304 100268 78360 100324
rect 78428 100268 78484 100324
rect 78552 100268 78608 100324
rect 77808 100144 77864 100200
rect 77932 100144 77988 100200
rect 78056 100144 78112 100200
rect 78180 100144 78236 100200
rect 78304 100144 78360 100200
rect 78428 100144 78484 100200
rect 78552 100144 78608 100200
rect 77808 100020 77864 100076
rect 77932 100020 77988 100076
rect 78056 100020 78112 100076
rect 78180 100020 78236 100076
rect 78304 100020 78360 100076
rect 78428 100020 78484 100076
rect 78552 100020 78608 100076
rect 77808 99896 77864 99952
rect 77932 99896 77988 99952
rect 78056 99896 78112 99952
rect 78180 99896 78236 99952
rect 78304 99896 78360 99952
rect 78428 99896 78484 99952
rect 78552 99896 78608 99952
rect 77808 99772 77864 99828
rect 77932 99772 77988 99828
rect 78056 99772 78112 99828
rect 78180 99772 78236 99828
rect 78304 99772 78360 99828
rect 78428 99772 78484 99828
rect 78552 99772 78608 99828
rect 77808 99648 77864 99704
rect 77932 99648 77988 99704
rect 78056 99648 78112 99704
rect 78180 99648 78236 99704
rect 78304 99648 78360 99704
rect 78428 99648 78484 99704
rect 78552 99648 78608 99704
rect 77808 99524 77864 99580
rect 77932 99524 77988 99580
rect 78056 99524 78112 99580
rect 78180 99524 78236 99580
rect 78304 99524 78360 99580
rect 78428 99524 78484 99580
rect 78552 99524 78608 99580
rect 77808 99400 77864 99456
rect 77932 99400 77988 99456
rect 78056 99400 78112 99456
rect 78180 99400 78236 99456
rect 78304 99400 78360 99456
rect 78428 99400 78484 99456
rect 78552 99400 78608 99456
rect 77808 99276 77864 99332
rect 77932 99276 77988 99332
rect 78056 99276 78112 99332
rect 78180 99276 78236 99332
rect 78304 99276 78360 99332
rect 78428 99276 78484 99332
rect 78552 99276 78608 99332
rect 77808 99152 77864 99208
rect 77932 99152 77988 99208
rect 78056 99152 78112 99208
rect 78180 99152 78236 99208
rect 78304 99152 78360 99208
rect 78428 99152 78484 99208
rect 78552 99152 78608 99208
rect 77808 99028 77864 99084
rect 77932 99028 77988 99084
rect 78056 99028 78112 99084
rect 78180 99028 78236 99084
rect 78304 99028 78360 99084
rect 78428 99028 78484 99084
rect 78552 99028 78608 99084
rect 77808 98904 77864 98960
rect 77932 98904 77988 98960
rect 78056 98904 78112 98960
rect 78180 98904 78236 98960
rect 78304 98904 78360 98960
rect 78428 98904 78484 98960
rect 78552 98904 78608 98960
rect 70074 98052 70130 98108
rect 70074 97928 70130 97984
rect 70074 97804 70130 97860
rect 70074 97680 70130 97736
rect 70074 97556 70130 97612
rect 70074 97432 70130 97488
rect 70074 97308 70130 97364
rect 70074 97184 70130 97240
rect 70074 97060 70130 97116
rect 70074 96936 70130 96992
rect 70074 96812 70130 96868
rect 70074 96688 70130 96744
rect 70074 96564 70130 96620
rect 70074 96440 70130 96496
rect 70074 96316 70130 96372
rect 70074 96192 70130 96248
rect 77808 98058 77864 98114
rect 77932 98058 77988 98114
rect 78056 98058 78112 98114
rect 78180 98058 78236 98114
rect 78304 98058 78360 98114
rect 78428 98058 78484 98114
rect 78552 98058 78608 98114
rect 77808 97934 77864 97990
rect 77932 97934 77988 97990
rect 78056 97934 78112 97990
rect 78180 97934 78236 97990
rect 78304 97934 78360 97990
rect 78428 97934 78484 97990
rect 78552 97934 78608 97990
rect 77808 97810 77864 97866
rect 77932 97810 77988 97866
rect 78056 97810 78112 97866
rect 78180 97810 78236 97866
rect 78304 97810 78360 97866
rect 78428 97810 78484 97866
rect 78552 97810 78608 97866
rect 77808 97686 77864 97742
rect 77932 97686 77988 97742
rect 78056 97686 78112 97742
rect 78180 97686 78236 97742
rect 78304 97686 78360 97742
rect 78428 97686 78484 97742
rect 78552 97686 78608 97742
rect 77808 97562 77864 97618
rect 77932 97562 77988 97618
rect 78056 97562 78112 97618
rect 78180 97562 78236 97618
rect 78304 97562 78360 97618
rect 78428 97562 78484 97618
rect 78552 97562 78608 97618
rect 77808 97438 77864 97494
rect 77932 97438 77988 97494
rect 78056 97438 78112 97494
rect 78180 97438 78236 97494
rect 78304 97438 78360 97494
rect 78428 97438 78484 97494
rect 78552 97438 78608 97494
rect 77808 97314 77864 97370
rect 77932 97314 77988 97370
rect 78056 97314 78112 97370
rect 78180 97314 78236 97370
rect 78304 97314 78360 97370
rect 78428 97314 78484 97370
rect 78552 97314 78608 97370
rect 77808 97190 77864 97246
rect 77932 97190 77988 97246
rect 78056 97190 78112 97246
rect 78180 97190 78236 97246
rect 78304 97190 78360 97246
rect 78428 97190 78484 97246
rect 78552 97190 78608 97246
rect 77808 97066 77864 97122
rect 77932 97066 77988 97122
rect 78056 97066 78112 97122
rect 78180 97066 78236 97122
rect 78304 97066 78360 97122
rect 78428 97066 78484 97122
rect 78552 97066 78608 97122
rect 77808 96942 77864 96998
rect 77932 96942 77988 96998
rect 78056 96942 78112 96998
rect 78180 96942 78236 96998
rect 78304 96942 78360 96998
rect 78428 96942 78484 96998
rect 78552 96942 78608 96998
rect 77808 96818 77864 96874
rect 77932 96818 77988 96874
rect 78056 96818 78112 96874
rect 78180 96818 78236 96874
rect 78304 96818 78360 96874
rect 78428 96818 78484 96874
rect 78552 96818 78608 96874
rect 77808 96694 77864 96750
rect 77932 96694 77988 96750
rect 78056 96694 78112 96750
rect 78180 96694 78236 96750
rect 78304 96694 78360 96750
rect 78428 96694 78484 96750
rect 78552 96694 78608 96750
rect 77808 96570 77864 96626
rect 77932 96570 77988 96626
rect 78056 96570 78112 96626
rect 78180 96570 78236 96626
rect 78304 96570 78360 96626
rect 78428 96570 78484 96626
rect 78552 96570 78608 96626
rect 77808 96446 77864 96502
rect 77932 96446 77988 96502
rect 78056 96446 78112 96502
rect 78180 96446 78236 96502
rect 78304 96446 78360 96502
rect 78428 96446 78484 96502
rect 78552 96446 78608 96502
rect 77808 96322 77864 96378
rect 77932 96322 77988 96378
rect 78056 96322 78112 96378
rect 78180 96322 78236 96378
rect 78304 96322 78360 96378
rect 78428 96322 78484 96378
rect 78552 96322 78608 96378
rect 77808 96198 77864 96254
rect 77932 96198 77988 96254
rect 78056 96198 78112 96254
rect 78180 96198 78236 96254
rect 78304 96198 78360 96254
rect 78428 96198 78484 96254
rect 78552 96198 78608 96254
rect 70074 95682 70130 95738
rect 70074 95558 70130 95614
rect 70074 95434 70130 95490
rect 70074 95310 70130 95366
rect 70074 95186 70130 95242
rect 70074 95062 70130 95118
rect 70074 94938 70130 94994
rect 70074 94814 70130 94870
rect 70074 94690 70130 94746
rect 70074 94566 70130 94622
rect 70074 94442 70130 94498
rect 70074 94318 70130 94374
rect 70074 94194 70130 94250
rect 70074 94070 70130 94126
rect 70074 93946 70130 94002
rect 70074 93822 70130 93878
rect 77808 95688 77864 95744
rect 77932 95688 77988 95744
rect 78056 95688 78112 95744
rect 78180 95688 78236 95744
rect 78304 95688 78360 95744
rect 78428 95688 78484 95744
rect 78552 95688 78608 95744
rect 77808 95564 77864 95620
rect 77932 95564 77988 95620
rect 78056 95564 78112 95620
rect 78180 95564 78236 95620
rect 78304 95564 78360 95620
rect 78428 95564 78484 95620
rect 78552 95564 78608 95620
rect 77808 95440 77864 95496
rect 77932 95440 77988 95496
rect 78056 95440 78112 95496
rect 78180 95440 78236 95496
rect 78304 95440 78360 95496
rect 78428 95440 78484 95496
rect 78552 95440 78608 95496
rect 77808 95316 77864 95372
rect 77932 95316 77988 95372
rect 78056 95316 78112 95372
rect 78180 95316 78236 95372
rect 78304 95316 78360 95372
rect 78428 95316 78484 95372
rect 78552 95316 78608 95372
rect 77808 95192 77864 95248
rect 77932 95192 77988 95248
rect 78056 95192 78112 95248
rect 78180 95192 78236 95248
rect 78304 95192 78360 95248
rect 78428 95192 78484 95248
rect 78552 95192 78608 95248
rect 77808 95068 77864 95124
rect 77932 95068 77988 95124
rect 78056 95068 78112 95124
rect 78180 95068 78236 95124
rect 78304 95068 78360 95124
rect 78428 95068 78484 95124
rect 78552 95068 78608 95124
rect 77808 94944 77864 95000
rect 77932 94944 77988 95000
rect 78056 94944 78112 95000
rect 78180 94944 78236 95000
rect 78304 94944 78360 95000
rect 78428 94944 78484 95000
rect 78552 94944 78608 95000
rect 77808 94820 77864 94876
rect 77932 94820 77988 94876
rect 78056 94820 78112 94876
rect 78180 94820 78236 94876
rect 78304 94820 78360 94876
rect 78428 94820 78484 94876
rect 78552 94820 78608 94876
rect 77808 94696 77864 94752
rect 77932 94696 77988 94752
rect 78056 94696 78112 94752
rect 78180 94696 78236 94752
rect 78304 94696 78360 94752
rect 78428 94696 78484 94752
rect 78552 94696 78608 94752
rect 77808 94572 77864 94628
rect 77932 94572 77988 94628
rect 78056 94572 78112 94628
rect 78180 94572 78236 94628
rect 78304 94572 78360 94628
rect 78428 94572 78484 94628
rect 78552 94572 78608 94628
rect 77808 94448 77864 94504
rect 77932 94448 77988 94504
rect 78056 94448 78112 94504
rect 78180 94448 78236 94504
rect 78304 94448 78360 94504
rect 78428 94448 78484 94504
rect 78552 94448 78608 94504
rect 77808 94324 77864 94380
rect 77932 94324 77988 94380
rect 78056 94324 78112 94380
rect 78180 94324 78236 94380
rect 78304 94324 78360 94380
rect 78428 94324 78484 94380
rect 78552 94324 78608 94380
rect 77808 94200 77864 94256
rect 77932 94200 77988 94256
rect 78056 94200 78112 94256
rect 78180 94200 78236 94256
rect 78304 94200 78360 94256
rect 78428 94200 78484 94256
rect 78552 94200 78608 94256
rect 77808 94076 77864 94132
rect 77932 94076 77988 94132
rect 78056 94076 78112 94132
rect 78180 94076 78236 94132
rect 78304 94076 78360 94132
rect 78428 94076 78484 94132
rect 78552 94076 78608 94132
rect 77808 93952 77864 94008
rect 77932 93952 77988 94008
rect 78056 93952 78112 94008
rect 78180 93952 78236 94008
rect 78304 93952 78360 94008
rect 78428 93952 78484 94008
rect 78552 93952 78608 94008
rect 77808 93828 77864 93884
rect 77932 93828 77988 93884
rect 78056 93828 78112 93884
rect 78180 93828 78236 93884
rect 78304 93828 78360 93884
rect 78428 93828 78484 93884
rect 78552 93828 78608 93884
rect 70074 93078 70130 93134
rect 70074 92954 70130 93010
rect 70074 92830 70130 92886
rect 70074 92706 70130 92762
rect 70074 92582 70130 92638
rect 70074 92458 70130 92514
rect 70074 92334 70130 92390
rect 70074 92210 70130 92266
rect 70074 92086 70130 92142
rect 70074 91962 70130 92018
rect 70074 91838 70130 91894
rect 70074 91714 70130 91770
rect 70074 91590 70130 91646
rect 70074 91466 70130 91522
rect 70074 91342 70130 91398
rect 77808 93084 77864 93140
rect 77932 93084 77988 93140
rect 78056 93084 78112 93140
rect 78180 93084 78236 93140
rect 78304 93084 78360 93140
rect 78428 93084 78484 93140
rect 78552 93084 78608 93140
rect 77808 92960 77864 93016
rect 77932 92960 77988 93016
rect 78056 92960 78112 93016
rect 78180 92960 78236 93016
rect 78304 92960 78360 93016
rect 78428 92960 78484 93016
rect 78552 92960 78608 93016
rect 77808 92836 77864 92892
rect 77932 92836 77988 92892
rect 78056 92836 78112 92892
rect 78180 92836 78236 92892
rect 78304 92836 78360 92892
rect 78428 92836 78484 92892
rect 78552 92836 78608 92892
rect 77808 92712 77864 92768
rect 77932 92712 77988 92768
rect 78056 92712 78112 92768
rect 78180 92712 78236 92768
rect 78304 92712 78360 92768
rect 78428 92712 78484 92768
rect 78552 92712 78608 92768
rect 77808 92588 77864 92644
rect 77932 92588 77988 92644
rect 78056 92588 78112 92644
rect 78180 92588 78236 92644
rect 78304 92588 78360 92644
rect 78428 92588 78484 92644
rect 78552 92588 78608 92644
rect 77808 92464 77864 92520
rect 77932 92464 77988 92520
rect 78056 92464 78112 92520
rect 78180 92464 78236 92520
rect 78304 92464 78360 92520
rect 78428 92464 78484 92520
rect 78552 92464 78608 92520
rect 77808 92340 77864 92396
rect 77932 92340 77988 92396
rect 78056 92340 78112 92396
rect 78180 92340 78236 92396
rect 78304 92340 78360 92396
rect 78428 92340 78484 92396
rect 78552 92340 78608 92396
rect 77808 92216 77864 92272
rect 77932 92216 77988 92272
rect 78056 92216 78112 92272
rect 78180 92216 78236 92272
rect 78304 92216 78360 92272
rect 78428 92216 78484 92272
rect 78552 92216 78608 92272
rect 77808 92092 77864 92148
rect 77932 92092 77988 92148
rect 78056 92092 78112 92148
rect 78180 92092 78236 92148
rect 78304 92092 78360 92148
rect 78428 92092 78484 92148
rect 78552 92092 78608 92148
rect 77808 91968 77864 92024
rect 77932 91968 77988 92024
rect 78056 91968 78112 92024
rect 78180 91968 78236 92024
rect 78304 91968 78360 92024
rect 78428 91968 78484 92024
rect 78552 91968 78608 92024
rect 77808 91844 77864 91900
rect 77932 91844 77988 91900
rect 78056 91844 78112 91900
rect 78180 91844 78236 91900
rect 78304 91844 78360 91900
rect 78428 91844 78484 91900
rect 78552 91844 78608 91900
rect 77808 91720 77864 91776
rect 77932 91720 77988 91776
rect 78056 91720 78112 91776
rect 78180 91720 78236 91776
rect 78304 91720 78360 91776
rect 78428 91720 78484 91776
rect 78552 91720 78608 91776
rect 77808 91596 77864 91652
rect 77932 91596 77988 91652
rect 78056 91596 78112 91652
rect 78180 91596 78236 91652
rect 78304 91596 78360 91652
rect 78428 91596 78484 91652
rect 78552 91596 78608 91652
rect 77808 91472 77864 91528
rect 77932 91472 77988 91528
rect 78056 91472 78112 91528
rect 78180 91472 78236 91528
rect 78304 91472 78360 91528
rect 78428 91472 78484 91528
rect 78552 91472 78608 91528
rect 77808 91348 77864 91404
rect 77932 91348 77988 91404
rect 78056 91348 78112 91404
rect 78180 91348 78236 91404
rect 78304 91348 78360 91404
rect 78428 91348 78484 91404
rect 78552 91348 78608 91404
rect 77748 86316 77804 86372
rect 77872 86316 77928 86372
rect 77996 86316 78052 86372
rect 78120 86316 78176 86372
rect 78244 86316 78300 86372
rect 78368 86316 78424 86372
rect 78492 86316 78548 86372
rect 77748 86192 77804 86248
rect 77872 86192 77928 86248
rect 77996 86192 78052 86248
rect 78120 86192 78176 86248
rect 78244 86192 78300 86248
rect 78368 86192 78424 86248
rect 78492 86192 78548 86248
rect 110548 943379 110604 943435
rect 79148 940796 79204 940852
rect 79272 940796 79328 940852
rect 79396 940796 79452 940852
rect 79520 940796 79576 940852
rect 79644 940796 79700 940852
rect 79768 940796 79824 940852
rect 79892 940796 79948 940852
rect 79148 940672 79204 940728
rect 79272 940672 79328 940728
rect 79396 940672 79452 940728
rect 79520 940672 79576 940728
rect 79644 940672 79700 940728
rect 79768 940672 79824 940728
rect 79892 940672 79948 940728
rect 79148 940548 79204 940604
rect 79272 940548 79328 940604
rect 79396 940548 79452 940604
rect 79520 940548 79576 940604
rect 79644 940548 79700 940604
rect 79768 940548 79824 940604
rect 79892 940548 79948 940604
rect 79148 940424 79204 940480
rect 79272 940424 79328 940480
rect 79396 940424 79452 940480
rect 79520 940424 79576 940480
rect 79644 940424 79700 940480
rect 79768 940424 79824 940480
rect 79892 940424 79948 940480
rect 79148 940300 79204 940356
rect 79272 940300 79328 940356
rect 79396 940300 79452 940356
rect 79520 940300 79576 940356
rect 79644 940300 79700 940356
rect 79768 940300 79824 940356
rect 79892 940300 79948 940356
rect 79148 940176 79204 940232
rect 79272 940176 79328 940232
rect 79396 940176 79452 940232
rect 79520 940176 79576 940232
rect 79644 940176 79700 940232
rect 79768 940176 79824 940232
rect 79892 940176 79948 940232
rect 79148 940052 79204 940108
rect 79272 940052 79328 940108
rect 79396 940052 79452 940108
rect 79520 940052 79576 940108
rect 79644 940052 79700 940108
rect 79768 940052 79824 940108
rect 79892 940052 79948 940108
rect 88207 942144 88263 942200
rect 88407 942144 88463 942200
rect 88207 941844 88263 941900
rect 88407 941844 88463 941900
rect 88207 941544 88263 941600
rect 88407 941544 88463 941600
rect 106207 940744 106263 940800
rect 106407 940744 106463 940800
rect 106207 940444 106263 940500
rect 106407 940444 106463 940500
rect 106207 940144 106263 940200
rect 106407 940144 106463 940200
rect 110546 940654 110602 940710
rect 110546 940354 110602 940410
rect 110546 940054 110602 940110
rect 117548 943379 117604 943435
rect 117546 940654 117602 940710
rect 117546 940354 117602 940410
rect 117546 940054 117602 940110
rect 124548 943379 124604 943435
rect 140406 942097 140462 942153
rect 140406 941797 140462 941853
rect 140406 941497 140462 941553
rect 124546 940654 124602 940710
rect 124546 940354 124602 940410
rect 124546 940054 124602 940110
rect 165548 943379 165604 943435
rect 160207 942144 160263 942200
rect 160407 942144 160463 942200
rect 160207 941844 160263 941900
rect 160407 941844 160463 941900
rect 160207 941544 160263 941600
rect 160407 941544 160463 941600
rect 140821 940660 140877 940716
rect 140821 940360 140877 940416
rect 140821 940060 140877 940116
rect 142207 940744 142263 940800
rect 142407 940744 142463 940800
rect 142207 940444 142263 940500
rect 142407 940444 142463 940500
rect 142207 940144 142263 940200
rect 142407 940144 142463 940200
rect 165546 940654 165602 940710
rect 165546 940354 165602 940410
rect 165546 940054 165602 940110
rect 172548 943379 172604 943435
rect 179548 943379 179604 943435
rect 172546 940654 172602 940710
rect 172546 940354 172602 940410
rect 172546 940054 172602 940110
rect 178207 940744 178263 940800
rect 178407 940744 178463 940800
rect 178207 940444 178263 940500
rect 178407 940444 178463 940500
rect 178207 940144 178263 940200
rect 178407 940144 178463 940200
rect 195406 942097 195462 942153
rect 195406 941797 195462 941853
rect 195406 941497 195462 941553
rect 179546 940654 179602 940710
rect 179546 940354 179602 940410
rect 179546 940054 179602 940110
rect 220548 943379 220604 943435
rect 195821 940660 195877 940716
rect 195821 940360 195877 940416
rect 195821 940060 195877 940116
rect 214207 940744 214263 940800
rect 214407 940744 214463 940800
rect 214207 940444 214263 940500
rect 214407 940444 214463 940500
rect 214207 940144 214263 940200
rect 214407 940144 214463 940200
rect 220546 940654 220602 940710
rect 220546 940354 220602 940410
rect 220546 940054 220602 940110
rect 227548 943379 227604 943435
rect 234548 943379 234604 943435
rect 227546 940654 227602 940710
rect 227546 940354 227602 940410
rect 227546 940054 227602 940110
rect 232207 942144 232263 942200
rect 232407 942144 232463 942200
rect 232207 941844 232263 941900
rect 232407 941844 232463 941900
rect 232207 941544 232263 941600
rect 232407 941544 232463 941600
rect 250406 942097 250462 942153
rect 250406 941797 250462 941853
rect 250406 941497 250462 941553
rect 234546 940654 234602 940710
rect 234546 940354 234602 940410
rect 234546 940054 234602 940110
rect 250207 940744 250263 940800
rect 250407 940744 250463 940800
rect 250207 940444 250263 940500
rect 250407 940444 250463 940500
rect 250207 940144 250263 940200
rect 250407 940144 250463 940200
rect 275548 943379 275604 943435
rect 250821 940660 250877 940716
rect 250821 940360 250877 940416
rect 250821 940060 250877 940116
rect 268207 942144 268263 942200
rect 268407 942144 268463 942200
rect 268207 941844 268263 941900
rect 268407 941844 268463 941900
rect 268207 941544 268263 941600
rect 268407 941544 268463 941600
rect 275546 940654 275602 940710
rect 275546 940354 275602 940410
rect 275546 940054 275602 940110
rect 282548 943379 282604 943435
rect 289548 943379 289604 943435
rect 282546 940654 282602 940710
rect 282546 940354 282602 940410
rect 282546 940054 282602 940110
rect 286207 940744 286263 940800
rect 286407 940744 286463 940800
rect 286207 940444 286263 940500
rect 286407 940444 286463 940500
rect 286207 940144 286263 940200
rect 286407 940144 286463 940200
rect 289546 940654 289602 940710
rect 289546 940354 289602 940410
rect 289546 940054 289602 940110
rect 304207 942144 304263 942200
rect 304407 942144 304463 942200
rect 304207 941844 304263 941900
rect 304407 941844 304463 941900
rect 304207 941544 304263 941600
rect 304407 941544 304463 941600
rect 305406 942097 305462 942153
rect 305406 941797 305462 941853
rect 305406 941497 305462 941553
rect 330548 943379 330604 943435
rect 305821 940660 305877 940716
rect 305821 940360 305877 940416
rect 305821 940060 305877 940116
rect 322207 940744 322263 940800
rect 322407 940744 322463 940800
rect 322207 940444 322263 940500
rect 322407 940444 322463 940500
rect 322207 940144 322263 940200
rect 322407 940144 322463 940200
rect 330546 940654 330602 940710
rect 330546 940354 330602 940410
rect 330546 940054 330602 940110
rect 337548 943379 337604 943435
rect 344548 943379 344604 943435
rect 337546 940654 337602 940710
rect 337546 940354 337602 940410
rect 337546 940054 337602 940110
rect 340207 942144 340263 942200
rect 340407 942144 340463 942200
rect 340207 941844 340263 941900
rect 340407 941844 340463 941900
rect 340207 941544 340263 941600
rect 340407 941544 340463 941600
rect 360406 942097 360462 942153
rect 360406 941797 360462 941853
rect 360406 941497 360462 941553
rect 344546 940654 344602 940710
rect 344546 940354 344602 940410
rect 344546 940054 344602 940110
rect 358207 940744 358263 940800
rect 358407 940744 358463 940800
rect 358207 940444 358263 940500
rect 358407 940444 358463 940500
rect 358207 940144 358263 940200
rect 358407 940144 358463 940200
rect 360821 940660 360877 940716
rect 360821 940360 360877 940416
rect 360821 940060 360877 940116
rect 376207 942144 376263 942200
rect 376407 942144 376463 942200
rect 376207 941844 376263 941900
rect 376407 941844 376463 941900
rect 376207 941544 376263 941600
rect 376407 941544 376463 941600
rect 381348 940736 381404 940792
rect 381472 940736 381528 940792
rect 381596 940736 381652 940792
rect 381720 940736 381776 940792
rect 381844 940736 381900 940792
rect 381968 940736 382024 940792
rect 382092 940736 382148 940792
rect 382216 940736 382272 940792
rect 382340 940736 382396 940792
rect 382464 940736 382520 940792
rect 382588 940736 382644 940792
rect 382712 940736 382768 940792
rect 382836 940736 382892 940792
rect 382960 940736 383016 940792
rect 383084 940736 383140 940792
rect 381348 940612 381404 940668
rect 381472 940612 381528 940668
rect 381596 940612 381652 940668
rect 381720 940612 381776 940668
rect 381844 940612 381900 940668
rect 381968 940612 382024 940668
rect 382092 940612 382148 940668
rect 382216 940612 382272 940668
rect 382340 940612 382396 940668
rect 382464 940612 382520 940668
rect 382588 940612 382644 940668
rect 382712 940612 382768 940668
rect 382836 940612 382892 940668
rect 382960 940612 383016 940668
rect 383084 940612 383140 940668
rect 381348 940488 381404 940544
rect 381472 940488 381528 940544
rect 381596 940488 381652 940544
rect 381720 940488 381776 940544
rect 381844 940488 381900 940544
rect 381968 940488 382024 940544
rect 382092 940488 382148 940544
rect 382216 940488 382272 940544
rect 382340 940488 382396 940544
rect 382464 940488 382520 940544
rect 382588 940488 382644 940544
rect 382712 940488 382768 940544
rect 382836 940488 382892 940544
rect 382960 940488 383016 940544
rect 383084 940488 383140 940544
rect 381348 940364 381404 940420
rect 381472 940364 381528 940420
rect 381596 940364 381652 940420
rect 381720 940364 381776 940420
rect 381844 940364 381900 940420
rect 381968 940364 382024 940420
rect 382092 940364 382148 940420
rect 382216 940364 382272 940420
rect 382340 940364 382396 940420
rect 382464 940364 382520 940420
rect 382588 940364 382644 940420
rect 382712 940364 382768 940420
rect 382836 940364 382892 940420
rect 382960 940364 383016 940420
rect 383084 940364 383140 940420
rect 381348 940240 381404 940296
rect 381472 940240 381528 940296
rect 381596 940240 381652 940296
rect 381720 940240 381776 940296
rect 381844 940240 381900 940296
rect 381968 940240 382024 940296
rect 382092 940240 382148 940296
rect 382216 940240 382272 940296
rect 382340 940240 382396 940296
rect 382464 940240 382520 940296
rect 382588 940240 382644 940296
rect 382712 940240 382768 940296
rect 382836 940240 382892 940296
rect 382960 940240 383016 940296
rect 383084 940240 383140 940296
rect 381348 940116 381404 940172
rect 381472 940116 381528 940172
rect 381596 940116 381652 940172
rect 381720 940116 381776 940172
rect 381844 940116 381900 940172
rect 381968 940116 382024 940172
rect 382092 940116 382148 940172
rect 382216 940116 382272 940172
rect 382340 940116 382396 940172
rect 382464 940116 382520 940172
rect 382588 940116 382644 940172
rect 382712 940116 382768 940172
rect 382836 940116 382892 940172
rect 382960 940116 383016 940172
rect 383084 940116 383140 940172
rect 381348 939992 381404 940048
rect 381472 939992 381528 940048
rect 381596 939992 381652 940048
rect 381720 939992 381776 940048
rect 381844 939992 381900 940048
rect 381968 939992 382024 940048
rect 382092 939992 382148 940048
rect 382216 939992 382272 940048
rect 382340 939992 382396 940048
rect 382464 939992 382520 940048
rect 382588 939992 382644 940048
rect 382712 939992 382768 940048
rect 382836 939992 382892 940048
rect 382960 939992 383016 940048
rect 383084 939992 383140 940048
rect 383828 940736 383884 940792
rect 383952 940736 384008 940792
rect 384076 940736 384132 940792
rect 384200 940736 384256 940792
rect 384324 940736 384380 940792
rect 384448 940736 384504 940792
rect 384572 940736 384628 940792
rect 384696 940736 384752 940792
rect 384820 940736 384876 940792
rect 384944 940736 385000 940792
rect 385068 940736 385124 940792
rect 385192 940736 385248 940792
rect 385316 940736 385372 940792
rect 385440 940736 385496 940792
rect 385564 940736 385620 940792
rect 385688 940736 385744 940792
rect 383828 940612 383884 940668
rect 383952 940612 384008 940668
rect 384076 940612 384132 940668
rect 384200 940612 384256 940668
rect 384324 940612 384380 940668
rect 384448 940612 384504 940668
rect 384572 940612 384628 940668
rect 384696 940612 384752 940668
rect 384820 940612 384876 940668
rect 384944 940612 385000 940668
rect 385068 940612 385124 940668
rect 385192 940612 385248 940668
rect 385316 940612 385372 940668
rect 385440 940612 385496 940668
rect 385564 940612 385620 940668
rect 385688 940612 385744 940668
rect 383828 940488 383884 940544
rect 383952 940488 384008 940544
rect 384076 940488 384132 940544
rect 384200 940488 384256 940544
rect 384324 940488 384380 940544
rect 384448 940488 384504 940544
rect 384572 940488 384628 940544
rect 384696 940488 384752 940544
rect 384820 940488 384876 940544
rect 384944 940488 385000 940544
rect 385068 940488 385124 940544
rect 385192 940488 385248 940544
rect 385316 940488 385372 940544
rect 385440 940488 385496 940544
rect 385564 940488 385620 940544
rect 385688 940488 385744 940544
rect 383828 940364 383884 940420
rect 383952 940364 384008 940420
rect 384076 940364 384132 940420
rect 384200 940364 384256 940420
rect 384324 940364 384380 940420
rect 384448 940364 384504 940420
rect 384572 940364 384628 940420
rect 384696 940364 384752 940420
rect 384820 940364 384876 940420
rect 384944 940364 385000 940420
rect 385068 940364 385124 940420
rect 385192 940364 385248 940420
rect 385316 940364 385372 940420
rect 385440 940364 385496 940420
rect 385564 940364 385620 940420
rect 385688 940364 385744 940420
rect 383828 940240 383884 940296
rect 383952 940240 384008 940296
rect 384076 940240 384132 940296
rect 384200 940240 384256 940296
rect 384324 940240 384380 940296
rect 384448 940240 384504 940296
rect 384572 940240 384628 940296
rect 384696 940240 384752 940296
rect 384820 940240 384876 940296
rect 384944 940240 385000 940296
rect 385068 940240 385124 940296
rect 385192 940240 385248 940296
rect 385316 940240 385372 940296
rect 385440 940240 385496 940296
rect 385564 940240 385620 940296
rect 385688 940240 385744 940296
rect 383828 940116 383884 940172
rect 383952 940116 384008 940172
rect 384076 940116 384132 940172
rect 384200 940116 384256 940172
rect 384324 940116 384380 940172
rect 384448 940116 384504 940172
rect 384572 940116 384628 940172
rect 384696 940116 384752 940172
rect 384820 940116 384876 940172
rect 384944 940116 385000 940172
rect 385068 940116 385124 940172
rect 385192 940116 385248 940172
rect 385316 940116 385372 940172
rect 385440 940116 385496 940172
rect 385564 940116 385620 940172
rect 385688 940116 385744 940172
rect 383828 939992 383884 940048
rect 383952 939992 384008 940048
rect 384076 939992 384132 940048
rect 384200 939992 384256 940048
rect 384324 939992 384380 940048
rect 384448 939992 384504 940048
rect 384572 939992 384628 940048
rect 384696 939992 384752 940048
rect 384820 939992 384876 940048
rect 384944 939992 385000 940048
rect 385068 939992 385124 940048
rect 385192 939992 385248 940048
rect 385316 939992 385372 940048
rect 385440 939992 385496 940048
rect 385564 939992 385620 940048
rect 385688 939992 385744 940048
rect 386198 940736 386254 940792
rect 386322 940736 386378 940792
rect 386446 940736 386502 940792
rect 386570 940736 386626 940792
rect 386694 940736 386750 940792
rect 386818 940736 386874 940792
rect 386942 940736 386998 940792
rect 387066 940736 387122 940792
rect 387190 940736 387246 940792
rect 387314 940736 387370 940792
rect 387438 940736 387494 940792
rect 387562 940736 387618 940792
rect 387686 940736 387742 940792
rect 387810 940736 387866 940792
rect 387934 940736 387990 940792
rect 388058 940736 388114 940792
rect 386198 940612 386254 940668
rect 386322 940612 386378 940668
rect 386446 940612 386502 940668
rect 386570 940612 386626 940668
rect 386694 940612 386750 940668
rect 386818 940612 386874 940668
rect 386942 940612 386998 940668
rect 387066 940612 387122 940668
rect 387190 940612 387246 940668
rect 387314 940612 387370 940668
rect 387438 940612 387494 940668
rect 387562 940612 387618 940668
rect 387686 940612 387742 940668
rect 387810 940612 387866 940668
rect 387934 940612 387990 940668
rect 388058 940612 388114 940668
rect 386198 940488 386254 940544
rect 386322 940488 386378 940544
rect 386446 940488 386502 940544
rect 386570 940488 386626 940544
rect 386694 940488 386750 940544
rect 386818 940488 386874 940544
rect 386942 940488 386998 940544
rect 387066 940488 387122 940544
rect 387190 940488 387246 940544
rect 387314 940488 387370 940544
rect 387438 940488 387494 940544
rect 387562 940488 387618 940544
rect 387686 940488 387742 940544
rect 387810 940488 387866 940544
rect 387934 940488 387990 940544
rect 388058 940488 388114 940544
rect 386198 940364 386254 940420
rect 386322 940364 386378 940420
rect 386446 940364 386502 940420
rect 386570 940364 386626 940420
rect 386694 940364 386750 940420
rect 386818 940364 386874 940420
rect 386942 940364 386998 940420
rect 387066 940364 387122 940420
rect 387190 940364 387246 940420
rect 387314 940364 387370 940420
rect 387438 940364 387494 940420
rect 387562 940364 387618 940420
rect 387686 940364 387742 940420
rect 387810 940364 387866 940420
rect 387934 940364 387990 940420
rect 388058 940364 388114 940420
rect 386198 940240 386254 940296
rect 386322 940240 386378 940296
rect 386446 940240 386502 940296
rect 386570 940240 386626 940296
rect 386694 940240 386750 940296
rect 386818 940240 386874 940296
rect 386942 940240 386998 940296
rect 387066 940240 387122 940296
rect 387190 940240 387246 940296
rect 387314 940240 387370 940296
rect 387438 940240 387494 940296
rect 387562 940240 387618 940296
rect 387686 940240 387742 940296
rect 387810 940240 387866 940296
rect 387934 940240 387990 940296
rect 388058 940240 388114 940296
rect 386198 940116 386254 940172
rect 386322 940116 386378 940172
rect 386446 940116 386502 940172
rect 386570 940116 386626 940172
rect 386694 940116 386750 940172
rect 386818 940116 386874 940172
rect 386942 940116 386998 940172
rect 387066 940116 387122 940172
rect 387190 940116 387246 940172
rect 387314 940116 387370 940172
rect 387438 940116 387494 940172
rect 387562 940116 387618 940172
rect 387686 940116 387742 940172
rect 387810 940116 387866 940172
rect 387934 940116 387990 940172
rect 388058 940116 388114 940172
rect 386198 939992 386254 940048
rect 386322 939992 386378 940048
rect 386446 939992 386502 940048
rect 386570 939992 386626 940048
rect 386694 939992 386750 940048
rect 386818 939992 386874 940048
rect 386942 939992 386998 940048
rect 387066 939992 387122 940048
rect 387190 939992 387246 940048
rect 387314 939992 387370 940048
rect 387438 939992 387494 940048
rect 387562 939992 387618 940048
rect 387686 939992 387742 940048
rect 387810 939992 387866 940048
rect 387934 939992 387990 940048
rect 388058 939992 388114 940048
rect 388904 940736 388960 940792
rect 389028 940736 389084 940792
rect 389152 940736 389208 940792
rect 389276 940736 389332 940792
rect 389400 940736 389456 940792
rect 389524 940736 389580 940792
rect 389648 940736 389704 940792
rect 389772 940736 389828 940792
rect 389896 940736 389952 940792
rect 390020 940736 390076 940792
rect 390144 940736 390200 940792
rect 390268 940736 390324 940792
rect 390392 940736 390448 940792
rect 390516 940736 390572 940792
rect 390640 940736 390696 940792
rect 390764 940736 390820 940792
rect 388904 940612 388960 940668
rect 389028 940612 389084 940668
rect 389152 940612 389208 940668
rect 389276 940612 389332 940668
rect 389400 940612 389456 940668
rect 389524 940612 389580 940668
rect 389648 940612 389704 940668
rect 389772 940612 389828 940668
rect 389896 940612 389952 940668
rect 390020 940612 390076 940668
rect 390144 940612 390200 940668
rect 390268 940612 390324 940668
rect 390392 940612 390448 940668
rect 390516 940612 390572 940668
rect 390640 940612 390696 940668
rect 390764 940612 390820 940668
rect 388904 940488 388960 940544
rect 389028 940488 389084 940544
rect 389152 940488 389208 940544
rect 389276 940488 389332 940544
rect 389400 940488 389456 940544
rect 389524 940488 389580 940544
rect 389648 940488 389704 940544
rect 389772 940488 389828 940544
rect 389896 940488 389952 940544
rect 390020 940488 390076 940544
rect 390144 940488 390200 940544
rect 390268 940488 390324 940544
rect 390392 940488 390448 940544
rect 390516 940488 390572 940544
rect 390640 940488 390696 940544
rect 390764 940488 390820 940544
rect 388904 940364 388960 940420
rect 389028 940364 389084 940420
rect 389152 940364 389208 940420
rect 389276 940364 389332 940420
rect 389400 940364 389456 940420
rect 389524 940364 389580 940420
rect 389648 940364 389704 940420
rect 389772 940364 389828 940420
rect 389896 940364 389952 940420
rect 390020 940364 390076 940420
rect 390144 940364 390200 940420
rect 390268 940364 390324 940420
rect 390392 940364 390448 940420
rect 390516 940364 390572 940420
rect 390640 940364 390696 940420
rect 390764 940364 390820 940420
rect 388904 940240 388960 940296
rect 389028 940240 389084 940296
rect 389152 940240 389208 940296
rect 389276 940240 389332 940296
rect 389400 940240 389456 940296
rect 389524 940240 389580 940296
rect 389648 940240 389704 940296
rect 389772 940240 389828 940296
rect 389896 940240 389952 940296
rect 390020 940240 390076 940296
rect 390144 940240 390200 940296
rect 390268 940240 390324 940296
rect 390392 940240 390448 940296
rect 390516 940240 390572 940296
rect 390640 940240 390696 940296
rect 390764 940240 390820 940296
rect 388904 940116 388960 940172
rect 389028 940116 389084 940172
rect 389152 940116 389208 940172
rect 389276 940116 389332 940172
rect 389400 940116 389456 940172
rect 389524 940116 389580 940172
rect 389648 940116 389704 940172
rect 389772 940116 389828 940172
rect 389896 940116 389952 940172
rect 390020 940116 390076 940172
rect 390144 940116 390200 940172
rect 390268 940116 390324 940172
rect 390392 940116 390448 940172
rect 390516 940116 390572 940172
rect 390640 940116 390696 940172
rect 390764 940116 390820 940172
rect 388904 939992 388960 940048
rect 389028 939992 389084 940048
rect 389152 939992 389208 940048
rect 389276 939992 389332 940048
rect 389400 939992 389456 940048
rect 389524 939992 389580 940048
rect 389648 939992 389704 940048
rect 389772 939992 389828 940048
rect 389896 939992 389952 940048
rect 390020 939992 390076 940048
rect 390144 939992 390200 940048
rect 390268 939992 390324 940048
rect 390392 939992 390448 940048
rect 390516 939992 390572 940048
rect 390640 939992 390696 940048
rect 390764 939992 390820 940048
rect 391274 940736 391330 940792
rect 391398 940736 391454 940792
rect 391522 940736 391578 940792
rect 391646 940736 391702 940792
rect 391770 940736 391826 940792
rect 391894 940736 391950 940792
rect 392018 940736 392074 940792
rect 392142 940736 392198 940792
rect 392266 940736 392322 940792
rect 392390 940736 392446 940792
rect 392514 940736 392570 940792
rect 392638 940736 392694 940792
rect 392762 940736 392818 940792
rect 392886 940736 392942 940792
rect 393010 940736 393066 940792
rect 393134 940736 393190 940792
rect 391274 940612 391330 940668
rect 391398 940612 391454 940668
rect 391522 940612 391578 940668
rect 391646 940612 391702 940668
rect 391770 940612 391826 940668
rect 391894 940612 391950 940668
rect 392018 940612 392074 940668
rect 392142 940612 392198 940668
rect 392266 940612 392322 940668
rect 392390 940612 392446 940668
rect 392514 940612 392570 940668
rect 392638 940612 392694 940668
rect 392762 940612 392818 940668
rect 392886 940612 392942 940668
rect 393010 940612 393066 940668
rect 393134 940612 393190 940668
rect 391274 940488 391330 940544
rect 391398 940488 391454 940544
rect 391522 940488 391578 940544
rect 391646 940488 391702 940544
rect 391770 940488 391826 940544
rect 391894 940488 391950 940544
rect 392018 940488 392074 940544
rect 392142 940488 392198 940544
rect 392266 940488 392322 940544
rect 392390 940488 392446 940544
rect 392514 940488 392570 940544
rect 392638 940488 392694 940544
rect 392762 940488 392818 940544
rect 392886 940488 392942 940544
rect 393010 940488 393066 940544
rect 393134 940488 393190 940544
rect 391274 940364 391330 940420
rect 391398 940364 391454 940420
rect 391522 940364 391578 940420
rect 391646 940364 391702 940420
rect 391770 940364 391826 940420
rect 391894 940364 391950 940420
rect 392018 940364 392074 940420
rect 392142 940364 392198 940420
rect 392266 940364 392322 940420
rect 392390 940364 392446 940420
rect 392514 940364 392570 940420
rect 392638 940364 392694 940420
rect 392762 940364 392818 940420
rect 392886 940364 392942 940420
rect 393010 940364 393066 940420
rect 393134 940364 393190 940420
rect 391274 940240 391330 940296
rect 391398 940240 391454 940296
rect 391522 940240 391578 940296
rect 391646 940240 391702 940296
rect 391770 940240 391826 940296
rect 391894 940240 391950 940296
rect 392018 940240 392074 940296
rect 392142 940240 392198 940296
rect 392266 940240 392322 940296
rect 392390 940240 392446 940296
rect 392514 940240 392570 940296
rect 392638 940240 392694 940296
rect 392762 940240 392818 940296
rect 392886 940240 392942 940296
rect 393010 940240 393066 940296
rect 393134 940240 393190 940296
rect 391274 940116 391330 940172
rect 391398 940116 391454 940172
rect 391522 940116 391578 940172
rect 391646 940116 391702 940172
rect 391770 940116 391826 940172
rect 391894 940116 391950 940172
rect 392018 940116 392074 940172
rect 392142 940116 392198 940172
rect 392266 940116 392322 940172
rect 392390 940116 392446 940172
rect 392514 940116 392570 940172
rect 392638 940116 392694 940172
rect 392762 940116 392818 940172
rect 392886 940116 392942 940172
rect 393010 940116 393066 940172
rect 393134 940116 393190 940172
rect 391274 939992 391330 940048
rect 391398 939992 391454 940048
rect 391522 939992 391578 940048
rect 391646 939992 391702 940048
rect 391770 939992 391826 940048
rect 391894 939992 391950 940048
rect 392018 939992 392074 940048
rect 392142 939992 392198 940048
rect 392266 939992 392322 940048
rect 392390 939992 392446 940048
rect 392514 939992 392570 940048
rect 392638 939992 392694 940048
rect 392762 939992 392818 940048
rect 392886 939992 392942 940048
rect 393010 939992 393066 940048
rect 393134 939992 393190 940048
rect 440548 943379 440604 943435
rect 393878 940736 393934 940792
rect 394002 940736 394058 940792
rect 394126 940736 394182 940792
rect 394250 940736 394306 940792
rect 394374 940736 394430 940792
rect 394498 940736 394554 940792
rect 394622 940736 394678 940792
rect 394746 940736 394802 940792
rect 394870 940736 394926 940792
rect 394994 940736 395050 940792
rect 395118 940736 395174 940792
rect 395242 940736 395298 940792
rect 395366 940736 395422 940792
rect 395490 940736 395546 940792
rect 395614 940736 395670 940792
rect 393878 940612 393934 940668
rect 394002 940612 394058 940668
rect 394126 940612 394182 940668
rect 394250 940612 394306 940668
rect 394374 940612 394430 940668
rect 394498 940612 394554 940668
rect 394622 940612 394678 940668
rect 394746 940612 394802 940668
rect 394870 940612 394926 940668
rect 394994 940612 395050 940668
rect 395118 940612 395174 940668
rect 395242 940612 395298 940668
rect 395366 940612 395422 940668
rect 395490 940612 395546 940668
rect 395614 940612 395670 940668
rect 393878 940488 393934 940544
rect 394002 940488 394058 940544
rect 394126 940488 394182 940544
rect 394250 940488 394306 940544
rect 394374 940488 394430 940544
rect 394498 940488 394554 940544
rect 394622 940488 394678 940544
rect 394746 940488 394802 940544
rect 394870 940488 394926 940544
rect 394994 940488 395050 940544
rect 395118 940488 395174 940544
rect 395242 940488 395298 940544
rect 395366 940488 395422 940544
rect 395490 940488 395546 940544
rect 395614 940488 395670 940544
rect 393878 940364 393934 940420
rect 394002 940364 394058 940420
rect 394126 940364 394182 940420
rect 394250 940364 394306 940420
rect 394374 940364 394430 940420
rect 394498 940364 394554 940420
rect 394622 940364 394678 940420
rect 394746 940364 394802 940420
rect 394870 940364 394926 940420
rect 394994 940364 395050 940420
rect 395118 940364 395174 940420
rect 395242 940364 395298 940420
rect 395366 940364 395422 940420
rect 395490 940364 395546 940420
rect 395614 940364 395670 940420
rect 393878 940240 393934 940296
rect 394002 940240 394058 940296
rect 394126 940240 394182 940296
rect 394250 940240 394306 940296
rect 394374 940240 394430 940296
rect 394498 940240 394554 940296
rect 394622 940240 394678 940296
rect 394746 940240 394802 940296
rect 394870 940240 394926 940296
rect 394994 940240 395050 940296
rect 395118 940240 395174 940296
rect 395242 940240 395298 940296
rect 395366 940240 395422 940296
rect 395490 940240 395546 940296
rect 395614 940240 395670 940296
rect 393878 940116 393934 940172
rect 394002 940116 394058 940172
rect 394126 940116 394182 940172
rect 394250 940116 394306 940172
rect 394374 940116 394430 940172
rect 394498 940116 394554 940172
rect 394622 940116 394678 940172
rect 394746 940116 394802 940172
rect 394870 940116 394926 940172
rect 394994 940116 395050 940172
rect 395118 940116 395174 940172
rect 395242 940116 395298 940172
rect 395366 940116 395422 940172
rect 395490 940116 395546 940172
rect 395614 940116 395670 940172
rect 393878 939992 393934 940048
rect 394002 939992 394058 940048
rect 394126 939992 394182 940048
rect 394250 939992 394306 940048
rect 394374 939992 394430 940048
rect 394498 939992 394554 940048
rect 394622 939992 394678 940048
rect 394746 939992 394802 940048
rect 394870 939992 394926 940048
rect 394994 939992 395050 940048
rect 395118 939992 395174 940048
rect 395242 939992 395298 940048
rect 395366 939992 395422 940048
rect 395490 939992 395546 940048
rect 395614 939992 395670 940048
rect 412207 942144 412263 942200
rect 412407 942144 412463 942200
rect 412207 941844 412263 941900
rect 412407 941844 412463 941900
rect 412207 941544 412263 941600
rect 412407 941544 412463 941600
rect 430207 940744 430263 940800
rect 430407 940744 430463 940800
rect 430207 940444 430263 940500
rect 430407 940444 430463 940500
rect 430207 940144 430263 940200
rect 430407 940144 430463 940200
rect 440546 940654 440602 940710
rect 440546 940354 440602 940410
rect 440546 940054 440602 940110
rect 447548 943379 447604 943435
rect 454548 943379 454604 943435
rect 447546 940654 447602 940710
rect 447546 940354 447602 940410
rect 447546 940054 447602 940110
rect 448207 942144 448263 942200
rect 448407 942144 448463 942200
rect 448207 941844 448263 941900
rect 448407 941844 448463 941900
rect 448207 941544 448263 941600
rect 448407 941544 448463 941600
rect 470406 942097 470462 942153
rect 470406 941797 470462 941853
rect 470406 941497 470462 941553
rect 454546 940654 454602 940710
rect 454546 940354 454602 940410
rect 454546 940054 454602 940110
rect 466207 940744 466263 940800
rect 466407 940744 466463 940800
rect 466207 940444 466263 940500
rect 466407 940444 466463 940500
rect 466207 940144 466263 940200
rect 466407 940144 466463 940200
rect 495548 943379 495604 943435
rect 470821 940660 470877 940716
rect 470821 940360 470877 940416
rect 470821 940060 470877 940116
rect 484207 942144 484263 942200
rect 484407 942144 484463 942200
rect 484207 941844 484263 941900
rect 484407 941844 484463 941900
rect 484207 941544 484263 941600
rect 484407 941544 484463 941600
rect 502548 943379 502604 943435
rect 495546 940654 495602 940710
rect 495546 940354 495602 940410
rect 495546 940054 495602 940110
rect 502207 940744 502263 940800
rect 502407 940744 502463 940800
rect 502546 940654 502602 940710
rect 502207 940444 502263 940500
rect 502407 940444 502463 940500
rect 502546 940354 502602 940410
rect 502207 940144 502263 940200
rect 502407 940144 502463 940200
rect 502546 940054 502602 940110
rect 509548 943379 509604 943435
rect 509546 940654 509602 940710
rect 509546 940354 509602 940410
rect 509546 940054 509602 940110
rect 520207 942144 520263 942200
rect 520407 942144 520463 942200
rect 520207 941844 520263 941900
rect 520407 941844 520463 941900
rect 520207 941544 520263 941600
rect 520407 941544 520463 941600
rect 525406 942097 525462 942153
rect 525406 941797 525462 941853
rect 525406 941497 525462 941553
rect 550548 943379 550604 943435
rect 525821 940660 525877 940716
rect 525821 940360 525877 940416
rect 525821 940060 525877 940116
rect 538207 940744 538263 940800
rect 538407 940744 538463 940800
rect 538207 940444 538263 940500
rect 538407 940444 538463 940500
rect 538207 940144 538263 940200
rect 538407 940144 538463 940200
rect 557548 943379 557604 943435
rect 550546 940654 550602 940710
rect 550546 940354 550602 940410
rect 550546 940054 550602 940110
rect 556207 942144 556263 942200
rect 556407 942144 556463 942200
rect 556207 941844 556263 941900
rect 556407 941844 556463 941900
rect 556207 941544 556263 941600
rect 556407 941544 556463 941600
rect 557546 940654 557602 940710
rect 557546 940354 557602 940410
rect 557546 940054 557602 940110
rect 564548 943379 564604 943435
rect 580406 942097 580462 942153
rect 580406 941797 580462 941853
rect 580406 941497 580462 941553
rect 564546 940654 564602 940710
rect 564546 940354 564602 940410
rect 564546 940054 564602 940110
rect 574207 940744 574263 940800
rect 574407 940744 574463 940800
rect 574207 940444 574263 940500
rect 574407 940444 574463 940500
rect 574207 940144 574263 940200
rect 574407 940144 574463 940200
rect 580821 940660 580877 940716
rect 580821 940360 580877 940416
rect 580821 940060 580877 940116
rect 592207 942144 592263 942200
rect 592407 942144 592463 942200
rect 592207 941844 592263 941900
rect 592407 941844 592463 941900
rect 592207 941544 592263 941600
rect 592407 941544 592463 941600
rect 601348 940736 601404 940792
rect 601472 940736 601528 940792
rect 601596 940736 601652 940792
rect 601720 940736 601776 940792
rect 601844 940736 601900 940792
rect 601968 940736 602024 940792
rect 602092 940736 602148 940792
rect 602216 940736 602272 940792
rect 602340 940736 602396 940792
rect 602464 940736 602520 940792
rect 602588 940736 602644 940792
rect 602712 940736 602768 940792
rect 602836 940736 602892 940792
rect 602960 940736 603016 940792
rect 603084 940736 603140 940792
rect 601348 940612 601404 940668
rect 601472 940612 601528 940668
rect 601596 940612 601652 940668
rect 601720 940612 601776 940668
rect 601844 940612 601900 940668
rect 601968 940612 602024 940668
rect 602092 940612 602148 940668
rect 602216 940612 602272 940668
rect 602340 940612 602396 940668
rect 602464 940612 602520 940668
rect 602588 940612 602644 940668
rect 602712 940612 602768 940668
rect 602836 940612 602892 940668
rect 602960 940612 603016 940668
rect 603084 940612 603140 940668
rect 601348 940488 601404 940544
rect 601472 940488 601528 940544
rect 601596 940488 601652 940544
rect 601720 940488 601776 940544
rect 601844 940488 601900 940544
rect 601968 940488 602024 940544
rect 602092 940488 602148 940544
rect 602216 940488 602272 940544
rect 602340 940488 602396 940544
rect 602464 940488 602520 940544
rect 602588 940488 602644 940544
rect 602712 940488 602768 940544
rect 602836 940488 602892 940544
rect 602960 940488 603016 940544
rect 603084 940488 603140 940544
rect 601348 940364 601404 940420
rect 601472 940364 601528 940420
rect 601596 940364 601652 940420
rect 601720 940364 601776 940420
rect 601844 940364 601900 940420
rect 601968 940364 602024 940420
rect 602092 940364 602148 940420
rect 602216 940364 602272 940420
rect 602340 940364 602396 940420
rect 602464 940364 602520 940420
rect 602588 940364 602644 940420
rect 602712 940364 602768 940420
rect 602836 940364 602892 940420
rect 602960 940364 603016 940420
rect 603084 940364 603140 940420
rect 601348 940240 601404 940296
rect 601472 940240 601528 940296
rect 601596 940240 601652 940296
rect 601720 940240 601776 940296
rect 601844 940240 601900 940296
rect 601968 940240 602024 940296
rect 602092 940240 602148 940296
rect 602216 940240 602272 940296
rect 602340 940240 602396 940296
rect 602464 940240 602520 940296
rect 602588 940240 602644 940296
rect 602712 940240 602768 940296
rect 602836 940240 602892 940296
rect 602960 940240 603016 940296
rect 603084 940240 603140 940296
rect 601348 940116 601404 940172
rect 601472 940116 601528 940172
rect 601596 940116 601652 940172
rect 601720 940116 601776 940172
rect 601844 940116 601900 940172
rect 601968 940116 602024 940172
rect 602092 940116 602148 940172
rect 602216 940116 602272 940172
rect 602340 940116 602396 940172
rect 602464 940116 602520 940172
rect 602588 940116 602644 940172
rect 602712 940116 602768 940172
rect 602836 940116 602892 940172
rect 602960 940116 603016 940172
rect 603084 940116 603140 940172
rect 601348 939992 601404 940048
rect 601472 939992 601528 940048
rect 601596 939992 601652 940048
rect 601720 939992 601776 940048
rect 601844 939992 601900 940048
rect 601968 939992 602024 940048
rect 602092 939992 602148 940048
rect 602216 939992 602272 940048
rect 602340 939992 602396 940048
rect 602464 939992 602520 940048
rect 602588 939992 602644 940048
rect 602712 939992 602768 940048
rect 602836 939992 602892 940048
rect 602960 939992 603016 940048
rect 603084 939992 603140 940048
rect 603828 940736 603884 940792
rect 603952 940736 604008 940792
rect 604076 940736 604132 940792
rect 604200 940736 604256 940792
rect 604324 940736 604380 940792
rect 604448 940736 604504 940792
rect 604572 940736 604628 940792
rect 604696 940736 604752 940792
rect 604820 940736 604876 940792
rect 604944 940736 605000 940792
rect 605068 940736 605124 940792
rect 605192 940736 605248 940792
rect 605316 940736 605372 940792
rect 605440 940736 605496 940792
rect 605564 940736 605620 940792
rect 605688 940736 605744 940792
rect 603828 940612 603884 940668
rect 603952 940612 604008 940668
rect 604076 940612 604132 940668
rect 604200 940612 604256 940668
rect 604324 940612 604380 940668
rect 604448 940612 604504 940668
rect 604572 940612 604628 940668
rect 604696 940612 604752 940668
rect 604820 940612 604876 940668
rect 604944 940612 605000 940668
rect 605068 940612 605124 940668
rect 605192 940612 605248 940668
rect 605316 940612 605372 940668
rect 605440 940612 605496 940668
rect 605564 940612 605620 940668
rect 605688 940612 605744 940668
rect 603828 940488 603884 940544
rect 603952 940488 604008 940544
rect 604076 940488 604132 940544
rect 604200 940488 604256 940544
rect 604324 940488 604380 940544
rect 604448 940488 604504 940544
rect 604572 940488 604628 940544
rect 604696 940488 604752 940544
rect 604820 940488 604876 940544
rect 604944 940488 605000 940544
rect 605068 940488 605124 940544
rect 605192 940488 605248 940544
rect 605316 940488 605372 940544
rect 605440 940488 605496 940544
rect 605564 940488 605620 940544
rect 605688 940488 605744 940544
rect 603828 940364 603884 940420
rect 603952 940364 604008 940420
rect 604076 940364 604132 940420
rect 604200 940364 604256 940420
rect 604324 940364 604380 940420
rect 604448 940364 604504 940420
rect 604572 940364 604628 940420
rect 604696 940364 604752 940420
rect 604820 940364 604876 940420
rect 604944 940364 605000 940420
rect 605068 940364 605124 940420
rect 605192 940364 605248 940420
rect 605316 940364 605372 940420
rect 605440 940364 605496 940420
rect 605564 940364 605620 940420
rect 605688 940364 605744 940420
rect 603828 940240 603884 940296
rect 603952 940240 604008 940296
rect 604076 940240 604132 940296
rect 604200 940240 604256 940296
rect 604324 940240 604380 940296
rect 604448 940240 604504 940296
rect 604572 940240 604628 940296
rect 604696 940240 604752 940296
rect 604820 940240 604876 940296
rect 604944 940240 605000 940296
rect 605068 940240 605124 940296
rect 605192 940240 605248 940296
rect 605316 940240 605372 940296
rect 605440 940240 605496 940296
rect 605564 940240 605620 940296
rect 605688 940240 605744 940296
rect 603828 940116 603884 940172
rect 603952 940116 604008 940172
rect 604076 940116 604132 940172
rect 604200 940116 604256 940172
rect 604324 940116 604380 940172
rect 604448 940116 604504 940172
rect 604572 940116 604628 940172
rect 604696 940116 604752 940172
rect 604820 940116 604876 940172
rect 604944 940116 605000 940172
rect 605068 940116 605124 940172
rect 605192 940116 605248 940172
rect 605316 940116 605372 940172
rect 605440 940116 605496 940172
rect 605564 940116 605620 940172
rect 605688 940116 605744 940172
rect 603828 939992 603884 940048
rect 603952 939992 604008 940048
rect 604076 939992 604132 940048
rect 604200 939992 604256 940048
rect 604324 939992 604380 940048
rect 604448 939992 604504 940048
rect 604572 939992 604628 940048
rect 604696 939992 604752 940048
rect 604820 939992 604876 940048
rect 604944 939992 605000 940048
rect 605068 939992 605124 940048
rect 605192 939992 605248 940048
rect 605316 939992 605372 940048
rect 605440 939992 605496 940048
rect 605564 939992 605620 940048
rect 605688 939992 605744 940048
rect 606198 940736 606254 940792
rect 606322 940736 606378 940792
rect 606446 940736 606502 940792
rect 606570 940736 606626 940792
rect 606694 940736 606750 940792
rect 606818 940736 606874 940792
rect 606942 940736 606998 940792
rect 607066 940736 607122 940792
rect 607190 940736 607246 940792
rect 607314 940736 607370 940792
rect 607438 940736 607494 940792
rect 607562 940736 607618 940792
rect 607686 940736 607742 940792
rect 607810 940736 607866 940792
rect 607934 940736 607990 940792
rect 608058 940736 608114 940792
rect 606198 940612 606254 940668
rect 606322 940612 606378 940668
rect 606446 940612 606502 940668
rect 606570 940612 606626 940668
rect 606694 940612 606750 940668
rect 606818 940612 606874 940668
rect 606942 940612 606998 940668
rect 607066 940612 607122 940668
rect 607190 940612 607246 940668
rect 607314 940612 607370 940668
rect 607438 940612 607494 940668
rect 607562 940612 607618 940668
rect 607686 940612 607742 940668
rect 607810 940612 607866 940668
rect 607934 940612 607990 940668
rect 608058 940612 608114 940668
rect 606198 940488 606254 940544
rect 606322 940488 606378 940544
rect 606446 940488 606502 940544
rect 606570 940488 606626 940544
rect 606694 940488 606750 940544
rect 606818 940488 606874 940544
rect 606942 940488 606998 940544
rect 607066 940488 607122 940544
rect 607190 940488 607246 940544
rect 607314 940488 607370 940544
rect 607438 940488 607494 940544
rect 607562 940488 607618 940544
rect 607686 940488 607742 940544
rect 607810 940488 607866 940544
rect 607934 940488 607990 940544
rect 608058 940488 608114 940544
rect 606198 940364 606254 940420
rect 606322 940364 606378 940420
rect 606446 940364 606502 940420
rect 606570 940364 606626 940420
rect 606694 940364 606750 940420
rect 606818 940364 606874 940420
rect 606942 940364 606998 940420
rect 607066 940364 607122 940420
rect 607190 940364 607246 940420
rect 607314 940364 607370 940420
rect 607438 940364 607494 940420
rect 607562 940364 607618 940420
rect 607686 940364 607742 940420
rect 607810 940364 607866 940420
rect 607934 940364 607990 940420
rect 608058 940364 608114 940420
rect 606198 940240 606254 940296
rect 606322 940240 606378 940296
rect 606446 940240 606502 940296
rect 606570 940240 606626 940296
rect 606694 940240 606750 940296
rect 606818 940240 606874 940296
rect 606942 940240 606998 940296
rect 607066 940240 607122 940296
rect 607190 940240 607246 940296
rect 607314 940240 607370 940296
rect 607438 940240 607494 940296
rect 607562 940240 607618 940296
rect 607686 940240 607742 940296
rect 607810 940240 607866 940296
rect 607934 940240 607990 940296
rect 608058 940240 608114 940296
rect 606198 940116 606254 940172
rect 606322 940116 606378 940172
rect 606446 940116 606502 940172
rect 606570 940116 606626 940172
rect 606694 940116 606750 940172
rect 606818 940116 606874 940172
rect 606942 940116 606998 940172
rect 607066 940116 607122 940172
rect 607190 940116 607246 940172
rect 607314 940116 607370 940172
rect 607438 940116 607494 940172
rect 607562 940116 607618 940172
rect 607686 940116 607742 940172
rect 607810 940116 607866 940172
rect 607934 940116 607990 940172
rect 608058 940116 608114 940172
rect 606198 939992 606254 940048
rect 606322 939992 606378 940048
rect 606446 939992 606502 940048
rect 606570 939992 606626 940048
rect 606694 939992 606750 940048
rect 606818 939992 606874 940048
rect 606942 939992 606998 940048
rect 607066 939992 607122 940048
rect 607190 939992 607246 940048
rect 607314 939992 607370 940048
rect 607438 939992 607494 940048
rect 607562 939992 607618 940048
rect 607686 939992 607742 940048
rect 607810 939992 607866 940048
rect 607934 939992 607990 940048
rect 608058 939992 608114 940048
rect 608904 940736 608960 940792
rect 609028 940736 609084 940792
rect 609152 940736 609208 940792
rect 609276 940736 609332 940792
rect 609400 940736 609456 940792
rect 609524 940736 609580 940792
rect 609648 940736 609704 940792
rect 609772 940736 609828 940792
rect 609896 940736 609952 940792
rect 610020 940736 610076 940792
rect 610144 940736 610200 940792
rect 610268 940736 610324 940792
rect 610392 940736 610448 940792
rect 610516 940736 610572 940792
rect 610640 940736 610696 940792
rect 610764 940736 610820 940792
rect 608904 940612 608960 940668
rect 609028 940612 609084 940668
rect 609152 940612 609208 940668
rect 609276 940612 609332 940668
rect 609400 940612 609456 940668
rect 609524 940612 609580 940668
rect 609648 940612 609704 940668
rect 609772 940612 609828 940668
rect 609896 940612 609952 940668
rect 610020 940612 610076 940668
rect 610144 940612 610200 940668
rect 610268 940612 610324 940668
rect 610392 940612 610448 940668
rect 610516 940612 610572 940668
rect 610640 940612 610696 940668
rect 610764 940612 610820 940668
rect 608904 940488 608960 940544
rect 609028 940488 609084 940544
rect 609152 940488 609208 940544
rect 609276 940488 609332 940544
rect 609400 940488 609456 940544
rect 609524 940488 609580 940544
rect 609648 940488 609704 940544
rect 609772 940488 609828 940544
rect 609896 940488 609952 940544
rect 610020 940488 610076 940544
rect 610144 940488 610200 940544
rect 610268 940488 610324 940544
rect 610392 940488 610448 940544
rect 610516 940488 610572 940544
rect 610640 940488 610696 940544
rect 610764 940488 610820 940544
rect 608904 940364 608960 940420
rect 609028 940364 609084 940420
rect 609152 940364 609208 940420
rect 609276 940364 609332 940420
rect 609400 940364 609456 940420
rect 609524 940364 609580 940420
rect 609648 940364 609704 940420
rect 609772 940364 609828 940420
rect 609896 940364 609952 940420
rect 610020 940364 610076 940420
rect 610144 940364 610200 940420
rect 610268 940364 610324 940420
rect 610392 940364 610448 940420
rect 610516 940364 610572 940420
rect 610640 940364 610696 940420
rect 610764 940364 610820 940420
rect 608904 940240 608960 940296
rect 609028 940240 609084 940296
rect 609152 940240 609208 940296
rect 609276 940240 609332 940296
rect 609400 940240 609456 940296
rect 609524 940240 609580 940296
rect 609648 940240 609704 940296
rect 609772 940240 609828 940296
rect 609896 940240 609952 940296
rect 610020 940240 610076 940296
rect 610144 940240 610200 940296
rect 610268 940240 610324 940296
rect 610392 940240 610448 940296
rect 610516 940240 610572 940296
rect 610640 940240 610696 940296
rect 610764 940240 610820 940296
rect 608904 940116 608960 940172
rect 609028 940116 609084 940172
rect 609152 940116 609208 940172
rect 609276 940116 609332 940172
rect 609400 940116 609456 940172
rect 609524 940116 609580 940172
rect 609648 940116 609704 940172
rect 609772 940116 609828 940172
rect 609896 940116 609952 940172
rect 610020 940116 610076 940172
rect 610144 940116 610200 940172
rect 610268 940116 610324 940172
rect 610392 940116 610448 940172
rect 610516 940116 610572 940172
rect 610640 940116 610696 940172
rect 610764 940116 610820 940172
rect 608904 939992 608960 940048
rect 609028 939992 609084 940048
rect 609152 939992 609208 940048
rect 609276 939992 609332 940048
rect 609400 939992 609456 940048
rect 609524 939992 609580 940048
rect 609648 939992 609704 940048
rect 609772 939992 609828 940048
rect 609896 939992 609952 940048
rect 610020 939992 610076 940048
rect 610144 939992 610200 940048
rect 610268 939992 610324 940048
rect 610392 939992 610448 940048
rect 610516 939992 610572 940048
rect 610640 939992 610696 940048
rect 610764 939992 610820 940048
rect 611274 940736 611330 940792
rect 611398 940736 611454 940792
rect 611522 940736 611578 940792
rect 611646 940736 611702 940792
rect 611770 940736 611826 940792
rect 611894 940736 611950 940792
rect 612018 940736 612074 940792
rect 612142 940736 612198 940792
rect 612266 940736 612322 940792
rect 612390 940736 612446 940792
rect 612514 940736 612570 940792
rect 612638 940736 612694 940792
rect 612762 940736 612818 940792
rect 612886 940736 612942 940792
rect 613010 940736 613066 940792
rect 613134 940736 613190 940792
rect 611274 940612 611330 940668
rect 611398 940612 611454 940668
rect 611522 940612 611578 940668
rect 611646 940612 611702 940668
rect 611770 940612 611826 940668
rect 611894 940612 611950 940668
rect 612018 940612 612074 940668
rect 612142 940612 612198 940668
rect 612266 940612 612322 940668
rect 612390 940612 612446 940668
rect 612514 940612 612570 940668
rect 612638 940612 612694 940668
rect 612762 940612 612818 940668
rect 612886 940612 612942 940668
rect 613010 940612 613066 940668
rect 613134 940612 613190 940668
rect 611274 940488 611330 940544
rect 611398 940488 611454 940544
rect 611522 940488 611578 940544
rect 611646 940488 611702 940544
rect 611770 940488 611826 940544
rect 611894 940488 611950 940544
rect 612018 940488 612074 940544
rect 612142 940488 612198 940544
rect 612266 940488 612322 940544
rect 612390 940488 612446 940544
rect 612514 940488 612570 940544
rect 612638 940488 612694 940544
rect 612762 940488 612818 940544
rect 612886 940488 612942 940544
rect 613010 940488 613066 940544
rect 613134 940488 613190 940544
rect 611274 940364 611330 940420
rect 611398 940364 611454 940420
rect 611522 940364 611578 940420
rect 611646 940364 611702 940420
rect 611770 940364 611826 940420
rect 611894 940364 611950 940420
rect 612018 940364 612074 940420
rect 612142 940364 612198 940420
rect 612266 940364 612322 940420
rect 612390 940364 612446 940420
rect 612514 940364 612570 940420
rect 612638 940364 612694 940420
rect 612762 940364 612818 940420
rect 612886 940364 612942 940420
rect 613010 940364 613066 940420
rect 613134 940364 613190 940420
rect 611274 940240 611330 940296
rect 611398 940240 611454 940296
rect 611522 940240 611578 940296
rect 611646 940240 611702 940296
rect 611770 940240 611826 940296
rect 611894 940240 611950 940296
rect 612018 940240 612074 940296
rect 612142 940240 612198 940296
rect 612266 940240 612322 940296
rect 612390 940240 612446 940296
rect 612514 940240 612570 940296
rect 612638 940240 612694 940296
rect 612762 940240 612818 940296
rect 612886 940240 612942 940296
rect 613010 940240 613066 940296
rect 613134 940240 613190 940296
rect 611274 940116 611330 940172
rect 611398 940116 611454 940172
rect 611522 940116 611578 940172
rect 611646 940116 611702 940172
rect 611770 940116 611826 940172
rect 611894 940116 611950 940172
rect 612018 940116 612074 940172
rect 612142 940116 612198 940172
rect 612266 940116 612322 940172
rect 612390 940116 612446 940172
rect 612514 940116 612570 940172
rect 612638 940116 612694 940172
rect 612762 940116 612818 940172
rect 612886 940116 612942 940172
rect 613010 940116 613066 940172
rect 613134 940116 613190 940172
rect 611274 939992 611330 940048
rect 611398 939992 611454 940048
rect 611522 939992 611578 940048
rect 611646 939992 611702 940048
rect 611770 939992 611826 940048
rect 611894 939992 611950 940048
rect 612018 939992 612074 940048
rect 612142 939992 612198 940048
rect 612266 939992 612322 940048
rect 612390 939992 612446 940048
rect 612514 939992 612570 940048
rect 612638 939992 612694 940048
rect 612762 939992 612818 940048
rect 612886 939992 612942 940048
rect 613010 939992 613066 940048
rect 613134 939992 613190 940048
rect 660548 943379 660604 943435
rect 613878 940736 613934 940792
rect 614002 940736 614058 940792
rect 614126 940736 614182 940792
rect 614250 940736 614306 940792
rect 614374 940736 614430 940792
rect 614498 940736 614554 940792
rect 614622 940736 614678 940792
rect 614746 940736 614802 940792
rect 614870 940736 614926 940792
rect 614994 940736 615050 940792
rect 615118 940736 615174 940792
rect 615242 940736 615298 940792
rect 615366 940736 615422 940792
rect 615490 940736 615546 940792
rect 615614 940736 615670 940792
rect 613878 940612 613934 940668
rect 614002 940612 614058 940668
rect 614126 940612 614182 940668
rect 614250 940612 614306 940668
rect 614374 940612 614430 940668
rect 614498 940612 614554 940668
rect 614622 940612 614678 940668
rect 614746 940612 614802 940668
rect 614870 940612 614926 940668
rect 614994 940612 615050 940668
rect 615118 940612 615174 940668
rect 615242 940612 615298 940668
rect 615366 940612 615422 940668
rect 615490 940612 615546 940668
rect 615614 940612 615670 940668
rect 613878 940488 613934 940544
rect 614002 940488 614058 940544
rect 614126 940488 614182 940544
rect 614250 940488 614306 940544
rect 614374 940488 614430 940544
rect 614498 940488 614554 940544
rect 614622 940488 614678 940544
rect 614746 940488 614802 940544
rect 614870 940488 614926 940544
rect 614994 940488 615050 940544
rect 615118 940488 615174 940544
rect 615242 940488 615298 940544
rect 615366 940488 615422 940544
rect 615490 940488 615546 940544
rect 615614 940488 615670 940544
rect 613878 940364 613934 940420
rect 614002 940364 614058 940420
rect 614126 940364 614182 940420
rect 614250 940364 614306 940420
rect 614374 940364 614430 940420
rect 614498 940364 614554 940420
rect 614622 940364 614678 940420
rect 614746 940364 614802 940420
rect 614870 940364 614926 940420
rect 614994 940364 615050 940420
rect 615118 940364 615174 940420
rect 615242 940364 615298 940420
rect 615366 940364 615422 940420
rect 615490 940364 615546 940420
rect 615614 940364 615670 940420
rect 613878 940240 613934 940296
rect 614002 940240 614058 940296
rect 614126 940240 614182 940296
rect 614250 940240 614306 940296
rect 614374 940240 614430 940296
rect 614498 940240 614554 940296
rect 614622 940240 614678 940296
rect 614746 940240 614802 940296
rect 614870 940240 614926 940296
rect 614994 940240 615050 940296
rect 615118 940240 615174 940296
rect 615242 940240 615298 940296
rect 615366 940240 615422 940296
rect 615490 940240 615546 940296
rect 615614 940240 615670 940296
rect 613878 940116 613934 940172
rect 614002 940116 614058 940172
rect 614126 940116 614182 940172
rect 614250 940116 614306 940172
rect 614374 940116 614430 940172
rect 614498 940116 614554 940172
rect 614622 940116 614678 940172
rect 614746 940116 614802 940172
rect 614870 940116 614926 940172
rect 614994 940116 615050 940172
rect 615118 940116 615174 940172
rect 615242 940116 615298 940172
rect 615366 940116 615422 940172
rect 615490 940116 615546 940172
rect 615614 940116 615670 940172
rect 613878 939992 613934 940048
rect 614002 939992 614058 940048
rect 614126 939992 614182 940048
rect 614250 939992 614306 940048
rect 614374 939992 614430 940048
rect 614498 939992 614554 940048
rect 614622 939992 614678 940048
rect 614746 939992 614802 940048
rect 614870 939992 614926 940048
rect 614994 939992 615050 940048
rect 615118 939992 615174 940048
rect 615242 939992 615298 940048
rect 615366 939992 615422 940048
rect 615490 939992 615546 940048
rect 615614 939992 615670 940048
rect 628207 942144 628263 942200
rect 628407 942144 628463 942200
rect 628207 941844 628263 941900
rect 628407 941844 628463 941900
rect 628207 941544 628263 941600
rect 628407 941544 628463 941600
rect 646207 940744 646263 940800
rect 646407 940744 646463 940800
rect 646207 940444 646263 940500
rect 646407 940444 646463 940500
rect 646207 940144 646263 940200
rect 646407 940144 646463 940200
rect 667548 943379 667604 943435
rect 660546 940654 660602 940710
rect 660546 940354 660602 940410
rect 660546 940054 660602 940110
rect 664207 942144 664263 942200
rect 664407 942144 664463 942200
rect 664207 941844 664263 941900
rect 664407 941844 664463 941900
rect 664207 941544 664263 941600
rect 664407 941544 664463 941600
rect 667546 940654 667602 940710
rect 667546 940354 667602 940410
rect 667546 940054 667602 940110
rect 674548 943379 674604 943435
rect 690406 942097 690462 942153
rect 690406 941797 690462 941853
rect 690406 941497 690462 941553
rect 674546 940654 674602 940710
rect 674546 940354 674602 940410
rect 674546 940054 674602 940110
rect 682207 940744 682263 940800
rect 682407 940744 682463 940800
rect 682207 940444 682263 940500
rect 682407 940444 682463 940500
rect 682207 940144 682263 940200
rect 682407 940144 682463 940200
rect 699452 942136 699508 942192
rect 699576 942136 699632 942192
rect 699700 942136 699756 942192
rect 699824 942136 699880 942192
rect 699948 942136 700004 942192
rect 700072 942136 700128 942192
rect 700196 942136 700252 942192
rect 699452 942012 699508 942068
rect 699576 942012 699632 942068
rect 699700 942012 699756 942068
rect 699824 942012 699880 942068
rect 699948 942012 700004 942068
rect 700072 942012 700128 942068
rect 700196 942012 700252 942068
rect 699452 941888 699508 941944
rect 699576 941888 699632 941944
rect 699700 941888 699756 941944
rect 699824 941888 699880 941944
rect 699948 941888 700004 941944
rect 700072 941888 700128 941944
rect 700196 941888 700252 941944
rect 699452 941764 699508 941820
rect 699576 941764 699632 941820
rect 699700 941764 699756 941820
rect 699824 941764 699880 941820
rect 699948 941764 700004 941820
rect 700072 941764 700128 941820
rect 700196 941764 700252 941820
rect 699452 941640 699508 941696
rect 699576 941640 699632 941696
rect 699700 941640 699756 941696
rect 699824 941640 699880 941696
rect 699948 941640 700004 941696
rect 700072 941640 700128 941696
rect 700196 941640 700252 941696
rect 699452 941516 699508 941572
rect 699576 941516 699632 941572
rect 699700 941516 699756 941572
rect 699824 941516 699880 941572
rect 699948 941516 700004 941572
rect 700072 941516 700128 941572
rect 700196 941516 700252 941572
rect 699452 941392 699508 941448
rect 699576 941392 699632 941448
rect 699700 941392 699756 941448
rect 699824 941392 699880 941448
rect 699948 941392 700004 941448
rect 700072 941392 700128 941448
rect 700196 941392 700252 941448
rect 690821 940660 690877 940716
rect 690821 940360 690877 940416
rect 690821 940060 690877 940116
rect 698052 940736 698108 940792
rect 698176 940736 698232 940792
rect 698300 940736 698356 940792
rect 698424 940736 698480 940792
rect 698548 940736 698604 940792
rect 698672 940736 698728 940792
rect 698796 940736 698852 940792
rect 698052 940612 698108 940668
rect 698176 940612 698232 940668
rect 698300 940612 698356 940668
rect 698424 940612 698480 940668
rect 698548 940612 698604 940668
rect 698672 940612 698728 940668
rect 698796 940612 698852 940668
rect 698052 940488 698108 940544
rect 698176 940488 698232 940544
rect 698300 940488 698356 940544
rect 698424 940488 698480 940544
rect 698548 940488 698604 940544
rect 698672 940488 698728 940544
rect 698796 940488 698852 940544
rect 698052 940364 698108 940420
rect 698176 940364 698232 940420
rect 698300 940364 698356 940420
rect 698424 940364 698480 940420
rect 698548 940364 698604 940420
rect 698672 940364 698728 940420
rect 698796 940364 698852 940420
rect 698052 940240 698108 940296
rect 698176 940240 698232 940296
rect 698300 940240 698356 940296
rect 698424 940240 698480 940296
rect 698548 940240 698604 940296
rect 698672 940240 698728 940296
rect 698796 940240 698852 940296
rect 698052 940116 698108 940172
rect 698176 940116 698232 940172
rect 698300 940116 698356 940172
rect 698424 940116 698480 940172
rect 698548 940116 698604 940172
rect 698672 940116 698728 940172
rect 698796 940116 698852 940172
rect 698052 939992 698108 940048
rect 698176 939992 698232 940048
rect 698300 939992 698356 940048
rect 698424 939992 698480 940048
rect 698548 939992 698604 940048
rect 698672 939992 698728 940048
rect 698796 939992 698852 940048
rect 79300 929566 79356 929622
rect 79600 929566 79656 929622
rect 79900 929566 79956 929622
rect 79300 922566 79356 922622
rect 79600 922566 79656 922622
rect 79900 922566 79956 922622
rect 79300 915566 79356 915622
rect 79600 915566 79656 915622
rect 79900 915566 79956 915622
rect 79200 896373 79256 896429
rect 79500 896373 79556 896429
rect 79800 896373 79856 896429
rect 79200 896173 79256 896229
rect 79500 896173 79556 896229
rect 79800 896173 79856 896229
rect 79200 860373 79256 860429
rect 79500 860373 79556 860429
rect 79800 860373 79856 860429
rect 79200 860173 79256 860229
rect 79500 860173 79556 860229
rect 79800 860173 79856 860229
rect 79200 824373 79256 824429
rect 79500 824373 79556 824429
rect 79800 824373 79856 824429
rect 79200 824173 79256 824229
rect 79500 824173 79556 824229
rect 79800 824173 79856 824229
rect 79208 802614 79264 802670
rect 79332 802614 79388 802670
rect 79456 802614 79512 802670
rect 79580 802614 79636 802670
rect 79704 802614 79760 802670
rect 79828 802614 79884 802670
rect 79952 802614 80008 802670
rect 79208 802490 79264 802546
rect 79332 802490 79388 802546
rect 79456 802490 79512 802546
rect 79580 802490 79636 802546
rect 79704 802490 79760 802546
rect 79828 802490 79884 802546
rect 79952 802490 80008 802546
rect 79208 802366 79264 802422
rect 79332 802366 79388 802422
rect 79456 802366 79512 802422
rect 79580 802366 79636 802422
rect 79704 802366 79760 802422
rect 79828 802366 79884 802422
rect 79952 802366 80008 802422
rect 79208 802242 79264 802298
rect 79332 802242 79388 802298
rect 79456 802242 79512 802298
rect 79580 802242 79636 802298
rect 79704 802242 79760 802298
rect 79828 802242 79884 802298
rect 79952 802242 80008 802298
rect 79208 802118 79264 802174
rect 79332 802118 79388 802174
rect 79456 802118 79512 802174
rect 79580 802118 79636 802174
rect 79704 802118 79760 802174
rect 79828 802118 79884 802174
rect 79952 802118 80008 802174
rect 79208 801994 79264 802050
rect 79332 801994 79388 802050
rect 79456 801994 79512 802050
rect 79580 801994 79636 802050
rect 79704 801994 79760 802050
rect 79828 801994 79884 802050
rect 79952 801994 80008 802050
rect 79208 801870 79264 801926
rect 79332 801870 79388 801926
rect 79456 801870 79512 801926
rect 79580 801870 79636 801926
rect 79704 801870 79760 801926
rect 79828 801870 79884 801926
rect 79952 801870 80008 801926
rect 79208 801746 79264 801802
rect 79332 801746 79388 801802
rect 79456 801746 79512 801802
rect 79580 801746 79636 801802
rect 79704 801746 79760 801802
rect 79828 801746 79884 801802
rect 79952 801746 80008 801802
rect 79208 801622 79264 801678
rect 79332 801622 79388 801678
rect 79456 801622 79512 801678
rect 79580 801622 79636 801678
rect 79704 801622 79760 801678
rect 79828 801622 79884 801678
rect 79952 801622 80008 801678
rect 79208 801498 79264 801554
rect 79332 801498 79388 801554
rect 79456 801498 79512 801554
rect 79580 801498 79636 801554
rect 79704 801498 79760 801554
rect 79828 801498 79884 801554
rect 79952 801498 80008 801554
rect 79208 801374 79264 801430
rect 79332 801374 79388 801430
rect 79456 801374 79512 801430
rect 79580 801374 79636 801430
rect 79704 801374 79760 801430
rect 79828 801374 79884 801430
rect 79952 801374 80008 801430
rect 79208 801250 79264 801306
rect 79332 801250 79388 801306
rect 79456 801250 79512 801306
rect 79580 801250 79636 801306
rect 79704 801250 79760 801306
rect 79828 801250 79884 801306
rect 79952 801250 80008 801306
rect 79208 801126 79264 801182
rect 79332 801126 79388 801182
rect 79456 801126 79512 801182
rect 79580 801126 79636 801182
rect 79704 801126 79760 801182
rect 79828 801126 79884 801182
rect 79952 801126 80008 801182
rect 79208 801002 79264 801058
rect 79332 801002 79388 801058
rect 79456 801002 79512 801058
rect 79580 801002 79636 801058
rect 79704 801002 79760 801058
rect 79828 801002 79884 801058
rect 79952 801002 80008 801058
rect 79208 800878 79264 800934
rect 79332 800878 79388 800934
rect 79456 800878 79512 800934
rect 79580 800878 79636 800934
rect 79704 800878 79760 800934
rect 79828 800878 79884 800934
rect 79952 800878 80008 800934
rect 79208 800134 79264 800190
rect 79332 800134 79388 800190
rect 79456 800134 79512 800190
rect 79580 800134 79636 800190
rect 79704 800134 79760 800190
rect 79828 800134 79884 800190
rect 79952 800134 80008 800190
rect 79208 800010 79264 800066
rect 79332 800010 79388 800066
rect 79456 800010 79512 800066
rect 79580 800010 79636 800066
rect 79704 800010 79760 800066
rect 79828 800010 79884 800066
rect 79952 800010 80008 800066
rect 79208 799886 79264 799942
rect 79332 799886 79388 799942
rect 79456 799886 79512 799942
rect 79580 799886 79636 799942
rect 79704 799886 79760 799942
rect 79828 799886 79884 799942
rect 79952 799886 80008 799942
rect 79208 799762 79264 799818
rect 79332 799762 79388 799818
rect 79456 799762 79512 799818
rect 79580 799762 79636 799818
rect 79704 799762 79760 799818
rect 79828 799762 79884 799818
rect 79952 799762 80008 799818
rect 79208 799638 79264 799694
rect 79332 799638 79388 799694
rect 79456 799638 79512 799694
rect 79580 799638 79636 799694
rect 79704 799638 79760 799694
rect 79828 799638 79884 799694
rect 79952 799638 80008 799694
rect 79208 799514 79264 799570
rect 79332 799514 79388 799570
rect 79456 799514 79512 799570
rect 79580 799514 79636 799570
rect 79704 799514 79760 799570
rect 79828 799514 79884 799570
rect 79952 799514 80008 799570
rect 79208 799390 79264 799446
rect 79332 799390 79388 799446
rect 79456 799390 79512 799446
rect 79580 799390 79636 799446
rect 79704 799390 79760 799446
rect 79828 799390 79884 799446
rect 79952 799390 80008 799446
rect 79208 799266 79264 799322
rect 79332 799266 79388 799322
rect 79456 799266 79512 799322
rect 79580 799266 79636 799322
rect 79704 799266 79760 799322
rect 79828 799266 79884 799322
rect 79952 799266 80008 799322
rect 79208 799142 79264 799198
rect 79332 799142 79388 799198
rect 79456 799142 79512 799198
rect 79580 799142 79636 799198
rect 79704 799142 79760 799198
rect 79828 799142 79884 799198
rect 79952 799142 80008 799198
rect 79208 799018 79264 799074
rect 79332 799018 79388 799074
rect 79456 799018 79512 799074
rect 79580 799018 79636 799074
rect 79704 799018 79760 799074
rect 79828 799018 79884 799074
rect 79952 799018 80008 799074
rect 79208 798894 79264 798950
rect 79332 798894 79388 798950
rect 79456 798894 79512 798950
rect 79580 798894 79636 798950
rect 79704 798894 79760 798950
rect 79828 798894 79884 798950
rect 79952 798894 80008 798950
rect 79208 798770 79264 798826
rect 79332 798770 79388 798826
rect 79456 798770 79512 798826
rect 79580 798770 79636 798826
rect 79704 798770 79760 798826
rect 79828 798770 79884 798826
rect 79952 798770 80008 798826
rect 79208 798646 79264 798702
rect 79332 798646 79388 798702
rect 79456 798646 79512 798702
rect 79580 798646 79636 798702
rect 79704 798646 79760 798702
rect 79828 798646 79884 798702
rect 79952 798646 80008 798702
rect 79208 798522 79264 798578
rect 79332 798522 79388 798578
rect 79456 798522 79512 798578
rect 79580 798522 79636 798578
rect 79704 798522 79760 798578
rect 79828 798522 79884 798578
rect 79952 798522 80008 798578
rect 79208 798398 79264 798454
rect 79332 798398 79388 798454
rect 79456 798398 79512 798454
rect 79580 798398 79636 798454
rect 79704 798398 79760 798454
rect 79828 798398 79884 798454
rect 79952 798398 80008 798454
rect 79208 798274 79264 798330
rect 79332 798274 79388 798330
rect 79456 798274 79512 798330
rect 79580 798274 79636 798330
rect 79704 798274 79760 798330
rect 79828 798274 79884 798330
rect 79952 798274 80008 798330
rect 79208 797764 79264 797820
rect 79332 797764 79388 797820
rect 79456 797764 79512 797820
rect 79580 797764 79636 797820
rect 79704 797764 79760 797820
rect 79828 797764 79884 797820
rect 79952 797764 80008 797820
rect 79208 797640 79264 797696
rect 79332 797640 79388 797696
rect 79456 797640 79512 797696
rect 79580 797640 79636 797696
rect 79704 797640 79760 797696
rect 79828 797640 79884 797696
rect 79952 797640 80008 797696
rect 79208 797516 79264 797572
rect 79332 797516 79388 797572
rect 79456 797516 79512 797572
rect 79580 797516 79636 797572
rect 79704 797516 79760 797572
rect 79828 797516 79884 797572
rect 79952 797516 80008 797572
rect 79208 797392 79264 797448
rect 79332 797392 79388 797448
rect 79456 797392 79512 797448
rect 79580 797392 79636 797448
rect 79704 797392 79760 797448
rect 79828 797392 79884 797448
rect 79952 797392 80008 797448
rect 79208 797268 79264 797324
rect 79332 797268 79388 797324
rect 79456 797268 79512 797324
rect 79580 797268 79636 797324
rect 79704 797268 79760 797324
rect 79828 797268 79884 797324
rect 79952 797268 80008 797324
rect 79208 797144 79264 797200
rect 79332 797144 79388 797200
rect 79456 797144 79512 797200
rect 79580 797144 79636 797200
rect 79704 797144 79760 797200
rect 79828 797144 79884 797200
rect 79952 797144 80008 797200
rect 79208 797020 79264 797076
rect 79332 797020 79388 797076
rect 79456 797020 79512 797076
rect 79580 797020 79636 797076
rect 79704 797020 79760 797076
rect 79828 797020 79884 797076
rect 79952 797020 80008 797076
rect 79208 796896 79264 796952
rect 79332 796896 79388 796952
rect 79456 796896 79512 796952
rect 79580 796896 79636 796952
rect 79704 796896 79760 796952
rect 79828 796896 79884 796952
rect 79952 796896 80008 796952
rect 79208 796772 79264 796828
rect 79332 796772 79388 796828
rect 79456 796772 79512 796828
rect 79580 796772 79636 796828
rect 79704 796772 79760 796828
rect 79828 796772 79884 796828
rect 79952 796772 80008 796828
rect 79208 796648 79264 796704
rect 79332 796648 79388 796704
rect 79456 796648 79512 796704
rect 79580 796648 79636 796704
rect 79704 796648 79760 796704
rect 79828 796648 79884 796704
rect 79952 796648 80008 796704
rect 79208 796524 79264 796580
rect 79332 796524 79388 796580
rect 79456 796524 79512 796580
rect 79580 796524 79636 796580
rect 79704 796524 79760 796580
rect 79828 796524 79884 796580
rect 79952 796524 80008 796580
rect 79208 796400 79264 796456
rect 79332 796400 79388 796456
rect 79456 796400 79512 796456
rect 79580 796400 79636 796456
rect 79704 796400 79760 796456
rect 79828 796400 79884 796456
rect 79952 796400 80008 796456
rect 79208 796276 79264 796332
rect 79332 796276 79388 796332
rect 79456 796276 79512 796332
rect 79580 796276 79636 796332
rect 79704 796276 79760 796332
rect 79828 796276 79884 796332
rect 79952 796276 80008 796332
rect 79208 796152 79264 796208
rect 79332 796152 79388 796208
rect 79456 796152 79512 796208
rect 79580 796152 79636 796208
rect 79704 796152 79760 796208
rect 79828 796152 79884 796208
rect 79952 796152 80008 796208
rect 79208 796028 79264 796084
rect 79332 796028 79388 796084
rect 79456 796028 79512 796084
rect 79580 796028 79636 796084
rect 79704 796028 79760 796084
rect 79828 796028 79884 796084
rect 79952 796028 80008 796084
rect 79208 795904 79264 795960
rect 79332 795904 79388 795960
rect 79456 795904 79512 795960
rect 79580 795904 79636 795960
rect 79704 795904 79760 795960
rect 79828 795904 79884 795960
rect 79952 795904 80008 795960
rect 79208 795058 79264 795114
rect 79332 795058 79388 795114
rect 79456 795058 79512 795114
rect 79580 795058 79636 795114
rect 79704 795058 79760 795114
rect 79828 795058 79884 795114
rect 79952 795058 80008 795114
rect 79208 794934 79264 794990
rect 79332 794934 79388 794990
rect 79456 794934 79512 794990
rect 79580 794934 79636 794990
rect 79704 794934 79760 794990
rect 79828 794934 79884 794990
rect 79952 794934 80008 794990
rect 79208 794810 79264 794866
rect 79332 794810 79388 794866
rect 79456 794810 79512 794866
rect 79580 794810 79636 794866
rect 79704 794810 79760 794866
rect 79828 794810 79884 794866
rect 79952 794810 80008 794866
rect 79208 794686 79264 794742
rect 79332 794686 79388 794742
rect 79456 794686 79512 794742
rect 79580 794686 79636 794742
rect 79704 794686 79760 794742
rect 79828 794686 79884 794742
rect 79952 794686 80008 794742
rect 79208 794562 79264 794618
rect 79332 794562 79388 794618
rect 79456 794562 79512 794618
rect 79580 794562 79636 794618
rect 79704 794562 79760 794618
rect 79828 794562 79884 794618
rect 79952 794562 80008 794618
rect 79208 794438 79264 794494
rect 79332 794438 79388 794494
rect 79456 794438 79512 794494
rect 79580 794438 79636 794494
rect 79704 794438 79760 794494
rect 79828 794438 79884 794494
rect 79952 794438 80008 794494
rect 79208 794314 79264 794370
rect 79332 794314 79388 794370
rect 79456 794314 79512 794370
rect 79580 794314 79636 794370
rect 79704 794314 79760 794370
rect 79828 794314 79884 794370
rect 79952 794314 80008 794370
rect 79208 794190 79264 794246
rect 79332 794190 79388 794246
rect 79456 794190 79512 794246
rect 79580 794190 79636 794246
rect 79704 794190 79760 794246
rect 79828 794190 79884 794246
rect 79952 794190 80008 794246
rect 79208 794066 79264 794122
rect 79332 794066 79388 794122
rect 79456 794066 79512 794122
rect 79580 794066 79636 794122
rect 79704 794066 79760 794122
rect 79828 794066 79884 794122
rect 79952 794066 80008 794122
rect 79208 793942 79264 793998
rect 79332 793942 79388 793998
rect 79456 793942 79512 793998
rect 79580 793942 79636 793998
rect 79704 793942 79760 793998
rect 79828 793942 79884 793998
rect 79952 793942 80008 793998
rect 79208 793818 79264 793874
rect 79332 793818 79388 793874
rect 79456 793818 79512 793874
rect 79580 793818 79636 793874
rect 79704 793818 79760 793874
rect 79828 793818 79884 793874
rect 79952 793818 80008 793874
rect 79208 793694 79264 793750
rect 79332 793694 79388 793750
rect 79456 793694 79512 793750
rect 79580 793694 79636 793750
rect 79704 793694 79760 793750
rect 79828 793694 79884 793750
rect 79952 793694 80008 793750
rect 79208 793570 79264 793626
rect 79332 793570 79388 793626
rect 79456 793570 79512 793626
rect 79580 793570 79636 793626
rect 79704 793570 79760 793626
rect 79828 793570 79884 793626
rect 79952 793570 80008 793626
rect 79208 793446 79264 793502
rect 79332 793446 79388 793502
rect 79456 793446 79512 793502
rect 79580 793446 79636 793502
rect 79704 793446 79760 793502
rect 79828 793446 79884 793502
rect 79952 793446 80008 793502
rect 79208 793322 79264 793378
rect 79332 793322 79388 793378
rect 79456 793322 79512 793378
rect 79580 793322 79636 793378
rect 79704 793322 79760 793378
rect 79828 793322 79884 793378
rect 79952 793322 80008 793378
rect 79208 793198 79264 793254
rect 79332 793198 79388 793254
rect 79456 793198 79512 793254
rect 79580 793198 79636 793254
rect 79704 793198 79760 793254
rect 79828 793198 79884 793254
rect 79952 793198 80008 793254
rect 79208 792688 79264 792744
rect 79332 792688 79388 792744
rect 79456 792688 79512 792744
rect 79580 792688 79636 792744
rect 79704 792688 79760 792744
rect 79828 792688 79884 792744
rect 79952 792688 80008 792744
rect 79208 792564 79264 792620
rect 79332 792564 79388 792620
rect 79456 792564 79512 792620
rect 79580 792564 79636 792620
rect 79704 792564 79760 792620
rect 79828 792564 79884 792620
rect 79952 792564 80008 792620
rect 79208 792440 79264 792496
rect 79332 792440 79388 792496
rect 79456 792440 79512 792496
rect 79580 792440 79636 792496
rect 79704 792440 79760 792496
rect 79828 792440 79884 792496
rect 79952 792440 80008 792496
rect 79208 792316 79264 792372
rect 79332 792316 79388 792372
rect 79456 792316 79512 792372
rect 79580 792316 79636 792372
rect 79704 792316 79760 792372
rect 79828 792316 79884 792372
rect 79952 792316 80008 792372
rect 79208 792192 79264 792248
rect 79332 792192 79388 792248
rect 79456 792192 79512 792248
rect 79580 792192 79636 792248
rect 79704 792192 79760 792248
rect 79828 792192 79884 792248
rect 79952 792192 80008 792248
rect 79208 792068 79264 792124
rect 79332 792068 79388 792124
rect 79456 792068 79512 792124
rect 79580 792068 79636 792124
rect 79704 792068 79760 792124
rect 79828 792068 79884 792124
rect 79952 792068 80008 792124
rect 79208 791944 79264 792000
rect 79332 791944 79388 792000
rect 79456 791944 79512 792000
rect 79580 791944 79636 792000
rect 79704 791944 79760 792000
rect 79828 791944 79884 792000
rect 79952 791944 80008 792000
rect 79208 791820 79264 791876
rect 79332 791820 79388 791876
rect 79456 791820 79512 791876
rect 79580 791820 79636 791876
rect 79704 791820 79760 791876
rect 79828 791820 79884 791876
rect 79952 791820 80008 791876
rect 79208 791696 79264 791752
rect 79332 791696 79388 791752
rect 79456 791696 79512 791752
rect 79580 791696 79636 791752
rect 79704 791696 79760 791752
rect 79828 791696 79884 791752
rect 79952 791696 80008 791752
rect 79208 791572 79264 791628
rect 79332 791572 79388 791628
rect 79456 791572 79512 791628
rect 79580 791572 79636 791628
rect 79704 791572 79760 791628
rect 79828 791572 79884 791628
rect 79952 791572 80008 791628
rect 79208 791448 79264 791504
rect 79332 791448 79388 791504
rect 79456 791448 79512 791504
rect 79580 791448 79636 791504
rect 79704 791448 79760 791504
rect 79828 791448 79884 791504
rect 79952 791448 80008 791504
rect 79208 791324 79264 791380
rect 79332 791324 79388 791380
rect 79456 791324 79512 791380
rect 79580 791324 79636 791380
rect 79704 791324 79760 791380
rect 79828 791324 79884 791380
rect 79952 791324 80008 791380
rect 79208 791200 79264 791256
rect 79332 791200 79388 791256
rect 79456 791200 79512 791256
rect 79580 791200 79636 791256
rect 79704 791200 79760 791256
rect 79828 791200 79884 791256
rect 79952 791200 80008 791256
rect 79208 791076 79264 791132
rect 79332 791076 79388 791132
rect 79456 791076 79512 791132
rect 79580 791076 79636 791132
rect 79704 791076 79760 791132
rect 79828 791076 79884 791132
rect 79952 791076 80008 791132
rect 79208 790952 79264 791008
rect 79332 790952 79388 791008
rect 79456 790952 79512 791008
rect 79580 790952 79636 791008
rect 79704 790952 79760 791008
rect 79828 790952 79884 791008
rect 79952 790952 80008 791008
rect 79208 790828 79264 790884
rect 79332 790828 79388 790884
rect 79456 790828 79512 790884
rect 79580 790828 79636 790884
rect 79704 790828 79760 790884
rect 79828 790828 79884 790884
rect 79952 790828 80008 790884
rect 79208 790084 79264 790140
rect 79332 790084 79388 790140
rect 79456 790084 79512 790140
rect 79580 790084 79636 790140
rect 79704 790084 79760 790140
rect 79828 790084 79884 790140
rect 79952 790084 80008 790140
rect 79208 789960 79264 790016
rect 79332 789960 79388 790016
rect 79456 789960 79512 790016
rect 79580 789960 79636 790016
rect 79704 789960 79760 790016
rect 79828 789960 79884 790016
rect 79952 789960 80008 790016
rect 79208 789836 79264 789892
rect 79332 789836 79388 789892
rect 79456 789836 79512 789892
rect 79580 789836 79636 789892
rect 79704 789836 79760 789892
rect 79828 789836 79884 789892
rect 79952 789836 80008 789892
rect 79208 789712 79264 789768
rect 79332 789712 79388 789768
rect 79456 789712 79512 789768
rect 79580 789712 79636 789768
rect 79704 789712 79760 789768
rect 79828 789712 79884 789768
rect 79952 789712 80008 789768
rect 79208 789588 79264 789644
rect 79332 789588 79388 789644
rect 79456 789588 79512 789644
rect 79580 789588 79636 789644
rect 79704 789588 79760 789644
rect 79828 789588 79884 789644
rect 79952 789588 80008 789644
rect 79208 789464 79264 789520
rect 79332 789464 79388 789520
rect 79456 789464 79512 789520
rect 79580 789464 79636 789520
rect 79704 789464 79760 789520
rect 79828 789464 79884 789520
rect 79952 789464 80008 789520
rect 79208 789340 79264 789396
rect 79332 789340 79388 789396
rect 79456 789340 79512 789396
rect 79580 789340 79636 789396
rect 79704 789340 79760 789396
rect 79828 789340 79884 789396
rect 79952 789340 80008 789396
rect 79208 789216 79264 789272
rect 79332 789216 79388 789272
rect 79456 789216 79512 789272
rect 79580 789216 79636 789272
rect 79704 789216 79760 789272
rect 79828 789216 79884 789272
rect 79952 789216 80008 789272
rect 79208 789092 79264 789148
rect 79332 789092 79388 789148
rect 79456 789092 79512 789148
rect 79580 789092 79636 789148
rect 79704 789092 79760 789148
rect 79828 789092 79884 789148
rect 79952 789092 80008 789148
rect 79208 788968 79264 789024
rect 79332 788968 79388 789024
rect 79456 788968 79512 789024
rect 79580 788968 79636 789024
rect 79704 788968 79760 789024
rect 79828 788968 79884 789024
rect 79952 788968 80008 789024
rect 79208 788844 79264 788900
rect 79332 788844 79388 788900
rect 79456 788844 79512 788900
rect 79580 788844 79636 788900
rect 79704 788844 79760 788900
rect 79828 788844 79884 788900
rect 79952 788844 80008 788900
rect 79208 788720 79264 788776
rect 79332 788720 79388 788776
rect 79456 788720 79512 788776
rect 79580 788720 79636 788776
rect 79704 788720 79760 788776
rect 79828 788720 79884 788776
rect 79952 788720 80008 788776
rect 79208 788596 79264 788652
rect 79332 788596 79388 788652
rect 79456 788596 79512 788652
rect 79580 788596 79636 788652
rect 79704 788596 79760 788652
rect 79828 788596 79884 788652
rect 79952 788596 80008 788652
rect 79208 788472 79264 788528
rect 79332 788472 79388 788528
rect 79456 788472 79512 788528
rect 79580 788472 79636 788528
rect 79704 788472 79760 788528
rect 79828 788472 79884 788528
rect 79952 788472 80008 788528
rect 79208 788348 79264 788404
rect 79332 788348 79388 788404
rect 79456 788348 79512 788404
rect 79580 788348 79636 788404
rect 79704 788348 79760 788404
rect 79828 788348 79884 788404
rect 79952 788348 80008 788404
rect 79284 781992 79340 782048
rect 79584 781992 79640 782048
rect 79884 781992 79940 782048
rect 79300 765566 79356 765622
rect 79600 765566 79656 765622
rect 79900 765566 79956 765622
rect 79300 758566 79356 758622
rect 79600 758566 79656 758622
rect 79900 758566 79956 758622
rect 79200 752373 79256 752429
rect 79500 752373 79556 752429
rect 79800 752373 79856 752429
rect 79200 752173 79256 752229
rect 79500 752173 79556 752229
rect 79800 752173 79856 752229
rect 79300 751566 79356 751622
rect 79600 751566 79656 751622
rect 79900 751566 79956 751622
rect 79284 740992 79340 741048
rect 79584 740992 79640 741048
rect 79884 740992 79940 741048
rect 79300 724566 79356 724622
rect 79600 724566 79656 724622
rect 79900 724566 79956 724622
rect 79300 717566 79356 717622
rect 79600 717566 79656 717622
rect 79900 717566 79956 717622
rect 79200 716373 79256 716429
rect 79500 716373 79556 716429
rect 79800 716373 79856 716429
rect 79200 716173 79256 716229
rect 79500 716173 79556 716229
rect 79800 716173 79856 716229
rect 79300 710566 79356 710622
rect 79600 710566 79656 710622
rect 79900 710566 79956 710622
rect 79284 699992 79340 700048
rect 79584 699992 79640 700048
rect 79884 699992 79940 700048
rect 79300 683566 79356 683622
rect 79600 683566 79656 683622
rect 79900 683566 79956 683622
rect 79200 680373 79256 680429
rect 79500 680373 79556 680429
rect 79800 680373 79856 680429
rect 79200 680173 79256 680229
rect 79500 680173 79556 680229
rect 79800 680173 79856 680229
rect 79300 676566 79356 676622
rect 79600 676566 79656 676622
rect 79900 676566 79956 676622
rect 79300 669566 79356 669622
rect 79600 669566 79656 669622
rect 79900 669566 79956 669622
rect 79284 658992 79340 659048
rect 79584 658992 79640 659048
rect 79884 658992 79940 659048
rect 79200 644373 79256 644429
rect 79500 644373 79556 644429
rect 79800 644373 79856 644429
rect 79200 644173 79256 644229
rect 79500 644173 79556 644229
rect 79800 644173 79856 644229
rect 79300 642566 79356 642622
rect 79600 642566 79656 642622
rect 79900 642566 79956 642622
rect 79300 635566 79356 635622
rect 79600 635566 79656 635622
rect 79900 635566 79956 635622
rect 79300 628566 79356 628622
rect 79600 628566 79656 628622
rect 79900 628566 79956 628622
rect 79284 617992 79340 618048
rect 79584 617992 79640 618048
rect 79884 617992 79940 618048
rect 79200 608373 79256 608429
rect 79500 608373 79556 608429
rect 79800 608373 79856 608429
rect 79200 608173 79256 608229
rect 79500 608173 79556 608229
rect 79800 608173 79856 608229
rect 79300 601566 79356 601622
rect 79600 601566 79656 601622
rect 79900 601566 79956 601622
rect 79300 594566 79356 594622
rect 79600 594566 79656 594622
rect 79900 594566 79956 594622
rect 79300 587566 79356 587622
rect 79600 587566 79656 587622
rect 79900 587566 79956 587622
rect 79284 576992 79340 577048
rect 79584 576992 79640 577048
rect 79884 576992 79940 577048
rect 79200 572373 79256 572429
rect 79500 572373 79556 572429
rect 79800 572373 79856 572429
rect 79200 572173 79256 572229
rect 79500 572173 79556 572229
rect 79800 572173 79856 572229
rect 79300 560566 79356 560622
rect 79600 560566 79656 560622
rect 79900 560566 79956 560622
rect 79300 553566 79356 553622
rect 79600 553566 79656 553622
rect 79900 553566 79956 553622
rect 79300 546566 79356 546622
rect 79600 546566 79656 546622
rect 79900 546566 79956 546622
rect 79200 536373 79256 536429
rect 79500 536373 79556 536429
rect 79800 536373 79856 536429
rect 79200 536173 79256 536229
rect 79500 536173 79556 536229
rect 79800 536173 79856 536229
rect 79284 535992 79340 536048
rect 79584 535992 79640 536048
rect 79884 535992 79940 536048
rect 79300 519566 79356 519622
rect 79600 519566 79656 519622
rect 79900 519566 79956 519622
rect 79300 512566 79356 512622
rect 79600 512566 79656 512622
rect 79900 512566 79956 512622
rect 79300 505566 79356 505622
rect 79600 505566 79656 505622
rect 79900 505566 79956 505622
rect 79200 500373 79256 500429
rect 79500 500373 79556 500429
rect 79800 500373 79856 500429
rect 79200 500173 79256 500229
rect 79500 500173 79556 500229
rect 79800 500173 79856 500229
rect 79208 433614 79264 433670
rect 79332 433614 79388 433670
rect 79456 433614 79512 433670
rect 79580 433614 79636 433670
rect 79704 433614 79760 433670
rect 79828 433614 79884 433670
rect 79952 433614 80008 433670
rect 79208 433490 79264 433546
rect 79332 433490 79388 433546
rect 79456 433490 79512 433546
rect 79580 433490 79636 433546
rect 79704 433490 79760 433546
rect 79828 433490 79884 433546
rect 79952 433490 80008 433546
rect 79208 433366 79264 433422
rect 79332 433366 79388 433422
rect 79456 433366 79512 433422
rect 79580 433366 79636 433422
rect 79704 433366 79760 433422
rect 79828 433366 79884 433422
rect 79952 433366 80008 433422
rect 79208 433242 79264 433298
rect 79332 433242 79388 433298
rect 79456 433242 79512 433298
rect 79580 433242 79636 433298
rect 79704 433242 79760 433298
rect 79828 433242 79884 433298
rect 79952 433242 80008 433298
rect 79208 433118 79264 433174
rect 79332 433118 79388 433174
rect 79456 433118 79512 433174
rect 79580 433118 79636 433174
rect 79704 433118 79760 433174
rect 79828 433118 79884 433174
rect 79952 433118 80008 433174
rect 79208 432994 79264 433050
rect 79332 432994 79388 433050
rect 79456 432994 79512 433050
rect 79580 432994 79636 433050
rect 79704 432994 79760 433050
rect 79828 432994 79884 433050
rect 79952 432994 80008 433050
rect 79208 432870 79264 432926
rect 79332 432870 79388 432926
rect 79456 432870 79512 432926
rect 79580 432870 79636 432926
rect 79704 432870 79760 432926
rect 79828 432870 79884 432926
rect 79952 432870 80008 432926
rect 79208 432746 79264 432802
rect 79332 432746 79388 432802
rect 79456 432746 79512 432802
rect 79580 432746 79636 432802
rect 79704 432746 79760 432802
rect 79828 432746 79884 432802
rect 79952 432746 80008 432802
rect 79208 432622 79264 432678
rect 79332 432622 79388 432678
rect 79456 432622 79512 432678
rect 79580 432622 79636 432678
rect 79704 432622 79760 432678
rect 79828 432622 79884 432678
rect 79952 432622 80008 432678
rect 79208 432498 79264 432554
rect 79332 432498 79388 432554
rect 79456 432498 79512 432554
rect 79580 432498 79636 432554
rect 79704 432498 79760 432554
rect 79828 432498 79884 432554
rect 79952 432498 80008 432554
rect 79208 432374 79264 432430
rect 79332 432374 79388 432430
rect 79456 432374 79512 432430
rect 79580 432374 79636 432430
rect 79704 432374 79760 432430
rect 79828 432374 79884 432430
rect 79952 432374 80008 432430
rect 79208 432250 79264 432306
rect 79332 432250 79388 432306
rect 79456 432250 79512 432306
rect 79580 432250 79636 432306
rect 79704 432250 79760 432306
rect 79828 432250 79884 432306
rect 79952 432250 80008 432306
rect 79208 432126 79264 432182
rect 79332 432126 79388 432182
rect 79456 432126 79512 432182
rect 79580 432126 79636 432182
rect 79704 432126 79760 432182
rect 79828 432126 79884 432182
rect 79952 432126 80008 432182
rect 79208 432002 79264 432058
rect 79332 432002 79388 432058
rect 79456 432002 79512 432058
rect 79580 432002 79636 432058
rect 79704 432002 79760 432058
rect 79828 432002 79884 432058
rect 79952 432002 80008 432058
rect 79208 431878 79264 431934
rect 79332 431878 79388 431934
rect 79456 431878 79512 431934
rect 79580 431878 79636 431934
rect 79704 431878 79760 431934
rect 79828 431878 79884 431934
rect 79952 431878 80008 431934
rect 79208 431134 79264 431190
rect 79332 431134 79388 431190
rect 79456 431134 79512 431190
rect 79580 431134 79636 431190
rect 79704 431134 79760 431190
rect 79828 431134 79884 431190
rect 79952 431134 80008 431190
rect 79208 431010 79264 431066
rect 79332 431010 79388 431066
rect 79456 431010 79512 431066
rect 79580 431010 79636 431066
rect 79704 431010 79760 431066
rect 79828 431010 79884 431066
rect 79952 431010 80008 431066
rect 79208 430886 79264 430942
rect 79332 430886 79388 430942
rect 79456 430886 79512 430942
rect 79580 430886 79636 430942
rect 79704 430886 79760 430942
rect 79828 430886 79884 430942
rect 79952 430886 80008 430942
rect 79208 430762 79264 430818
rect 79332 430762 79388 430818
rect 79456 430762 79512 430818
rect 79580 430762 79636 430818
rect 79704 430762 79760 430818
rect 79828 430762 79884 430818
rect 79952 430762 80008 430818
rect 79208 430638 79264 430694
rect 79332 430638 79388 430694
rect 79456 430638 79512 430694
rect 79580 430638 79636 430694
rect 79704 430638 79760 430694
rect 79828 430638 79884 430694
rect 79952 430638 80008 430694
rect 79208 430514 79264 430570
rect 79332 430514 79388 430570
rect 79456 430514 79512 430570
rect 79580 430514 79636 430570
rect 79704 430514 79760 430570
rect 79828 430514 79884 430570
rect 79952 430514 80008 430570
rect 79208 430390 79264 430446
rect 79332 430390 79388 430446
rect 79456 430390 79512 430446
rect 79580 430390 79636 430446
rect 79704 430390 79760 430446
rect 79828 430390 79884 430446
rect 79952 430390 80008 430446
rect 79208 430266 79264 430322
rect 79332 430266 79388 430322
rect 79456 430266 79512 430322
rect 79580 430266 79636 430322
rect 79704 430266 79760 430322
rect 79828 430266 79884 430322
rect 79952 430266 80008 430322
rect 79208 430142 79264 430198
rect 79332 430142 79388 430198
rect 79456 430142 79512 430198
rect 79580 430142 79636 430198
rect 79704 430142 79760 430198
rect 79828 430142 79884 430198
rect 79952 430142 80008 430198
rect 79208 430018 79264 430074
rect 79332 430018 79388 430074
rect 79456 430018 79512 430074
rect 79580 430018 79636 430074
rect 79704 430018 79760 430074
rect 79828 430018 79884 430074
rect 79952 430018 80008 430074
rect 79208 429894 79264 429950
rect 79332 429894 79388 429950
rect 79456 429894 79512 429950
rect 79580 429894 79636 429950
rect 79704 429894 79760 429950
rect 79828 429894 79884 429950
rect 79952 429894 80008 429950
rect 79208 429770 79264 429826
rect 79332 429770 79388 429826
rect 79456 429770 79512 429826
rect 79580 429770 79636 429826
rect 79704 429770 79760 429826
rect 79828 429770 79884 429826
rect 79952 429770 80008 429826
rect 79208 429646 79264 429702
rect 79332 429646 79388 429702
rect 79456 429646 79512 429702
rect 79580 429646 79636 429702
rect 79704 429646 79760 429702
rect 79828 429646 79884 429702
rect 79952 429646 80008 429702
rect 79208 429522 79264 429578
rect 79332 429522 79388 429578
rect 79456 429522 79512 429578
rect 79580 429522 79636 429578
rect 79704 429522 79760 429578
rect 79828 429522 79884 429578
rect 79952 429522 80008 429578
rect 79208 429398 79264 429454
rect 79332 429398 79388 429454
rect 79456 429398 79512 429454
rect 79580 429398 79636 429454
rect 79704 429398 79760 429454
rect 79828 429398 79884 429454
rect 79952 429398 80008 429454
rect 79208 429274 79264 429330
rect 79332 429274 79388 429330
rect 79456 429274 79512 429330
rect 79580 429274 79636 429330
rect 79704 429274 79760 429330
rect 79828 429274 79884 429330
rect 79952 429274 80008 429330
rect 79208 428764 79264 428820
rect 79332 428764 79388 428820
rect 79456 428764 79512 428820
rect 79580 428764 79636 428820
rect 79704 428764 79760 428820
rect 79828 428764 79884 428820
rect 79952 428764 80008 428820
rect 79208 428640 79264 428696
rect 79332 428640 79388 428696
rect 79456 428640 79512 428696
rect 79580 428640 79636 428696
rect 79704 428640 79760 428696
rect 79828 428640 79884 428696
rect 79952 428640 80008 428696
rect 79208 428516 79264 428572
rect 79332 428516 79388 428572
rect 79456 428516 79512 428572
rect 79580 428516 79636 428572
rect 79704 428516 79760 428572
rect 79828 428516 79884 428572
rect 79952 428516 80008 428572
rect 79208 428392 79264 428448
rect 79332 428392 79388 428448
rect 79456 428392 79512 428448
rect 79580 428392 79636 428448
rect 79704 428392 79760 428448
rect 79828 428392 79884 428448
rect 79952 428392 80008 428448
rect 79208 428268 79264 428324
rect 79332 428268 79388 428324
rect 79456 428268 79512 428324
rect 79580 428268 79636 428324
rect 79704 428268 79760 428324
rect 79828 428268 79884 428324
rect 79952 428268 80008 428324
rect 79208 428144 79264 428200
rect 79332 428144 79388 428200
rect 79456 428144 79512 428200
rect 79580 428144 79636 428200
rect 79704 428144 79760 428200
rect 79828 428144 79884 428200
rect 79952 428144 80008 428200
rect 79208 428020 79264 428076
rect 79332 428020 79388 428076
rect 79456 428020 79512 428076
rect 79580 428020 79636 428076
rect 79704 428020 79760 428076
rect 79828 428020 79884 428076
rect 79952 428020 80008 428076
rect 79208 427896 79264 427952
rect 79332 427896 79388 427952
rect 79456 427896 79512 427952
rect 79580 427896 79636 427952
rect 79704 427896 79760 427952
rect 79828 427896 79884 427952
rect 79952 427896 80008 427952
rect 79208 427772 79264 427828
rect 79332 427772 79388 427828
rect 79456 427772 79512 427828
rect 79580 427772 79636 427828
rect 79704 427772 79760 427828
rect 79828 427772 79884 427828
rect 79952 427772 80008 427828
rect 79208 427648 79264 427704
rect 79332 427648 79388 427704
rect 79456 427648 79512 427704
rect 79580 427648 79636 427704
rect 79704 427648 79760 427704
rect 79828 427648 79884 427704
rect 79952 427648 80008 427704
rect 79208 427524 79264 427580
rect 79332 427524 79388 427580
rect 79456 427524 79512 427580
rect 79580 427524 79636 427580
rect 79704 427524 79760 427580
rect 79828 427524 79884 427580
rect 79952 427524 80008 427580
rect 79208 427400 79264 427456
rect 79332 427400 79388 427456
rect 79456 427400 79512 427456
rect 79580 427400 79636 427456
rect 79704 427400 79760 427456
rect 79828 427400 79884 427456
rect 79952 427400 80008 427456
rect 79208 427276 79264 427332
rect 79332 427276 79388 427332
rect 79456 427276 79512 427332
rect 79580 427276 79636 427332
rect 79704 427276 79760 427332
rect 79828 427276 79884 427332
rect 79952 427276 80008 427332
rect 79208 427152 79264 427208
rect 79332 427152 79388 427208
rect 79456 427152 79512 427208
rect 79580 427152 79636 427208
rect 79704 427152 79760 427208
rect 79828 427152 79884 427208
rect 79952 427152 80008 427208
rect 79208 427028 79264 427084
rect 79332 427028 79388 427084
rect 79456 427028 79512 427084
rect 79580 427028 79636 427084
rect 79704 427028 79760 427084
rect 79828 427028 79884 427084
rect 79952 427028 80008 427084
rect 79208 426904 79264 426960
rect 79332 426904 79388 426960
rect 79456 426904 79512 426960
rect 79580 426904 79636 426960
rect 79704 426904 79760 426960
rect 79828 426904 79884 426960
rect 79952 426904 80008 426960
rect 79208 426058 79264 426114
rect 79332 426058 79388 426114
rect 79456 426058 79512 426114
rect 79580 426058 79636 426114
rect 79704 426058 79760 426114
rect 79828 426058 79884 426114
rect 79952 426058 80008 426114
rect 79208 425934 79264 425990
rect 79332 425934 79388 425990
rect 79456 425934 79512 425990
rect 79580 425934 79636 425990
rect 79704 425934 79760 425990
rect 79828 425934 79884 425990
rect 79952 425934 80008 425990
rect 79208 425810 79264 425866
rect 79332 425810 79388 425866
rect 79456 425810 79512 425866
rect 79580 425810 79636 425866
rect 79704 425810 79760 425866
rect 79828 425810 79884 425866
rect 79952 425810 80008 425866
rect 79208 425686 79264 425742
rect 79332 425686 79388 425742
rect 79456 425686 79512 425742
rect 79580 425686 79636 425742
rect 79704 425686 79760 425742
rect 79828 425686 79884 425742
rect 79952 425686 80008 425742
rect 79208 425562 79264 425618
rect 79332 425562 79388 425618
rect 79456 425562 79512 425618
rect 79580 425562 79636 425618
rect 79704 425562 79760 425618
rect 79828 425562 79884 425618
rect 79952 425562 80008 425618
rect 79208 425438 79264 425494
rect 79332 425438 79388 425494
rect 79456 425438 79512 425494
rect 79580 425438 79636 425494
rect 79704 425438 79760 425494
rect 79828 425438 79884 425494
rect 79952 425438 80008 425494
rect 79208 425314 79264 425370
rect 79332 425314 79388 425370
rect 79456 425314 79512 425370
rect 79580 425314 79636 425370
rect 79704 425314 79760 425370
rect 79828 425314 79884 425370
rect 79952 425314 80008 425370
rect 79208 425190 79264 425246
rect 79332 425190 79388 425246
rect 79456 425190 79512 425246
rect 79580 425190 79636 425246
rect 79704 425190 79760 425246
rect 79828 425190 79884 425246
rect 79952 425190 80008 425246
rect 79208 425066 79264 425122
rect 79332 425066 79388 425122
rect 79456 425066 79512 425122
rect 79580 425066 79636 425122
rect 79704 425066 79760 425122
rect 79828 425066 79884 425122
rect 79952 425066 80008 425122
rect 79208 424942 79264 424998
rect 79332 424942 79388 424998
rect 79456 424942 79512 424998
rect 79580 424942 79636 424998
rect 79704 424942 79760 424998
rect 79828 424942 79884 424998
rect 79952 424942 80008 424998
rect 79208 424818 79264 424874
rect 79332 424818 79388 424874
rect 79456 424818 79512 424874
rect 79580 424818 79636 424874
rect 79704 424818 79760 424874
rect 79828 424818 79884 424874
rect 79952 424818 80008 424874
rect 79208 424694 79264 424750
rect 79332 424694 79388 424750
rect 79456 424694 79512 424750
rect 79580 424694 79636 424750
rect 79704 424694 79760 424750
rect 79828 424694 79884 424750
rect 79952 424694 80008 424750
rect 79208 424570 79264 424626
rect 79332 424570 79388 424626
rect 79456 424570 79512 424626
rect 79580 424570 79636 424626
rect 79704 424570 79760 424626
rect 79828 424570 79884 424626
rect 79952 424570 80008 424626
rect 79208 424446 79264 424502
rect 79332 424446 79388 424502
rect 79456 424446 79512 424502
rect 79580 424446 79636 424502
rect 79704 424446 79760 424502
rect 79828 424446 79884 424502
rect 79952 424446 80008 424502
rect 79208 424322 79264 424378
rect 79332 424322 79388 424378
rect 79456 424322 79512 424378
rect 79580 424322 79636 424378
rect 79704 424322 79760 424378
rect 79828 424322 79884 424378
rect 79952 424322 80008 424378
rect 79208 424198 79264 424254
rect 79332 424198 79388 424254
rect 79456 424198 79512 424254
rect 79580 424198 79636 424254
rect 79704 424198 79760 424254
rect 79828 424198 79884 424254
rect 79952 424198 80008 424254
rect 79208 423688 79264 423744
rect 79332 423688 79388 423744
rect 79456 423688 79512 423744
rect 79580 423688 79636 423744
rect 79704 423688 79760 423744
rect 79828 423688 79884 423744
rect 79952 423688 80008 423744
rect 79208 423564 79264 423620
rect 79332 423564 79388 423620
rect 79456 423564 79512 423620
rect 79580 423564 79636 423620
rect 79704 423564 79760 423620
rect 79828 423564 79884 423620
rect 79952 423564 80008 423620
rect 79208 423440 79264 423496
rect 79332 423440 79388 423496
rect 79456 423440 79512 423496
rect 79580 423440 79636 423496
rect 79704 423440 79760 423496
rect 79828 423440 79884 423496
rect 79952 423440 80008 423496
rect 79208 423316 79264 423372
rect 79332 423316 79388 423372
rect 79456 423316 79512 423372
rect 79580 423316 79636 423372
rect 79704 423316 79760 423372
rect 79828 423316 79884 423372
rect 79952 423316 80008 423372
rect 79208 423192 79264 423248
rect 79332 423192 79388 423248
rect 79456 423192 79512 423248
rect 79580 423192 79636 423248
rect 79704 423192 79760 423248
rect 79828 423192 79884 423248
rect 79952 423192 80008 423248
rect 79208 423068 79264 423124
rect 79332 423068 79388 423124
rect 79456 423068 79512 423124
rect 79580 423068 79636 423124
rect 79704 423068 79760 423124
rect 79828 423068 79884 423124
rect 79952 423068 80008 423124
rect 79208 422944 79264 423000
rect 79332 422944 79388 423000
rect 79456 422944 79512 423000
rect 79580 422944 79636 423000
rect 79704 422944 79760 423000
rect 79828 422944 79884 423000
rect 79952 422944 80008 423000
rect 79208 422820 79264 422876
rect 79332 422820 79388 422876
rect 79456 422820 79512 422876
rect 79580 422820 79636 422876
rect 79704 422820 79760 422876
rect 79828 422820 79884 422876
rect 79952 422820 80008 422876
rect 79208 422696 79264 422752
rect 79332 422696 79388 422752
rect 79456 422696 79512 422752
rect 79580 422696 79636 422752
rect 79704 422696 79760 422752
rect 79828 422696 79884 422752
rect 79952 422696 80008 422752
rect 79208 422572 79264 422628
rect 79332 422572 79388 422628
rect 79456 422572 79512 422628
rect 79580 422572 79636 422628
rect 79704 422572 79760 422628
rect 79828 422572 79884 422628
rect 79952 422572 80008 422628
rect 79208 422448 79264 422504
rect 79332 422448 79388 422504
rect 79456 422448 79512 422504
rect 79580 422448 79636 422504
rect 79704 422448 79760 422504
rect 79828 422448 79884 422504
rect 79952 422448 80008 422504
rect 79208 422324 79264 422380
rect 79332 422324 79388 422380
rect 79456 422324 79512 422380
rect 79580 422324 79636 422380
rect 79704 422324 79760 422380
rect 79828 422324 79884 422380
rect 79952 422324 80008 422380
rect 79208 422200 79264 422256
rect 79332 422200 79388 422256
rect 79456 422200 79512 422256
rect 79580 422200 79636 422256
rect 79704 422200 79760 422256
rect 79828 422200 79884 422256
rect 79952 422200 80008 422256
rect 79208 422076 79264 422132
rect 79332 422076 79388 422132
rect 79456 422076 79512 422132
rect 79580 422076 79636 422132
rect 79704 422076 79760 422132
rect 79828 422076 79884 422132
rect 79952 422076 80008 422132
rect 79208 421952 79264 422008
rect 79332 421952 79388 422008
rect 79456 421952 79512 422008
rect 79580 421952 79636 422008
rect 79704 421952 79760 422008
rect 79828 421952 79884 422008
rect 79952 421952 80008 422008
rect 79208 421828 79264 421884
rect 79332 421828 79388 421884
rect 79456 421828 79512 421884
rect 79580 421828 79636 421884
rect 79704 421828 79760 421884
rect 79828 421828 79884 421884
rect 79952 421828 80008 421884
rect 79208 421084 79264 421140
rect 79332 421084 79388 421140
rect 79456 421084 79512 421140
rect 79580 421084 79636 421140
rect 79704 421084 79760 421140
rect 79828 421084 79884 421140
rect 79952 421084 80008 421140
rect 79208 420960 79264 421016
rect 79332 420960 79388 421016
rect 79456 420960 79512 421016
rect 79580 420960 79636 421016
rect 79704 420960 79760 421016
rect 79828 420960 79884 421016
rect 79952 420960 80008 421016
rect 79208 420836 79264 420892
rect 79332 420836 79388 420892
rect 79456 420836 79512 420892
rect 79580 420836 79636 420892
rect 79704 420836 79760 420892
rect 79828 420836 79884 420892
rect 79952 420836 80008 420892
rect 79208 420712 79264 420768
rect 79332 420712 79388 420768
rect 79456 420712 79512 420768
rect 79580 420712 79636 420768
rect 79704 420712 79760 420768
rect 79828 420712 79884 420768
rect 79952 420712 80008 420768
rect 79208 420588 79264 420644
rect 79332 420588 79388 420644
rect 79456 420588 79512 420644
rect 79580 420588 79636 420644
rect 79704 420588 79760 420644
rect 79828 420588 79884 420644
rect 79952 420588 80008 420644
rect 79208 420464 79264 420520
rect 79332 420464 79388 420520
rect 79456 420464 79512 420520
rect 79580 420464 79636 420520
rect 79704 420464 79760 420520
rect 79828 420464 79884 420520
rect 79952 420464 80008 420520
rect 79208 420340 79264 420396
rect 79332 420340 79388 420396
rect 79456 420340 79512 420396
rect 79580 420340 79636 420396
rect 79704 420340 79760 420396
rect 79828 420340 79884 420396
rect 79952 420340 80008 420396
rect 79208 420216 79264 420272
rect 79332 420216 79388 420272
rect 79456 420216 79512 420272
rect 79580 420216 79636 420272
rect 79704 420216 79760 420272
rect 79828 420216 79884 420272
rect 79952 420216 80008 420272
rect 79208 420092 79264 420148
rect 79332 420092 79388 420148
rect 79456 420092 79512 420148
rect 79580 420092 79636 420148
rect 79704 420092 79760 420148
rect 79828 420092 79884 420148
rect 79952 420092 80008 420148
rect 79208 419968 79264 420024
rect 79332 419968 79388 420024
rect 79456 419968 79512 420024
rect 79580 419968 79636 420024
rect 79704 419968 79760 420024
rect 79828 419968 79884 420024
rect 79952 419968 80008 420024
rect 79208 419844 79264 419900
rect 79332 419844 79388 419900
rect 79456 419844 79512 419900
rect 79580 419844 79636 419900
rect 79704 419844 79760 419900
rect 79828 419844 79884 419900
rect 79952 419844 80008 419900
rect 79208 419720 79264 419776
rect 79332 419720 79388 419776
rect 79456 419720 79512 419776
rect 79580 419720 79636 419776
rect 79704 419720 79760 419776
rect 79828 419720 79884 419776
rect 79952 419720 80008 419776
rect 79208 419596 79264 419652
rect 79332 419596 79388 419652
rect 79456 419596 79512 419652
rect 79580 419596 79636 419652
rect 79704 419596 79760 419652
rect 79828 419596 79884 419652
rect 79952 419596 80008 419652
rect 79208 419472 79264 419528
rect 79332 419472 79388 419528
rect 79456 419472 79512 419528
rect 79580 419472 79636 419528
rect 79704 419472 79760 419528
rect 79828 419472 79884 419528
rect 79952 419472 80008 419528
rect 79208 419348 79264 419404
rect 79332 419348 79388 419404
rect 79456 419348 79512 419404
rect 79580 419348 79636 419404
rect 79704 419348 79760 419404
rect 79828 419348 79884 419404
rect 79952 419348 80008 419404
rect 79284 412992 79340 413048
rect 79584 412992 79640 413048
rect 79884 412992 79940 413048
rect 79300 396566 79356 396622
rect 79600 396566 79656 396622
rect 79900 396566 79956 396622
rect 79200 392373 79256 392429
rect 79500 392373 79556 392429
rect 79800 392373 79856 392429
rect 79200 392173 79256 392229
rect 79500 392173 79556 392229
rect 79800 392173 79856 392229
rect 79300 389566 79356 389622
rect 79600 389566 79656 389622
rect 79900 389566 79956 389622
rect 79300 382566 79356 382622
rect 79600 382566 79656 382622
rect 79900 382566 79956 382622
rect 79284 371992 79340 372048
rect 79584 371992 79640 372048
rect 79884 371992 79940 372048
rect 79200 356373 79256 356429
rect 79500 356373 79556 356429
rect 79800 356373 79856 356429
rect 79200 356173 79256 356229
rect 79500 356173 79556 356229
rect 79800 356173 79856 356229
rect 79300 355566 79356 355622
rect 79600 355566 79656 355622
rect 79900 355566 79956 355622
rect 79300 348566 79356 348622
rect 79600 348566 79656 348622
rect 79900 348566 79956 348622
rect 79300 341566 79356 341622
rect 79600 341566 79656 341622
rect 79900 341566 79956 341622
rect 698044 922378 698100 922434
rect 698344 922378 698400 922434
rect 698644 922378 698700 922434
rect 698044 915378 698100 915434
rect 698344 915378 698400 915434
rect 698644 915378 698700 915434
rect 698044 908378 698100 908434
rect 698344 908378 698400 908434
rect 698644 908378 698700 908434
rect 698144 896373 698200 896429
rect 698444 896373 698500 896429
rect 698744 896373 698800 896429
rect 698144 896173 698200 896229
rect 698444 896173 698500 896229
rect 698744 896173 698800 896229
rect 698060 891952 698116 892008
rect 698360 891952 698416 892008
rect 698660 891952 698716 892008
rect 698144 860373 698200 860429
rect 698444 860373 698500 860429
rect 698744 860373 698800 860429
rect 698144 860173 698200 860229
rect 698444 860173 698500 860229
rect 698744 860173 698800 860229
rect 698044 836378 698100 836434
rect 698344 836378 698400 836434
rect 698644 836378 698700 836434
rect 698044 829378 698100 829434
rect 698344 829378 698400 829434
rect 698644 829378 698700 829434
rect 698144 824373 698200 824429
rect 698444 824373 698500 824429
rect 698744 824373 698800 824429
rect 698144 824173 698200 824229
rect 698444 824173 698500 824229
rect 698744 824173 698800 824229
rect 698044 822378 698100 822434
rect 698344 822378 698400 822434
rect 698644 822378 698700 822434
rect 698060 805952 698116 806008
rect 698360 805952 698416 806008
rect 698660 805952 698716 806008
rect 698144 752373 698200 752429
rect 698444 752373 698500 752429
rect 698744 752373 698800 752429
rect 698144 752173 698200 752229
rect 698444 752173 698500 752229
rect 698744 752173 698800 752229
rect 698044 750378 698100 750434
rect 698344 750378 698400 750434
rect 698644 750378 698700 750434
rect 698044 743378 698100 743434
rect 698344 743378 698400 743434
rect 698644 743378 698700 743434
rect 698044 736378 698100 736434
rect 698344 736378 698400 736434
rect 698644 736378 698700 736434
rect 698060 719952 698116 720008
rect 698360 719952 698416 720008
rect 698660 719952 698716 720008
rect 698144 716373 698200 716429
rect 698444 716373 698500 716429
rect 698744 716373 698800 716429
rect 698144 716173 698200 716229
rect 698444 716173 698500 716229
rect 698744 716173 698800 716229
rect 698044 707378 698100 707434
rect 698344 707378 698400 707434
rect 698644 707378 698700 707434
rect 698044 700378 698100 700434
rect 698344 700378 698400 700434
rect 698644 700378 698700 700434
rect 698044 693378 698100 693434
rect 698344 693378 698400 693434
rect 698644 693378 698700 693434
rect 698144 680373 698200 680429
rect 698444 680373 698500 680429
rect 698744 680373 698800 680429
rect 698144 680173 698200 680229
rect 698444 680173 698500 680229
rect 698744 680173 698800 680229
rect 698060 676952 698116 677008
rect 698360 676952 698416 677008
rect 698660 676952 698716 677008
rect 698044 664378 698100 664434
rect 698344 664378 698400 664434
rect 698644 664378 698700 664434
rect 698044 657378 698100 657434
rect 698344 657378 698400 657434
rect 698644 657378 698700 657434
rect 698044 650378 698100 650434
rect 698344 650378 698400 650434
rect 698644 650378 698700 650434
rect 698144 644373 698200 644429
rect 698444 644373 698500 644429
rect 698744 644373 698800 644429
rect 698144 644173 698200 644229
rect 698444 644173 698500 644229
rect 698744 644173 698800 644229
rect 698060 633952 698116 634008
rect 698360 633952 698416 634008
rect 698660 633952 698716 634008
rect 698044 621378 698100 621434
rect 698344 621378 698400 621434
rect 698644 621378 698700 621434
rect 698044 614378 698100 614434
rect 698344 614378 698400 614434
rect 698644 614378 698700 614434
rect 698144 608373 698200 608429
rect 698444 608373 698500 608429
rect 698744 608373 698800 608429
rect 698144 608173 698200 608229
rect 698444 608173 698500 608229
rect 698744 608173 698800 608229
rect 698044 607378 698100 607434
rect 698344 607378 698400 607434
rect 698644 607378 698700 607434
rect 698060 590952 698116 591008
rect 698360 590952 698416 591008
rect 698660 590952 698716 591008
rect 698044 578378 698100 578434
rect 698344 578378 698400 578434
rect 698644 578378 698700 578434
rect 698144 572373 698200 572429
rect 698444 572373 698500 572429
rect 698744 572373 698800 572429
rect 698144 572173 698200 572229
rect 698444 572173 698500 572229
rect 698744 572173 698800 572229
rect 698044 571378 698100 571434
rect 698344 571378 698400 571434
rect 698644 571378 698700 571434
rect 698044 564378 698100 564434
rect 698344 564378 698400 564434
rect 698644 564378 698700 564434
rect 698060 547952 698116 548008
rect 698360 547952 698416 548008
rect 698660 547952 698716 548008
rect 698144 536373 698200 536429
rect 698444 536373 698500 536429
rect 698744 536373 698800 536429
rect 698144 536173 698200 536229
rect 698444 536173 698500 536229
rect 698744 536173 698800 536229
rect 698044 535378 698100 535434
rect 698344 535378 698400 535434
rect 698644 535378 698700 535434
rect 698044 528378 698100 528434
rect 698344 528378 698400 528434
rect 698644 528378 698700 528434
rect 698044 521378 698100 521434
rect 698344 521378 698400 521434
rect 698644 521378 698700 521434
rect 698060 504952 698116 505008
rect 698360 504952 698416 505008
rect 698660 504952 698716 505008
rect 698144 500373 698200 500429
rect 698444 500373 698500 500429
rect 698744 500373 698800 500429
rect 698144 500173 698200 500229
rect 698444 500173 698500 500229
rect 698744 500173 698800 500229
rect 698144 464373 698200 464429
rect 698444 464373 698500 464429
rect 698744 464373 698800 464429
rect 698144 464173 698200 464229
rect 698444 464173 698500 464229
rect 698744 464173 698800 464229
rect 697992 453596 698048 453652
rect 698116 453596 698172 453652
rect 698240 453596 698296 453652
rect 698364 453596 698420 453652
rect 698488 453596 698544 453652
rect 698612 453596 698668 453652
rect 698736 453596 698792 453652
rect 697992 453472 698048 453528
rect 698116 453472 698172 453528
rect 698240 453472 698296 453528
rect 698364 453472 698420 453528
rect 698488 453472 698544 453528
rect 698612 453472 698668 453528
rect 698736 453472 698792 453528
rect 697992 453348 698048 453404
rect 698116 453348 698172 453404
rect 698240 453348 698296 453404
rect 698364 453348 698420 453404
rect 698488 453348 698544 453404
rect 698612 453348 698668 453404
rect 698736 453348 698792 453404
rect 697992 453224 698048 453280
rect 698116 453224 698172 453280
rect 698240 453224 698296 453280
rect 698364 453224 698420 453280
rect 698488 453224 698544 453280
rect 698612 453224 698668 453280
rect 698736 453224 698792 453280
rect 697992 453100 698048 453156
rect 698116 453100 698172 453156
rect 698240 453100 698296 453156
rect 698364 453100 698420 453156
rect 698488 453100 698544 453156
rect 698612 453100 698668 453156
rect 698736 453100 698792 453156
rect 697992 452976 698048 453032
rect 698116 452976 698172 453032
rect 698240 452976 698296 453032
rect 698364 452976 698420 453032
rect 698488 452976 698544 453032
rect 698612 452976 698668 453032
rect 698736 452976 698792 453032
rect 697992 452852 698048 452908
rect 698116 452852 698172 452908
rect 698240 452852 698296 452908
rect 698364 452852 698420 452908
rect 698488 452852 698544 452908
rect 698612 452852 698668 452908
rect 698736 452852 698792 452908
rect 697992 452728 698048 452784
rect 698116 452728 698172 452784
rect 698240 452728 698296 452784
rect 698364 452728 698420 452784
rect 698488 452728 698544 452784
rect 698612 452728 698668 452784
rect 698736 452728 698792 452784
rect 697992 452604 698048 452660
rect 698116 452604 698172 452660
rect 698240 452604 698296 452660
rect 698364 452604 698420 452660
rect 698488 452604 698544 452660
rect 698612 452604 698668 452660
rect 698736 452604 698792 452660
rect 697992 452480 698048 452536
rect 698116 452480 698172 452536
rect 698240 452480 698296 452536
rect 698364 452480 698420 452536
rect 698488 452480 698544 452536
rect 698612 452480 698668 452536
rect 698736 452480 698792 452536
rect 697992 452356 698048 452412
rect 698116 452356 698172 452412
rect 698240 452356 698296 452412
rect 698364 452356 698420 452412
rect 698488 452356 698544 452412
rect 698612 452356 698668 452412
rect 698736 452356 698792 452412
rect 697992 452232 698048 452288
rect 698116 452232 698172 452288
rect 698240 452232 698296 452288
rect 698364 452232 698420 452288
rect 698488 452232 698544 452288
rect 698612 452232 698668 452288
rect 698736 452232 698792 452288
rect 697992 452108 698048 452164
rect 698116 452108 698172 452164
rect 698240 452108 698296 452164
rect 698364 452108 698420 452164
rect 698488 452108 698544 452164
rect 698612 452108 698668 452164
rect 698736 452108 698792 452164
rect 697992 451984 698048 452040
rect 698116 451984 698172 452040
rect 698240 451984 698296 452040
rect 698364 451984 698420 452040
rect 698488 451984 698544 452040
rect 698612 451984 698668 452040
rect 698736 451984 698792 452040
rect 697992 451860 698048 451916
rect 698116 451860 698172 451916
rect 698240 451860 698296 451916
rect 698364 451860 698420 451916
rect 698488 451860 698544 451916
rect 698612 451860 698668 451916
rect 698736 451860 698792 451916
rect 697992 451116 698048 451172
rect 698116 451116 698172 451172
rect 698240 451116 698296 451172
rect 698364 451116 698420 451172
rect 698488 451116 698544 451172
rect 698612 451116 698668 451172
rect 698736 451116 698792 451172
rect 697992 450992 698048 451048
rect 698116 450992 698172 451048
rect 698240 450992 698296 451048
rect 698364 450992 698420 451048
rect 698488 450992 698544 451048
rect 698612 450992 698668 451048
rect 698736 450992 698792 451048
rect 697992 450868 698048 450924
rect 698116 450868 698172 450924
rect 698240 450868 698296 450924
rect 698364 450868 698420 450924
rect 698488 450868 698544 450924
rect 698612 450868 698668 450924
rect 698736 450868 698792 450924
rect 697992 450744 698048 450800
rect 698116 450744 698172 450800
rect 698240 450744 698296 450800
rect 698364 450744 698420 450800
rect 698488 450744 698544 450800
rect 698612 450744 698668 450800
rect 698736 450744 698792 450800
rect 697992 450620 698048 450676
rect 698116 450620 698172 450676
rect 698240 450620 698296 450676
rect 698364 450620 698420 450676
rect 698488 450620 698544 450676
rect 698612 450620 698668 450676
rect 698736 450620 698792 450676
rect 697992 450496 698048 450552
rect 698116 450496 698172 450552
rect 698240 450496 698296 450552
rect 698364 450496 698420 450552
rect 698488 450496 698544 450552
rect 698612 450496 698668 450552
rect 698736 450496 698792 450552
rect 697992 450372 698048 450428
rect 698116 450372 698172 450428
rect 698240 450372 698296 450428
rect 698364 450372 698420 450428
rect 698488 450372 698544 450428
rect 698612 450372 698668 450428
rect 698736 450372 698792 450428
rect 697992 450248 698048 450304
rect 698116 450248 698172 450304
rect 698240 450248 698296 450304
rect 698364 450248 698420 450304
rect 698488 450248 698544 450304
rect 698612 450248 698668 450304
rect 698736 450248 698792 450304
rect 697992 450124 698048 450180
rect 698116 450124 698172 450180
rect 698240 450124 698296 450180
rect 698364 450124 698420 450180
rect 698488 450124 698544 450180
rect 698612 450124 698668 450180
rect 698736 450124 698792 450180
rect 697992 450000 698048 450056
rect 698116 450000 698172 450056
rect 698240 450000 698296 450056
rect 698364 450000 698420 450056
rect 698488 450000 698544 450056
rect 698612 450000 698668 450056
rect 698736 450000 698792 450056
rect 697992 449876 698048 449932
rect 698116 449876 698172 449932
rect 698240 449876 698296 449932
rect 698364 449876 698420 449932
rect 698488 449876 698544 449932
rect 698612 449876 698668 449932
rect 698736 449876 698792 449932
rect 697992 449752 698048 449808
rect 698116 449752 698172 449808
rect 698240 449752 698296 449808
rect 698364 449752 698420 449808
rect 698488 449752 698544 449808
rect 698612 449752 698668 449808
rect 698736 449752 698792 449808
rect 697992 449628 698048 449684
rect 698116 449628 698172 449684
rect 698240 449628 698296 449684
rect 698364 449628 698420 449684
rect 698488 449628 698544 449684
rect 698612 449628 698668 449684
rect 698736 449628 698792 449684
rect 697992 449504 698048 449560
rect 698116 449504 698172 449560
rect 698240 449504 698296 449560
rect 698364 449504 698420 449560
rect 698488 449504 698544 449560
rect 698612 449504 698668 449560
rect 698736 449504 698792 449560
rect 697992 449380 698048 449436
rect 698116 449380 698172 449436
rect 698240 449380 698296 449436
rect 698364 449380 698420 449436
rect 698488 449380 698544 449436
rect 698612 449380 698668 449436
rect 698736 449380 698792 449436
rect 697992 449256 698048 449312
rect 698116 449256 698172 449312
rect 698240 449256 698296 449312
rect 698364 449256 698420 449312
rect 698488 449256 698544 449312
rect 698612 449256 698668 449312
rect 698736 449256 698792 449312
rect 697992 448746 698048 448802
rect 698116 448746 698172 448802
rect 698240 448746 698296 448802
rect 698364 448746 698420 448802
rect 698488 448746 698544 448802
rect 698612 448746 698668 448802
rect 698736 448746 698792 448802
rect 697992 448622 698048 448678
rect 698116 448622 698172 448678
rect 698240 448622 698296 448678
rect 698364 448622 698420 448678
rect 698488 448622 698544 448678
rect 698612 448622 698668 448678
rect 698736 448622 698792 448678
rect 697992 448498 698048 448554
rect 698116 448498 698172 448554
rect 698240 448498 698296 448554
rect 698364 448498 698420 448554
rect 698488 448498 698544 448554
rect 698612 448498 698668 448554
rect 698736 448498 698792 448554
rect 697992 448374 698048 448430
rect 698116 448374 698172 448430
rect 698240 448374 698296 448430
rect 698364 448374 698420 448430
rect 698488 448374 698544 448430
rect 698612 448374 698668 448430
rect 698736 448374 698792 448430
rect 697992 448250 698048 448306
rect 698116 448250 698172 448306
rect 698240 448250 698296 448306
rect 698364 448250 698420 448306
rect 698488 448250 698544 448306
rect 698612 448250 698668 448306
rect 698736 448250 698792 448306
rect 697992 448126 698048 448182
rect 698116 448126 698172 448182
rect 698240 448126 698296 448182
rect 698364 448126 698420 448182
rect 698488 448126 698544 448182
rect 698612 448126 698668 448182
rect 698736 448126 698792 448182
rect 697992 448002 698048 448058
rect 698116 448002 698172 448058
rect 698240 448002 698296 448058
rect 698364 448002 698420 448058
rect 698488 448002 698544 448058
rect 698612 448002 698668 448058
rect 698736 448002 698792 448058
rect 697992 447878 698048 447934
rect 698116 447878 698172 447934
rect 698240 447878 698296 447934
rect 698364 447878 698420 447934
rect 698488 447878 698544 447934
rect 698612 447878 698668 447934
rect 698736 447878 698792 447934
rect 697992 447754 698048 447810
rect 698116 447754 698172 447810
rect 698240 447754 698296 447810
rect 698364 447754 698420 447810
rect 698488 447754 698544 447810
rect 698612 447754 698668 447810
rect 698736 447754 698792 447810
rect 697992 447630 698048 447686
rect 698116 447630 698172 447686
rect 698240 447630 698296 447686
rect 698364 447630 698420 447686
rect 698488 447630 698544 447686
rect 698612 447630 698668 447686
rect 698736 447630 698792 447686
rect 697992 447506 698048 447562
rect 698116 447506 698172 447562
rect 698240 447506 698296 447562
rect 698364 447506 698420 447562
rect 698488 447506 698544 447562
rect 698612 447506 698668 447562
rect 698736 447506 698792 447562
rect 697992 447382 698048 447438
rect 698116 447382 698172 447438
rect 698240 447382 698296 447438
rect 698364 447382 698420 447438
rect 698488 447382 698544 447438
rect 698612 447382 698668 447438
rect 698736 447382 698792 447438
rect 697992 447258 698048 447314
rect 698116 447258 698172 447314
rect 698240 447258 698296 447314
rect 698364 447258 698420 447314
rect 698488 447258 698544 447314
rect 698612 447258 698668 447314
rect 698736 447258 698792 447314
rect 697992 447134 698048 447190
rect 698116 447134 698172 447190
rect 698240 447134 698296 447190
rect 698364 447134 698420 447190
rect 698488 447134 698544 447190
rect 698612 447134 698668 447190
rect 698736 447134 698792 447190
rect 697992 447010 698048 447066
rect 698116 447010 698172 447066
rect 698240 447010 698296 447066
rect 698364 447010 698420 447066
rect 698488 447010 698544 447066
rect 698612 447010 698668 447066
rect 698736 447010 698792 447066
rect 697992 446886 698048 446942
rect 698116 446886 698172 446942
rect 698240 446886 698296 446942
rect 698364 446886 698420 446942
rect 698488 446886 698544 446942
rect 698612 446886 698668 446942
rect 698736 446886 698792 446942
rect 697992 446040 698048 446096
rect 698116 446040 698172 446096
rect 698240 446040 698296 446096
rect 698364 446040 698420 446096
rect 698488 446040 698544 446096
rect 698612 446040 698668 446096
rect 698736 446040 698792 446096
rect 697992 445916 698048 445972
rect 698116 445916 698172 445972
rect 698240 445916 698296 445972
rect 698364 445916 698420 445972
rect 698488 445916 698544 445972
rect 698612 445916 698668 445972
rect 698736 445916 698792 445972
rect 697992 445792 698048 445848
rect 698116 445792 698172 445848
rect 698240 445792 698296 445848
rect 698364 445792 698420 445848
rect 698488 445792 698544 445848
rect 698612 445792 698668 445848
rect 698736 445792 698792 445848
rect 697992 445668 698048 445724
rect 698116 445668 698172 445724
rect 698240 445668 698296 445724
rect 698364 445668 698420 445724
rect 698488 445668 698544 445724
rect 698612 445668 698668 445724
rect 698736 445668 698792 445724
rect 697992 445544 698048 445600
rect 698116 445544 698172 445600
rect 698240 445544 698296 445600
rect 698364 445544 698420 445600
rect 698488 445544 698544 445600
rect 698612 445544 698668 445600
rect 698736 445544 698792 445600
rect 697992 445420 698048 445476
rect 698116 445420 698172 445476
rect 698240 445420 698296 445476
rect 698364 445420 698420 445476
rect 698488 445420 698544 445476
rect 698612 445420 698668 445476
rect 698736 445420 698792 445476
rect 697992 445296 698048 445352
rect 698116 445296 698172 445352
rect 698240 445296 698296 445352
rect 698364 445296 698420 445352
rect 698488 445296 698544 445352
rect 698612 445296 698668 445352
rect 698736 445296 698792 445352
rect 697992 445172 698048 445228
rect 698116 445172 698172 445228
rect 698240 445172 698296 445228
rect 698364 445172 698420 445228
rect 698488 445172 698544 445228
rect 698612 445172 698668 445228
rect 698736 445172 698792 445228
rect 697992 445048 698048 445104
rect 698116 445048 698172 445104
rect 698240 445048 698296 445104
rect 698364 445048 698420 445104
rect 698488 445048 698544 445104
rect 698612 445048 698668 445104
rect 698736 445048 698792 445104
rect 697992 444924 698048 444980
rect 698116 444924 698172 444980
rect 698240 444924 698296 444980
rect 698364 444924 698420 444980
rect 698488 444924 698544 444980
rect 698612 444924 698668 444980
rect 698736 444924 698792 444980
rect 697992 444800 698048 444856
rect 698116 444800 698172 444856
rect 698240 444800 698296 444856
rect 698364 444800 698420 444856
rect 698488 444800 698544 444856
rect 698612 444800 698668 444856
rect 698736 444800 698792 444856
rect 697992 444676 698048 444732
rect 698116 444676 698172 444732
rect 698240 444676 698296 444732
rect 698364 444676 698420 444732
rect 698488 444676 698544 444732
rect 698612 444676 698668 444732
rect 698736 444676 698792 444732
rect 697992 444552 698048 444608
rect 698116 444552 698172 444608
rect 698240 444552 698296 444608
rect 698364 444552 698420 444608
rect 698488 444552 698544 444608
rect 698612 444552 698668 444608
rect 698736 444552 698792 444608
rect 697992 444428 698048 444484
rect 698116 444428 698172 444484
rect 698240 444428 698296 444484
rect 698364 444428 698420 444484
rect 698488 444428 698544 444484
rect 698612 444428 698668 444484
rect 698736 444428 698792 444484
rect 697992 444304 698048 444360
rect 698116 444304 698172 444360
rect 698240 444304 698296 444360
rect 698364 444304 698420 444360
rect 698488 444304 698544 444360
rect 698612 444304 698668 444360
rect 698736 444304 698792 444360
rect 697992 444180 698048 444236
rect 698116 444180 698172 444236
rect 698240 444180 698296 444236
rect 698364 444180 698420 444236
rect 698488 444180 698544 444236
rect 698612 444180 698668 444236
rect 698736 444180 698792 444236
rect 697992 443670 698048 443726
rect 698116 443670 698172 443726
rect 698240 443670 698296 443726
rect 698364 443670 698420 443726
rect 698488 443670 698544 443726
rect 698612 443670 698668 443726
rect 698736 443670 698792 443726
rect 697992 443546 698048 443602
rect 698116 443546 698172 443602
rect 698240 443546 698296 443602
rect 698364 443546 698420 443602
rect 698488 443546 698544 443602
rect 698612 443546 698668 443602
rect 698736 443546 698792 443602
rect 697992 443422 698048 443478
rect 698116 443422 698172 443478
rect 698240 443422 698296 443478
rect 698364 443422 698420 443478
rect 698488 443422 698544 443478
rect 698612 443422 698668 443478
rect 698736 443422 698792 443478
rect 697992 443298 698048 443354
rect 698116 443298 698172 443354
rect 698240 443298 698296 443354
rect 698364 443298 698420 443354
rect 698488 443298 698544 443354
rect 698612 443298 698668 443354
rect 698736 443298 698792 443354
rect 697992 443174 698048 443230
rect 698116 443174 698172 443230
rect 698240 443174 698296 443230
rect 698364 443174 698420 443230
rect 698488 443174 698544 443230
rect 698612 443174 698668 443230
rect 698736 443174 698792 443230
rect 697992 443050 698048 443106
rect 698116 443050 698172 443106
rect 698240 443050 698296 443106
rect 698364 443050 698420 443106
rect 698488 443050 698544 443106
rect 698612 443050 698668 443106
rect 698736 443050 698792 443106
rect 697992 442926 698048 442982
rect 698116 442926 698172 442982
rect 698240 442926 698296 442982
rect 698364 442926 698420 442982
rect 698488 442926 698544 442982
rect 698612 442926 698668 442982
rect 698736 442926 698792 442982
rect 697992 442802 698048 442858
rect 698116 442802 698172 442858
rect 698240 442802 698296 442858
rect 698364 442802 698420 442858
rect 698488 442802 698544 442858
rect 698612 442802 698668 442858
rect 698736 442802 698792 442858
rect 697992 442678 698048 442734
rect 698116 442678 698172 442734
rect 698240 442678 698296 442734
rect 698364 442678 698420 442734
rect 698488 442678 698544 442734
rect 698612 442678 698668 442734
rect 698736 442678 698792 442734
rect 697992 442554 698048 442610
rect 698116 442554 698172 442610
rect 698240 442554 698296 442610
rect 698364 442554 698420 442610
rect 698488 442554 698544 442610
rect 698612 442554 698668 442610
rect 698736 442554 698792 442610
rect 697992 442430 698048 442486
rect 698116 442430 698172 442486
rect 698240 442430 698296 442486
rect 698364 442430 698420 442486
rect 698488 442430 698544 442486
rect 698612 442430 698668 442486
rect 698736 442430 698792 442486
rect 697992 442306 698048 442362
rect 698116 442306 698172 442362
rect 698240 442306 698296 442362
rect 698364 442306 698420 442362
rect 698488 442306 698544 442362
rect 698612 442306 698668 442362
rect 698736 442306 698792 442362
rect 697992 442182 698048 442238
rect 698116 442182 698172 442238
rect 698240 442182 698296 442238
rect 698364 442182 698420 442238
rect 698488 442182 698544 442238
rect 698612 442182 698668 442238
rect 698736 442182 698792 442238
rect 697992 442058 698048 442114
rect 698116 442058 698172 442114
rect 698240 442058 698296 442114
rect 698364 442058 698420 442114
rect 698488 442058 698544 442114
rect 698612 442058 698668 442114
rect 698736 442058 698792 442114
rect 697992 441934 698048 441990
rect 698116 441934 698172 441990
rect 698240 441934 698296 441990
rect 698364 441934 698420 441990
rect 698488 441934 698544 441990
rect 698612 441934 698668 441990
rect 698736 441934 698792 441990
rect 697992 441810 698048 441866
rect 698116 441810 698172 441866
rect 698240 441810 698296 441866
rect 698364 441810 698420 441866
rect 698488 441810 698544 441866
rect 698612 441810 698668 441866
rect 698736 441810 698792 441866
rect 697992 441066 698048 441122
rect 698116 441066 698172 441122
rect 698240 441066 698296 441122
rect 698364 441066 698420 441122
rect 698488 441066 698544 441122
rect 698612 441066 698668 441122
rect 698736 441066 698792 441122
rect 697992 440942 698048 440998
rect 698116 440942 698172 440998
rect 698240 440942 698296 440998
rect 698364 440942 698420 440998
rect 698488 440942 698544 440998
rect 698612 440942 698668 440998
rect 698736 440942 698792 440998
rect 697992 440818 698048 440874
rect 698116 440818 698172 440874
rect 698240 440818 698296 440874
rect 698364 440818 698420 440874
rect 698488 440818 698544 440874
rect 698612 440818 698668 440874
rect 698736 440818 698792 440874
rect 697992 440694 698048 440750
rect 698116 440694 698172 440750
rect 698240 440694 698296 440750
rect 698364 440694 698420 440750
rect 698488 440694 698544 440750
rect 698612 440694 698668 440750
rect 698736 440694 698792 440750
rect 697992 440570 698048 440626
rect 698116 440570 698172 440626
rect 698240 440570 698296 440626
rect 698364 440570 698420 440626
rect 698488 440570 698544 440626
rect 698612 440570 698668 440626
rect 698736 440570 698792 440626
rect 697992 440446 698048 440502
rect 698116 440446 698172 440502
rect 698240 440446 698296 440502
rect 698364 440446 698420 440502
rect 698488 440446 698544 440502
rect 698612 440446 698668 440502
rect 698736 440446 698792 440502
rect 697992 440322 698048 440378
rect 698116 440322 698172 440378
rect 698240 440322 698296 440378
rect 698364 440322 698420 440378
rect 698488 440322 698544 440378
rect 698612 440322 698668 440378
rect 698736 440322 698792 440378
rect 697992 440198 698048 440254
rect 698116 440198 698172 440254
rect 698240 440198 698296 440254
rect 698364 440198 698420 440254
rect 698488 440198 698544 440254
rect 698612 440198 698668 440254
rect 698736 440198 698792 440254
rect 697992 440074 698048 440130
rect 698116 440074 698172 440130
rect 698240 440074 698296 440130
rect 698364 440074 698420 440130
rect 698488 440074 698544 440130
rect 698612 440074 698668 440130
rect 698736 440074 698792 440130
rect 697992 439950 698048 440006
rect 698116 439950 698172 440006
rect 698240 439950 698296 440006
rect 698364 439950 698420 440006
rect 698488 439950 698544 440006
rect 698612 439950 698668 440006
rect 698736 439950 698792 440006
rect 697992 439826 698048 439882
rect 698116 439826 698172 439882
rect 698240 439826 698296 439882
rect 698364 439826 698420 439882
rect 698488 439826 698544 439882
rect 698612 439826 698668 439882
rect 698736 439826 698792 439882
rect 697992 439702 698048 439758
rect 698116 439702 698172 439758
rect 698240 439702 698296 439758
rect 698364 439702 698420 439758
rect 698488 439702 698544 439758
rect 698612 439702 698668 439758
rect 698736 439702 698792 439758
rect 697992 439578 698048 439634
rect 698116 439578 698172 439634
rect 698240 439578 698296 439634
rect 698364 439578 698420 439634
rect 698488 439578 698544 439634
rect 698612 439578 698668 439634
rect 698736 439578 698792 439634
rect 697992 439454 698048 439510
rect 698116 439454 698172 439510
rect 698240 439454 698296 439510
rect 698364 439454 698420 439510
rect 698488 439454 698544 439510
rect 698612 439454 698668 439510
rect 698736 439454 698792 439510
rect 697992 439330 698048 439386
rect 698116 439330 698172 439386
rect 698240 439330 698296 439386
rect 698364 439330 698420 439386
rect 698488 439330 698544 439386
rect 698612 439330 698668 439386
rect 698736 439330 698792 439386
rect 698144 428373 698200 428429
rect 698444 428373 698500 428429
rect 698744 428373 698800 428429
rect 698144 428173 698200 428229
rect 698444 428173 698500 428229
rect 698744 428173 698800 428229
rect 697992 410596 698048 410652
rect 698116 410596 698172 410652
rect 698240 410596 698296 410652
rect 698364 410596 698420 410652
rect 698488 410596 698544 410652
rect 698612 410596 698668 410652
rect 698736 410596 698792 410652
rect 697992 410472 698048 410528
rect 698116 410472 698172 410528
rect 698240 410472 698296 410528
rect 698364 410472 698420 410528
rect 698488 410472 698544 410528
rect 698612 410472 698668 410528
rect 698736 410472 698792 410528
rect 697992 410348 698048 410404
rect 698116 410348 698172 410404
rect 698240 410348 698296 410404
rect 698364 410348 698420 410404
rect 698488 410348 698544 410404
rect 698612 410348 698668 410404
rect 698736 410348 698792 410404
rect 697992 410224 698048 410280
rect 698116 410224 698172 410280
rect 698240 410224 698296 410280
rect 698364 410224 698420 410280
rect 698488 410224 698544 410280
rect 698612 410224 698668 410280
rect 698736 410224 698792 410280
rect 697992 410100 698048 410156
rect 698116 410100 698172 410156
rect 698240 410100 698296 410156
rect 698364 410100 698420 410156
rect 698488 410100 698544 410156
rect 698612 410100 698668 410156
rect 698736 410100 698792 410156
rect 697992 409976 698048 410032
rect 698116 409976 698172 410032
rect 698240 409976 698296 410032
rect 698364 409976 698420 410032
rect 698488 409976 698544 410032
rect 698612 409976 698668 410032
rect 698736 409976 698792 410032
rect 697992 409852 698048 409908
rect 698116 409852 698172 409908
rect 698240 409852 698296 409908
rect 698364 409852 698420 409908
rect 698488 409852 698544 409908
rect 698612 409852 698668 409908
rect 698736 409852 698792 409908
rect 697992 409728 698048 409784
rect 698116 409728 698172 409784
rect 698240 409728 698296 409784
rect 698364 409728 698420 409784
rect 698488 409728 698544 409784
rect 698612 409728 698668 409784
rect 698736 409728 698792 409784
rect 697992 409604 698048 409660
rect 698116 409604 698172 409660
rect 698240 409604 698296 409660
rect 698364 409604 698420 409660
rect 698488 409604 698544 409660
rect 698612 409604 698668 409660
rect 698736 409604 698792 409660
rect 697992 409480 698048 409536
rect 698116 409480 698172 409536
rect 698240 409480 698296 409536
rect 698364 409480 698420 409536
rect 698488 409480 698544 409536
rect 698612 409480 698668 409536
rect 698736 409480 698792 409536
rect 697992 409356 698048 409412
rect 698116 409356 698172 409412
rect 698240 409356 698296 409412
rect 698364 409356 698420 409412
rect 698488 409356 698544 409412
rect 698612 409356 698668 409412
rect 698736 409356 698792 409412
rect 697992 409232 698048 409288
rect 698116 409232 698172 409288
rect 698240 409232 698296 409288
rect 698364 409232 698420 409288
rect 698488 409232 698544 409288
rect 698612 409232 698668 409288
rect 698736 409232 698792 409288
rect 697992 409108 698048 409164
rect 698116 409108 698172 409164
rect 698240 409108 698296 409164
rect 698364 409108 698420 409164
rect 698488 409108 698544 409164
rect 698612 409108 698668 409164
rect 698736 409108 698792 409164
rect 697992 408984 698048 409040
rect 698116 408984 698172 409040
rect 698240 408984 698296 409040
rect 698364 408984 698420 409040
rect 698488 408984 698544 409040
rect 698612 408984 698668 409040
rect 698736 408984 698792 409040
rect 697992 408860 698048 408916
rect 698116 408860 698172 408916
rect 698240 408860 698296 408916
rect 698364 408860 698420 408916
rect 698488 408860 698544 408916
rect 698612 408860 698668 408916
rect 698736 408860 698792 408916
rect 697992 408116 698048 408172
rect 698116 408116 698172 408172
rect 698240 408116 698296 408172
rect 698364 408116 698420 408172
rect 698488 408116 698544 408172
rect 698612 408116 698668 408172
rect 698736 408116 698792 408172
rect 697992 407992 698048 408048
rect 698116 407992 698172 408048
rect 698240 407992 698296 408048
rect 698364 407992 698420 408048
rect 698488 407992 698544 408048
rect 698612 407992 698668 408048
rect 698736 407992 698792 408048
rect 697992 407868 698048 407924
rect 698116 407868 698172 407924
rect 698240 407868 698296 407924
rect 698364 407868 698420 407924
rect 698488 407868 698544 407924
rect 698612 407868 698668 407924
rect 698736 407868 698792 407924
rect 697992 407744 698048 407800
rect 698116 407744 698172 407800
rect 698240 407744 698296 407800
rect 698364 407744 698420 407800
rect 698488 407744 698544 407800
rect 698612 407744 698668 407800
rect 698736 407744 698792 407800
rect 697992 407620 698048 407676
rect 698116 407620 698172 407676
rect 698240 407620 698296 407676
rect 698364 407620 698420 407676
rect 698488 407620 698544 407676
rect 698612 407620 698668 407676
rect 698736 407620 698792 407676
rect 697992 407496 698048 407552
rect 698116 407496 698172 407552
rect 698240 407496 698296 407552
rect 698364 407496 698420 407552
rect 698488 407496 698544 407552
rect 698612 407496 698668 407552
rect 698736 407496 698792 407552
rect 697992 407372 698048 407428
rect 698116 407372 698172 407428
rect 698240 407372 698296 407428
rect 698364 407372 698420 407428
rect 698488 407372 698544 407428
rect 698612 407372 698668 407428
rect 698736 407372 698792 407428
rect 697992 407248 698048 407304
rect 698116 407248 698172 407304
rect 698240 407248 698296 407304
rect 698364 407248 698420 407304
rect 698488 407248 698544 407304
rect 698612 407248 698668 407304
rect 698736 407248 698792 407304
rect 697992 407124 698048 407180
rect 698116 407124 698172 407180
rect 698240 407124 698296 407180
rect 698364 407124 698420 407180
rect 698488 407124 698544 407180
rect 698612 407124 698668 407180
rect 698736 407124 698792 407180
rect 697992 407000 698048 407056
rect 698116 407000 698172 407056
rect 698240 407000 698296 407056
rect 698364 407000 698420 407056
rect 698488 407000 698544 407056
rect 698612 407000 698668 407056
rect 698736 407000 698792 407056
rect 697992 406876 698048 406932
rect 698116 406876 698172 406932
rect 698240 406876 698296 406932
rect 698364 406876 698420 406932
rect 698488 406876 698544 406932
rect 698612 406876 698668 406932
rect 698736 406876 698792 406932
rect 697992 406752 698048 406808
rect 698116 406752 698172 406808
rect 698240 406752 698296 406808
rect 698364 406752 698420 406808
rect 698488 406752 698544 406808
rect 698612 406752 698668 406808
rect 698736 406752 698792 406808
rect 697992 406628 698048 406684
rect 698116 406628 698172 406684
rect 698240 406628 698296 406684
rect 698364 406628 698420 406684
rect 698488 406628 698544 406684
rect 698612 406628 698668 406684
rect 698736 406628 698792 406684
rect 697992 406504 698048 406560
rect 698116 406504 698172 406560
rect 698240 406504 698296 406560
rect 698364 406504 698420 406560
rect 698488 406504 698544 406560
rect 698612 406504 698668 406560
rect 698736 406504 698792 406560
rect 697992 406380 698048 406436
rect 698116 406380 698172 406436
rect 698240 406380 698296 406436
rect 698364 406380 698420 406436
rect 698488 406380 698544 406436
rect 698612 406380 698668 406436
rect 698736 406380 698792 406436
rect 697992 406256 698048 406312
rect 698116 406256 698172 406312
rect 698240 406256 698296 406312
rect 698364 406256 698420 406312
rect 698488 406256 698544 406312
rect 698612 406256 698668 406312
rect 698736 406256 698792 406312
rect 697992 405746 698048 405802
rect 698116 405746 698172 405802
rect 698240 405746 698296 405802
rect 698364 405746 698420 405802
rect 698488 405746 698544 405802
rect 698612 405746 698668 405802
rect 698736 405746 698792 405802
rect 697992 405622 698048 405678
rect 698116 405622 698172 405678
rect 698240 405622 698296 405678
rect 698364 405622 698420 405678
rect 698488 405622 698544 405678
rect 698612 405622 698668 405678
rect 698736 405622 698792 405678
rect 697992 405498 698048 405554
rect 698116 405498 698172 405554
rect 698240 405498 698296 405554
rect 698364 405498 698420 405554
rect 698488 405498 698544 405554
rect 698612 405498 698668 405554
rect 698736 405498 698792 405554
rect 697992 405374 698048 405430
rect 698116 405374 698172 405430
rect 698240 405374 698296 405430
rect 698364 405374 698420 405430
rect 698488 405374 698544 405430
rect 698612 405374 698668 405430
rect 698736 405374 698792 405430
rect 697992 405250 698048 405306
rect 698116 405250 698172 405306
rect 698240 405250 698296 405306
rect 698364 405250 698420 405306
rect 698488 405250 698544 405306
rect 698612 405250 698668 405306
rect 698736 405250 698792 405306
rect 697992 405126 698048 405182
rect 698116 405126 698172 405182
rect 698240 405126 698296 405182
rect 698364 405126 698420 405182
rect 698488 405126 698544 405182
rect 698612 405126 698668 405182
rect 698736 405126 698792 405182
rect 697992 405002 698048 405058
rect 698116 405002 698172 405058
rect 698240 405002 698296 405058
rect 698364 405002 698420 405058
rect 698488 405002 698544 405058
rect 698612 405002 698668 405058
rect 698736 405002 698792 405058
rect 697992 404878 698048 404934
rect 698116 404878 698172 404934
rect 698240 404878 698296 404934
rect 698364 404878 698420 404934
rect 698488 404878 698544 404934
rect 698612 404878 698668 404934
rect 698736 404878 698792 404934
rect 697992 404754 698048 404810
rect 698116 404754 698172 404810
rect 698240 404754 698296 404810
rect 698364 404754 698420 404810
rect 698488 404754 698544 404810
rect 698612 404754 698668 404810
rect 698736 404754 698792 404810
rect 697992 404630 698048 404686
rect 698116 404630 698172 404686
rect 698240 404630 698296 404686
rect 698364 404630 698420 404686
rect 698488 404630 698544 404686
rect 698612 404630 698668 404686
rect 698736 404630 698792 404686
rect 697992 404506 698048 404562
rect 698116 404506 698172 404562
rect 698240 404506 698296 404562
rect 698364 404506 698420 404562
rect 698488 404506 698544 404562
rect 698612 404506 698668 404562
rect 698736 404506 698792 404562
rect 697992 404382 698048 404438
rect 698116 404382 698172 404438
rect 698240 404382 698296 404438
rect 698364 404382 698420 404438
rect 698488 404382 698544 404438
rect 698612 404382 698668 404438
rect 698736 404382 698792 404438
rect 697992 404258 698048 404314
rect 698116 404258 698172 404314
rect 698240 404258 698296 404314
rect 698364 404258 698420 404314
rect 698488 404258 698544 404314
rect 698612 404258 698668 404314
rect 698736 404258 698792 404314
rect 697992 404134 698048 404190
rect 698116 404134 698172 404190
rect 698240 404134 698296 404190
rect 698364 404134 698420 404190
rect 698488 404134 698544 404190
rect 698612 404134 698668 404190
rect 698736 404134 698792 404190
rect 697992 404010 698048 404066
rect 698116 404010 698172 404066
rect 698240 404010 698296 404066
rect 698364 404010 698420 404066
rect 698488 404010 698544 404066
rect 698612 404010 698668 404066
rect 698736 404010 698792 404066
rect 697992 403886 698048 403942
rect 698116 403886 698172 403942
rect 698240 403886 698296 403942
rect 698364 403886 698420 403942
rect 698488 403886 698544 403942
rect 698612 403886 698668 403942
rect 698736 403886 698792 403942
rect 697992 403040 698048 403096
rect 698116 403040 698172 403096
rect 698240 403040 698296 403096
rect 698364 403040 698420 403096
rect 698488 403040 698544 403096
rect 698612 403040 698668 403096
rect 698736 403040 698792 403096
rect 697992 402916 698048 402972
rect 698116 402916 698172 402972
rect 698240 402916 698296 402972
rect 698364 402916 698420 402972
rect 698488 402916 698544 402972
rect 698612 402916 698668 402972
rect 698736 402916 698792 402972
rect 697992 402792 698048 402848
rect 698116 402792 698172 402848
rect 698240 402792 698296 402848
rect 698364 402792 698420 402848
rect 698488 402792 698544 402848
rect 698612 402792 698668 402848
rect 698736 402792 698792 402848
rect 697992 402668 698048 402724
rect 698116 402668 698172 402724
rect 698240 402668 698296 402724
rect 698364 402668 698420 402724
rect 698488 402668 698544 402724
rect 698612 402668 698668 402724
rect 698736 402668 698792 402724
rect 697992 402544 698048 402600
rect 698116 402544 698172 402600
rect 698240 402544 698296 402600
rect 698364 402544 698420 402600
rect 698488 402544 698544 402600
rect 698612 402544 698668 402600
rect 698736 402544 698792 402600
rect 697992 402420 698048 402476
rect 698116 402420 698172 402476
rect 698240 402420 698296 402476
rect 698364 402420 698420 402476
rect 698488 402420 698544 402476
rect 698612 402420 698668 402476
rect 698736 402420 698792 402476
rect 697992 402296 698048 402352
rect 698116 402296 698172 402352
rect 698240 402296 698296 402352
rect 698364 402296 698420 402352
rect 698488 402296 698544 402352
rect 698612 402296 698668 402352
rect 698736 402296 698792 402352
rect 697992 402172 698048 402228
rect 698116 402172 698172 402228
rect 698240 402172 698296 402228
rect 698364 402172 698420 402228
rect 698488 402172 698544 402228
rect 698612 402172 698668 402228
rect 698736 402172 698792 402228
rect 697992 402048 698048 402104
rect 698116 402048 698172 402104
rect 698240 402048 698296 402104
rect 698364 402048 698420 402104
rect 698488 402048 698544 402104
rect 698612 402048 698668 402104
rect 698736 402048 698792 402104
rect 697992 401924 698048 401980
rect 698116 401924 698172 401980
rect 698240 401924 698296 401980
rect 698364 401924 698420 401980
rect 698488 401924 698544 401980
rect 698612 401924 698668 401980
rect 698736 401924 698792 401980
rect 697992 401800 698048 401856
rect 698116 401800 698172 401856
rect 698240 401800 698296 401856
rect 698364 401800 698420 401856
rect 698488 401800 698544 401856
rect 698612 401800 698668 401856
rect 698736 401800 698792 401856
rect 697992 401676 698048 401732
rect 698116 401676 698172 401732
rect 698240 401676 698296 401732
rect 698364 401676 698420 401732
rect 698488 401676 698544 401732
rect 698612 401676 698668 401732
rect 698736 401676 698792 401732
rect 697992 401552 698048 401608
rect 698116 401552 698172 401608
rect 698240 401552 698296 401608
rect 698364 401552 698420 401608
rect 698488 401552 698544 401608
rect 698612 401552 698668 401608
rect 698736 401552 698792 401608
rect 697992 401428 698048 401484
rect 698116 401428 698172 401484
rect 698240 401428 698296 401484
rect 698364 401428 698420 401484
rect 698488 401428 698544 401484
rect 698612 401428 698668 401484
rect 698736 401428 698792 401484
rect 697992 401304 698048 401360
rect 698116 401304 698172 401360
rect 698240 401304 698296 401360
rect 698364 401304 698420 401360
rect 698488 401304 698544 401360
rect 698612 401304 698668 401360
rect 698736 401304 698792 401360
rect 697992 401180 698048 401236
rect 698116 401180 698172 401236
rect 698240 401180 698296 401236
rect 698364 401180 698420 401236
rect 698488 401180 698544 401236
rect 698612 401180 698668 401236
rect 698736 401180 698792 401236
rect 697992 400670 698048 400726
rect 698116 400670 698172 400726
rect 698240 400670 698296 400726
rect 698364 400670 698420 400726
rect 698488 400670 698544 400726
rect 698612 400670 698668 400726
rect 698736 400670 698792 400726
rect 697992 400546 698048 400602
rect 698116 400546 698172 400602
rect 698240 400546 698296 400602
rect 698364 400546 698420 400602
rect 698488 400546 698544 400602
rect 698612 400546 698668 400602
rect 698736 400546 698792 400602
rect 697992 400422 698048 400478
rect 698116 400422 698172 400478
rect 698240 400422 698296 400478
rect 698364 400422 698420 400478
rect 698488 400422 698544 400478
rect 698612 400422 698668 400478
rect 698736 400422 698792 400478
rect 697992 400298 698048 400354
rect 698116 400298 698172 400354
rect 698240 400298 698296 400354
rect 698364 400298 698420 400354
rect 698488 400298 698544 400354
rect 698612 400298 698668 400354
rect 698736 400298 698792 400354
rect 697992 400174 698048 400230
rect 698116 400174 698172 400230
rect 698240 400174 698296 400230
rect 698364 400174 698420 400230
rect 698488 400174 698544 400230
rect 698612 400174 698668 400230
rect 698736 400174 698792 400230
rect 697992 400050 698048 400106
rect 698116 400050 698172 400106
rect 698240 400050 698296 400106
rect 698364 400050 698420 400106
rect 698488 400050 698544 400106
rect 698612 400050 698668 400106
rect 698736 400050 698792 400106
rect 697992 399926 698048 399982
rect 698116 399926 698172 399982
rect 698240 399926 698296 399982
rect 698364 399926 698420 399982
rect 698488 399926 698544 399982
rect 698612 399926 698668 399982
rect 698736 399926 698792 399982
rect 697992 399802 698048 399858
rect 698116 399802 698172 399858
rect 698240 399802 698296 399858
rect 698364 399802 698420 399858
rect 698488 399802 698544 399858
rect 698612 399802 698668 399858
rect 698736 399802 698792 399858
rect 697992 399678 698048 399734
rect 698116 399678 698172 399734
rect 698240 399678 698296 399734
rect 698364 399678 698420 399734
rect 698488 399678 698544 399734
rect 698612 399678 698668 399734
rect 698736 399678 698792 399734
rect 697992 399554 698048 399610
rect 698116 399554 698172 399610
rect 698240 399554 698296 399610
rect 698364 399554 698420 399610
rect 698488 399554 698544 399610
rect 698612 399554 698668 399610
rect 698736 399554 698792 399610
rect 697992 399430 698048 399486
rect 698116 399430 698172 399486
rect 698240 399430 698296 399486
rect 698364 399430 698420 399486
rect 698488 399430 698544 399486
rect 698612 399430 698668 399486
rect 698736 399430 698792 399486
rect 697992 399306 698048 399362
rect 698116 399306 698172 399362
rect 698240 399306 698296 399362
rect 698364 399306 698420 399362
rect 698488 399306 698544 399362
rect 698612 399306 698668 399362
rect 698736 399306 698792 399362
rect 697992 399182 698048 399238
rect 698116 399182 698172 399238
rect 698240 399182 698296 399238
rect 698364 399182 698420 399238
rect 698488 399182 698544 399238
rect 698612 399182 698668 399238
rect 698736 399182 698792 399238
rect 697992 399058 698048 399114
rect 698116 399058 698172 399114
rect 698240 399058 698296 399114
rect 698364 399058 698420 399114
rect 698488 399058 698544 399114
rect 698612 399058 698668 399114
rect 698736 399058 698792 399114
rect 697992 398934 698048 398990
rect 698116 398934 698172 398990
rect 698240 398934 698296 398990
rect 698364 398934 698420 398990
rect 698488 398934 698544 398990
rect 698612 398934 698668 398990
rect 698736 398934 698792 398990
rect 697992 398810 698048 398866
rect 698116 398810 698172 398866
rect 698240 398810 698296 398866
rect 698364 398810 698420 398866
rect 698488 398810 698544 398866
rect 698612 398810 698668 398866
rect 698736 398810 698792 398866
rect 697992 398066 698048 398122
rect 698116 398066 698172 398122
rect 698240 398066 698296 398122
rect 698364 398066 698420 398122
rect 698488 398066 698544 398122
rect 698612 398066 698668 398122
rect 698736 398066 698792 398122
rect 697992 397942 698048 397998
rect 698116 397942 698172 397998
rect 698240 397942 698296 397998
rect 698364 397942 698420 397998
rect 698488 397942 698544 397998
rect 698612 397942 698668 397998
rect 698736 397942 698792 397998
rect 697992 397818 698048 397874
rect 698116 397818 698172 397874
rect 698240 397818 698296 397874
rect 698364 397818 698420 397874
rect 698488 397818 698544 397874
rect 698612 397818 698668 397874
rect 698736 397818 698792 397874
rect 697992 397694 698048 397750
rect 698116 397694 698172 397750
rect 698240 397694 698296 397750
rect 698364 397694 698420 397750
rect 698488 397694 698544 397750
rect 698612 397694 698668 397750
rect 698736 397694 698792 397750
rect 697992 397570 698048 397626
rect 698116 397570 698172 397626
rect 698240 397570 698296 397626
rect 698364 397570 698420 397626
rect 698488 397570 698544 397626
rect 698612 397570 698668 397626
rect 698736 397570 698792 397626
rect 697992 397446 698048 397502
rect 698116 397446 698172 397502
rect 698240 397446 698296 397502
rect 698364 397446 698420 397502
rect 698488 397446 698544 397502
rect 698612 397446 698668 397502
rect 698736 397446 698792 397502
rect 697992 397322 698048 397378
rect 698116 397322 698172 397378
rect 698240 397322 698296 397378
rect 698364 397322 698420 397378
rect 698488 397322 698544 397378
rect 698612 397322 698668 397378
rect 698736 397322 698792 397378
rect 697992 397198 698048 397254
rect 698116 397198 698172 397254
rect 698240 397198 698296 397254
rect 698364 397198 698420 397254
rect 698488 397198 698544 397254
rect 698612 397198 698668 397254
rect 698736 397198 698792 397254
rect 697992 397074 698048 397130
rect 698116 397074 698172 397130
rect 698240 397074 698296 397130
rect 698364 397074 698420 397130
rect 698488 397074 698544 397130
rect 698612 397074 698668 397130
rect 698736 397074 698792 397130
rect 697992 396950 698048 397006
rect 698116 396950 698172 397006
rect 698240 396950 698296 397006
rect 698364 396950 698420 397006
rect 698488 396950 698544 397006
rect 698612 396950 698668 397006
rect 698736 396950 698792 397006
rect 697992 396826 698048 396882
rect 698116 396826 698172 396882
rect 698240 396826 698296 396882
rect 698364 396826 698420 396882
rect 698488 396826 698544 396882
rect 698612 396826 698668 396882
rect 698736 396826 698792 396882
rect 697992 396702 698048 396758
rect 698116 396702 698172 396758
rect 698240 396702 698296 396758
rect 698364 396702 698420 396758
rect 698488 396702 698544 396758
rect 698612 396702 698668 396758
rect 698736 396702 698792 396758
rect 697992 396578 698048 396634
rect 698116 396578 698172 396634
rect 698240 396578 698296 396634
rect 698364 396578 698420 396634
rect 698488 396578 698544 396634
rect 698612 396578 698668 396634
rect 698736 396578 698792 396634
rect 697992 396454 698048 396510
rect 698116 396454 698172 396510
rect 698240 396454 698296 396510
rect 698364 396454 698420 396510
rect 698488 396454 698544 396510
rect 698612 396454 698668 396510
rect 698736 396454 698792 396510
rect 697992 396330 698048 396386
rect 698116 396330 698172 396386
rect 698240 396330 698296 396386
rect 698364 396330 698420 396386
rect 698488 396330 698544 396386
rect 698612 396330 698668 396386
rect 698736 396330 698792 396386
rect 698144 392373 698200 392429
rect 698444 392373 698500 392429
rect 698744 392373 698800 392429
rect 698144 392173 698200 392229
rect 698444 392173 698500 392229
rect 698744 392173 698800 392229
rect 698044 363378 698100 363434
rect 698344 363378 698400 363434
rect 698644 363378 698700 363434
rect 698144 356373 698200 356429
rect 698444 356373 698500 356429
rect 698744 356373 698800 356429
rect 698144 356173 698200 356229
rect 698444 356173 698500 356229
rect 698744 356173 698800 356229
rect 698044 349378 698100 349434
rect 698344 349378 698400 349434
rect 698644 349378 698700 349434
rect 79208 330984 79264 331040
rect 79332 330984 79388 331040
rect 79456 330984 79512 331040
rect 79580 330984 79636 331040
rect 79704 330984 79760 331040
rect 79828 330984 79884 331040
rect 79952 330984 80008 331040
rect 79208 330860 79264 330916
rect 79332 330860 79388 330916
rect 79456 330860 79512 330916
rect 79580 330860 79636 330916
rect 79704 330860 79760 330916
rect 79828 330860 79884 330916
rect 79952 330860 80008 330916
rect 79208 330736 79264 330792
rect 79332 330736 79388 330792
rect 79456 330736 79512 330792
rect 79580 330736 79636 330792
rect 79704 330736 79760 330792
rect 79828 330736 79884 330792
rect 79952 330736 80008 330792
rect 79208 330612 79264 330668
rect 79332 330612 79388 330668
rect 79456 330612 79512 330668
rect 79580 330612 79636 330668
rect 79704 330612 79760 330668
rect 79828 330612 79884 330668
rect 79952 330612 80008 330668
rect 79208 330488 79264 330544
rect 79332 330488 79388 330544
rect 79456 330488 79512 330544
rect 79580 330488 79636 330544
rect 79704 330488 79760 330544
rect 79828 330488 79884 330544
rect 79952 330488 80008 330544
rect 79208 330364 79264 330420
rect 79332 330364 79388 330420
rect 79456 330364 79512 330420
rect 79580 330364 79636 330420
rect 79704 330364 79760 330420
rect 79828 330364 79884 330420
rect 79952 330364 80008 330420
rect 79208 330240 79264 330296
rect 79332 330240 79388 330296
rect 79456 330240 79512 330296
rect 79580 330240 79636 330296
rect 79704 330240 79760 330296
rect 79828 330240 79884 330296
rect 79952 330240 80008 330296
rect 106207 330832 106263 330888
rect 106407 330832 106463 330888
rect 106207 330532 106263 330588
rect 106407 330532 106463 330588
rect 106207 330232 106263 330288
rect 106407 330232 106463 330288
rect 88207 329432 88263 329488
rect 88407 329432 88463 329488
rect 88207 329132 88263 329188
rect 88407 329132 88463 329188
rect 88207 328832 88263 328888
rect 88407 328832 88463 328888
rect 142207 330832 142263 330888
rect 142407 330832 142463 330888
rect 142207 330532 142263 330588
rect 142407 330532 142463 330588
rect 142207 330232 142263 330288
rect 142407 330232 142463 330288
rect 158178 330984 158234 331040
rect 158302 330984 158358 331040
rect 158426 330984 158482 331040
rect 158550 330984 158606 331040
rect 158178 330860 158234 330916
rect 158302 330860 158358 330916
rect 158426 330860 158482 330916
rect 158550 330860 158606 330916
rect 158178 330736 158234 330792
rect 158302 330736 158358 330792
rect 158426 330736 158482 330792
rect 158550 330736 158606 330792
rect 158178 330612 158234 330668
rect 158302 330612 158358 330668
rect 158426 330612 158482 330668
rect 158550 330612 158606 330668
rect 158178 330488 158234 330544
rect 158302 330488 158358 330544
rect 158426 330488 158482 330544
rect 158550 330488 158606 330544
rect 158178 330364 158234 330420
rect 158302 330364 158358 330420
rect 158426 330364 158482 330420
rect 158550 330364 158606 330420
rect 158178 330240 158234 330296
rect 158302 330240 158358 330296
rect 158426 330240 158482 330296
rect 158550 330240 158606 330296
rect 124207 329432 124263 329488
rect 124407 329432 124463 329488
rect 124207 329132 124263 329188
rect 124407 329132 124463 329188
rect 124207 328832 124263 328888
rect 124407 328832 124463 328888
rect 157158 329584 157214 329640
rect 157282 329584 157338 329640
rect 157406 329584 157462 329640
rect 157530 329584 157586 329640
rect 157158 329460 157214 329516
rect 157282 329460 157338 329516
rect 157406 329460 157462 329516
rect 157530 329460 157586 329516
rect 157158 329336 157214 329392
rect 157282 329336 157338 329392
rect 157406 329336 157462 329392
rect 157530 329336 157586 329392
rect 157158 329212 157214 329268
rect 157282 329212 157338 329268
rect 157406 329212 157462 329268
rect 157530 329212 157586 329268
rect 157158 329088 157214 329144
rect 157282 329088 157338 329144
rect 157406 329088 157462 329144
rect 157530 329088 157586 329144
rect 157158 328964 157214 329020
rect 157282 328964 157338 329020
rect 157406 328964 157462 329020
rect 157530 328964 157586 329020
rect 157158 328840 157214 328896
rect 157282 328840 157338 328896
rect 157406 328840 157462 328896
rect 157530 328840 157586 328896
rect 79300 314566 79356 314622
rect 79600 314566 79656 314622
rect 79900 314566 79956 314622
rect 157210 318368 157266 318424
rect 157510 318368 157566 318424
rect 157210 316970 157266 317026
rect 157510 316970 157566 317026
rect 157210 315572 157266 315628
rect 157510 315572 157566 315628
rect 79300 307566 79356 307622
rect 79600 307566 79656 307622
rect 79900 307566 79956 307622
rect 79208 307130 79264 307186
rect 79332 307130 79388 307186
rect 79456 307130 79512 307186
rect 79580 307130 79636 307186
rect 79704 307130 79760 307186
rect 79828 307130 79884 307186
rect 79952 307130 80008 307186
rect 79208 307006 79264 307062
rect 79332 307006 79388 307062
rect 79456 307006 79512 307062
rect 79580 307006 79636 307062
rect 79704 307006 79760 307062
rect 79828 307006 79884 307062
rect 79952 307006 80008 307062
rect 79208 306882 79264 306938
rect 79332 306882 79388 306938
rect 79456 306882 79512 306938
rect 79580 306882 79636 306938
rect 79704 306882 79760 306938
rect 79828 306882 79884 306938
rect 79952 306882 80008 306938
rect 79208 306758 79264 306814
rect 79332 306758 79388 306814
rect 79456 306758 79512 306814
rect 79580 306758 79636 306814
rect 79704 306758 79760 306814
rect 79828 306758 79884 306814
rect 79952 306758 80008 306814
rect 79208 306634 79264 306690
rect 79332 306634 79388 306690
rect 79456 306634 79512 306690
rect 79580 306634 79636 306690
rect 79704 306634 79760 306690
rect 79828 306634 79884 306690
rect 79952 306634 80008 306690
rect 79208 306510 79264 306566
rect 79332 306510 79388 306566
rect 79456 306510 79512 306566
rect 79580 306510 79636 306566
rect 79704 306510 79760 306566
rect 79828 306510 79884 306566
rect 79952 306510 80008 306566
rect 79208 306386 79264 306442
rect 79332 306386 79388 306442
rect 79456 306386 79512 306442
rect 79580 306386 79636 306442
rect 79704 306386 79760 306442
rect 79828 306386 79884 306442
rect 79952 306386 80008 306442
rect 116220 307130 116276 307186
rect 116344 307130 116400 307186
rect 116220 307006 116276 307062
rect 116344 307006 116400 307062
rect 116220 306882 116276 306938
rect 116344 306882 116400 306938
rect 116220 306758 116276 306814
rect 116344 306758 116400 306814
rect 116220 306634 116276 306690
rect 116344 306634 116400 306690
rect 116220 306510 116276 306566
rect 116344 306510 116400 306566
rect 116220 306386 116276 306442
rect 116344 306386 116400 306442
rect 114625 305730 114681 305786
rect 114749 305730 114805 305786
rect 114625 305606 114681 305662
rect 114749 305606 114805 305662
rect 114625 305482 114681 305538
rect 114749 305482 114805 305538
rect 114625 305358 114681 305414
rect 114749 305358 114805 305414
rect 114625 305234 114681 305290
rect 114749 305234 114805 305290
rect 114625 305110 114681 305166
rect 114749 305110 114805 305166
rect 114625 304986 114681 305042
rect 114749 304986 114805 305042
rect 119410 307130 119466 307186
rect 119534 307130 119590 307186
rect 119410 307006 119466 307062
rect 119534 307006 119590 307062
rect 119410 306882 119466 306938
rect 119534 306882 119590 306938
rect 119410 306758 119466 306814
rect 119534 306758 119590 306814
rect 119410 306634 119466 306690
rect 119534 306634 119590 306690
rect 119410 306510 119466 306566
rect 119534 306510 119590 306566
rect 119410 306386 119466 306442
rect 119534 306386 119590 306442
rect 117815 305730 117871 305786
rect 117939 305730 117995 305786
rect 117815 305606 117871 305662
rect 117939 305606 117995 305662
rect 117815 305482 117871 305538
rect 117939 305482 117995 305538
rect 117815 305358 117871 305414
rect 117939 305358 117995 305414
rect 117815 305234 117871 305290
rect 117939 305234 117995 305290
rect 117815 305110 117871 305166
rect 117939 305110 117995 305166
rect 117815 304986 117871 305042
rect 117939 304986 117995 305042
rect 122600 307130 122656 307186
rect 122724 307130 122780 307186
rect 122600 307006 122656 307062
rect 122724 307006 122780 307062
rect 122600 306882 122656 306938
rect 122724 306882 122780 306938
rect 122600 306758 122656 306814
rect 122724 306758 122780 306814
rect 122600 306634 122656 306690
rect 122724 306634 122780 306690
rect 122600 306510 122656 306566
rect 122724 306510 122780 306566
rect 122600 306386 122656 306442
rect 122724 306386 122780 306442
rect 121005 305730 121061 305786
rect 121129 305730 121185 305786
rect 121005 305606 121061 305662
rect 121129 305606 121185 305662
rect 121005 305482 121061 305538
rect 121129 305482 121185 305538
rect 121005 305358 121061 305414
rect 121129 305358 121185 305414
rect 121005 305234 121061 305290
rect 121129 305234 121185 305290
rect 121005 305110 121061 305166
rect 121129 305110 121185 305166
rect 121005 304986 121061 305042
rect 121129 304986 121185 305042
rect 124195 305730 124251 305786
rect 124319 305730 124375 305786
rect 124195 305606 124251 305662
rect 124319 305606 124375 305662
rect 124195 305482 124251 305538
rect 124319 305482 124375 305538
rect 124195 305358 124251 305414
rect 124319 305358 124375 305414
rect 124195 305234 124251 305290
rect 124319 305234 124375 305290
rect 124195 305110 124251 305166
rect 124319 305110 124375 305166
rect 124195 304986 124251 305042
rect 124319 304986 124375 305042
rect 157210 314174 157266 314230
rect 157510 314174 157566 314230
rect 178207 330832 178263 330888
rect 178407 330832 178463 330888
rect 178207 330532 178263 330588
rect 178407 330532 178463 330588
rect 178207 330232 178263 330288
rect 178407 330232 178463 330288
rect 160207 329432 160263 329488
rect 160407 329432 160463 329488
rect 160207 329132 160263 329188
rect 160407 329132 160463 329188
rect 160207 328832 160263 328888
rect 160407 328832 160463 328888
rect 214207 330832 214263 330888
rect 214407 330832 214463 330888
rect 214207 330532 214263 330588
rect 214407 330532 214463 330588
rect 214207 330232 214263 330288
rect 214407 330232 214463 330288
rect 196207 329432 196263 329488
rect 196407 329432 196463 329488
rect 196207 329132 196263 329188
rect 196407 329132 196463 329188
rect 196207 328832 196263 328888
rect 196407 328832 196463 328888
rect 250207 330832 250263 330888
rect 250407 330832 250463 330888
rect 250207 330532 250263 330588
rect 250407 330532 250463 330588
rect 250207 330232 250263 330288
rect 250407 330232 250463 330288
rect 232207 329432 232263 329488
rect 232407 329432 232463 329488
rect 232207 329132 232263 329188
rect 232407 329132 232463 329188
rect 232207 328832 232263 328888
rect 232407 328832 232463 328888
rect 286207 330832 286263 330888
rect 286407 330832 286463 330888
rect 286207 330532 286263 330588
rect 286407 330532 286463 330588
rect 286207 330232 286263 330288
rect 286407 330232 286463 330288
rect 268207 329432 268263 329488
rect 268407 329432 268463 329488
rect 268207 329132 268263 329188
rect 268407 329132 268463 329188
rect 268207 328832 268263 328888
rect 268407 328832 268463 328888
rect 322207 330832 322263 330888
rect 322407 330832 322463 330888
rect 322207 330532 322263 330588
rect 322407 330532 322463 330588
rect 322207 330232 322263 330288
rect 322407 330232 322463 330288
rect 304207 329432 304263 329488
rect 304407 329432 304463 329488
rect 304207 329132 304263 329188
rect 304407 329132 304463 329188
rect 304207 328832 304263 328888
rect 304407 328832 304463 328888
rect 358207 330832 358263 330888
rect 358407 330832 358463 330888
rect 358207 330532 358263 330588
rect 358407 330532 358463 330588
rect 358207 330232 358263 330288
rect 358407 330232 358463 330288
rect 340207 329432 340263 329488
rect 340407 329432 340463 329488
rect 340207 329132 340263 329188
rect 340407 329132 340463 329188
rect 340207 328832 340263 328888
rect 340407 328832 340463 328888
rect 376207 329432 376263 329488
rect 376407 329432 376463 329488
rect 376207 329132 376263 329188
rect 376407 329132 376463 329188
rect 376207 328832 376263 328888
rect 376407 328832 376463 328888
rect 381310 330984 381366 331040
rect 381434 330984 381490 331040
rect 381558 330984 381614 331040
rect 381682 330984 381738 331040
rect 381310 330860 381366 330916
rect 381434 330860 381490 330916
rect 381558 330860 381614 330916
rect 381682 330860 381738 330916
rect 381310 330736 381366 330792
rect 381434 330736 381490 330792
rect 381558 330736 381614 330792
rect 381682 330736 381738 330792
rect 381310 330612 381366 330668
rect 381434 330612 381490 330668
rect 381558 330612 381614 330668
rect 381682 330612 381738 330668
rect 381310 330488 381366 330544
rect 381434 330488 381490 330544
rect 381558 330488 381614 330544
rect 381682 330488 381738 330544
rect 381310 330364 381366 330420
rect 381434 330364 381490 330420
rect 381558 330364 381614 330420
rect 381682 330364 381738 330420
rect 381310 330240 381366 330296
rect 381434 330240 381490 330296
rect 381558 330240 381614 330296
rect 381682 330240 381738 330296
rect 158230 317669 158286 317725
rect 158530 317669 158586 317725
rect 158230 316271 158286 316327
rect 158530 316271 158586 316327
rect 158230 314873 158286 314929
rect 158530 314873 158586 314929
rect 158178 307070 158234 307126
rect 158302 307070 158358 307126
rect 158426 307070 158482 307126
rect 158550 307070 158606 307126
rect 158178 306946 158234 307002
rect 158302 306946 158358 307002
rect 158426 306946 158482 307002
rect 158550 306946 158606 307002
rect 158178 306822 158234 306878
rect 158302 306822 158358 306878
rect 158426 306822 158482 306878
rect 158550 306822 158606 306878
rect 158178 306698 158234 306754
rect 158302 306698 158358 306754
rect 158426 306698 158482 306754
rect 158550 306698 158606 306754
rect 158178 306574 158234 306630
rect 158302 306574 158358 306630
rect 158426 306574 158482 306630
rect 158550 306574 158606 306630
rect 158178 306450 158234 306506
rect 158302 306450 158358 306506
rect 158426 306450 158482 306506
rect 158550 306450 158606 306506
rect 158178 306326 158234 306382
rect 158302 306326 158358 306382
rect 158426 306326 158482 306382
rect 158550 306326 158606 306382
rect 394207 330832 394263 330888
rect 394407 330832 394463 330888
rect 394207 330532 394263 330588
rect 394407 330532 394463 330588
rect 394207 330232 394263 330288
rect 394407 330232 394463 330288
rect 381382 317671 381438 317727
rect 381682 317671 381738 317727
rect 381382 316273 381438 316329
rect 381682 316273 381738 316329
rect 381382 314875 381438 314931
rect 381682 314875 381738 314931
rect 381310 307070 381366 307126
rect 381434 307070 381490 307126
rect 381558 307070 381614 307126
rect 381682 307070 381738 307126
rect 381310 306946 381366 307002
rect 381434 306946 381490 307002
rect 381558 306946 381614 307002
rect 381682 306946 381738 307002
rect 381310 306822 381366 306878
rect 381434 306822 381490 306878
rect 381558 306822 381614 306878
rect 381682 306822 381738 306878
rect 381310 306698 381366 306754
rect 381434 306698 381490 306754
rect 381558 306698 381614 306754
rect 381682 306698 381738 306754
rect 381310 306574 381366 306630
rect 381434 306574 381490 306630
rect 381558 306574 381614 306630
rect 381682 306574 381738 306630
rect 381310 306450 381366 306506
rect 381434 306450 381490 306506
rect 381558 306450 381614 306506
rect 381682 306450 381738 306506
rect 381310 306326 381366 306382
rect 381434 306326 381490 306382
rect 381558 306326 381614 306382
rect 381682 306326 381738 306382
rect 382330 329584 382386 329640
rect 382454 329584 382510 329640
rect 382578 329584 382634 329640
rect 382702 329584 382758 329640
rect 382330 329460 382386 329516
rect 382454 329460 382510 329516
rect 382578 329460 382634 329516
rect 382702 329460 382758 329516
rect 382330 329336 382386 329392
rect 382454 329336 382510 329392
rect 382578 329336 382634 329392
rect 382702 329336 382758 329392
rect 382330 329212 382386 329268
rect 382454 329212 382510 329268
rect 382578 329212 382634 329268
rect 382702 329212 382758 329268
rect 382330 329088 382386 329144
rect 382454 329088 382510 329144
rect 382578 329088 382634 329144
rect 382702 329088 382758 329144
rect 382330 328964 382386 329020
rect 382454 328964 382510 329020
rect 382578 328964 382634 329020
rect 382702 328964 382758 329020
rect 382330 328840 382386 328896
rect 382454 328840 382510 328896
rect 382578 328840 382634 328896
rect 382702 328840 382758 328896
rect 430207 330832 430263 330888
rect 430407 330832 430463 330888
rect 430207 330532 430263 330588
rect 430407 330532 430463 330588
rect 430207 330232 430263 330288
rect 430407 330232 430463 330288
rect 412207 329432 412263 329488
rect 412407 329432 412463 329488
rect 412207 329132 412263 329188
rect 412407 329132 412463 329188
rect 412207 328832 412263 328888
rect 412407 328832 412463 328888
rect 466207 330832 466263 330888
rect 466407 330832 466463 330888
rect 466207 330532 466263 330588
rect 466407 330532 466463 330588
rect 466207 330232 466263 330288
rect 466407 330232 466463 330288
rect 448207 329432 448263 329488
rect 448407 329432 448463 329488
rect 448207 329132 448263 329188
rect 448407 329132 448463 329188
rect 448207 328832 448263 328888
rect 448407 328832 448463 328888
rect 502207 330832 502263 330888
rect 502407 330832 502463 330888
rect 502207 330532 502263 330588
rect 502407 330532 502463 330588
rect 502207 330232 502263 330288
rect 502407 330232 502463 330288
rect 484207 329432 484263 329488
rect 484407 329432 484463 329488
rect 484207 329132 484263 329188
rect 484407 329132 484463 329188
rect 484207 328832 484263 328888
rect 484407 328832 484463 328888
rect 538207 330832 538263 330888
rect 538407 330832 538463 330888
rect 538207 330532 538263 330588
rect 538407 330532 538463 330588
rect 538207 330232 538263 330288
rect 538407 330232 538463 330288
rect 520207 329432 520263 329488
rect 520407 329432 520463 329488
rect 520207 329132 520263 329188
rect 520407 329132 520463 329188
rect 520207 328832 520263 328888
rect 520407 328832 520463 328888
rect 574207 330832 574263 330888
rect 574407 330832 574463 330888
rect 574207 330532 574263 330588
rect 574407 330532 574463 330588
rect 574207 330232 574263 330288
rect 574407 330232 574463 330288
rect 556207 329432 556263 329488
rect 556407 329432 556463 329488
rect 556207 329132 556263 329188
rect 556407 329132 556463 329188
rect 556207 328832 556263 328888
rect 556407 328832 556463 328888
rect 610207 330832 610263 330888
rect 610407 330832 610463 330888
rect 610207 330532 610263 330588
rect 610407 330532 610463 330588
rect 610207 330232 610263 330288
rect 610407 330232 610463 330288
rect 592207 329432 592263 329488
rect 592407 329432 592463 329488
rect 592207 329132 592263 329188
rect 592407 329132 592463 329188
rect 592207 328832 592263 328888
rect 592407 328832 592463 328888
rect 646207 330832 646263 330888
rect 646407 330832 646463 330888
rect 646207 330532 646263 330588
rect 646407 330532 646463 330588
rect 646207 330232 646263 330288
rect 646407 330232 646463 330288
rect 628207 329432 628263 329488
rect 628407 329432 628463 329488
rect 628207 329132 628263 329188
rect 628407 329132 628463 329188
rect 628207 328832 628263 328888
rect 628407 328832 628463 328888
rect 682207 330832 682263 330888
rect 682407 330832 682463 330888
rect 682207 330532 682263 330588
rect 682407 330532 682463 330588
rect 682207 330232 682263 330288
rect 682407 330232 682463 330288
rect 698060 332952 698116 333008
rect 698360 332952 698416 333008
rect 698660 332952 698716 333008
rect 698052 330984 698108 331040
rect 698176 330984 698232 331040
rect 698300 330984 698356 331040
rect 698424 330984 698480 331040
rect 698548 330984 698604 331040
rect 698672 330984 698728 331040
rect 698796 330984 698852 331040
rect 698052 330860 698108 330916
rect 698176 330860 698232 330916
rect 698300 330860 698356 330916
rect 698424 330860 698480 330916
rect 698548 330860 698604 330916
rect 698672 330860 698728 330916
rect 698796 330860 698852 330916
rect 698052 330736 698108 330792
rect 698176 330736 698232 330792
rect 698300 330736 698356 330792
rect 698424 330736 698480 330792
rect 698548 330736 698604 330792
rect 698672 330736 698728 330792
rect 698796 330736 698852 330792
rect 698052 330612 698108 330668
rect 698176 330612 698232 330668
rect 698300 330612 698356 330668
rect 698424 330612 698480 330668
rect 698548 330612 698604 330668
rect 698672 330612 698728 330668
rect 698796 330612 698852 330668
rect 698052 330488 698108 330544
rect 698176 330488 698232 330544
rect 698300 330488 698356 330544
rect 698424 330488 698480 330544
rect 698548 330488 698604 330544
rect 698672 330488 698728 330544
rect 698796 330488 698852 330544
rect 698052 330364 698108 330420
rect 698176 330364 698232 330420
rect 698300 330364 698356 330420
rect 698424 330364 698480 330420
rect 698548 330364 698604 330420
rect 698672 330364 698728 330420
rect 698796 330364 698852 330420
rect 698052 330240 698108 330296
rect 698176 330240 698232 330296
rect 698300 330240 698356 330296
rect 698424 330240 698480 330296
rect 698548 330240 698604 330296
rect 698672 330240 698728 330296
rect 698796 330240 698852 330296
rect 664207 329432 664263 329488
rect 664407 329432 664463 329488
rect 664207 329132 664263 329188
rect 664407 329132 664463 329188
rect 664207 328832 664263 328888
rect 664407 328832 664463 328888
rect 382402 318370 382458 318426
rect 382702 318370 382758 318426
rect 382402 316972 382458 317028
rect 382702 316972 382758 317028
rect 382402 315574 382458 315630
rect 382702 315574 382758 315630
rect 698044 320378 698100 320434
rect 698344 320378 698400 320434
rect 698644 320378 698700 320434
rect 382402 314176 382458 314232
rect 382702 314176 382758 314232
rect 157158 305670 157214 305726
rect 157282 305670 157338 305726
rect 157406 305670 157462 305726
rect 157530 305670 157586 305726
rect 157158 305546 157214 305602
rect 157282 305546 157338 305602
rect 157406 305546 157462 305602
rect 157530 305546 157586 305602
rect 157158 305422 157214 305478
rect 157282 305422 157338 305478
rect 157406 305422 157462 305478
rect 157530 305422 157586 305478
rect 157158 305298 157214 305354
rect 157282 305298 157338 305354
rect 157406 305298 157462 305354
rect 157530 305298 157586 305354
rect 157158 305174 157214 305230
rect 157282 305174 157338 305230
rect 157406 305174 157462 305230
rect 157530 305174 157586 305230
rect 157158 305050 157214 305106
rect 157282 305050 157338 305106
rect 157406 305050 157462 305106
rect 157530 305050 157586 305106
rect 157158 304926 157214 304982
rect 157282 304926 157338 304982
rect 157406 304926 157462 304982
rect 157530 304926 157586 304982
rect 382330 305670 382386 305726
rect 382454 305670 382510 305726
rect 382578 305670 382634 305726
rect 382702 305670 382758 305726
rect 382330 305546 382386 305602
rect 382454 305546 382510 305602
rect 382578 305546 382634 305602
rect 382702 305546 382758 305602
rect 382330 305422 382386 305478
rect 382454 305422 382510 305478
rect 382578 305422 382634 305478
rect 382702 305422 382758 305478
rect 382330 305298 382386 305354
rect 382454 305298 382510 305354
rect 382578 305298 382634 305354
rect 382702 305298 382758 305354
rect 382330 305174 382386 305230
rect 382454 305174 382510 305230
rect 382578 305174 382634 305230
rect 382702 305174 382758 305230
rect 382330 305050 382386 305106
rect 382454 305050 382510 305106
rect 382578 305050 382634 305106
rect 382702 305050 382758 305106
rect 382330 304926 382386 304982
rect 382454 304926 382510 304982
rect 382578 304926 382634 304982
rect 382702 304926 382758 304982
rect 390220 307130 390276 307186
rect 390344 307130 390400 307186
rect 390220 307006 390276 307062
rect 390344 307006 390400 307062
rect 390220 306882 390276 306938
rect 390344 306882 390400 306938
rect 390220 306758 390276 306814
rect 390344 306758 390400 306814
rect 390220 306634 390276 306690
rect 390344 306634 390400 306690
rect 390220 306510 390276 306566
rect 390344 306510 390400 306566
rect 390220 306386 390276 306442
rect 390344 306386 390400 306442
rect 388625 305730 388681 305786
rect 388749 305730 388805 305786
rect 388625 305606 388681 305662
rect 388749 305606 388805 305662
rect 388625 305482 388681 305538
rect 388749 305482 388805 305538
rect 388625 305358 388681 305414
rect 388749 305358 388805 305414
rect 388625 305234 388681 305290
rect 388749 305234 388805 305290
rect 388625 305110 388681 305166
rect 388749 305110 388805 305166
rect 388625 304986 388681 305042
rect 388749 304986 388805 305042
rect 393410 307130 393466 307186
rect 393534 307130 393590 307186
rect 393410 307006 393466 307062
rect 393534 307006 393590 307062
rect 393410 306882 393466 306938
rect 393534 306882 393590 306938
rect 393410 306758 393466 306814
rect 393534 306758 393590 306814
rect 393410 306634 393466 306690
rect 393534 306634 393590 306690
rect 393410 306510 393466 306566
rect 393534 306510 393590 306566
rect 393410 306386 393466 306442
rect 393534 306386 393590 306442
rect 391815 305730 391871 305786
rect 391939 305730 391995 305786
rect 391815 305606 391871 305662
rect 391939 305606 391995 305662
rect 391815 305482 391871 305538
rect 391939 305482 391995 305538
rect 391815 305358 391871 305414
rect 391939 305358 391995 305414
rect 391815 305234 391871 305290
rect 391939 305234 391995 305290
rect 391815 305110 391871 305166
rect 391939 305110 391995 305166
rect 391815 304986 391871 305042
rect 391939 304986 391995 305042
rect 396600 307130 396656 307186
rect 396724 307130 396780 307186
rect 396600 307006 396656 307062
rect 396724 307006 396780 307062
rect 396600 306882 396656 306938
rect 396724 306882 396780 306938
rect 396600 306758 396656 306814
rect 396724 306758 396780 306814
rect 396600 306634 396656 306690
rect 396724 306634 396780 306690
rect 396600 306510 396656 306566
rect 396724 306510 396780 306566
rect 396600 306386 396656 306442
rect 396724 306386 396780 306442
rect 395005 305730 395061 305786
rect 395129 305730 395185 305786
rect 395005 305606 395061 305662
rect 395129 305606 395185 305662
rect 395005 305482 395061 305538
rect 395129 305482 395185 305538
rect 395005 305358 395061 305414
rect 395129 305358 395185 305414
rect 395005 305234 395061 305290
rect 395129 305234 395185 305290
rect 395005 305110 395061 305166
rect 395129 305110 395185 305166
rect 395005 304986 395061 305042
rect 395129 304986 395185 305042
rect 398195 305730 398251 305786
rect 398319 305730 398375 305786
rect 398195 305606 398251 305662
rect 398319 305606 398375 305662
rect 398195 305482 398251 305538
rect 398319 305482 398375 305538
rect 398195 305358 398251 305414
rect 398319 305358 398375 305414
rect 398195 305234 398251 305290
rect 398319 305234 398375 305290
rect 398195 305110 398251 305166
rect 398319 305110 398375 305166
rect 398195 304986 398251 305042
rect 398319 304986 398375 305042
rect 490220 307130 490276 307186
rect 490344 307130 490400 307186
rect 490220 307006 490276 307062
rect 490344 307006 490400 307062
rect 490220 306882 490276 306938
rect 490344 306882 490400 306938
rect 490220 306758 490276 306814
rect 490344 306758 490400 306814
rect 490220 306634 490276 306690
rect 490344 306634 490400 306690
rect 490220 306510 490276 306566
rect 490344 306510 490400 306566
rect 490220 306386 490276 306442
rect 490344 306386 490400 306442
rect 488625 305730 488681 305786
rect 488749 305730 488805 305786
rect 488625 305606 488681 305662
rect 488749 305606 488805 305662
rect 488625 305482 488681 305538
rect 488749 305482 488805 305538
rect 488625 305358 488681 305414
rect 488749 305358 488805 305414
rect 488625 305234 488681 305290
rect 488749 305234 488805 305290
rect 488625 305110 488681 305166
rect 488749 305110 488805 305166
rect 488625 304986 488681 305042
rect 488749 304986 488805 305042
rect 493410 307130 493466 307186
rect 493534 307130 493590 307186
rect 493410 307006 493466 307062
rect 493534 307006 493590 307062
rect 493410 306882 493466 306938
rect 493534 306882 493590 306938
rect 493410 306758 493466 306814
rect 493534 306758 493590 306814
rect 493410 306634 493466 306690
rect 493534 306634 493590 306690
rect 493410 306510 493466 306566
rect 493534 306510 493590 306566
rect 493410 306386 493466 306442
rect 493534 306386 493590 306442
rect 491815 305730 491871 305786
rect 491939 305730 491995 305786
rect 491815 305606 491871 305662
rect 491939 305606 491995 305662
rect 491815 305482 491871 305538
rect 491939 305482 491995 305538
rect 491815 305358 491871 305414
rect 491939 305358 491995 305414
rect 491815 305234 491871 305290
rect 491939 305234 491995 305290
rect 491815 305110 491871 305166
rect 491939 305110 491995 305166
rect 491815 304986 491871 305042
rect 491939 304986 491995 305042
rect 496600 307130 496656 307186
rect 496724 307130 496780 307186
rect 496600 307006 496656 307062
rect 496724 307006 496780 307062
rect 496600 306882 496656 306938
rect 496724 306882 496780 306938
rect 496600 306758 496656 306814
rect 496724 306758 496780 306814
rect 496600 306634 496656 306690
rect 496724 306634 496780 306690
rect 496600 306510 496656 306566
rect 496724 306510 496780 306566
rect 496600 306386 496656 306442
rect 496724 306386 496780 306442
rect 495005 305730 495061 305786
rect 495129 305730 495185 305786
rect 495005 305606 495061 305662
rect 495129 305606 495185 305662
rect 495005 305482 495061 305538
rect 495129 305482 495185 305538
rect 495005 305358 495061 305414
rect 495129 305358 495185 305414
rect 495005 305234 495061 305290
rect 495129 305234 495185 305290
rect 495005 305110 495061 305166
rect 495129 305110 495185 305166
rect 495005 304986 495061 305042
rect 495129 304986 495185 305042
rect 498195 305730 498251 305786
rect 498319 305730 498375 305786
rect 498195 305606 498251 305662
rect 498319 305606 498375 305662
rect 498195 305482 498251 305538
rect 498319 305482 498375 305538
rect 498195 305358 498251 305414
rect 498319 305358 498375 305414
rect 498195 305234 498251 305290
rect 498319 305234 498375 305290
rect 498195 305110 498251 305166
rect 498319 305110 498375 305166
rect 498195 304986 498251 305042
rect 498319 304986 498375 305042
rect 590910 307070 590966 307126
rect 591034 307070 591090 307126
rect 591158 307070 591214 307126
rect 591282 307070 591338 307126
rect 591406 307070 591462 307126
rect 591530 307070 591586 307126
rect 591654 307070 591710 307126
rect 590910 306946 590966 307002
rect 591034 306946 591090 307002
rect 591158 306946 591214 307002
rect 591282 306946 591338 307002
rect 591406 306946 591462 307002
rect 591530 306946 591586 307002
rect 591654 306946 591710 307002
rect 590910 306822 590966 306878
rect 591034 306822 591090 306878
rect 591158 306822 591214 306878
rect 591282 306822 591338 306878
rect 591406 306822 591462 306878
rect 591530 306822 591586 306878
rect 591654 306822 591710 306878
rect 590910 306698 590966 306754
rect 591034 306698 591090 306754
rect 591158 306698 591214 306754
rect 591282 306698 591338 306754
rect 591406 306698 591462 306754
rect 591530 306698 591586 306754
rect 591654 306698 591710 306754
rect 590910 306574 590966 306630
rect 591034 306574 591090 306630
rect 591158 306574 591214 306630
rect 591282 306574 591338 306630
rect 591406 306574 591462 306630
rect 591530 306574 591586 306630
rect 591654 306574 591710 306630
rect 590910 306450 590966 306506
rect 591034 306450 591090 306506
rect 591158 306450 591214 306506
rect 591282 306450 591338 306506
rect 591406 306450 591462 306506
rect 591530 306450 591586 306506
rect 591654 306450 591710 306506
rect 590910 306326 590966 306382
rect 591034 306326 591090 306382
rect 591158 306326 591214 306382
rect 591282 306326 591338 306382
rect 591406 306326 591462 306382
rect 591530 306326 591586 306382
rect 591654 306326 591710 306382
rect 79300 300566 79356 300622
rect 79600 300566 79656 300622
rect 79900 300566 79956 300622
rect 79284 289992 79340 290048
rect 79584 289992 79640 290048
rect 79884 289992 79940 290048
rect 79208 283316 79264 283372
rect 79332 283316 79388 283372
rect 79456 283316 79512 283372
rect 79580 283316 79636 283372
rect 79704 283316 79760 283372
rect 79828 283316 79884 283372
rect 79952 283316 80008 283372
rect 79208 283192 79264 283248
rect 79332 283192 79388 283248
rect 79456 283192 79512 283248
rect 79580 283192 79636 283248
rect 79704 283192 79760 283248
rect 79828 283192 79884 283248
rect 79952 283192 80008 283248
rect 79208 283068 79264 283124
rect 79332 283068 79388 283124
rect 79456 283068 79512 283124
rect 79580 283068 79636 283124
rect 79704 283068 79760 283124
rect 79828 283068 79884 283124
rect 79952 283068 80008 283124
rect 79208 282944 79264 283000
rect 79332 282944 79388 283000
rect 79456 282944 79512 283000
rect 79580 282944 79636 283000
rect 79704 282944 79760 283000
rect 79828 282944 79884 283000
rect 79952 282944 80008 283000
rect 79208 282820 79264 282876
rect 79332 282820 79388 282876
rect 79456 282820 79512 282876
rect 79580 282820 79636 282876
rect 79704 282820 79760 282876
rect 79828 282820 79884 282876
rect 79952 282820 80008 282876
rect 79208 282696 79264 282752
rect 79332 282696 79388 282752
rect 79456 282696 79512 282752
rect 79580 282696 79636 282752
rect 79704 282696 79760 282752
rect 79828 282696 79884 282752
rect 79952 282696 80008 282752
rect 79208 282572 79264 282628
rect 79332 282572 79388 282628
rect 79456 282572 79512 282628
rect 79580 282572 79636 282628
rect 79704 282572 79760 282628
rect 79828 282572 79884 282628
rect 79952 282572 80008 282628
rect 99294 283256 99350 283312
rect 99418 283256 99474 283312
rect 99294 283132 99350 283188
rect 99418 283132 99474 283188
rect 99294 283008 99350 283064
rect 99418 283008 99474 283064
rect 99294 282884 99350 282940
rect 99418 282884 99474 282940
rect 99294 282760 99350 282816
rect 99418 282760 99474 282816
rect 99294 282636 99350 282692
rect 99418 282636 99474 282692
rect 99294 282512 99350 282568
rect 99418 282512 99474 282568
rect 94294 281856 94350 281912
rect 94418 281856 94474 281912
rect 94294 281732 94350 281788
rect 94418 281732 94474 281788
rect 94294 281608 94350 281664
rect 94418 281608 94474 281664
rect 94294 281484 94350 281540
rect 94418 281484 94474 281540
rect 94294 281360 94350 281416
rect 94418 281360 94474 281416
rect 94294 281236 94350 281292
rect 94418 281236 94474 281292
rect 94294 281112 94350 281168
rect 94418 281112 94474 281168
rect 109294 283256 109350 283312
rect 109418 283256 109474 283312
rect 109294 283132 109350 283188
rect 109418 283132 109474 283188
rect 109294 283008 109350 283064
rect 109418 283008 109474 283064
rect 109294 282884 109350 282940
rect 109418 282884 109474 282940
rect 109294 282760 109350 282816
rect 109418 282760 109474 282816
rect 109294 282636 109350 282692
rect 109418 282636 109474 282692
rect 109294 282512 109350 282568
rect 109418 282512 109474 282568
rect 104294 281856 104350 281912
rect 104418 281856 104474 281912
rect 104294 281732 104350 281788
rect 104418 281732 104474 281788
rect 104294 281608 104350 281664
rect 104418 281608 104474 281664
rect 104294 281484 104350 281540
rect 104418 281484 104474 281540
rect 104294 281360 104350 281416
rect 104418 281360 104474 281416
rect 104294 281236 104350 281292
rect 104418 281236 104474 281292
rect 104294 281112 104350 281168
rect 104418 281112 104474 281168
rect 119294 283256 119350 283312
rect 119418 283256 119474 283312
rect 119294 283132 119350 283188
rect 119418 283132 119474 283188
rect 119294 283008 119350 283064
rect 119418 283008 119474 283064
rect 119294 282884 119350 282940
rect 119418 282884 119474 282940
rect 119294 282760 119350 282816
rect 119418 282760 119474 282816
rect 119294 282636 119350 282692
rect 119418 282636 119474 282692
rect 119294 282512 119350 282568
rect 119418 282512 119474 282568
rect 114294 281856 114350 281912
rect 114418 281856 114474 281912
rect 114294 281732 114350 281788
rect 114418 281732 114474 281788
rect 114294 281608 114350 281664
rect 114418 281608 114474 281664
rect 114294 281484 114350 281540
rect 114418 281484 114474 281540
rect 114294 281360 114350 281416
rect 114418 281360 114474 281416
rect 114294 281236 114350 281292
rect 114418 281236 114474 281292
rect 114294 281112 114350 281168
rect 114418 281112 114474 281168
rect 129294 283256 129350 283312
rect 129418 283256 129474 283312
rect 129294 283132 129350 283188
rect 129418 283132 129474 283188
rect 129294 283008 129350 283064
rect 129418 283008 129474 283064
rect 129294 282884 129350 282940
rect 129418 282884 129474 282940
rect 129294 282760 129350 282816
rect 129418 282760 129474 282816
rect 129294 282636 129350 282692
rect 129418 282636 129474 282692
rect 129294 282512 129350 282568
rect 129418 282512 129474 282568
rect 124294 281856 124350 281912
rect 124418 281856 124474 281912
rect 124294 281732 124350 281788
rect 124418 281732 124474 281788
rect 124294 281608 124350 281664
rect 124418 281608 124474 281664
rect 124294 281484 124350 281540
rect 124418 281484 124474 281540
rect 124294 281360 124350 281416
rect 124418 281360 124474 281416
rect 124294 281236 124350 281292
rect 124418 281236 124474 281292
rect 124294 281112 124350 281168
rect 124418 281112 124474 281168
rect 139294 283256 139350 283312
rect 139418 283256 139474 283312
rect 139294 283132 139350 283188
rect 139418 283132 139474 283188
rect 139294 283008 139350 283064
rect 139418 283008 139474 283064
rect 139294 282884 139350 282940
rect 139418 282884 139474 282940
rect 139294 282760 139350 282816
rect 139418 282760 139474 282816
rect 139294 282636 139350 282692
rect 139418 282636 139474 282692
rect 139294 282512 139350 282568
rect 139418 282512 139474 282568
rect 134294 281856 134350 281912
rect 134418 281856 134474 281912
rect 134294 281732 134350 281788
rect 134418 281732 134474 281788
rect 134294 281608 134350 281664
rect 134418 281608 134474 281664
rect 134294 281484 134350 281540
rect 134418 281484 134474 281540
rect 134294 281360 134350 281416
rect 134418 281360 134474 281416
rect 134294 281236 134350 281292
rect 134418 281236 134474 281292
rect 134294 281112 134350 281168
rect 134418 281112 134474 281168
rect 149294 283256 149350 283312
rect 149418 283256 149474 283312
rect 149294 283132 149350 283188
rect 149418 283132 149474 283188
rect 149294 283008 149350 283064
rect 149418 283008 149474 283064
rect 149294 282884 149350 282940
rect 149418 282884 149474 282940
rect 149294 282760 149350 282816
rect 149418 282760 149474 282816
rect 149294 282636 149350 282692
rect 149418 282636 149474 282692
rect 149294 282512 149350 282568
rect 149418 282512 149474 282568
rect 144294 281856 144350 281912
rect 144418 281856 144474 281912
rect 144294 281732 144350 281788
rect 144418 281732 144474 281788
rect 144294 281608 144350 281664
rect 144418 281608 144474 281664
rect 144294 281484 144350 281540
rect 144418 281484 144474 281540
rect 144294 281360 144350 281416
rect 144418 281360 144474 281416
rect 144294 281236 144350 281292
rect 144418 281236 144474 281292
rect 144294 281112 144350 281168
rect 144418 281112 144474 281168
rect 159294 283256 159350 283312
rect 159418 283256 159474 283312
rect 159294 283132 159350 283188
rect 159418 283132 159474 283188
rect 159294 283008 159350 283064
rect 159418 283008 159474 283064
rect 159294 282884 159350 282940
rect 159418 282884 159474 282940
rect 159294 282760 159350 282816
rect 159418 282760 159474 282816
rect 159294 282636 159350 282692
rect 159418 282636 159474 282692
rect 159294 282512 159350 282568
rect 159418 282512 159474 282568
rect 154294 281856 154350 281912
rect 154418 281856 154474 281912
rect 154294 281732 154350 281788
rect 154418 281732 154474 281788
rect 154294 281608 154350 281664
rect 154418 281608 154474 281664
rect 154294 281484 154350 281540
rect 154418 281484 154474 281540
rect 154294 281360 154350 281416
rect 154418 281360 154474 281416
rect 154294 281236 154350 281292
rect 154418 281236 154474 281292
rect 154294 281112 154350 281168
rect 154418 281112 154474 281168
rect 169294 283256 169350 283312
rect 169418 283256 169474 283312
rect 169294 283132 169350 283188
rect 169418 283132 169474 283188
rect 169294 283008 169350 283064
rect 169418 283008 169474 283064
rect 169294 282884 169350 282940
rect 169418 282884 169474 282940
rect 169294 282760 169350 282816
rect 169418 282760 169474 282816
rect 169294 282636 169350 282692
rect 169418 282636 169474 282692
rect 169294 282512 169350 282568
rect 169418 282512 169474 282568
rect 164294 281856 164350 281912
rect 164418 281856 164474 281912
rect 164294 281732 164350 281788
rect 164418 281732 164474 281788
rect 164294 281608 164350 281664
rect 164418 281608 164474 281664
rect 164294 281484 164350 281540
rect 164418 281484 164474 281540
rect 164294 281360 164350 281416
rect 164418 281360 164474 281416
rect 164294 281236 164350 281292
rect 164418 281236 164474 281292
rect 164294 281112 164350 281168
rect 164418 281112 164474 281168
rect 179294 283256 179350 283312
rect 179418 283256 179474 283312
rect 179294 283132 179350 283188
rect 179418 283132 179474 283188
rect 179294 283008 179350 283064
rect 179418 283008 179474 283064
rect 179294 282884 179350 282940
rect 179418 282884 179474 282940
rect 179294 282760 179350 282816
rect 179418 282760 179474 282816
rect 179294 282636 179350 282692
rect 179418 282636 179474 282692
rect 179294 282512 179350 282568
rect 179418 282512 179474 282568
rect 174294 281856 174350 281912
rect 174418 281856 174474 281912
rect 174294 281732 174350 281788
rect 174418 281732 174474 281788
rect 174294 281608 174350 281664
rect 174418 281608 174474 281664
rect 174294 281484 174350 281540
rect 174418 281484 174474 281540
rect 174294 281360 174350 281416
rect 174418 281360 174474 281416
rect 174294 281236 174350 281292
rect 174418 281236 174474 281292
rect 174294 281112 174350 281168
rect 174418 281112 174474 281168
rect 189294 283256 189350 283312
rect 189418 283256 189474 283312
rect 189294 283132 189350 283188
rect 189418 283132 189474 283188
rect 189294 283008 189350 283064
rect 189418 283008 189474 283064
rect 189294 282884 189350 282940
rect 189418 282884 189474 282940
rect 189294 282760 189350 282816
rect 189418 282760 189474 282816
rect 189294 282636 189350 282692
rect 189418 282636 189474 282692
rect 189294 282512 189350 282568
rect 189418 282512 189474 282568
rect 184294 281856 184350 281912
rect 184418 281856 184474 281912
rect 184294 281732 184350 281788
rect 184418 281732 184474 281788
rect 184294 281608 184350 281664
rect 184418 281608 184474 281664
rect 184294 281484 184350 281540
rect 184418 281484 184474 281540
rect 184294 281360 184350 281416
rect 184418 281360 184474 281416
rect 184294 281236 184350 281292
rect 184418 281236 184474 281292
rect 184294 281112 184350 281168
rect 184418 281112 184474 281168
rect 199294 283256 199350 283312
rect 199418 283256 199474 283312
rect 199294 283132 199350 283188
rect 199418 283132 199474 283188
rect 199294 283008 199350 283064
rect 199418 283008 199474 283064
rect 199294 282884 199350 282940
rect 199418 282884 199474 282940
rect 199294 282760 199350 282816
rect 199418 282760 199474 282816
rect 199294 282636 199350 282692
rect 199418 282636 199474 282692
rect 199294 282512 199350 282568
rect 199418 282512 199474 282568
rect 194294 281856 194350 281912
rect 194418 281856 194474 281912
rect 194294 281732 194350 281788
rect 194418 281732 194474 281788
rect 194294 281608 194350 281664
rect 194418 281608 194474 281664
rect 194294 281484 194350 281540
rect 194418 281484 194474 281540
rect 194294 281360 194350 281416
rect 194418 281360 194474 281416
rect 194294 281236 194350 281292
rect 194418 281236 194474 281292
rect 194294 281112 194350 281168
rect 194418 281112 194474 281168
rect 209294 283256 209350 283312
rect 209418 283256 209474 283312
rect 209294 283132 209350 283188
rect 209418 283132 209474 283188
rect 209294 283008 209350 283064
rect 209418 283008 209474 283064
rect 209294 282884 209350 282940
rect 209418 282884 209474 282940
rect 209294 282760 209350 282816
rect 209418 282760 209474 282816
rect 209294 282636 209350 282692
rect 209418 282636 209474 282692
rect 209294 282512 209350 282568
rect 209418 282512 209474 282568
rect 204294 281856 204350 281912
rect 204418 281856 204474 281912
rect 204294 281732 204350 281788
rect 204418 281732 204474 281788
rect 204294 281608 204350 281664
rect 204418 281608 204474 281664
rect 204294 281484 204350 281540
rect 204418 281484 204474 281540
rect 204294 281360 204350 281416
rect 204418 281360 204474 281416
rect 204294 281236 204350 281292
rect 204418 281236 204474 281292
rect 204294 281112 204350 281168
rect 204418 281112 204474 281168
rect 219294 283256 219350 283312
rect 219418 283256 219474 283312
rect 219294 283132 219350 283188
rect 219418 283132 219474 283188
rect 219294 283008 219350 283064
rect 219418 283008 219474 283064
rect 219294 282884 219350 282940
rect 219418 282884 219474 282940
rect 219294 282760 219350 282816
rect 219418 282760 219474 282816
rect 219294 282636 219350 282692
rect 219418 282636 219474 282692
rect 219294 282512 219350 282568
rect 219418 282512 219474 282568
rect 214294 281856 214350 281912
rect 214418 281856 214474 281912
rect 214294 281732 214350 281788
rect 214418 281732 214474 281788
rect 214294 281608 214350 281664
rect 214418 281608 214474 281664
rect 214294 281484 214350 281540
rect 214418 281484 214474 281540
rect 214294 281360 214350 281416
rect 214418 281360 214474 281416
rect 214294 281236 214350 281292
rect 214418 281236 214474 281292
rect 214294 281112 214350 281168
rect 214418 281112 214474 281168
rect 229294 283256 229350 283312
rect 229418 283256 229474 283312
rect 229294 283132 229350 283188
rect 229418 283132 229474 283188
rect 229294 283008 229350 283064
rect 229418 283008 229474 283064
rect 229294 282884 229350 282940
rect 229418 282884 229474 282940
rect 229294 282760 229350 282816
rect 229418 282760 229474 282816
rect 229294 282636 229350 282692
rect 229418 282636 229474 282692
rect 229294 282512 229350 282568
rect 229418 282512 229474 282568
rect 224294 281856 224350 281912
rect 224418 281856 224474 281912
rect 224294 281732 224350 281788
rect 224418 281732 224474 281788
rect 224294 281608 224350 281664
rect 224418 281608 224474 281664
rect 224294 281484 224350 281540
rect 224418 281484 224474 281540
rect 224294 281360 224350 281416
rect 224418 281360 224474 281416
rect 224294 281236 224350 281292
rect 224418 281236 224474 281292
rect 224294 281112 224350 281168
rect 224418 281112 224474 281168
rect 239294 283256 239350 283312
rect 239418 283256 239474 283312
rect 239294 283132 239350 283188
rect 239418 283132 239474 283188
rect 239294 283008 239350 283064
rect 239418 283008 239474 283064
rect 239294 282884 239350 282940
rect 239418 282884 239474 282940
rect 239294 282760 239350 282816
rect 239418 282760 239474 282816
rect 239294 282636 239350 282692
rect 239418 282636 239474 282692
rect 239294 282512 239350 282568
rect 239418 282512 239474 282568
rect 234294 281856 234350 281912
rect 234418 281856 234474 281912
rect 234294 281732 234350 281788
rect 234418 281732 234474 281788
rect 234294 281608 234350 281664
rect 234418 281608 234474 281664
rect 234294 281484 234350 281540
rect 234418 281484 234474 281540
rect 234294 281360 234350 281416
rect 234418 281360 234474 281416
rect 234294 281236 234350 281292
rect 234418 281236 234474 281292
rect 234294 281112 234350 281168
rect 234418 281112 234474 281168
rect 249294 283256 249350 283312
rect 249418 283256 249474 283312
rect 249294 283132 249350 283188
rect 249418 283132 249474 283188
rect 249294 283008 249350 283064
rect 249418 283008 249474 283064
rect 249294 282884 249350 282940
rect 249418 282884 249474 282940
rect 249294 282760 249350 282816
rect 249418 282760 249474 282816
rect 249294 282636 249350 282692
rect 249418 282636 249474 282692
rect 249294 282512 249350 282568
rect 249418 282512 249474 282568
rect 244294 281856 244350 281912
rect 244418 281856 244474 281912
rect 244294 281732 244350 281788
rect 244418 281732 244474 281788
rect 244294 281608 244350 281664
rect 244418 281608 244474 281664
rect 244294 281484 244350 281540
rect 244418 281484 244474 281540
rect 244294 281360 244350 281416
rect 244418 281360 244474 281416
rect 244294 281236 244350 281292
rect 244418 281236 244474 281292
rect 244294 281112 244350 281168
rect 244418 281112 244474 281168
rect 259294 283256 259350 283312
rect 259418 283256 259474 283312
rect 259294 283132 259350 283188
rect 259418 283132 259474 283188
rect 259294 283008 259350 283064
rect 259418 283008 259474 283064
rect 259294 282884 259350 282940
rect 259418 282884 259474 282940
rect 259294 282760 259350 282816
rect 259418 282760 259474 282816
rect 259294 282636 259350 282692
rect 259418 282636 259474 282692
rect 259294 282512 259350 282568
rect 259418 282512 259474 282568
rect 254294 281856 254350 281912
rect 254418 281856 254474 281912
rect 254294 281732 254350 281788
rect 254418 281732 254474 281788
rect 254294 281608 254350 281664
rect 254418 281608 254474 281664
rect 254294 281484 254350 281540
rect 254418 281484 254474 281540
rect 254294 281360 254350 281416
rect 254418 281360 254474 281416
rect 254294 281236 254350 281292
rect 254418 281236 254474 281292
rect 254294 281112 254350 281168
rect 254418 281112 254474 281168
rect 269294 283256 269350 283312
rect 269418 283256 269474 283312
rect 269294 283132 269350 283188
rect 269418 283132 269474 283188
rect 269294 283008 269350 283064
rect 269418 283008 269474 283064
rect 269294 282884 269350 282940
rect 269418 282884 269474 282940
rect 269294 282760 269350 282816
rect 269418 282760 269474 282816
rect 269294 282636 269350 282692
rect 269418 282636 269474 282692
rect 269294 282512 269350 282568
rect 269418 282512 269474 282568
rect 264294 281856 264350 281912
rect 264418 281856 264474 281912
rect 264294 281732 264350 281788
rect 264418 281732 264474 281788
rect 264294 281608 264350 281664
rect 264418 281608 264474 281664
rect 264294 281484 264350 281540
rect 264418 281484 264474 281540
rect 264294 281360 264350 281416
rect 264418 281360 264474 281416
rect 264294 281236 264350 281292
rect 264418 281236 264474 281292
rect 264294 281112 264350 281168
rect 264418 281112 264474 281168
rect 279294 283256 279350 283312
rect 279418 283256 279474 283312
rect 279294 283132 279350 283188
rect 279418 283132 279474 283188
rect 279294 283008 279350 283064
rect 279418 283008 279474 283064
rect 279294 282884 279350 282940
rect 279418 282884 279474 282940
rect 279294 282760 279350 282816
rect 279418 282760 279474 282816
rect 279294 282636 279350 282692
rect 279418 282636 279474 282692
rect 279294 282512 279350 282568
rect 279418 282512 279474 282568
rect 274294 281856 274350 281912
rect 274418 281856 274474 281912
rect 274294 281732 274350 281788
rect 274418 281732 274474 281788
rect 274294 281608 274350 281664
rect 274418 281608 274474 281664
rect 274294 281484 274350 281540
rect 274418 281484 274474 281540
rect 274294 281360 274350 281416
rect 274418 281360 274474 281416
rect 274294 281236 274350 281292
rect 274418 281236 274474 281292
rect 274294 281112 274350 281168
rect 274418 281112 274474 281168
rect 289294 283256 289350 283312
rect 289418 283256 289474 283312
rect 289294 283132 289350 283188
rect 289418 283132 289474 283188
rect 289294 283008 289350 283064
rect 289418 283008 289474 283064
rect 289294 282884 289350 282940
rect 289418 282884 289474 282940
rect 289294 282760 289350 282816
rect 289418 282760 289474 282816
rect 289294 282636 289350 282692
rect 289418 282636 289474 282692
rect 289294 282512 289350 282568
rect 289418 282512 289474 282568
rect 284294 281856 284350 281912
rect 284418 281856 284474 281912
rect 284294 281732 284350 281788
rect 284418 281732 284474 281788
rect 284294 281608 284350 281664
rect 284418 281608 284474 281664
rect 284294 281484 284350 281540
rect 284418 281484 284474 281540
rect 284294 281360 284350 281416
rect 284418 281360 284474 281416
rect 284294 281236 284350 281292
rect 284418 281236 284474 281292
rect 284294 281112 284350 281168
rect 284418 281112 284474 281168
rect 299294 283256 299350 283312
rect 299418 283256 299474 283312
rect 299294 283132 299350 283188
rect 299418 283132 299474 283188
rect 299294 283008 299350 283064
rect 299418 283008 299474 283064
rect 299294 282884 299350 282940
rect 299418 282884 299474 282940
rect 299294 282760 299350 282816
rect 299418 282760 299474 282816
rect 299294 282636 299350 282692
rect 299418 282636 299474 282692
rect 299294 282512 299350 282568
rect 299418 282512 299474 282568
rect 294294 281856 294350 281912
rect 294418 281856 294474 281912
rect 294294 281732 294350 281788
rect 294418 281732 294474 281788
rect 294294 281608 294350 281664
rect 294418 281608 294474 281664
rect 294294 281484 294350 281540
rect 294418 281484 294474 281540
rect 294294 281360 294350 281416
rect 294418 281360 294474 281416
rect 294294 281236 294350 281292
rect 294418 281236 294474 281292
rect 294294 281112 294350 281168
rect 294418 281112 294474 281168
rect 309294 283256 309350 283312
rect 309418 283256 309474 283312
rect 309294 283132 309350 283188
rect 309418 283132 309474 283188
rect 309294 283008 309350 283064
rect 309418 283008 309474 283064
rect 309294 282884 309350 282940
rect 309418 282884 309474 282940
rect 309294 282760 309350 282816
rect 309418 282760 309474 282816
rect 309294 282636 309350 282692
rect 309418 282636 309474 282692
rect 309294 282512 309350 282568
rect 309418 282512 309474 282568
rect 304294 281856 304350 281912
rect 304418 281856 304474 281912
rect 304294 281732 304350 281788
rect 304418 281732 304474 281788
rect 304294 281608 304350 281664
rect 304418 281608 304474 281664
rect 304294 281484 304350 281540
rect 304418 281484 304474 281540
rect 304294 281360 304350 281416
rect 304418 281360 304474 281416
rect 304294 281236 304350 281292
rect 304418 281236 304474 281292
rect 304294 281112 304350 281168
rect 304418 281112 304474 281168
rect 319294 283256 319350 283312
rect 319418 283256 319474 283312
rect 319294 283132 319350 283188
rect 319418 283132 319474 283188
rect 319294 283008 319350 283064
rect 319418 283008 319474 283064
rect 319294 282884 319350 282940
rect 319418 282884 319474 282940
rect 319294 282760 319350 282816
rect 319418 282760 319474 282816
rect 319294 282636 319350 282692
rect 319418 282636 319474 282692
rect 319294 282512 319350 282568
rect 319418 282512 319474 282568
rect 314294 281856 314350 281912
rect 314418 281856 314474 281912
rect 314294 281732 314350 281788
rect 314418 281732 314474 281788
rect 314294 281608 314350 281664
rect 314418 281608 314474 281664
rect 314294 281484 314350 281540
rect 314418 281484 314474 281540
rect 314294 281360 314350 281416
rect 314418 281360 314474 281416
rect 314294 281236 314350 281292
rect 314418 281236 314474 281292
rect 314294 281112 314350 281168
rect 314418 281112 314474 281168
rect 329294 283256 329350 283312
rect 329418 283256 329474 283312
rect 329294 283132 329350 283188
rect 329418 283132 329474 283188
rect 329294 283008 329350 283064
rect 329418 283008 329474 283064
rect 329294 282884 329350 282940
rect 329418 282884 329474 282940
rect 329294 282760 329350 282816
rect 329418 282760 329474 282816
rect 329294 282636 329350 282692
rect 329418 282636 329474 282692
rect 329294 282512 329350 282568
rect 329418 282512 329474 282568
rect 324294 281856 324350 281912
rect 324418 281856 324474 281912
rect 324294 281732 324350 281788
rect 324418 281732 324474 281788
rect 324294 281608 324350 281664
rect 324418 281608 324474 281664
rect 324294 281484 324350 281540
rect 324418 281484 324474 281540
rect 324294 281360 324350 281416
rect 324418 281360 324474 281416
rect 324294 281236 324350 281292
rect 324418 281236 324474 281292
rect 324294 281112 324350 281168
rect 324418 281112 324474 281168
rect 339294 283256 339350 283312
rect 339418 283256 339474 283312
rect 339294 283132 339350 283188
rect 339418 283132 339474 283188
rect 339294 283008 339350 283064
rect 339418 283008 339474 283064
rect 339294 282884 339350 282940
rect 339418 282884 339474 282940
rect 339294 282760 339350 282816
rect 339418 282760 339474 282816
rect 339294 282636 339350 282692
rect 339418 282636 339474 282692
rect 339294 282512 339350 282568
rect 339418 282512 339474 282568
rect 334294 281856 334350 281912
rect 334418 281856 334474 281912
rect 334294 281732 334350 281788
rect 334418 281732 334474 281788
rect 334294 281608 334350 281664
rect 334418 281608 334474 281664
rect 334294 281484 334350 281540
rect 334418 281484 334474 281540
rect 334294 281360 334350 281416
rect 334418 281360 334474 281416
rect 334294 281236 334350 281292
rect 334418 281236 334474 281292
rect 334294 281112 334350 281168
rect 334418 281112 334474 281168
rect 349294 283256 349350 283312
rect 349418 283256 349474 283312
rect 349294 283132 349350 283188
rect 349418 283132 349474 283188
rect 349294 283008 349350 283064
rect 349418 283008 349474 283064
rect 349294 282884 349350 282940
rect 349418 282884 349474 282940
rect 349294 282760 349350 282816
rect 349418 282760 349474 282816
rect 349294 282636 349350 282692
rect 349418 282636 349474 282692
rect 349294 282512 349350 282568
rect 349418 282512 349474 282568
rect 344294 281856 344350 281912
rect 344418 281856 344474 281912
rect 344294 281732 344350 281788
rect 344418 281732 344474 281788
rect 344294 281608 344350 281664
rect 344418 281608 344474 281664
rect 344294 281484 344350 281540
rect 344418 281484 344474 281540
rect 344294 281360 344350 281416
rect 344418 281360 344474 281416
rect 344294 281236 344350 281292
rect 344418 281236 344474 281292
rect 344294 281112 344350 281168
rect 344418 281112 344474 281168
rect 359294 283256 359350 283312
rect 359418 283256 359474 283312
rect 359294 283132 359350 283188
rect 359418 283132 359474 283188
rect 359294 283008 359350 283064
rect 359418 283008 359474 283064
rect 359294 282884 359350 282940
rect 359418 282884 359474 282940
rect 359294 282760 359350 282816
rect 359418 282760 359474 282816
rect 359294 282636 359350 282692
rect 359418 282636 359474 282692
rect 359294 282512 359350 282568
rect 359418 282512 359474 282568
rect 354294 281856 354350 281912
rect 354418 281856 354474 281912
rect 354294 281732 354350 281788
rect 354418 281732 354474 281788
rect 354294 281608 354350 281664
rect 354418 281608 354474 281664
rect 354294 281484 354350 281540
rect 354418 281484 354474 281540
rect 354294 281360 354350 281416
rect 354418 281360 354474 281416
rect 354294 281236 354350 281292
rect 354418 281236 354474 281292
rect 354294 281112 354350 281168
rect 354418 281112 354474 281168
rect 369294 283256 369350 283312
rect 369418 283256 369474 283312
rect 369294 283132 369350 283188
rect 369418 283132 369474 283188
rect 369294 283008 369350 283064
rect 369418 283008 369474 283064
rect 369294 282884 369350 282940
rect 369418 282884 369474 282940
rect 369294 282760 369350 282816
rect 369418 282760 369474 282816
rect 369294 282636 369350 282692
rect 369418 282636 369474 282692
rect 369294 282512 369350 282568
rect 369418 282512 369474 282568
rect 364294 281856 364350 281912
rect 364418 281856 364474 281912
rect 364294 281732 364350 281788
rect 364418 281732 364474 281788
rect 364294 281608 364350 281664
rect 364418 281608 364474 281664
rect 364294 281484 364350 281540
rect 364418 281484 364474 281540
rect 364294 281360 364350 281416
rect 364418 281360 364474 281416
rect 364294 281236 364350 281292
rect 364418 281236 364474 281292
rect 364294 281112 364350 281168
rect 364418 281112 364474 281168
rect 379294 283256 379350 283312
rect 379418 283256 379474 283312
rect 379294 283132 379350 283188
rect 379418 283132 379474 283188
rect 379294 283008 379350 283064
rect 379418 283008 379474 283064
rect 379294 282884 379350 282940
rect 379418 282884 379474 282940
rect 379294 282760 379350 282816
rect 379418 282760 379474 282816
rect 379294 282636 379350 282692
rect 379418 282636 379474 282692
rect 379294 282512 379350 282568
rect 379418 282512 379474 282568
rect 374294 281856 374350 281912
rect 374418 281856 374474 281912
rect 374294 281732 374350 281788
rect 374418 281732 374474 281788
rect 374294 281608 374350 281664
rect 374418 281608 374474 281664
rect 374294 281484 374350 281540
rect 374418 281484 374474 281540
rect 374294 281360 374350 281416
rect 374418 281360 374474 281416
rect 374294 281236 374350 281292
rect 374418 281236 374474 281292
rect 374294 281112 374350 281168
rect 374418 281112 374474 281168
rect 389294 283256 389350 283312
rect 389418 283256 389474 283312
rect 389294 283132 389350 283188
rect 389418 283132 389474 283188
rect 389294 283008 389350 283064
rect 389418 283008 389474 283064
rect 389294 282884 389350 282940
rect 389418 282884 389474 282940
rect 389294 282760 389350 282816
rect 389418 282760 389474 282816
rect 389294 282636 389350 282692
rect 389418 282636 389474 282692
rect 389294 282512 389350 282568
rect 389418 282512 389474 282568
rect 384294 281856 384350 281912
rect 384418 281856 384474 281912
rect 384294 281732 384350 281788
rect 384418 281732 384474 281788
rect 384294 281608 384350 281664
rect 384418 281608 384474 281664
rect 384294 281484 384350 281540
rect 384418 281484 384474 281540
rect 384294 281360 384350 281416
rect 384418 281360 384474 281416
rect 384294 281236 384350 281292
rect 384418 281236 384474 281292
rect 384294 281112 384350 281168
rect 384418 281112 384474 281168
rect 399294 283256 399350 283312
rect 399418 283256 399474 283312
rect 399294 283132 399350 283188
rect 399418 283132 399474 283188
rect 399294 283008 399350 283064
rect 399418 283008 399474 283064
rect 399294 282884 399350 282940
rect 399418 282884 399474 282940
rect 399294 282760 399350 282816
rect 399418 282760 399474 282816
rect 399294 282636 399350 282692
rect 399418 282636 399474 282692
rect 399294 282512 399350 282568
rect 399418 282512 399474 282568
rect 394294 281856 394350 281912
rect 394418 281856 394474 281912
rect 394294 281732 394350 281788
rect 394418 281732 394474 281788
rect 394294 281608 394350 281664
rect 394418 281608 394474 281664
rect 394294 281484 394350 281540
rect 394418 281484 394474 281540
rect 394294 281360 394350 281416
rect 394418 281360 394474 281416
rect 394294 281236 394350 281292
rect 394418 281236 394474 281292
rect 394294 281112 394350 281168
rect 394418 281112 394474 281168
rect 409294 283256 409350 283312
rect 409418 283256 409474 283312
rect 409294 283132 409350 283188
rect 409418 283132 409474 283188
rect 409294 283008 409350 283064
rect 409418 283008 409474 283064
rect 409294 282884 409350 282940
rect 409418 282884 409474 282940
rect 409294 282760 409350 282816
rect 409418 282760 409474 282816
rect 409294 282636 409350 282692
rect 409418 282636 409474 282692
rect 409294 282512 409350 282568
rect 409418 282512 409474 282568
rect 404294 281856 404350 281912
rect 404418 281856 404474 281912
rect 404294 281732 404350 281788
rect 404418 281732 404474 281788
rect 404294 281608 404350 281664
rect 404418 281608 404474 281664
rect 404294 281484 404350 281540
rect 404418 281484 404474 281540
rect 404294 281360 404350 281416
rect 404418 281360 404474 281416
rect 404294 281236 404350 281292
rect 404418 281236 404474 281292
rect 404294 281112 404350 281168
rect 404418 281112 404474 281168
rect 419294 283256 419350 283312
rect 419418 283256 419474 283312
rect 419294 283132 419350 283188
rect 419418 283132 419474 283188
rect 419294 283008 419350 283064
rect 419418 283008 419474 283064
rect 419294 282884 419350 282940
rect 419418 282884 419474 282940
rect 419294 282760 419350 282816
rect 419418 282760 419474 282816
rect 419294 282636 419350 282692
rect 419418 282636 419474 282692
rect 419294 282512 419350 282568
rect 419418 282512 419474 282568
rect 414294 281856 414350 281912
rect 414418 281856 414474 281912
rect 414294 281732 414350 281788
rect 414418 281732 414474 281788
rect 414294 281608 414350 281664
rect 414418 281608 414474 281664
rect 414294 281484 414350 281540
rect 414418 281484 414474 281540
rect 414294 281360 414350 281416
rect 414418 281360 414474 281416
rect 414294 281236 414350 281292
rect 414418 281236 414474 281292
rect 414294 281112 414350 281168
rect 414418 281112 414474 281168
rect 429294 283256 429350 283312
rect 429418 283256 429474 283312
rect 429294 283132 429350 283188
rect 429418 283132 429474 283188
rect 429294 283008 429350 283064
rect 429418 283008 429474 283064
rect 429294 282884 429350 282940
rect 429418 282884 429474 282940
rect 429294 282760 429350 282816
rect 429418 282760 429474 282816
rect 429294 282636 429350 282692
rect 429418 282636 429474 282692
rect 429294 282512 429350 282568
rect 429418 282512 429474 282568
rect 424294 281856 424350 281912
rect 424418 281856 424474 281912
rect 424294 281732 424350 281788
rect 424418 281732 424474 281788
rect 424294 281608 424350 281664
rect 424418 281608 424474 281664
rect 424294 281484 424350 281540
rect 424418 281484 424474 281540
rect 424294 281360 424350 281416
rect 424418 281360 424474 281416
rect 424294 281236 424350 281292
rect 424418 281236 424474 281292
rect 424294 281112 424350 281168
rect 424418 281112 424474 281168
rect 439294 283256 439350 283312
rect 439418 283256 439474 283312
rect 439294 283132 439350 283188
rect 439418 283132 439474 283188
rect 439294 283008 439350 283064
rect 439418 283008 439474 283064
rect 439294 282884 439350 282940
rect 439418 282884 439474 282940
rect 439294 282760 439350 282816
rect 439418 282760 439474 282816
rect 439294 282636 439350 282692
rect 439418 282636 439474 282692
rect 439294 282512 439350 282568
rect 439418 282512 439474 282568
rect 434294 281856 434350 281912
rect 434418 281856 434474 281912
rect 434294 281732 434350 281788
rect 434418 281732 434474 281788
rect 434294 281608 434350 281664
rect 434418 281608 434474 281664
rect 434294 281484 434350 281540
rect 434418 281484 434474 281540
rect 434294 281360 434350 281416
rect 434418 281360 434474 281416
rect 434294 281236 434350 281292
rect 434418 281236 434474 281292
rect 434294 281112 434350 281168
rect 434418 281112 434474 281168
rect 449294 283256 449350 283312
rect 449418 283256 449474 283312
rect 449294 283132 449350 283188
rect 449418 283132 449474 283188
rect 449294 283008 449350 283064
rect 449418 283008 449474 283064
rect 449294 282884 449350 282940
rect 449418 282884 449474 282940
rect 449294 282760 449350 282816
rect 449418 282760 449474 282816
rect 449294 282636 449350 282692
rect 449418 282636 449474 282692
rect 449294 282512 449350 282568
rect 449418 282512 449474 282568
rect 444294 281856 444350 281912
rect 444418 281856 444474 281912
rect 444294 281732 444350 281788
rect 444418 281732 444474 281788
rect 444294 281608 444350 281664
rect 444418 281608 444474 281664
rect 444294 281484 444350 281540
rect 444418 281484 444474 281540
rect 444294 281360 444350 281416
rect 444418 281360 444474 281416
rect 444294 281236 444350 281292
rect 444418 281236 444474 281292
rect 444294 281112 444350 281168
rect 444418 281112 444474 281168
rect 459294 283256 459350 283312
rect 459418 283256 459474 283312
rect 459294 283132 459350 283188
rect 459418 283132 459474 283188
rect 459294 283008 459350 283064
rect 459418 283008 459474 283064
rect 459294 282884 459350 282940
rect 459418 282884 459474 282940
rect 459294 282760 459350 282816
rect 459418 282760 459474 282816
rect 459294 282636 459350 282692
rect 459418 282636 459474 282692
rect 459294 282512 459350 282568
rect 459418 282512 459474 282568
rect 454294 281856 454350 281912
rect 454418 281856 454474 281912
rect 454294 281732 454350 281788
rect 454418 281732 454474 281788
rect 454294 281608 454350 281664
rect 454418 281608 454474 281664
rect 454294 281484 454350 281540
rect 454418 281484 454474 281540
rect 454294 281360 454350 281416
rect 454418 281360 454474 281416
rect 454294 281236 454350 281292
rect 454418 281236 454474 281292
rect 454294 281112 454350 281168
rect 454418 281112 454474 281168
rect 469294 283256 469350 283312
rect 469418 283256 469474 283312
rect 469294 283132 469350 283188
rect 469418 283132 469474 283188
rect 469294 283008 469350 283064
rect 469418 283008 469474 283064
rect 469294 282884 469350 282940
rect 469418 282884 469474 282940
rect 469294 282760 469350 282816
rect 469418 282760 469474 282816
rect 469294 282636 469350 282692
rect 469418 282636 469474 282692
rect 469294 282512 469350 282568
rect 469418 282512 469474 282568
rect 464294 281856 464350 281912
rect 464418 281856 464474 281912
rect 464294 281732 464350 281788
rect 464418 281732 464474 281788
rect 464294 281608 464350 281664
rect 464418 281608 464474 281664
rect 464294 281484 464350 281540
rect 464418 281484 464474 281540
rect 464294 281360 464350 281416
rect 464418 281360 464474 281416
rect 464294 281236 464350 281292
rect 464418 281236 464474 281292
rect 464294 281112 464350 281168
rect 464418 281112 464474 281168
rect 479294 283256 479350 283312
rect 479418 283256 479474 283312
rect 479294 283132 479350 283188
rect 479418 283132 479474 283188
rect 479294 283008 479350 283064
rect 479418 283008 479474 283064
rect 479294 282884 479350 282940
rect 479418 282884 479474 282940
rect 479294 282760 479350 282816
rect 479418 282760 479474 282816
rect 479294 282636 479350 282692
rect 479418 282636 479474 282692
rect 479294 282512 479350 282568
rect 479418 282512 479474 282568
rect 474294 281856 474350 281912
rect 474418 281856 474474 281912
rect 474294 281732 474350 281788
rect 474418 281732 474474 281788
rect 474294 281608 474350 281664
rect 474418 281608 474474 281664
rect 474294 281484 474350 281540
rect 474418 281484 474474 281540
rect 474294 281360 474350 281416
rect 474418 281360 474474 281416
rect 474294 281236 474350 281292
rect 474418 281236 474474 281292
rect 474294 281112 474350 281168
rect 474418 281112 474474 281168
rect 489294 283256 489350 283312
rect 489418 283256 489474 283312
rect 489294 283132 489350 283188
rect 489418 283132 489474 283188
rect 489294 283008 489350 283064
rect 489418 283008 489474 283064
rect 489294 282884 489350 282940
rect 489418 282884 489474 282940
rect 489294 282760 489350 282816
rect 489418 282760 489474 282816
rect 489294 282636 489350 282692
rect 489418 282636 489474 282692
rect 489294 282512 489350 282568
rect 489418 282512 489474 282568
rect 484294 281856 484350 281912
rect 484418 281856 484474 281912
rect 484294 281732 484350 281788
rect 484418 281732 484474 281788
rect 484294 281608 484350 281664
rect 484418 281608 484474 281664
rect 484294 281484 484350 281540
rect 484418 281484 484474 281540
rect 484294 281360 484350 281416
rect 484418 281360 484474 281416
rect 484294 281236 484350 281292
rect 484418 281236 484474 281292
rect 484294 281112 484350 281168
rect 484418 281112 484474 281168
rect 499294 283256 499350 283312
rect 499418 283256 499474 283312
rect 499294 283132 499350 283188
rect 499418 283132 499474 283188
rect 499294 283008 499350 283064
rect 499418 283008 499474 283064
rect 499294 282884 499350 282940
rect 499418 282884 499474 282940
rect 499294 282760 499350 282816
rect 499418 282760 499474 282816
rect 499294 282636 499350 282692
rect 499418 282636 499474 282692
rect 499294 282512 499350 282568
rect 499418 282512 499474 282568
rect 494294 281856 494350 281912
rect 494418 281856 494474 281912
rect 494294 281732 494350 281788
rect 494418 281732 494474 281788
rect 494294 281608 494350 281664
rect 494418 281608 494474 281664
rect 494294 281484 494350 281540
rect 494418 281484 494474 281540
rect 494294 281360 494350 281416
rect 494418 281360 494474 281416
rect 494294 281236 494350 281292
rect 494418 281236 494474 281292
rect 494294 281112 494350 281168
rect 494418 281112 494474 281168
rect 509294 283256 509350 283312
rect 509418 283256 509474 283312
rect 509294 283132 509350 283188
rect 509418 283132 509474 283188
rect 509294 283008 509350 283064
rect 509418 283008 509474 283064
rect 509294 282884 509350 282940
rect 509418 282884 509474 282940
rect 509294 282760 509350 282816
rect 509418 282760 509474 282816
rect 509294 282636 509350 282692
rect 509418 282636 509474 282692
rect 509294 282512 509350 282568
rect 509418 282512 509474 282568
rect 504294 281856 504350 281912
rect 504418 281856 504474 281912
rect 504294 281732 504350 281788
rect 504418 281732 504474 281788
rect 504294 281608 504350 281664
rect 504418 281608 504474 281664
rect 504294 281484 504350 281540
rect 504418 281484 504474 281540
rect 504294 281360 504350 281416
rect 504418 281360 504474 281416
rect 504294 281236 504350 281292
rect 504418 281236 504474 281292
rect 504294 281112 504350 281168
rect 504418 281112 504474 281168
rect 519294 283256 519350 283312
rect 519418 283256 519474 283312
rect 519294 283132 519350 283188
rect 519418 283132 519474 283188
rect 519294 283008 519350 283064
rect 519418 283008 519474 283064
rect 519294 282884 519350 282940
rect 519418 282884 519474 282940
rect 519294 282760 519350 282816
rect 519418 282760 519474 282816
rect 519294 282636 519350 282692
rect 519418 282636 519474 282692
rect 519294 282512 519350 282568
rect 519418 282512 519474 282568
rect 514294 281856 514350 281912
rect 514418 281856 514474 281912
rect 514294 281732 514350 281788
rect 514418 281732 514474 281788
rect 514294 281608 514350 281664
rect 514418 281608 514474 281664
rect 514294 281484 514350 281540
rect 514418 281484 514474 281540
rect 514294 281360 514350 281416
rect 514418 281360 514474 281416
rect 514294 281236 514350 281292
rect 514418 281236 514474 281292
rect 514294 281112 514350 281168
rect 514418 281112 514474 281168
rect 529294 283256 529350 283312
rect 529418 283256 529474 283312
rect 529294 283132 529350 283188
rect 529418 283132 529474 283188
rect 529294 283008 529350 283064
rect 529418 283008 529474 283064
rect 529294 282884 529350 282940
rect 529418 282884 529474 282940
rect 529294 282760 529350 282816
rect 529418 282760 529474 282816
rect 529294 282636 529350 282692
rect 529418 282636 529474 282692
rect 529294 282512 529350 282568
rect 529418 282512 529474 282568
rect 524294 281856 524350 281912
rect 524418 281856 524474 281912
rect 524294 281732 524350 281788
rect 524418 281732 524474 281788
rect 524294 281608 524350 281664
rect 524418 281608 524474 281664
rect 524294 281484 524350 281540
rect 524418 281484 524474 281540
rect 524294 281360 524350 281416
rect 524418 281360 524474 281416
rect 524294 281236 524350 281292
rect 524418 281236 524474 281292
rect 524294 281112 524350 281168
rect 524418 281112 524474 281168
rect 539294 283256 539350 283312
rect 539418 283256 539474 283312
rect 539294 283132 539350 283188
rect 539418 283132 539474 283188
rect 539294 283008 539350 283064
rect 539418 283008 539474 283064
rect 539294 282884 539350 282940
rect 539418 282884 539474 282940
rect 539294 282760 539350 282816
rect 539418 282760 539474 282816
rect 539294 282636 539350 282692
rect 539418 282636 539474 282692
rect 539294 282512 539350 282568
rect 539418 282512 539474 282568
rect 534294 281856 534350 281912
rect 534418 281856 534474 281912
rect 534294 281732 534350 281788
rect 534418 281732 534474 281788
rect 534294 281608 534350 281664
rect 534418 281608 534474 281664
rect 534294 281484 534350 281540
rect 534418 281484 534474 281540
rect 534294 281360 534350 281416
rect 534418 281360 534474 281416
rect 534294 281236 534350 281292
rect 534418 281236 534474 281292
rect 534294 281112 534350 281168
rect 534418 281112 534474 281168
rect 549294 283256 549350 283312
rect 549418 283256 549474 283312
rect 549294 283132 549350 283188
rect 549418 283132 549474 283188
rect 549294 283008 549350 283064
rect 549418 283008 549474 283064
rect 549294 282884 549350 282940
rect 549418 282884 549474 282940
rect 549294 282760 549350 282816
rect 549418 282760 549474 282816
rect 549294 282636 549350 282692
rect 549418 282636 549474 282692
rect 549294 282512 549350 282568
rect 549418 282512 549474 282568
rect 544294 281856 544350 281912
rect 544418 281856 544474 281912
rect 544294 281732 544350 281788
rect 544418 281732 544474 281788
rect 544294 281608 544350 281664
rect 544418 281608 544474 281664
rect 544294 281484 544350 281540
rect 544418 281484 544474 281540
rect 544294 281360 544350 281416
rect 544418 281360 544474 281416
rect 544294 281236 544350 281292
rect 544418 281236 544474 281292
rect 544294 281112 544350 281168
rect 544418 281112 544474 281168
rect 590970 283316 591026 283372
rect 591094 283316 591150 283372
rect 591218 283316 591274 283372
rect 591342 283316 591398 283372
rect 591466 283316 591522 283372
rect 591590 283316 591646 283372
rect 591714 283316 591770 283372
rect 590970 283192 591026 283248
rect 591094 283192 591150 283248
rect 591218 283192 591274 283248
rect 591342 283192 591398 283248
rect 591466 283192 591522 283248
rect 591590 283192 591646 283248
rect 591714 283192 591770 283248
rect 590970 283068 591026 283124
rect 591094 283068 591150 283124
rect 591218 283068 591274 283124
rect 591342 283068 591398 283124
rect 591466 283068 591522 283124
rect 591590 283068 591646 283124
rect 591714 283068 591770 283124
rect 590970 282944 591026 283000
rect 591094 282944 591150 283000
rect 591218 282944 591274 283000
rect 591342 282944 591398 283000
rect 591466 282944 591522 283000
rect 591590 282944 591646 283000
rect 591714 282944 591770 283000
rect 590970 282820 591026 282876
rect 591094 282820 591150 282876
rect 591218 282820 591274 282876
rect 591342 282820 591398 282876
rect 591466 282820 591522 282876
rect 591590 282820 591646 282876
rect 591714 282820 591770 282876
rect 590970 282696 591026 282752
rect 591094 282696 591150 282752
rect 591218 282696 591274 282752
rect 591342 282696 591398 282752
rect 591466 282696 591522 282752
rect 591590 282696 591646 282752
rect 591714 282696 591770 282752
rect 590970 282572 591026 282628
rect 591094 282572 591150 282628
rect 591218 282572 591274 282628
rect 591342 282572 591398 282628
rect 591466 282572 591522 282628
rect 591590 282572 591646 282628
rect 591714 282572 591770 282628
rect 554294 281856 554350 281912
rect 554418 281856 554474 281912
rect 554294 281732 554350 281788
rect 554418 281732 554474 281788
rect 554294 281608 554350 281664
rect 554418 281608 554474 281664
rect 554294 281484 554350 281540
rect 554418 281484 554474 281540
rect 554294 281360 554350 281416
rect 554418 281360 554474 281416
rect 554294 281236 554350 281292
rect 554418 281236 554474 281292
rect 554294 281112 554350 281168
rect 554418 281112 554474 281168
rect 79300 273566 79356 273622
rect 79600 273566 79656 273622
rect 79900 273566 79956 273622
rect 79300 266566 79356 266622
rect 79600 266566 79656 266622
rect 79900 266566 79956 266622
rect 79300 259566 79356 259622
rect 79600 259566 79656 259622
rect 79900 259566 79956 259622
rect 79148 255316 79204 255372
rect 79272 255316 79328 255372
rect 79396 255316 79452 255372
rect 79520 255316 79576 255372
rect 79644 255316 79700 255372
rect 79768 255316 79824 255372
rect 79892 255316 79948 255372
rect 79148 255192 79204 255248
rect 79272 255192 79328 255248
rect 79396 255192 79452 255248
rect 79520 255192 79576 255248
rect 79644 255192 79700 255248
rect 79768 255192 79824 255248
rect 79892 255192 79948 255248
rect 79284 248992 79340 249048
rect 79584 248992 79640 249048
rect 79884 248992 79940 249048
rect 79300 232566 79356 232622
rect 79600 232566 79656 232622
rect 79900 232566 79956 232622
rect 79148 229316 79204 229372
rect 79272 229316 79328 229372
rect 79396 229316 79452 229372
rect 79520 229316 79576 229372
rect 79644 229316 79700 229372
rect 79768 229316 79824 229372
rect 79892 229316 79948 229372
rect 79148 229192 79204 229248
rect 79272 229192 79328 229248
rect 79396 229192 79452 229248
rect 79520 229192 79576 229248
rect 79644 229192 79700 229248
rect 79768 229192 79824 229248
rect 79892 229192 79948 229248
rect 79300 225566 79356 225622
rect 79600 225566 79656 225622
rect 79900 225566 79956 225622
rect 79300 218566 79356 218622
rect 79600 218566 79656 218622
rect 79900 218566 79956 218622
rect 79284 207992 79340 208048
rect 79584 207992 79640 208048
rect 79884 207992 79940 208048
rect 79148 203316 79204 203372
rect 79272 203316 79328 203372
rect 79396 203316 79452 203372
rect 79520 203316 79576 203372
rect 79644 203316 79700 203372
rect 79768 203316 79824 203372
rect 79892 203316 79948 203372
rect 79148 203192 79204 203248
rect 79272 203192 79328 203248
rect 79396 203192 79452 203248
rect 79520 203192 79576 203248
rect 79644 203192 79700 203248
rect 79768 203192 79824 203248
rect 79892 203192 79948 203248
rect 79300 191566 79356 191622
rect 79600 191566 79656 191622
rect 79900 191566 79956 191622
rect 79300 184566 79356 184622
rect 79600 184566 79656 184622
rect 79900 184566 79956 184622
rect 79300 177566 79356 177622
rect 79600 177566 79656 177622
rect 79900 177566 79956 177622
rect 79148 177316 79204 177372
rect 79272 177316 79328 177372
rect 79396 177316 79452 177372
rect 79520 177316 79576 177372
rect 79644 177316 79700 177372
rect 79768 177316 79824 177372
rect 79892 177316 79948 177372
rect 79148 177192 79204 177248
rect 79272 177192 79328 177248
rect 79396 177192 79452 177248
rect 79520 177192 79576 177248
rect 79644 177192 79700 177248
rect 79768 177192 79824 177248
rect 79892 177192 79948 177248
rect 79148 151316 79204 151372
rect 79272 151316 79328 151372
rect 79396 151316 79452 151372
rect 79520 151316 79576 151372
rect 79644 151316 79700 151372
rect 79768 151316 79824 151372
rect 79892 151316 79948 151372
rect 79148 151192 79204 151248
rect 79272 151192 79328 151248
rect 79396 151192 79452 151248
rect 79520 151192 79576 151248
rect 79644 151192 79700 151248
rect 79768 151192 79824 151248
rect 79892 151192 79948 151248
rect 79148 125316 79204 125372
rect 79272 125316 79328 125372
rect 79396 125316 79452 125372
rect 79520 125316 79576 125372
rect 79644 125316 79700 125372
rect 79768 125316 79824 125372
rect 79892 125316 79948 125372
rect 79148 125192 79204 125248
rect 79272 125192 79328 125248
rect 79396 125192 79452 125248
rect 79520 125192 79576 125248
rect 79644 125192 79700 125248
rect 79768 125192 79824 125248
rect 79892 125192 79948 125248
rect 79148 99316 79204 99372
rect 79272 99316 79328 99372
rect 79396 99316 79452 99372
rect 79520 99316 79576 99372
rect 79644 99316 79700 99372
rect 79768 99316 79824 99372
rect 79892 99316 79948 99372
rect 79148 99192 79204 99248
rect 79272 99192 79328 99248
rect 79396 99192 79452 99248
rect 79520 99192 79576 99248
rect 79644 99192 79700 99248
rect 79768 99192 79824 99248
rect 79892 99192 79948 99248
rect 590970 255316 591026 255372
rect 591094 255316 591150 255372
rect 591218 255316 591274 255372
rect 591342 255316 591398 255372
rect 591466 255316 591522 255372
rect 591590 255316 591646 255372
rect 591714 255316 591770 255372
rect 590970 255192 591026 255248
rect 591094 255192 591150 255248
rect 591218 255192 591274 255248
rect 591342 255192 591398 255248
rect 591466 255192 591522 255248
rect 591590 255192 591646 255248
rect 591714 255192 591770 255248
rect 590970 229316 591026 229372
rect 591094 229316 591150 229372
rect 591218 229316 591274 229372
rect 591342 229316 591398 229372
rect 591466 229316 591522 229372
rect 591590 229316 591646 229372
rect 591714 229316 591770 229372
rect 590970 229192 591026 229248
rect 591094 229192 591150 229248
rect 591218 229192 591274 229248
rect 591342 229192 591398 229248
rect 591466 229192 591522 229248
rect 591590 229192 591646 229248
rect 591714 229192 591770 229248
rect 590970 203316 591026 203372
rect 591094 203316 591150 203372
rect 591218 203316 591274 203372
rect 591342 203316 591398 203372
rect 591466 203316 591522 203372
rect 591590 203316 591646 203372
rect 591714 203316 591770 203372
rect 590970 203192 591026 203248
rect 591094 203192 591150 203248
rect 591218 203192 591274 203248
rect 591342 203192 591398 203248
rect 591466 203192 591522 203248
rect 591590 203192 591646 203248
rect 591714 203192 591770 203248
rect 590970 177316 591026 177372
rect 591094 177316 591150 177372
rect 591218 177316 591274 177372
rect 591342 177316 591398 177372
rect 591466 177316 591522 177372
rect 591590 177316 591646 177372
rect 591714 177316 591770 177372
rect 590970 177192 591026 177248
rect 591094 177192 591150 177248
rect 591218 177192 591274 177248
rect 591342 177192 591398 177248
rect 591466 177192 591522 177248
rect 591590 177192 591646 177248
rect 591714 177192 591770 177248
rect 590970 151316 591026 151372
rect 591094 151316 591150 151372
rect 591218 151316 591274 151372
rect 591342 151316 591398 151372
rect 591466 151316 591522 151372
rect 591590 151316 591646 151372
rect 591714 151316 591770 151372
rect 590970 151192 591026 151248
rect 591094 151192 591150 151248
rect 591218 151192 591274 151248
rect 591342 151192 591398 151248
rect 591466 151192 591522 151248
rect 591590 151192 591646 151248
rect 591714 151192 591770 151248
rect 590970 125316 591026 125372
rect 591094 125316 591150 125372
rect 591218 125316 591274 125372
rect 591342 125316 591398 125372
rect 591466 125316 591522 125372
rect 591590 125316 591646 125372
rect 591714 125316 591770 125372
rect 590970 125192 591026 125248
rect 591094 125192 591150 125248
rect 591218 125192 591274 125248
rect 591342 125192 591398 125248
rect 591466 125192 591522 125248
rect 591590 125192 591646 125248
rect 591714 125192 591770 125248
rect 590959 120081 591015 120137
rect 591259 120081 591315 120137
rect 591559 120081 591615 120137
rect 590959 116973 591015 117029
rect 591259 116973 591315 117029
rect 591559 116973 591615 117029
rect 590959 113865 591015 113921
rect 591259 113865 591315 113921
rect 591559 113865 591615 113921
rect 590970 99316 591026 99372
rect 591094 99316 591150 99372
rect 591218 99316 591274 99372
rect 591342 99316 591398 99372
rect 591466 99316 591522 99372
rect 591590 99316 591646 99372
rect 591714 99316 591770 99372
rect 590970 99192 591026 99248
rect 591094 99192 591150 99248
rect 591218 99192 591274 99248
rect 591342 99192 591398 99248
rect 591466 99192 591522 99248
rect 591590 99192 591646 99248
rect 591714 99192 591770 99248
rect 79208 79952 79264 80008
rect 79332 79952 79388 80008
rect 79456 79952 79512 80008
rect 79580 79952 79636 80008
rect 79704 79952 79760 80008
rect 79828 79952 79884 80008
rect 79952 79952 80008 80008
rect 79208 79828 79264 79884
rect 79332 79828 79388 79884
rect 79456 79828 79512 79884
rect 79580 79828 79636 79884
rect 79704 79828 79760 79884
rect 79828 79828 79884 79884
rect 79952 79828 80008 79884
rect 79208 79704 79264 79760
rect 79332 79704 79388 79760
rect 79456 79704 79512 79760
rect 79580 79704 79636 79760
rect 79704 79704 79760 79760
rect 79828 79704 79884 79760
rect 79952 79704 80008 79760
rect 79208 79580 79264 79636
rect 79332 79580 79388 79636
rect 79456 79580 79512 79636
rect 79580 79580 79636 79636
rect 79704 79580 79760 79636
rect 79828 79580 79884 79636
rect 79952 79580 80008 79636
rect 79208 79456 79264 79512
rect 79332 79456 79388 79512
rect 79456 79456 79512 79512
rect 79580 79456 79636 79512
rect 79704 79456 79760 79512
rect 79828 79456 79884 79512
rect 79952 79456 80008 79512
rect 79208 79332 79264 79388
rect 79332 79332 79388 79388
rect 79456 79332 79512 79388
rect 79580 79332 79636 79388
rect 79704 79332 79760 79388
rect 79828 79332 79884 79388
rect 79952 79332 80008 79388
rect 79208 79208 79264 79264
rect 79332 79208 79388 79264
rect 79456 79208 79512 79264
rect 79580 79208 79636 79264
rect 79704 79208 79760 79264
rect 79828 79208 79884 79264
rect 79952 79208 80008 79264
rect 77808 78552 77864 78608
rect 77932 78552 77988 78608
rect 78056 78552 78112 78608
rect 78180 78552 78236 78608
rect 78304 78552 78360 78608
rect 78428 78552 78484 78608
rect 78552 78552 78608 78608
rect 77808 78428 77864 78484
rect 77932 78428 77988 78484
rect 78056 78428 78112 78484
rect 78180 78428 78236 78484
rect 78304 78428 78360 78484
rect 78428 78428 78484 78484
rect 78552 78428 78608 78484
rect 77808 78304 77864 78360
rect 77932 78304 77988 78360
rect 78056 78304 78112 78360
rect 78180 78304 78236 78360
rect 78304 78304 78360 78360
rect 78428 78304 78484 78360
rect 78552 78304 78608 78360
rect 77808 78180 77864 78236
rect 77932 78180 77988 78236
rect 78056 78180 78112 78236
rect 78180 78180 78236 78236
rect 78304 78180 78360 78236
rect 78428 78180 78484 78236
rect 78552 78180 78608 78236
rect 77808 78056 77864 78112
rect 77932 78056 77988 78112
rect 78056 78056 78112 78112
rect 78180 78056 78236 78112
rect 78304 78056 78360 78112
rect 78428 78056 78484 78112
rect 78552 78056 78608 78112
rect 77808 77932 77864 77988
rect 77932 77932 77988 77988
rect 78056 77932 78112 77988
rect 78180 77932 78236 77988
rect 78304 77932 78360 77988
rect 78428 77932 78484 77988
rect 78552 77932 78608 77988
rect 77808 77808 77864 77864
rect 77932 77808 77988 77864
rect 78056 77808 78112 77864
rect 78180 77808 78236 77864
rect 78304 77808 78360 77864
rect 78428 77808 78484 77864
rect 78552 77808 78608 77864
rect 99294 79952 99350 80008
rect 99418 79952 99474 80008
rect 99294 79828 99350 79884
rect 99418 79828 99474 79884
rect 99294 79704 99350 79760
rect 99418 79704 99474 79760
rect 99294 79580 99350 79636
rect 99418 79580 99474 79636
rect 99294 79456 99350 79512
rect 99418 79456 99474 79512
rect 99294 79332 99350 79388
rect 99418 79332 99474 79388
rect 99294 79208 99350 79264
rect 99418 79208 99474 79264
rect 94294 78552 94350 78608
rect 94418 78552 94474 78608
rect 94294 78428 94350 78484
rect 94418 78428 94474 78484
rect 94294 78304 94350 78360
rect 94418 78304 94474 78360
rect 94294 78180 94350 78236
rect 94418 78180 94474 78236
rect 94294 78056 94350 78112
rect 94418 78056 94474 78112
rect 94294 77932 94350 77988
rect 94418 77932 94474 77988
rect 94294 77808 94350 77864
rect 94418 77808 94474 77864
rect 104294 78552 104350 78608
rect 104418 78552 104474 78608
rect 104294 78428 104350 78484
rect 104418 78428 104474 78484
rect 104294 78304 104350 78360
rect 104418 78304 104474 78360
rect 104294 78180 104350 78236
rect 104418 78180 104474 78236
rect 104294 78056 104350 78112
rect 104418 78056 104474 78112
rect 104294 77932 104350 77988
rect 104418 77932 104474 77988
rect 104294 77808 104350 77864
rect 104418 77808 104474 77864
rect 107330 79952 107386 80008
rect 107454 79952 107510 80008
rect 107578 79952 107634 80008
rect 107702 79952 107758 80008
rect 107826 79952 107882 80008
rect 107950 79952 108006 80008
rect 108074 79952 108130 80008
rect 108198 79952 108254 80008
rect 108322 79952 108378 80008
rect 108446 79952 108502 80008
rect 108570 79952 108626 80008
rect 108694 79952 108750 80008
rect 108818 79952 108874 80008
rect 108942 79952 108998 80008
rect 109066 79952 109122 80008
rect 107330 79828 107386 79884
rect 107454 79828 107510 79884
rect 107578 79828 107634 79884
rect 107702 79828 107758 79884
rect 107826 79828 107882 79884
rect 107950 79828 108006 79884
rect 108074 79828 108130 79884
rect 108198 79828 108254 79884
rect 108322 79828 108378 79884
rect 108446 79828 108502 79884
rect 108570 79828 108626 79884
rect 108694 79828 108750 79884
rect 108818 79828 108874 79884
rect 108942 79828 108998 79884
rect 109066 79828 109122 79884
rect 107330 79704 107386 79760
rect 107454 79704 107510 79760
rect 107578 79704 107634 79760
rect 107702 79704 107758 79760
rect 107826 79704 107882 79760
rect 107950 79704 108006 79760
rect 108074 79704 108130 79760
rect 108198 79704 108254 79760
rect 108322 79704 108378 79760
rect 108446 79704 108502 79760
rect 108570 79704 108626 79760
rect 108694 79704 108750 79760
rect 108818 79704 108874 79760
rect 108942 79704 108998 79760
rect 109066 79704 109122 79760
rect 107330 79580 107386 79636
rect 107454 79580 107510 79636
rect 107578 79580 107634 79636
rect 107702 79580 107758 79636
rect 107826 79580 107882 79636
rect 107950 79580 108006 79636
rect 108074 79580 108130 79636
rect 108198 79580 108254 79636
rect 108322 79580 108378 79636
rect 108446 79580 108502 79636
rect 108570 79580 108626 79636
rect 108694 79580 108750 79636
rect 108818 79580 108874 79636
rect 108942 79580 108998 79636
rect 109066 79580 109122 79636
rect 107330 79456 107386 79512
rect 107454 79456 107510 79512
rect 107578 79456 107634 79512
rect 107702 79456 107758 79512
rect 107826 79456 107882 79512
rect 107950 79456 108006 79512
rect 108074 79456 108130 79512
rect 108198 79456 108254 79512
rect 108322 79456 108378 79512
rect 108446 79456 108502 79512
rect 108570 79456 108626 79512
rect 108694 79456 108750 79512
rect 108818 79456 108874 79512
rect 108942 79456 108998 79512
rect 109066 79456 109122 79512
rect 107330 79332 107386 79388
rect 107454 79332 107510 79388
rect 107578 79332 107634 79388
rect 107702 79332 107758 79388
rect 107826 79332 107882 79388
rect 107950 79332 108006 79388
rect 108074 79332 108130 79388
rect 108198 79332 108254 79388
rect 108322 79332 108378 79388
rect 108446 79332 108502 79388
rect 108570 79332 108626 79388
rect 108694 79332 108750 79388
rect 108818 79332 108874 79388
rect 108942 79332 108998 79388
rect 109066 79332 109122 79388
rect 107330 79208 107386 79264
rect 107454 79208 107510 79264
rect 107578 79208 107634 79264
rect 107702 79208 107758 79264
rect 107826 79208 107882 79264
rect 107950 79208 108006 79264
rect 108074 79208 108130 79264
rect 108198 79208 108254 79264
rect 108322 79208 108378 79264
rect 108446 79208 108502 79264
rect 108570 79208 108626 79264
rect 108694 79208 108750 79264
rect 108818 79208 108874 79264
rect 108942 79208 108998 79264
rect 109066 79208 109122 79264
rect 109810 79952 109866 80008
rect 109934 79952 109990 80008
rect 110058 79952 110114 80008
rect 110182 79952 110238 80008
rect 110306 79952 110362 80008
rect 110430 79952 110486 80008
rect 110554 79952 110610 80008
rect 110678 79952 110734 80008
rect 110802 79952 110858 80008
rect 110926 79952 110982 80008
rect 111050 79952 111106 80008
rect 111174 79952 111230 80008
rect 111298 79952 111354 80008
rect 111422 79952 111478 80008
rect 111546 79952 111602 80008
rect 111670 79952 111726 80008
rect 109810 79828 109866 79884
rect 109934 79828 109990 79884
rect 110058 79828 110114 79884
rect 110182 79828 110238 79884
rect 110306 79828 110362 79884
rect 110430 79828 110486 79884
rect 110554 79828 110610 79884
rect 110678 79828 110734 79884
rect 110802 79828 110858 79884
rect 110926 79828 110982 79884
rect 111050 79828 111106 79884
rect 111174 79828 111230 79884
rect 111298 79828 111354 79884
rect 111422 79828 111478 79884
rect 111546 79828 111602 79884
rect 111670 79828 111726 79884
rect 109810 79704 109866 79760
rect 109934 79704 109990 79760
rect 110058 79704 110114 79760
rect 110182 79704 110238 79760
rect 110306 79704 110362 79760
rect 110430 79704 110486 79760
rect 110554 79704 110610 79760
rect 110678 79704 110734 79760
rect 110802 79704 110858 79760
rect 110926 79704 110982 79760
rect 111050 79704 111106 79760
rect 111174 79704 111230 79760
rect 111298 79704 111354 79760
rect 111422 79704 111478 79760
rect 111546 79704 111602 79760
rect 111670 79704 111726 79760
rect 109810 79580 109866 79636
rect 109934 79580 109990 79636
rect 110058 79580 110114 79636
rect 110182 79580 110238 79636
rect 110306 79580 110362 79636
rect 110430 79580 110486 79636
rect 110554 79580 110610 79636
rect 110678 79580 110734 79636
rect 110802 79580 110858 79636
rect 110926 79580 110982 79636
rect 111050 79580 111106 79636
rect 111174 79580 111230 79636
rect 111298 79580 111354 79636
rect 111422 79580 111478 79636
rect 111546 79580 111602 79636
rect 111670 79580 111726 79636
rect 109810 79456 109866 79512
rect 109934 79456 109990 79512
rect 110058 79456 110114 79512
rect 110182 79456 110238 79512
rect 110306 79456 110362 79512
rect 110430 79456 110486 79512
rect 110554 79456 110610 79512
rect 110678 79456 110734 79512
rect 110802 79456 110858 79512
rect 110926 79456 110982 79512
rect 111050 79456 111106 79512
rect 111174 79456 111230 79512
rect 111298 79456 111354 79512
rect 111422 79456 111478 79512
rect 111546 79456 111602 79512
rect 111670 79456 111726 79512
rect 109810 79332 109866 79388
rect 109934 79332 109990 79388
rect 110058 79332 110114 79388
rect 110182 79332 110238 79388
rect 110306 79332 110362 79388
rect 110430 79332 110486 79388
rect 110554 79332 110610 79388
rect 110678 79332 110734 79388
rect 110802 79332 110858 79388
rect 110926 79332 110982 79388
rect 111050 79332 111106 79388
rect 111174 79332 111230 79388
rect 111298 79332 111354 79388
rect 111422 79332 111478 79388
rect 111546 79332 111602 79388
rect 111670 79332 111726 79388
rect 109810 79208 109866 79264
rect 109934 79208 109990 79264
rect 110058 79208 110114 79264
rect 110182 79208 110238 79264
rect 110306 79208 110362 79264
rect 110430 79208 110486 79264
rect 110554 79208 110610 79264
rect 110678 79208 110734 79264
rect 110802 79208 110858 79264
rect 110926 79208 110982 79264
rect 111050 79208 111106 79264
rect 111174 79208 111230 79264
rect 111298 79208 111354 79264
rect 111422 79208 111478 79264
rect 111546 79208 111602 79264
rect 111670 79208 111726 79264
rect 112180 79952 112236 80008
rect 112304 79952 112360 80008
rect 112428 79952 112484 80008
rect 112552 79952 112608 80008
rect 112676 79952 112732 80008
rect 112800 79952 112856 80008
rect 112924 79952 112980 80008
rect 113048 79952 113104 80008
rect 113172 79952 113228 80008
rect 113296 79952 113352 80008
rect 113420 79952 113476 80008
rect 113544 79952 113600 80008
rect 113668 79952 113724 80008
rect 113792 79952 113848 80008
rect 113916 79952 113972 80008
rect 114040 79952 114096 80008
rect 112180 79828 112236 79884
rect 112304 79828 112360 79884
rect 112428 79828 112484 79884
rect 112552 79828 112608 79884
rect 112676 79828 112732 79884
rect 112800 79828 112856 79884
rect 112924 79828 112980 79884
rect 113048 79828 113104 79884
rect 113172 79828 113228 79884
rect 113296 79828 113352 79884
rect 113420 79828 113476 79884
rect 113544 79828 113600 79884
rect 113668 79828 113724 79884
rect 113792 79828 113848 79884
rect 113916 79828 113972 79884
rect 114040 79828 114096 79884
rect 112180 79704 112236 79760
rect 112304 79704 112360 79760
rect 112428 79704 112484 79760
rect 112552 79704 112608 79760
rect 112676 79704 112732 79760
rect 112800 79704 112856 79760
rect 112924 79704 112980 79760
rect 113048 79704 113104 79760
rect 113172 79704 113228 79760
rect 113296 79704 113352 79760
rect 113420 79704 113476 79760
rect 113544 79704 113600 79760
rect 113668 79704 113724 79760
rect 113792 79704 113848 79760
rect 113916 79704 113972 79760
rect 114040 79704 114096 79760
rect 112180 79580 112236 79636
rect 112304 79580 112360 79636
rect 112428 79580 112484 79636
rect 112552 79580 112608 79636
rect 112676 79580 112732 79636
rect 112800 79580 112856 79636
rect 112924 79580 112980 79636
rect 113048 79580 113104 79636
rect 113172 79580 113228 79636
rect 113296 79580 113352 79636
rect 113420 79580 113476 79636
rect 113544 79580 113600 79636
rect 113668 79580 113724 79636
rect 113792 79580 113848 79636
rect 113916 79580 113972 79636
rect 114040 79580 114096 79636
rect 112180 79456 112236 79512
rect 112304 79456 112360 79512
rect 112428 79456 112484 79512
rect 112552 79456 112608 79512
rect 112676 79456 112732 79512
rect 112800 79456 112856 79512
rect 112924 79456 112980 79512
rect 113048 79456 113104 79512
rect 113172 79456 113228 79512
rect 113296 79456 113352 79512
rect 113420 79456 113476 79512
rect 113544 79456 113600 79512
rect 113668 79456 113724 79512
rect 113792 79456 113848 79512
rect 113916 79456 113972 79512
rect 114040 79456 114096 79512
rect 112180 79332 112236 79388
rect 112304 79332 112360 79388
rect 112428 79332 112484 79388
rect 112552 79332 112608 79388
rect 112676 79332 112732 79388
rect 112800 79332 112856 79388
rect 112924 79332 112980 79388
rect 113048 79332 113104 79388
rect 113172 79332 113228 79388
rect 113296 79332 113352 79388
rect 113420 79332 113476 79388
rect 113544 79332 113600 79388
rect 113668 79332 113724 79388
rect 113792 79332 113848 79388
rect 113916 79332 113972 79388
rect 114040 79332 114096 79388
rect 112180 79208 112236 79264
rect 112304 79208 112360 79264
rect 112428 79208 112484 79264
rect 112552 79208 112608 79264
rect 112676 79208 112732 79264
rect 112800 79208 112856 79264
rect 112924 79208 112980 79264
rect 113048 79208 113104 79264
rect 113172 79208 113228 79264
rect 113296 79208 113352 79264
rect 113420 79208 113476 79264
rect 113544 79208 113600 79264
rect 113668 79208 113724 79264
rect 113792 79208 113848 79264
rect 113916 79208 113972 79264
rect 114040 79208 114096 79264
rect 114886 79952 114942 80008
rect 115010 79952 115066 80008
rect 115134 79952 115190 80008
rect 115258 79952 115314 80008
rect 115382 79952 115438 80008
rect 115506 79952 115562 80008
rect 115630 79952 115686 80008
rect 115754 79952 115810 80008
rect 115878 79952 115934 80008
rect 116002 79952 116058 80008
rect 116126 79952 116182 80008
rect 116250 79952 116306 80008
rect 116374 79952 116430 80008
rect 116498 79952 116554 80008
rect 116622 79952 116678 80008
rect 116746 79952 116802 80008
rect 114886 79828 114942 79884
rect 115010 79828 115066 79884
rect 115134 79828 115190 79884
rect 115258 79828 115314 79884
rect 115382 79828 115438 79884
rect 115506 79828 115562 79884
rect 115630 79828 115686 79884
rect 115754 79828 115810 79884
rect 115878 79828 115934 79884
rect 116002 79828 116058 79884
rect 116126 79828 116182 79884
rect 116250 79828 116306 79884
rect 116374 79828 116430 79884
rect 116498 79828 116554 79884
rect 116622 79828 116678 79884
rect 116746 79828 116802 79884
rect 114886 79704 114942 79760
rect 115010 79704 115066 79760
rect 115134 79704 115190 79760
rect 115258 79704 115314 79760
rect 115382 79704 115438 79760
rect 115506 79704 115562 79760
rect 115630 79704 115686 79760
rect 115754 79704 115810 79760
rect 115878 79704 115934 79760
rect 116002 79704 116058 79760
rect 116126 79704 116182 79760
rect 116250 79704 116306 79760
rect 116374 79704 116430 79760
rect 116498 79704 116554 79760
rect 116622 79704 116678 79760
rect 116746 79704 116802 79760
rect 114886 79580 114942 79636
rect 115010 79580 115066 79636
rect 115134 79580 115190 79636
rect 115258 79580 115314 79636
rect 115382 79580 115438 79636
rect 115506 79580 115562 79636
rect 115630 79580 115686 79636
rect 115754 79580 115810 79636
rect 115878 79580 115934 79636
rect 116002 79580 116058 79636
rect 116126 79580 116182 79636
rect 116250 79580 116306 79636
rect 116374 79580 116430 79636
rect 116498 79580 116554 79636
rect 116622 79580 116678 79636
rect 116746 79580 116802 79636
rect 114886 79456 114942 79512
rect 115010 79456 115066 79512
rect 115134 79456 115190 79512
rect 115258 79456 115314 79512
rect 115382 79456 115438 79512
rect 115506 79456 115562 79512
rect 115630 79456 115686 79512
rect 115754 79456 115810 79512
rect 115878 79456 115934 79512
rect 116002 79456 116058 79512
rect 116126 79456 116182 79512
rect 116250 79456 116306 79512
rect 116374 79456 116430 79512
rect 116498 79456 116554 79512
rect 116622 79456 116678 79512
rect 116746 79456 116802 79512
rect 114886 79332 114942 79388
rect 115010 79332 115066 79388
rect 115134 79332 115190 79388
rect 115258 79332 115314 79388
rect 115382 79332 115438 79388
rect 115506 79332 115562 79388
rect 115630 79332 115686 79388
rect 115754 79332 115810 79388
rect 115878 79332 115934 79388
rect 116002 79332 116058 79388
rect 116126 79332 116182 79388
rect 116250 79332 116306 79388
rect 116374 79332 116430 79388
rect 116498 79332 116554 79388
rect 116622 79332 116678 79388
rect 116746 79332 116802 79388
rect 114886 79208 114942 79264
rect 115010 79208 115066 79264
rect 115134 79208 115190 79264
rect 115258 79208 115314 79264
rect 115382 79208 115438 79264
rect 115506 79208 115562 79264
rect 115630 79208 115686 79264
rect 115754 79208 115810 79264
rect 115878 79208 115934 79264
rect 116002 79208 116058 79264
rect 116126 79208 116182 79264
rect 116250 79208 116306 79264
rect 116374 79208 116430 79264
rect 116498 79208 116554 79264
rect 116622 79208 116678 79264
rect 116746 79208 116802 79264
rect 117256 79952 117312 80008
rect 117380 79952 117436 80008
rect 117504 79952 117560 80008
rect 117628 79952 117684 80008
rect 117752 79952 117808 80008
rect 117876 79952 117932 80008
rect 118000 79952 118056 80008
rect 118124 79952 118180 80008
rect 118248 79952 118304 80008
rect 118372 79952 118428 80008
rect 118496 79952 118552 80008
rect 118620 79952 118676 80008
rect 118744 79952 118800 80008
rect 118868 79952 118924 80008
rect 118992 79952 119048 80008
rect 119116 79952 119172 80008
rect 117256 79828 117312 79884
rect 117380 79828 117436 79884
rect 117504 79828 117560 79884
rect 117628 79828 117684 79884
rect 117752 79828 117808 79884
rect 117876 79828 117932 79884
rect 118000 79828 118056 79884
rect 118124 79828 118180 79884
rect 118248 79828 118304 79884
rect 118372 79828 118428 79884
rect 118496 79828 118552 79884
rect 118620 79828 118676 79884
rect 118744 79828 118800 79884
rect 118868 79828 118924 79884
rect 118992 79828 119048 79884
rect 119116 79828 119172 79884
rect 117256 79704 117312 79760
rect 117380 79704 117436 79760
rect 117504 79704 117560 79760
rect 117628 79704 117684 79760
rect 117752 79704 117808 79760
rect 117876 79704 117932 79760
rect 118000 79704 118056 79760
rect 118124 79704 118180 79760
rect 118248 79704 118304 79760
rect 118372 79704 118428 79760
rect 118496 79704 118552 79760
rect 118620 79704 118676 79760
rect 118744 79704 118800 79760
rect 118868 79704 118924 79760
rect 118992 79704 119048 79760
rect 119116 79704 119172 79760
rect 117256 79580 117312 79636
rect 117380 79580 117436 79636
rect 117504 79580 117560 79636
rect 117628 79580 117684 79636
rect 117752 79580 117808 79636
rect 117876 79580 117932 79636
rect 118000 79580 118056 79636
rect 118124 79580 118180 79636
rect 118248 79580 118304 79636
rect 118372 79580 118428 79636
rect 118496 79580 118552 79636
rect 118620 79580 118676 79636
rect 118744 79580 118800 79636
rect 118868 79580 118924 79636
rect 118992 79580 119048 79636
rect 119116 79580 119172 79636
rect 117256 79456 117312 79512
rect 117380 79456 117436 79512
rect 117504 79456 117560 79512
rect 117628 79456 117684 79512
rect 117752 79456 117808 79512
rect 117876 79456 117932 79512
rect 118000 79456 118056 79512
rect 118124 79456 118180 79512
rect 118248 79456 118304 79512
rect 118372 79456 118428 79512
rect 118496 79456 118552 79512
rect 118620 79456 118676 79512
rect 118744 79456 118800 79512
rect 118868 79456 118924 79512
rect 118992 79456 119048 79512
rect 119116 79456 119172 79512
rect 117256 79332 117312 79388
rect 117380 79332 117436 79388
rect 117504 79332 117560 79388
rect 117628 79332 117684 79388
rect 117752 79332 117808 79388
rect 117876 79332 117932 79388
rect 118000 79332 118056 79388
rect 118124 79332 118180 79388
rect 118248 79332 118304 79388
rect 118372 79332 118428 79388
rect 118496 79332 118552 79388
rect 118620 79332 118676 79388
rect 118744 79332 118800 79388
rect 118868 79332 118924 79388
rect 118992 79332 119048 79388
rect 119116 79332 119172 79388
rect 117256 79208 117312 79264
rect 117380 79208 117436 79264
rect 117504 79208 117560 79264
rect 117628 79208 117684 79264
rect 117752 79208 117808 79264
rect 117876 79208 117932 79264
rect 118000 79208 118056 79264
rect 118124 79208 118180 79264
rect 118248 79208 118304 79264
rect 118372 79208 118428 79264
rect 118496 79208 118552 79264
rect 118620 79208 118676 79264
rect 118744 79208 118800 79264
rect 118868 79208 118924 79264
rect 118992 79208 119048 79264
rect 119116 79208 119172 79264
rect 119860 79952 119916 80008
rect 119984 79952 120040 80008
rect 120108 79952 120164 80008
rect 120232 79952 120288 80008
rect 120356 79952 120412 80008
rect 120480 79952 120536 80008
rect 120604 79952 120660 80008
rect 120728 79952 120784 80008
rect 120852 79952 120908 80008
rect 120976 79952 121032 80008
rect 121100 79952 121156 80008
rect 121224 79952 121280 80008
rect 121348 79952 121404 80008
rect 121472 79952 121528 80008
rect 121596 79952 121652 80008
rect 119860 79828 119916 79884
rect 119984 79828 120040 79884
rect 120108 79828 120164 79884
rect 120232 79828 120288 79884
rect 120356 79828 120412 79884
rect 120480 79828 120536 79884
rect 120604 79828 120660 79884
rect 120728 79828 120784 79884
rect 120852 79828 120908 79884
rect 120976 79828 121032 79884
rect 121100 79828 121156 79884
rect 121224 79828 121280 79884
rect 121348 79828 121404 79884
rect 121472 79828 121528 79884
rect 121596 79828 121652 79884
rect 119860 79704 119916 79760
rect 119984 79704 120040 79760
rect 120108 79704 120164 79760
rect 120232 79704 120288 79760
rect 120356 79704 120412 79760
rect 120480 79704 120536 79760
rect 120604 79704 120660 79760
rect 120728 79704 120784 79760
rect 120852 79704 120908 79760
rect 120976 79704 121032 79760
rect 121100 79704 121156 79760
rect 121224 79704 121280 79760
rect 121348 79704 121404 79760
rect 121472 79704 121528 79760
rect 121596 79704 121652 79760
rect 119860 79580 119916 79636
rect 119984 79580 120040 79636
rect 120108 79580 120164 79636
rect 120232 79580 120288 79636
rect 120356 79580 120412 79636
rect 120480 79580 120536 79636
rect 120604 79580 120660 79636
rect 120728 79580 120784 79636
rect 120852 79580 120908 79636
rect 120976 79580 121032 79636
rect 121100 79580 121156 79636
rect 121224 79580 121280 79636
rect 121348 79580 121404 79636
rect 121472 79580 121528 79636
rect 121596 79580 121652 79636
rect 119860 79456 119916 79512
rect 119984 79456 120040 79512
rect 120108 79456 120164 79512
rect 120232 79456 120288 79512
rect 120356 79456 120412 79512
rect 120480 79456 120536 79512
rect 120604 79456 120660 79512
rect 120728 79456 120784 79512
rect 120852 79456 120908 79512
rect 120976 79456 121032 79512
rect 121100 79456 121156 79512
rect 121224 79456 121280 79512
rect 121348 79456 121404 79512
rect 121472 79456 121528 79512
rect 121596 79456 121652 79512
rect 119860 79332 119916 79388
rect 119984 79332 120040 79388
rect 120108 79332 120164 79388
rect 120232 79332 120288 79388
rect 120356 79332 120412 79388
rect 120480 79332 120536 79388
rect 120604 79332 120660 79388
rect 120728 79332 120784 79388
rect 120852 79332 120908 79388
rect 120976 79332 121032 79388
rect 121100 79332 121156 79388
rect 121224 79332 121280 79388
rect 121348 79332 121404 79388
rect 121472 79332 121528 79388
rect 121596 79332 121652 79388
rect 119860 79208 119916 79264
rect 119984 79208 120040 79264
rect 120108 79208 120164 79264
rect 120232 79208 120288 79264
rect 120356 79208 120412 79264
rect 120480 79208 120536 79264
rect 120604 79208 120660 79264
rect 120728 79208 120784 79264
rect 120852 79208 120908 79264
rect 120976 79208 121032 79264
rect 121100 79208 121156 79264
rect 121224 79208 121280 79264
rect 121348 79208 121404 79264
rect 121472 79208 121528 79264
rect 121596 79208 121652 79264
rect 129294 79952 129350 80008
rect 129418 79952 129474 80008
rect 129294 79828 129350 79884
rect 129418 79828 129474 79884
rect 129294 79704 129350 79760
rect 129418 79704 129474 79760
rect 129294 79580 129350 79636
rect 129418 79580 129474 79636
rect 129294 79456 129350 79512
rect 129418 79456 129474 79512
rect 129294 79332 129350 79388
rect 129418 79332 129474 79388
rect 129294 79208 129350 79264
rect 129418 79208 129474 79264
rect 124294 78552 124350 78608
rect 124418 78552 124474 78608
rect 124294 78428 124350 78484
rect 124418 78428 124474 78484
rect 124294 78304 124350 78360
rect 124418 78304 124474 78360
rect 124294 78180 124350 78236
rect 124418 78180 124474 78236
rect 124294 78056 124350 78112
rect 124418 78056 124474 78112
rect 124294 77932 124350 77988
rect 124418 77932 124474 77988
rect 124294 77808 124350 77864
rect 124418 77808 124474 77864
rect 139294 79952 139350 80008
rect 139418 79952 139474 80008
rect 139294 79828 139350 79884
rect 139418 79828 139474 79884
rect 139294 79704 139350 79760
rect 139418 79704 139474 79760
rect 139294 79580 139350 79636
rect 139418 79580 139474 79636
rect 139294 79456 139350 79512
rect 139418 79456 139474 79512
rect 139294 79332 139350 79388
rect 139418 79332 139474 79388
rect 139294 79208 139350 79264
rect 139418 79208 139474 79264
rect 134294 78552 134350 78608
rect 134418 78552 134474 78608
rect 134294 78428 134350 78484
rect 134418 78428 134474 78484
rect 134294 78304 134350 78360
rect 134418 78304 134474 78360
rect 134294 78180 134350 78236
rect 134418 78180 134474 78236
rect 134294 78056 134350 78112
rect 134418 78056 134474 78112
rect 134294 77932 134350 77988
rect 134418 77932 134474 77988
rect 134294 77808 134350 77864
rect 134418 77808 134474 77864
rect 149294 79952 149350 80008
rect 149418 79952 149474 80008
rect 149294 79828 149350 79884
rect 149418 79828 149474 79884
rect 149294 79704 149350 79760
rect 149418 79704 149474 79760
rect 149294 79580 149350 79636
rect 149418 79580 149474 79636
rect 149294 79456 149350 79512
rect 149418 79456 149474 79512
rect 149294 79332 149350 79388
rect 149418 79332 149474 79388
rect 149294 79208 149350 79264
rect 149418 79208 149474 79264
rect 144294 78552 144350 78608
rect 144418 78552 144474 78608
rect 144294 78428 144350 78484
rect 144418 78428 144474 78484
rect 144294 78304 144350 78360
rect 144418 78304 144474 78360
rect 144294 78180 144350 78236
rect 144418 78180 144474 78236
rect 144294 78056 144350 78112
rect 144418 78056 144474 78112
rect 144294 77932 144350 77988
rect 144418 77932 144474 77988
rect 144294 77808 144350 77864
rect 144418 77808 144474 77864
rect 159294 79952 159350 80008
rect 159418 79952 159474 80008
rect 159294 79828 159350 79884
rect 159418 79828 159474 79884
rect 159294 79704 159350 79760
rect 159418 79704 159474 79760
rect 159294 79580 159350 79636
rect 159418 79580 159474 79636
rect 159294 79456 159350 79512
rect 159418 79456 159474 79512
rect 159294 79332 159350 79388
rect 159418 79332 159474 79388
rect 159294 79208 159350 79264
rect 159418 79208 159474 79264
rect 154294 78552 154350 78608
rect 154418 78552 154474 78608
rect 154294 78428 154350 78484
rect 154418 78428 154474 78484
rect 154294 78304 154350 78360
rect 154418 78304 154474 78360
rect 154294 78180 154350 78236
rect 154418 78180 154474 78236
rect 154294 78056 154350 78112
rect 154418 78056 154474 78112
rect 154294 77932 154350 77988
rect 154418 77932 154474 77988
rect 154294 77808 154350 77864
rect 154418 77808 154474 77864
rect 169294 79952 169350 80008
rect 169418 79952 169474 80008
rect 169294 79828 169350 79884
rect 169418 79828 169474 79884
rect 169294 79704 169350 79760
rect 169418 79704 169474 79760
rect 169294 79580 169350 79636
rect 169418 79580 169474 79636
rect 169294 79456 169350 79512
rect 169418 79456 169474 79512
rect 169294 79332 169350 79388
rect 169418 79332 169474 79388
rect 169294 79208 169350 79264
rect 169418 79208 169474 79264
rect 164294 78552 164350 78608
rect 164418 78552 164474 78608
rect 164294 78428 164350 78484
rect 164418 78428 164474 78484
rect 164294 78304 164350 78360
rect 164418 78304 164474 78360
rect 164294 78180 164350 78236
rect 164418 78180 164474 78236
rect 164294 78056 164350 78112
rect 164418 78056 164474 78112
rect 164294 77932 164350 77988
rect 164418 77932 164474 77988
rect 164294 77808 164350 77864
rect 164418 77808 164474 77864
rect 179294 79952 179350 80008
rect 179418 79952 179474 80008
rect 179294 79828 179350 79884
rect 179418 79828 179474 79884
rect 179294 79704 179350 79760
rect 179418 79704 179474 79760
rect 179294 79580 179350 79636
rect 179418 79580 179474 79636
rect 179294 79456 179350 79512
rect 179418 79456 179474 79512
rect 179294 79332 179350 79388
rect 179418 79332 179474 79388
rect 179294 79208 179350 79264
rect 179418 79208 179474 79264
rect 174294 78552 174350 78608
rect 174418 78552 174474 78608
rect 174294 78428 174350 78484
rect 174418 78428 174474 78484
rect 174294 78304 174350 78360
rect 174418 78304 174474 78360
rect 174294 78180 174350 78236
rect 174418 78180 174474 78236
rect 174294 78056 174350 78112
rect 174418 78056 174474 78112
rect 174294 77932 174350 77988
rect 174418 77932 174474 77988
rect 174294 77808 174350 77864
rect 174418 77808 174474 77864
rect 189294 79952 189350 80008
rect 189418 79952 189474 80008
rect 189294 79828 189350 79884
rect 189418 79828 189474 79884
rect 189294 79704 189350 79760
rect 189418 79704 189474 79760
rect 189294 79580 189350 79636
rect 189418 79580 189474 79636
rect 189294 79456 189350 79512
rect 189418 79456 189474 79512
rect 189294 79332 189350 79388
rect 189418 79332 189474 79388
rect 189294 79208 189350 79264
rect 189418 79208 189474 79264
rect 184294 78552 184350 78608
rect 184418 78552 184474 78608
rect 184294 78428 184350 78484
rect 184418 78428 184474 78484
rect 184294 78304 184350 78360
rect 184418 78304 184474 78360
rect 184294 78180 184350 78236
rect 184418 78180 184474 78236
rect 184294 78056 184350 78112
rect 184418 78056 184474 78112
rect 184294 77932 184350 77988
rect 184418 77932 184474 77988
rect 184294 77808 184350 77864
rect 184418 77808 184474 77864
rect 199294 79952 199350 80008
rect 199418 79952 199474 80008
rect 199294 79828 199350 79884
rect 199418 79828 199474 79884
rect 199294 79704 199350 79760
rect 199418 79704 199474 79760
rect 199294 79580 199350 79636
rect 199418 79580 199474 79636
rect 199294 79456 199350 79512
rect 199418 79456 199474 79512
rect 199294 79332 199350 79388
rect 199418 79332 199474 79388
rect 199294 79208 199350 79264
rect 199418 79208 199474 79264
rect 194294 78552 194350 78608
rect 194418 78552 194474 78608
rect 194294 78428 194350 78484
rect 194418 78428 194474 78484
rect 194294 78304 194350 78360
rect 194418 78304 194474 78360
rect 194294 78180 194350 78236
rect 194418 78180 194474 78236
rect 194294 78056 194350 78112
rect 194418 78056 194474 78112
rect 194294 77932 194350 77988
rect 194418 77932 194474 77988
rect 194294 77808 194350 77864
rect 194418 77808 194474 77864
rect 209294 79952 209350 80008
rect 209418 79952 209474 80008
rect 209294 79828 209350 79884
rect 209418 79828 209474 79884
rect 209294 79704 209350 79760
rect 209418 79704 209474 79760
rect 209294 79580 209350 79636
rect 209418 79580 209474 79636
rect 209294 79456 209350 79512
rect 209418 79456 209474 79512
rect 209294 79332 209350 79388
rect 209418 79332 209474 79388
rect 209294 79208 209350 79264
rect 209418 79208 209474 79264
rect 204294 78552 204350 78608
rect 204418 78552 204474 78608
rect 204294 78428 204350 78484
rect 204418 78428 204474 78484
rect 204294 78304 204350 78360
rect 204418 78304 204474 78360
rect 204294 78180 204350 78236
rect 204418 78180 204474 78236
rect 204294 78056 204350 78112
rect 204418 78056 204474 78112
rect 204294 77932 204350 77988
rect 204418 77932 204474 77988
rect 204294 77808 204350 77864
rect 204418 77808 204474 77864
rect 219294 79952 219350 80008
rect 219418 79952 219474 80008
rect 219294 79828 219350 79884
rect 219418 79828 219474 79884
rect 219294 79704 219350 79760
rect 219418 79704 219474 79760
rect 219294 79580 219350 79636
rect 219418 79580 219474 79636
rect 219294 79456 219350 79512
rect 219418 79456 219474 79512
rect 219294 79332 219350 79388
rect 219418 79332 219474 79388
rect 219294 79208 219350 79264
rect 219418 79208 219474 79264
rect 214294 78552 214350 78608
rect 214418 78552 214474 78608
rect 214294 78428 214350 78484
rect 214418 78428 214474 78484
rect 214294 78304 214350 78360
rect 214418 78304 214474 78360
rect 214294 78180 214350 78236
rect 214418 78180 214474 78236
rect 214294 78056 214350 78112
rect 214418 78056 214474 78112
rect 214294 77932 214350 77988
rect 214418 77932 214474 77988
rect 214294 77808 214350 77864
rect 214418 77808 214474 77864
rect 229294 79952 229350 80008
rect 229418 79952 229474 80008
rect 229294 79828 229350 79884
rect 229418 79828 229474 79884
rect 229294 79704 229350 79760
rect 229418 79704 229474 79760
rect 229294 79580 229350 79636
rect 229418 79580 229474 79636
rect 229294 79456 229350 79512
rect 229418 79456 229474 79512
rect 229294 79332 229350 79388
rect 229418 79332 229474 79388
rect 229294 79208 229350 79264
rect 229418 79208 229474 79264
rect 224294 78552 224350 78608
rect 224418 78552 224474 78608
rect 224294 78428 224350 78484
rect 224418 78428 224474 78484
rect 224294 78304 224350 78360
rect 224418 78304 224474 78360
rect 224294 78180 224350 78236
rect 224418 78180 224474 78236
rect 224294 78056 224350 78112
rect 224418 78056 224474 78112
rect 224294 77932 224350 77988
rect 224418 77932 224474 77988
rect 224294 77808 224350 77864
rect 224418 77808 224474 77864
rect 239294 79952 239350 80008
rect 239418 79952 239474 80008
rect 239294 79828 239350 79884
rect 239418 79828 239474 79884
rect 239294 79704 239350 79760
rect 239418 79704 239474 79760
rect 239294 79580 239350 79636
rect 239418 79580 239474 79636
rect 239294 79456 239350 79512
rect 239418 79456 239474 79512
rect 239294 79332 239350 79388
rect 239418 79332 239474 79388
rect 239294 79208 239350 79264
rect 239418 79208 239474 79264
rect 234294 78552 234350 78608
rect 234418 78552 234474 78608
rect 234294 78428 234350 78484
rect 234418 78428 234474 78484
rect 234294 78304 234350 78360
rect 234418 78304 234474 78360
rect 234294 78180 234350 78236
rect 234418 78180 234474 78236
rect 234294 78056 234350 78112
rect 234418 78056 234474 78112
rect 234294 77932 234350 77988
rect 234418 77932 234474 77988
rect 234294 77808 234350 77864
rect 234418 77808 234474 77864
rect 249294 79952 249350 80008
rect 249418 79952 249474 80008
rect 249294 79828 249350 79884
rect 249418 79828 249474 79884
rect 249294 79704 249350 79760
rect 249418 79704 249474 79760
rect 249294 79580 249350 79636
rect 249418 79580 249474 79636
rect 249294 79456 249350 79512
rect 249418 79456 249474 79512
rect 249294 79332 249350 79388
rect 249418 79332 249474 79388
rect 249294 79208 249350 79264
rect 249418 79208 249474 79264
rect 244294 78552 244350 78608
rect 244418 78552 244474 78608
rect 244294 78428 244350 78484
rect 244418 78428 244474 78484
rect 244294 78304 244350 78360
rect 244418 78304 244474 78360
rect 244294 78180 244350 78236
rect 244418 78180 244474 78236
rect 244294 78056 244350 78112
rect 244418 78056 244474 78112
rect 244294 77932 244350 77988
rect 244418 77932 244474 77988
rect 244294 77808 244350 77864
rect 244418 77808 244474 77864
rect 259294 79952 259350 80008
rect 259418 79952 259474 80008
rect 259294 79828 259350 79884
rect 259418 79828 259474 79884
rect 259294 79704 259350 79760
rect 259418 79704 259474 79760
rect 259294 79580 259350 79636
rect 259418 79580 259474 79636
rect 259294 79456 259350 79512
rect 259418 79456 259474 79512
rect 259294 79332 259350 79388
rect 259418 79332 259474 79388
rect 259294 79208 259350 79264
rect 259418 79208 259474 79264
rect 254294 78552 254350 78608
rect 254418 78552 254474 78608
rect 254294 78428 254350 78484
rect 254418 78428 254474 78484
rect 254294 78304 254350 78360
rect 254418 78304 254474 78360
rect 254294 78180 254350 78236
rect 254418 78180 254474 78236
rect 254294 78056 254350 78112
rect 254418 78056 254474 78112
rect 254294 77932 254350 77988
rect 254418 77932 254474 77988
rect 254294 77808 254350 77864
rect 254418 77808 254474 77864
rect 269294 79952 269350 80008
rect 269418 79952 269474 80008
rect 269294 79828 269350 79884
rect 269418 79828 269474 79884
rect 269294 79704 269350 79760
rect 269418 79704 269474 79760
rect 269294 79580 269350 79636
rect 269418 79580 269474 79636
rect 269294 79456 269350 79512
rect 269418 79456 269474 79512
rect 269294 79332 269350 79388
rect 269418 79332 269474 79388
rect 269294 79208 269350 79264
rect 269418 79208 269474 79264
rect 272330 79952 272386 80008
rect 272454 79952 272510 80008
rect 272578 79952 272634 80008
rect 272702 79952 272758 80008
rect 272826 79952 272882 80008
rect 272950 79952 273006 80008
rect 273074 79952 273130 80008
rect 273198 79952 273254 80008
rect 273322 79952 273378 80008
rect 273446 79952 273502 80008
rect 273570 79952 273626 80008
rect 273694 79952 273750 80008
rect 273818 79952 273874 80008
rect 273942 79952 273998 80008
rect 274066 79952 274122 80008
rect 272330 79828 272386 79884
rect 272454 79828 272510 79884
rect 272578 79828 272634 79884
rect 272702 79828 272758 79884
rect 272826 79828 272882 79884
rect 272950 79828 273006 79884
rect 273074 79828 273130 79884
rect 273198 79828 273254 79884
rect 273322 79828 273378 79884
rect 273446 79828 273502 79884
rect 273570 79828 273626 79884
rect 273694 79828 273750 79884
rect 273818 79828 273874 79884
rect 273942 79828 273998 79884
rect 274066 79828 274122 79884
rect 272330 79704 272386 79760
rect 272454 79704 272510 79760
rect 272578 79704 272634 79760
rect 272702 79704 272758 79760
rect 272826 79704 272882 79760
rect 272950 79704 273006 79760
rect 273074 79704 273130 79760
rect 273198 79704 273254 79760
rect 273322 79704 273378 79760
rect 273446 79704 273502 79760
rect 273570 79704 273626 79760
rect 273694 79704 273750 79760
rect 273818 79704 273874 79760
rect 273942 79704 273998 79760
rect 274066 79704 274122 79760
rect 272330 79580 272386 79636
rect 272454 79580 272510 79636
rect 272578 79580 272634 79636
rect 272702 79580 272758 79636
rect 272826 79580 272882 79636
rect 272950 79580 273006 79636
rect 273074 79580 273130 79636
rect 273198 79580 273254 79636
rect 273322 79580 273378 79636
rect 273446 79580 273502 79636
rect 273570 79580 273626 79636
rect 273694 79580 273750 79636
rect 273818 79580 273874 79636
rect 273942 79580 273998 79636
rect 274066 79580 274122 79636
rect 272330 79456 272386 79512
rect 272454 79456 272510 79512
rect 272578 79456 272634 79512
rect 272702 79456 272758 79512
rect 272826 79456 272882 79512
rect 272950 79456 273006 79512
rect 273074 79456 273130 79512
rect 273198 79456 273254 79512
rect 273322 79456 273378 79512
rect 273446 79456 273502 79512
rect 273570 79456 273626 79512
rect 273694 79456 273750 79512
rect 273818 79456 273874 79512
rect 273942 79456 273998 79512
rect 274066 79456 274122 79512
rect 272330 79332 272386 79388
rect 272454 79332 272510 79388
rect 272578 79332 272634 79388
rect 272702 79332 272758 79388
rect 272826 79332 272882 79388
rect 272950 79332 273006 79388
rect 273074 79332 273130 79388
rect 273198 79332 273254 79388
rect 273322 79332 273378 79388
rect 273446 79332 273502 79388
rect 273570 79332 273626 79388
rect 273694 79332 273750 79388
rect 273818 79332 273874 79388
rect 273942 79332 273998 79388
rect 274066 79332 274122 79388
rect 272330 79208 272386 79264
rect 272454 79208 272510 79264
rect 272578 79208 272634 79264
rect 272702 79208 272758 79264
rect 272826 79208 272882 79264
rect 272950 79208 273006 79264
rect 273074 79208 273130 79264
rect 273198 79208 273254 79264
rect 273322 79208 273378 79264
rect 273446 79208 273502 79264
rect 273570 79208 273626 79264
rect 273694 79208 273750 79264
rect 273818 79208 273874 79264
rect 273942 79208 273998 79264
rect 274066 79208 274122 79264
rect 264294 78552 264350 78608
rect 264418 78552 264474 78608
rect 264294 78428 264350 78484
rect 264418 78428 264474 78484
rect 264294 78304 264350 78360
rect 264418 78304 264474 78360
rect 264294 78180 264350 78236
rect 264418 78180 264474 78236
rect 264294 78056 264350 78112
rect 264418 78056 264474 78112
rect 264294 77932 264350 77988
rect 264418 77932 264474 77988
rect 264294 77808 264350 77864
rect 264418 77808 264474 77864
rect 274810 79952 274866 80008
rect 274934 79952 274990 80008
rect 275058 79952 275114 80008
rect 275182 79952 275238 80008
rect 275306 79952 275362 80008
rect 275430 79952 275486 80008
rect 275554 79952 275610 80008
rect 275678 79952 275734 80008
rect 275802 79952 275858 80008
rect 275926 79952 275982 80008
rect 276050 79952 276106 80008
rect 276174 79952 276230 80008
rect 276298 79952 276354 80008
rect 276422 79952 276478 80008
rect 276546 79952 276602 80008
rect 276670 79952 276726 80008
rect 274810 79828 274866 79884
rect 274934 79828 274990 79884
rect 275058 79828 275114 79884
rect 275182 79828 275238 79884
rect 275306 79828 275362 79884
rect 275430 79828 275486 79884
rect 275554 79828 275610 79884
rect 275678 79828 275734 79884
rect 275802 79828 275858 79884
rect 275926 79828 275982 79884
rect 276050 79828 276106 79884
rect 276174 79828 276230 79884
rect 276298 79828 276354 79884
rect 276422 79828 276478 79884
rect 276546 79828 276602 79884
rect 276670 79828 276726 79884
rect 274810 79704 274866 79760
rect 274934 79704 274990 79760
rect 275058 79704 275114 79760
rect 275182 79704 275238 79760
rect 275306 79704 275362 79760
rect 275430 79704 275486 79760
rect 275554 79704 275610 79760
rect 275678 79704 275734 79760
rect 275802 79704 275858 79760
rect 275926 79704 275982 79760
rect 276050 79704 276106 79760
rect 276174 79704 276230 79760
rect 276298 79704 276354 79760
rect 276422 79704 276478 79760
rect 276546 79704 276602 79760
rect 276670 79704 276726 79760
rect 274810 79580 274866 79636
rect 274934 79580 274990 79636
rect 275058 79580 275114 79636
rect 275182 79580 275238 79636
rect 275306 79580 275362 79636
rect 275430 79580 275486 79636
rect 275554 79580 275610 79636
rect 275678 79580 275734 79636
rect 275802 79580 275858 79636
rect 275926 79580 275982 79636
rect 276050 79580 276106 79636
rect 276174 79580 276230 79636
rect 276298 79580 276354 79636
rect 276422 79580 276478 79636
rect 276546 79580 276602 79636
rect 276670 79580 276726 79636
rect 274810 79456 274866 79512
rect 274934 79456 274990 79512
rect 275058 79456 275114 79512
rect 275182 79456 275238 79512
rect 275306 79456 275362 79512
rect 275430 79456 275486 79512
rect 275554 79456 275610 79512
rect 275678 79456 275734 79512
rect 275802 79456 275858 79512
rect 275926 79456 275982 79512
rect 276050 79456 276106 79512
rect 276174 79456 276230 79512
rect 276298 79456 276354 79512
rect 276422 79456 276478 79512
rect 276546 79456 276602 79512
rect 276670 79456 276726 79512
rect 274810 79332 274866 79388
rect 274934 79332 274990 79388
rect 275058 79332 275114 79388
rect 275182 79332 275238 79388
rect 275306 79332 275362 79388
rect 275430 79332 275486 79388
rect 275554 79332 275610 79388
rect 275678 79332 275734 79388
rect 275802 79332 275858 79388
rect 275926 79332 275982 79388
rect 276050 79332 276106 79388
rect 276174 79332 276230 79388
rect 276298 79332 276354 79388
rect 276422 79332 276478 79388
rect 276546 79332 276602 79388
rect 276670 79332 276726 79388
rect 274810 79208 274866 79264
rect 274934 79208 274990 79264
rect 275058 79208 275114 79264
rect 275182 79208 275238 79264
rect 275306 79208 275362 79264
rect 275430 79208 275486 79264
rect 275554 79208 275610 79264
rect 275678 79208 275734 79264
rect 275802 79208 275858 79264
rect 275926 79208 275982 79264
rect 276050 79208 276106 79264
rect 276174 79208 276230 79264
rect 276298 79208 276354 79264
rect 276422 79208 276478 79264
rect 276546 79208 276602 79264
rect 276670 79208 276726 79264
rect 277180 79952 277236 80008
rect 277304 79952 277360 80008
rect 277428 79952 277484 80008
rect 277552 79952 277608 80008
rect 277676 79952 277732 80008
rect 277800 79952 277856 80008
rect 277924 79952 277980 80008
rect 278048 79952 278104 80008
rect 278172 79952 278228 80008
rect 278296 79952 278352 80008
rect 278420 79952 278476 80008
rect 278544 79952 278600 80008
rect 278668 79952 278724 80008
rect 278792 79952 278848 80008
rect 278916 79952 278972 80008
rect 279040 79952 279096 80008
rect 277180 79828 277236 79884
rect 277304 79828 277360 79884
rect 277428 79828 277484 79884
rect 277552 79828 277608 79884
rect 277676 79828 277732 79884
rect 277800 79828 277856 79884
rect 277924 79828 277980 79884
rect 278048 79828 278104 79884
rect 278172 79828 278228 79884
rect 278296 79828 278352 79884
rect 278420 79828 278476 79884
rect 278544 79828 278600 79884
rect 278668 79828 278724 79884
rect 278792 79828 278848 79884
rect 278916 79828 278972 79884
rect 279040 79828 279096 79884
rect 277180 79704 277236 79760
rect 277304 79704 277360 79760
rect 277428 79704 277484 79760
rect 277552 79704 277608 79760
rect 277676 79704 277732 79760
rect 277800 79704 277856 79760
rect 277924 79704 277980 79760
rect 278048 79704 278104 79760
rect 278172 79704 278228 79760
rect 278296 79704 278352 79760
rect 278420 79704 278476 79760
rect 278544 79704 278600 79760
rect 278668 79704 278724 79760
rect 278792 79704 278848 79760
rect 278916 79704 278972 79760
rect 279040 79704 279096 79760
rect 277180 79580 277236 79636
rect 277304 79580 277360 79636
rect 277428 79580 277484 79636
rect 277552 79580 277608 79636
rect 277676 79580 277732 79636
rect 277800 79580 277856 79636
rect 277924 79580 277980 79636
rect 278048 79580 278104 79636
rect 278172 79580 278228 79636
rect 278296 79580 278352 79636
rect 278420 79580 278476 79636
rect 278544 79580 278600 79636
rect 278668 79580 278724 79636
rect 278792 79580 278848 79636
rect 278916 79580 278972 79636
rect 279040 79580 279096 79636
rect 277180 79456 277236 79512
rect 277304 79456 277360 79512
rect 277428 79456 277484 79512
rect 277552 79456 277608 79512
rect 277676 79456 277732 79512
rect 277800 79456 277856 79512
rect 277924 79456 277980 79512
rect 278048 79456 278104 79512
rect 278172 79456 278228 79512
rect 278296 79456 278352 79512
rect 278420 79456 278476 79512
rect 278544 79456 278600 79512
rect 278668 79456 278724 79512
rect 278792 79456 278848 79512
rect 278916 79456 278972 79512
rect 279040 79456 279096 79512
rect 277180 79332 277236 79388
rect 277304 79332 277360 79388
rect 277428 79332 277484 79388
rect 277552 79332 277608 79388
rect 277676 79332 277732 79388
rect 277800 79332 277856 79388
rect 277924 79332 277980 79388
rect 278048 79332 278104 79388
rect 278172 79332 278228 79388
rect 278296 79332 278352 79388
rect 278420 79332 278476 79388
rect 278544 79332 278600 79388
rect 278668 79332 278724 79388
rect 278792 79332 278848 79388
rect 278916 79332 278972 79388
rect 279040 79332 279096 79388
rect 277180 79208 277236 79264
rect 277304 79208 277360 79264
rect 277428 79208 277484 79264
rect 277552 79208 277608 79264
rect 277676 79208 277732 79264
rect 277800 79208 277856 79264
rect 277924 79208 277980 79264
rect 278048 79208 278104 79264
rect 278172 79208 278228 79264
rect 278296 79208 278352 79264
rect 278420 79208 278476 79264
rect 278544 79208 278600 79264
rect 278668 79208 278724 79264
rect 278792 79208 278848 79264
rect 278916 79208 278972 79264
rect 279040 79208 279096 79264
rect 279886 79952 279942 80008
rect 280010 79952 280066 80008
rect 280134 79952 280190 80008
rect 280258 79952 280314 80008
rect 280382 79952 280438 80008
rect 280506 79952 280562 80008
rect 280630 79952 280686 80008
rect 280754 79952 280810 80008
rect 280878 79952 280934 80008
rect 281002 79952 281058 80008
rect 281126 79952 281182 80008
rect 281250 79952 281306 80008
rect 281374 79952 281430 80008
rect 281498 79952 281554 80008
rect 281622 79952 281678 80008
rect 281746 79952 281802 80008
rect 279886 79828 279942 79884
rect 280010 79828 280066 79884
rect 280134 79828 280190 79884
rect 280258 79828 280314 79884
rect 280382 79828 280438 79884
rect 280506 79828 280562 79884
rect 280630 79828 280686 79884
rect 280754 79828 280810 79884
rect 280878 79828 280934 79884
rect 281002 79828 281058 79884
rect 281126 79828 281182 79884
rect 281250 79828 281306 79884
rect 281374 79828 281430 79884
rect 281498 79828 281554 79884
rect 281622 79828 281678 79884
rect 281746 79828 281802 79884
rect 279886 79704 279942 79760
rect 280010 79704 280066 79760
rect 280134 79704 280190 79760
rect 280258 79704 280314 79760
rect 280382 79704 280438 79760
rect 280506 79704 280562 79760
rect 280630 79704 280686 79760
rect 280754 79704 280810 79760
rect 280878 79704 280934 79760
rect 281002 79704 281058 79760
rect 281126 79704 281182 79760
rect 281250 79704 281306 79760
rect 281374 79704 281430 79760
rect 281498 79704 281554 79760
rect 281622 79704 281678 79760
rect 281746 79704 281802 79760
rect 279886 79580 279942 79636
rect 280010 79580 280066 79636
rect 280134 79580 280190 79636
rect 280258 79580 280314 79636
rect 280382 79580 280438 79636
rect 280506 79580 280562 79636
rect 280630 79580 280686 79636
rect 280754 79580 280810 79636
rect 280878 79580 280934 79636
rect 281002 79580 281058 79636
rect 281126 79580 281182 79636
rect 281250 79580 281306 79636
rect 281374 79580 281430 79636
rect 281498 79580 281554 79636
rect 281622 79580 281678 79636
rect 281746 79580 281802 79636
rect 279886 79456 279942 79512
rect 280010 79456 280066 79512
rect 280134 79456 280190 79512
rect 280258 79456 280314 79512
rect 280382 79456 280438 79512
rect 280506 79456 280562 79512
rect 280630 79456 280686 79512
rect 280754 79456 280810 79512
rect 280878 79456 280934 79512
rect 281002 79456 281058 79512
rect 281126 79456 281182 79512
rect 281250 79456 281306 79512
rect 281374 79456 281430 79512
rect 281498 79456 281554 79512
rect 281622 79456 281678 79512
rect 281746 79456 281802 79512
rect 279886 79332 279942 79388
rect 280010 79332 280066 79388
rect 280134 79332 280190 79388
rect 280258 79332 280314 79388
rect 280382 79332 280438 79388
rect 280506 79332 280562 79388
rect 280630 79332 280686 79388
rect 280754 79332 280810 79388
rect 280878 79332 280934 79388
rect 281002 79332 281058 79388
rect 281126 79332 281182 79388
rect 281250 79332 281306 79388
rect 281374 79332 281430 79388
rect 281498 79332 281554 79388
rect 281622 79332 281678 79388
rect 281746 79332 281802 79388
rect 279886 79208 279942 79264
rect 280010 79208 280066 79264
rect 280134 79208 280190 79264
rect 280258 79208 280314 79264
rect 280382 79208 280438 79264
rect 280506 79208 280562 79264
rect 280630 79208 280686 79264
rect 280754 79208 280810 79264
rect 280878 79208 280934 79264
rect 281002 79208 281058 79264
rect 281126 79208 281182 79264
rect 281250 79208 281306 79264
rect 281374 79208 281430 79264
rect 281498 79208 281554 79264
rect 281622 79208 281678 79264
rect 281746 79208 281802 79264
rect 282256 79952 282312 80008
rect 282380 79952 282436 80008
rect 282504 79952 282560 80008
rect 282628 79952 282684 80008
rect 282752 79952 282808 80008
rect 282876 79952 282932 80008
rect 283000 79952 283056 80008
rect 283124 79952 283180 80008
rect 283248 79952 283304 80008
rect 283372 79952 283428 80008
rect 283496 79952 283552 80008
rect 283620 79952 283676 80008
rect 283744 79952 283800 80008
rect 283868 79952 283924 80008
rect 283992 79952 284048 80008
rect 284116 79952 284172 80008
rect 282256 79828 282312 79884
rect 282380 79828 282436 79884
rect 282504 79828 282560 79884
rect 282628 79828 282684 79884
rect 282752 79828 282808 79884
rect 282876 79828 282932 79884
rect 283000 79828 283056 79884
rect 283124 79828 283180 79884
rect 283248 79828 283304 79884
rect 283372 79828 283428 79884
rect 283496 79828 283552 79884
rect 283620 79828 283676 79884
rect 283744 79828 283800 79884
rect 283868 79828 283924 79884
rect 283992 79828 284048 79884
rect 284116 79828 284172 79884
rect 282256 79704 282312 79760
rect 282380 79704 282436 79760
rect 282504 79704 282560 79760
rect 282628 79704 282684 79760
rect 282752 79704 282808 79760
rect 282876 79704 282932 79760
rect 283000 79704 283056 79760
rect 283124 79704 283180 79760
rect 283248 79704 283304 79760
rect 283372 79704 283428 79760
rect 283496 79704 283552 79760
rect 283620 79704 283676 79760
rect 283744 79704 283800 79760
rect 283868 79704 283924 79760
rect 283992 79704 284048 79760
rect 284116 79704 284172 79760
rect 282256 79580 282312 79636
rect 282380 79580 282436 79636
rect 282504 79580 282560 79636
rect 282628 79580 282684 79636
rect 282752 79580 282808 79636
rect 282876 79580 282932 79636
rect 283000 79580 283056 79636
rect 283124 79580 283180 79636
rect 283248 79580 283304 79636
rect 283372 79580 283428 79636
rect 283496 79580 283552 79636
rect 283620 79580 283676 79636
rect 283744 79580 283800 79636
rect 283868 79580 283924 79636
rect 283992 79580 284048 79636
rect 284116 79580 284172 79636
rect 282256 79456 282312 79512
rect 282380 79456 282436 79512
rect 282504 79456 282560 79512
rect 282628 79456 282684 79512
rect 282752 79456 282808 79512
rect 282876 79456 282932 79512
rect 283000 79456 283056 79512
rect 283124 79456 283180 79512
rect 283248 79456 283304 79512
rect 283372 79456 283428 79512
rect 283496 79456 283552 79512
rect 283620 79456 283676 79512
rect 283744 79456 283800 79512
rect 283868 79456 283924 79512
rect 283992 79456 284048 79512
rect 284116 79456 284172 79512
rect 282256 79332 282312 79388
rect 282380 79332 282436 79388
rect 282504 79332 282560 79388
rect 282628 79332 282684 79388
rect 282752 79332 282808 79388
rect 282876 79332 282932 79388
rect 283000 79332 283056 79388
rect 283124 79332 283180 79388
rect 283248 79332 283304 79388
rect 283372 79332 283428 79388
rect 283496 79332 283552 79388
rect 283620 79332 283676 79388
rect 283744 79332 283800 79388
rect 283868 79332 283924 79388
rect 283992 79332 284048 79388
rect 284116 79332 284172 79388
rect 282256 79208 282312 79264
rect 282380 79208 282436 79264
rect 282504 79208 282560 79264
rect 282628 79208 282684 79264
rect 282752 79208 282808 79264
rect 282876 79208 282932 79264
rect 283000 79208 283056 79264
rect 283124 79208 283180 79264
rect 283248 79208 283304 79264
rect 283372 79208 283428 79264
rect 283496 79208 283552 79264
rect 283620 79208 283676 79264
rect 283744 79208 283800 79264
rect 283868 79208 283924 79264
rect 283992 79208 284048 79264
rect 284116 79208 284172 79264
rect 284860 79952 284916 80008
rect 284984 79952 285040 80008
rect 285108 79952 285164 80008
rect 285232 79952 285288 80008
rect 285356 79952 285412 80008
rect 285480 79952 285536 80008
rect 285604 79952 285660 80008
rect 285728 79952 285784 80008
rect 285852 79952 285908 80008
rect 285976 79952 286032 80008
rect 286100 79952 286156 80008
rect 286224 79952 286280 80008
rect 286348 79952 286404 80008
rect 286472 79952 286528 80008
rect 286596 79952 286652 80008
rect 284860 79828 284916 79884
rect 284984 79828 285040 79884
rect 285108 79828 285164 79884
rect 285232 79828 285288 79884
rect 285356 79828 285412 79884
rect 285480 79828 285536 79884
rect 285604 79828 285660 79884
rect 285728 79828 285784 79884
rect 285852 79828 285908 79884
rect 285976 79828 286032 79884
rect 286100 79828 286156 79884
rect 286224 79828 286280 79884
rect 286348 79828 286404 79884
rect 286472 79828 286528 79884
rect 286596 79828 286652 79884
rect 284860 79704 284916 79760
rect 284984 79704 285040 79760
rect 285108 79704 285164 79760
rect 285232 79704 285288 79760
rect 285356 79704 285412 79760
rect 285480 79704 285536 79760
rect 285604 79704 285660 79760
rect 285728 79704 285784 79760
rect 285852 79704 285908 79760
rect 285976 79704 286032 79760
rect 286100 79704 286156 79760
rect 286224 79704 286280 79760
rect 286348 79704 286404 79760
rect 286472 79704 286528 79760
rect 286596 79704 286652 79760
rect 284860 79580 284916 79636
rect 284984 79580 285040 79636
rect 285108 79580 285164 79636
rect 285232 79580 285288 79636
rect 285356 79580 285412 79636
rect 285480 79580 285536 79636
rect 285604 79580 285660 79636
rect 285728 79580 285784 79636
rect 285852 79580 285908 79636
rect 285976 79580 286032 79636
rect 286100 79580 286156 79636
rect 286224 79580 286280 79636
rect 286348 79580 286404 79636
rect 286472 79580 286528 79636
rect 286596 79580 286652 79636
rect 284860 79456 284916 79512
rect 284984 79456 285040 79512
rect 285108 79456 285164 79512
rect 285232 79456 285288 79512
rect 285356 79456 285412 79512
rect 285480 79456 285536 79512
rect 285604 79456 285660 79512
rect 285728 79456 285784 79512
rect 285852 79456 285908 79512
rect 285976 79456 286032 79512
rect 286100 79456 286156 79512
rect 286224 79456 286280 79512
rect 286348 79456 286404 79512
rect 286472 79456 286528 79512
rect 286596 79456 286652 79512
rect 284860 79332 284916 79388
rect 284984 79332 285040 79388
rect 285108 79332 285164 79388
rect 285232 79332 285288 79388
rect 285356 79332 285412 79388
rect 285480 79332 285536 79388
rect 285604 79332 285660 79388
rect 285728 79332 285784 79388
rect 285852 79332 285908 79388
rect 285976 79332 286032 79388
rect 286100 79332 286156 79388
rect 286224 79332 286280 79388
rect 286348 79332 286404 79388
rect 286472 79332 286528 79388
rect 286596 79332 286652 79388
rect 284860 79208 284916 79264
rect 284984 79208 285040 79264
rect 285108 79208 285164 79264
rect 285232 79208 285288 79264
rect 285356 79208 285412 79264
rect 285480 79208 285536 79264
rect 285604 79208 285660 79264
rect 285728 79208 285784 79264
rect 285852 79208 285908 79264
rect 285976 79208 286032 79264
rect 286100 79208 286156 79264
rect 286224 79208 286280 79264
rect 286348 79208 286404 79264
rect 286472 79208 286528 79264
rect 286596 79208 286652 79264
rect 289294 79952 289350 80008
rect 289418 79952 289474 80008
rect 289294 79828 289350 79884
rect 289418 79828 289474 79884
rect 289294 79704 289350 79760
rect 289418 79704 289474 79760
rect 289294 79580 289350 79636
rect 289418 79580 289474 79636
rect 289294 79456 289350 79512
rect 289418 79456 289474 79512
rect 289294 79332 289350 79388
rect 289418 79332 289474 79388
rect 289294 79208 289350 79264
rect 289418 79208 289474 79264
rect 299294 79952 299350 80008
rect 299418 79952 299474 80008
rect 299294 79828 299350 79884
rect 299418 79828 299474 79884
rect 299294 79704 299350 79760
rect 299418 79704 299474 79760
rect 299294 79580 299350 79636
rect 299418 79580 299474 79636
rect 299294 79456 299350 79512
rect 299418 79456 299474 79512
rect 299294 79332 299350 79388
rect 299418 79332 299474 79388
rect 299294 79208 299350 79264
rect 299418 79208 299474 79264
rect 294294 78552 294350 78608
rect 294418 78552 294474 78608
rect 294294 78428 294350 78484
rect 294418 78428 294474 78484
rect 294294 78304 294350 78360
rect 294418 78304 294474 78360
rect 294294 78180 294350 78236
rect 294418 78180 294474 78236
rect 294294 78056 294350 78112
rect 294418 78056 294474 78112
rect 294294 77932 294350 77988
rect 294418 77932 294474 77988
rect 294294 77808 294350 77864
rect 294418 77808 294474 77864
rect 309294 79952 309350 80008
rect 309418 79952 309474 80008
rect 309294 79828 309350 79884
rect 309418 79828 309474 79884
rect 309294 79704 309350 79760
rect 309418 79704 309474 79760
rect 309294 79580 309350 79636
rect 309418 79580 309474 79636
rect 309294 79456 309350 79512
rect 309418 79456 309474 79512
rect 309294 79332 309350 79388
rect 309418 79332 309474 79388
rect 309294 79208 309350 79264
rect 309418 79208 309474 79264
rect 304294 78552 304350 78608
rect 304418 78552 304474 78608
rect 304294 78428 304350 78484
rect 304418 78428 304474 78484
rect 304294 78304 304350 78360
rect 304418 78304 304474 78360
rect 304294 78180 304350 78236
rect 304418 78180 304474 78236
rect 304294 78056 304350 78112
rect 304418 78056 304474 78112
rect 304294 77932 304350 77988
rect 304418 77932 304474 77988
rect 304294 77808 304350 77864
rect 304418 77808 304474 77864
rect 319294 79952 319350 80008
rect 319418 79952 319474 80008
rect 319294 79828 319350 79884
rect 319418 79828 319474 79884
rect 319294 79704 319350 79760
rect 319418 79704 319474 79760
rect 319294 79580 319350 79636
rect 319418 79580 319474 79636
rect 319294 79456 319350 79512
rect 319418 79456 319474 79512
rect 319294 79332 319350 79388
rect 319418 79332 319474 79388
rect 319294 79208 319350 79264
rect 319418 79208 319474 79264
rect 314294 78552 314350 78608
rect 314418 78552 314474 78608
rect 314294 78428 314350 78484
rect 314418 78428 314474 78484
rect 314294 78304 314350 78360
rect 314418 78304 314474 78360
rect 314294 78180 314350 78236
rect 314418 78180 314474 78236
rect 314294 78056 314350 78112
rect 314418 78056 314474 78112
rect 314294 77932 314350 77988
rect 314418 77932 314474 77988
rect 314294 77808 314350 77864
rect 314418 77808 314474 77864
rect 329294 79952 329350 80008
rect 329418 79952 329474 80008
rect 329294 79828 329350 79884
rect 329418 79828 329474 79884
rect 329294 79704 329350 79760
rect 329418 79704 329474 79760
rect 329294 79580 329350 79636
rect 329418 79580 329474 79636
rect 329294 79456 329350 79512
rect 329418 79456 329474 79512
rect 329294 79332 329350 79388
rect 329418 79332 329474 79388
rect 329294 79208 329350 79264
rect 329418 79208 329474 79264
rect 324294 78552 324350 78608
rect 324418 78552 324474 78608
rect 324294 78428 324350 78484
rect 324418 78428 324474 78484
rect 324294 78304 324350 78360
rect 324418 78304 324474 78360
rect 324294 78180 324350 78236
rect 324418 78180 324474 78236
rect 324294 78056 324350 78112
rect 324418 78056 324474 78112
rect 324294 77932 324350 77988
rect 324418 77932 324474 77988
rect 324294 77808 324350 77864
rect 324418 77808 324474 77864
rect 339294 79952 339350 80008
rect 339418 79952 339474 80008
rect 339294 79828 339350 79884
rect 339418 79828 339474 79884
rect 339294 79704 339350 79760
rect 339418 79704 339474 79760
rect 339294 79580 339350 79636
rect 339418 79580 339474 79636
rect 339294 79456 339350 79512
rect 339418 79456 339474 79512
rect 339294 79332 339350 79388
rect 339418 79332 339474 79388
rect 339294 79208 339350 79264
rect 339418 79208 339474 79264
rect 334294 78552 334350 78608
rect 334418 78552 334474 78608
rect 334294 78428 334350 78484
rect 334418 78428 334474 78484
rect 334294 78304 334350 78360
rect 334418 78304 334474 78360
rect 334294 78180 334350 78236
rect 334418 78180 334474 78236
rect 334294 78056 334350 78112
rect 334418 78056 334474 78112
rect 334294 77932 334350 77988
rect 334418 77932 334474 77988
rect 334294 77808 334350 77864
rect 334418 77808 334474 77864
rect 349294 79952 349350 80008
rect 349418 79952 349474 80008
rect 349294 79828 349350 79884
rect 349418 79828 349474 79884
rect 349294 79704 349350 79760
rect 349418 79704 349474 79760
rect 349294 79580 349350 79636
rect 349418 79580 349474 79636
rect 349294 79456 349350 79512
rect 349418 79456 349474 79512
rect 349294 79332 349350 79388
rect 349418 79332 349474 79388
rect 349294 79208 349350 79264
rect 349418 79208 349474 79264
rect 344294 78552 344350 78608
rect 344418 78552 344474 78608
rect 344294 78428 344350 78484
rect 344418 78428 344474 78484
rect 344294 78304 344350 78360
rect 344418 78304 344474 78360
rect 344294 78180 344350 78236
rect 344418 78180 344474 78236
rect 344294 78056 344350 78112
rect 344418 78056 344474 78112
rect 344294 77932 344350 77988
rect 344418 77932 344474 77988
rect 344294 77808 344350 77864
rect 344418 77808 344474 77864
rect 359294 79952 359350 80008
rect 359418 79952 359474 80008
rect 359294 79828 359350 79884
rect 359418 79828 359474 79884
rect 359294 79704 359350 79760
rect 359418 79704 359474 79760
rect 359294 79580 359350 79636
rect 359418 79580 359474 79636
rect 359294 79456 359350 79512
rect 359418 79456 359474 79512
rect 359294 79332 359350 79388
rect 359418 79332 359474 79388
rect 359294 79208 359350 79264
rect 359418 79208 359474 79264
rect 354294 78552 354350 78608
rect 354418 78552 354474 78608
rect 354294 78428 354350 78484
rect 354418 78428 354474 78484
rect 354294 78304 354350 78360
rect 354418 78304 354474 78360
rect 354294 78180 354350 78236
rect 354418 78180 354474 78236
rect 354294 78056 354350 78112
rect 354418 78056 354474 78112
rect 354294 77932 354350 77988
rect 354418 77932 354474 77988
rect 354294 77808 354350 77864
rect 354418 77808 354474 77864
rect 369294 79952 369350 80008
rect 369418 79952 369474 80008
rect 369294 79828 369350 79884
rect 369418 79828 369474 79884
rect 369294 79704 369350 79760
rect 369418 79704 369474 79760
rect 369294 79580 369350 79636
rect 369418 79580 369474 79636
rect 369294 79456 369350 79512
rect 369418 79456 369474 79512
rect 369294 79332 369350 79388
rect 369418 79332 369474 79388
rect 369294 79208 369350 79264
rect 369418 79208 369474 79264
rect 364294 78552 364350 78608
rect 364418 78552 364474 78608
rect 364294 78428 364350 78484
rect 364418 78428 364474 78484
rect 364294 78304 364350 78360
rect 364418 78304 364474 78360
rect 364294 78180 364350 78236
rect 364418 78180 364474 78236
rect 364294 78056 364350 78112
rect 364418 78056 364474 78112
rect 364294 77932 364350 77988
rect 364418 77932 364474 77988
rect 364294 77808 364350 77864
rect 364418 77808 364474 77864
rect 379294 79952 379350 80008
rect 379418 79952 379474 80008
rect 379294 79828 379350 79884
rect 379418 79828 379474 79884
rect 379294 79704 379350 79760
rect 379418 79704 379474 79760
rect 379294 79580 379350 79636
rect 379418 79580 379474 79636
rect 379294 79456 379350 79512
rect 379418 79456 379474 79512
rect 379294 79332 379350 79388
rect 379418 79332 379474 79388
rect 379294 79208 379350 79264
rect 379418 79208 379474 79264
rect 374294 78552 374350 78608
rect 374418 78552 374474 78608
rect 374294 78428 374350 78484
rect 374418 78428 374474 78484
rect 374294 78304 374350 78360
rect 374418 78304 374474 78360
rect 374294 78180 374350 78236
rect 374418 78180 374474 78236
rect 374294 78056 374350 78112
rect 374418 78056 374474 78112
rect 374294 77932 374350 77988
rect 374418 77932 374474 77988
rect 374294 77808 374350 77864
rect 374418 77808 374474 77864
rect 389294 79952 389350 80008
rect 389418 79952 389474 80008
rect 389294 79828 389350 79884
rect 389418 79828 389474 79884
rect 389294 79704 389350 79760
rect 389418 79704 389474 79760
rect 389294 79580 389350 79636
rect 389418 79580 389474 79636
rect 389294 79456 389350 79512
rect 389418 79456 389474 79512
rect 389294 79332 389350 79388
rect 389418 79332 389474 79388
rect 389294 79208 389350 79264
rect 389418 79208 389474 79264
rect 384294 78552 384350 78608
rect 384418 78552 384474 78608
rect 384294 78428 384350 78484
rect 384418 78428 384474 78484
rect 384294 78304 384350 78360
rect 384418 78304 384474 78360
rect 384294 78180 384350 78236
rect 384418 78180 384474 78236
rect 384294 78056 384350 78112
rect 384418 78056 384474 78112
rect 384294 77932 384350 77988
rect 384418 77932 384474 77988
rect 384294 77808 384350 77864
rect 384418 77808 384474 77864
rect 399294 79952 399350 80008
rect 399418 79952 399474 80008
rect 399294 79828 399350 79884
rect 399418 79828 399474 79884
rect 399294 79704 399350 79760
rect 399418 79704 399474 79760
rect 399294 79580 399350 79636
rect 399418 79580 399474 79636
rect 399294 79456 399350 79512
rect 399418 79456 399474 79512
rect 399294 79332 399350 79388
rect 399418 79332 399474 79388
rect 399294 79208 399350 79264
rect 399418 79208 399474 79264
rect 394294 78552 394350 78608
rect 394418 78552 394474 78608
rect 394294 78428 394350 78484
rect 394418 78428 394474 78484
rect 394294 78304 394350 78360
rect 394418 78304 394474 78360
rect 394294 78180 394350 78236
rect 394418 78180 394474 78236
rect 394294 78056 394350 78112
rect 394418 78056 394474 78112
rect 394294 77932 394350 77988
rect 394418 77932 394474 77988
rect 394294 77808 394350 77864
rect 394418 77808 394474 77864
rect 409294 79952 409350 80008
rect 409418 79952 409474 80008
rect 409294 79828 409350 79884
rect 409418 79828 409474 79884
rect 409294 79704 409350 79760
rect 409418 79704 409474 79760
rect 409294 79580 409350 79636
rect 409418 79580 409474 79636
rect 409294 79456 409350 79512
rect 409418 79456 409474 79512
rect 409294 79332 409350 79388
rect 409418 79332 409474 79388
rect 409294 79208 409350 79264
rect 409418 79208 409474 79264
rect 404294 78552 404350 78608
rect 404418 78552 404474 78608
rect 404294 78428 404350 78484
rect 404418 78428 404474 78484
rect 404294 78304 404350 78360
rect 404418 78304 404474 78360
rect 404294 78180 404350 78236
rect 404418 78180 404474 78236
rect 404294 78056 404350 78112
rect 404418 78056 404474 78112
rect 404294 77932 404350 77988
rect 404418 77932 404474 77988
rect 404294 77808 404350 77864
rect 404418 77808 404474 77864
rect 419294 79952 419350 80008
rect 419418 79952 419474 80008
rect 419294 79828 419350 79884
rect 419418 79828 419474 79884
rect 419294 79704 419350 79760
rect 419418 79704 419474 79760
rect 419294 79580 419350 79636
rect 419418 79580 419474 79636
rect 419294 79456 419350 79512
rect 419418 79456 419474 79512
rect 419294 79332 419350 79388
rect 419418 79332 419474 79388
rect 419294 79208 419350 79264
rect 419418 79208 419474 79264
rect 414294 78552 414350 78608
rect 414418 78552 414474 78608
rect 414294 78428 414350 78484
rect 414418 78428 414474 78484
rect 414294 78304 414350 78360
rect 414418 78304 414474 78360
rect 414294 78180 414350 78236
rect 414418 78180 414474 78236
rect 414294 78056 414350 78112
rect 414418 78056 414474 78112
rect 414294 77932 414350 77988
rect 414418 77932 414474 77988
rect 414294 77808 414350 77864
rect 414418 77808 414474 77864
rect 429294 79952 429350 80008
rect 429418 79952 429474 80008
rect 429294 79828 429350 79884
rect 429418 79828 429474 79884
rect 429294 79704 429350 79760
rect 429418 79704 429474 79760
rect 429294 79580 429350 79636
rect 429418 79580 429474 79636
rect 429294 79456 429350 79512
rect 429418 79456 429474 79512
rect 429294 79332 429350 79388
rect 429418 79332 429474 79388
rect 429294 79208 429350 79264
rect 429418 79208 429474 79264
rect 424294 78552 424350 78608
rect 424418 78552 424474 78608
rect 424294 78428 424350 78484
rect 424418 78428 424474 78484
rect 424294 78304 424350 78360
rect 424418 78304 424474 78360
rect 424294 78180 424350 78236
rect 424418 78180 424474 78236
rect 424294 78056 424350 78112
rect 424418 78056 424474 78112
rect 424294 77932 424350 77988
rect 424418 77932 424474 77988
rect 424294 77808 424350 77864
rect 424418 77808 424474 77864
rect 439294 79952 439350 80008
rect 439418 79952 439474 80008
rect 439294 79828 439350 79884
rect 439418 79828 439474 79884
rect 439294 79704 439350 79760
rect 439418 79704 439474 79760
rect 439294 79580 439350 79636
rect 439418 79580 439474 79636
rect 439294 79456 439350 79512
rect 439418 79456 439474 79512
rect 439294 79332 439350 79388
rect 439418 79332 439474 79388
rect 439294 79208 439350 79264
rect 439418 79208 439474 79264
rect 434294 78552 434350 78608
rect 434418 78552 434474 78608
rect 434294 78428 434350 78484
rect 434418 78428 434474 78484
rect 434294 78304 434350 78360
rect 434418 78304 434474 78360
rect 434294 78180 434350 78236
rect 434418 78180 434474 78236
rect 434294 78056 434350 78112
rect 434418 78056 434474 78112
rect 434294 77932 434350 77988
rect 434418 77932 434474 77988
rect 434294 77808 434350 77864
rect 434418 77808 434474 77864
rect 449294 79952 449350 80008
rect 449418 79952 449474 80008
rect 449294 79828 449350 79884
rect 449418 79828 449474 79884
rect 449294 79704 449350 79760
rect 449418 79704 449474 79760
rect 449294 79580 449350 79636
rect 449418 79580 449474 79636
rect 449294 79456 449350 79512
rect 449418 79456 449474 79512
rect 449294 79332 449350 79388
rect 449418 79332 449474 79388
rect 449294 79208 449350 79264
rect 449418 79208 449474 79264
rect 444294 78552 444350 78608
rect 444418 78552 444474 78608
rect 444294 78428 444350 78484
rect 444418 78428 444474 78484
rect 444294 78304 444350 78360
rect 444418 78304 444474 78360
rect 444294 78180 444350 78236
rect 444418 78180 444474 78236
rect 444294 78056 444350 78112
rect 444418 78056 444474 78112
rect 444294 77932 444350 77988
rect 444418 77932 444474 77988
rect 444294 77808 444350 77864
rect 444418 77808 444474 77864
rect 459294 79952 459350 80008
rect 459418 79952 459474 80008
rect 459294 79828 459350 79884
rect 459418 79828 459474 79884
rect 459294 79704 459350 79760
rect 459418 79704 459474 79760
rect 459294 79580 459350 79636
rect 459418 79580 459474 79636
rect 459294 79456 459350 79512
rect 459418 79456 459474 79512
rect 459294 79332 459350 79388
rect 459418 79332 459474 79388
rect 459294 79208 459350 79264
rect 459418 79208 459474 79264
rect 454294 78552 454350 78608
rect 454418 78552 454474 78608
rect 454294 78428 454350 78484
rect 454418 78428 454474 78484
rect 454294 78304 454350 78360
rect 454418 78304 454474 78360
rect 454294 78180 454350 78236
rect 454418 78180 454474 78236
rect 454294 78056 454350 78112
rect 454418 78056 454474 78112
rect 454294 77932 454350 77988
rect 454418 77932 454474 77988
rect 454294 77808 454350 77864
rect 454418 77808 454474 77864
rect 469294 79952 469350 80008
rect 469418 79952 469474 80008
rect 469294 79828 469350 79884
rect 469418 79828 469474 79884
rect 469294 79704 469350 79760
rect 469418 79704 469474 79760
rect 469294 79580 469350 79636
rect 469418 79580 469474 79636
rect 469294 79456 469350 79512
rect 469418 79456 469474 79512
rect 469294 79332 469350 79388
rect 469418 79332 469474 79388
rect 469294 79208 469350 79264
rect 469418 79208 469474 79264
rect 464294 78552 464350 78608
rect 464418 78552 464474 78608
rect 464294 78428 464350 78484
rect 464418 78428 464474 78484
rect 464294 78304 464350 78360
rect 464418 78304 464474 78360
rect 464294 78180 464350 78236
rect 464418 78180 464474 78236
rect 464294 78056 464350 78112
rect 464418 78056 464474 78112
rect 464294 77932 464350 77988
rect 464418 77932 464474 77988
rect 464294 77808 464350 77864
rect 464418 77808 464474 77864
rect 479294 79952 479350 80008
rect 479418 79952 479474 80008
rect 479294 79828 479350 79884
rect 479418 79828 479474 79884
rect 479294 79704 479350 79760
rect 479418 79704 479474 79760
rect 479294 79580 479350 79636
rect 479418 79580 479474 79636
rect 479294 79456 479350 79512
rect 479418 79456 479474 79512
rect 479294 79332 479350 79388
rect 479418 79332 479474 79388
rect 479294 79208 479350 79264
rect 479418 79208 479474 79264
rect 474294 78552 474350 78608
rect 474418 78552 474474 78608
rect 474294 78428 474350 78484
rect 474418 78428 474474 78484
rect 474294 78304 474350 78360
rect 474418 78304 474474 78360
rect 474294 78180 474350 78236
rect 474418 78180 474474 78236
rect 474294 78056 474350 78112
rect 474418 78056 474474 78112
rect 474294 77932 474350 77988
rect 474418 77932 474474 77988
rect 474294 77808 474350 77864
rect 474418 77808 474474 77864
rect 489294 79952 489350 80008
rect 489418 79952 489474 80008
rect 489294 79828 489350 79884
rect 489418 79828 489474 79884
rect 489294 79704 489350 79760
rect 489418 79704 489474 79760
rect 489294 79580 489350 79636
rect 489418 79580 489474 79636
rect 489294 79456 489350 79512
rect 489418 79456 489474 79512
rect 489294 79332 489350 79388
rect 489418 79332 489474 79388
rect 489294 79208 489350 79264
rect 489418 79208 489474 79264
rect 484294 78552 484350 78608
rect 484418 78552 484474 78608
rect 484294 78428 484350 78484
rect 484418 78428 484474 78484
rect 484294 78304 484350 78360
rect 484418 78304 484474 78360
rect 484294 78180 484350 78236
rect 484418 78180 484474 78236
rect 484294 78056 484350 78112
rect 484418 78056 484474 78112
rect 484294 77932 484350 77988
rect 484418 77932 484474 77988
rect 484294 77808 484350 77864
rect 484418 77808 484474 77864
rect 499294 79952 499350 80008
rect 499418 79952 499474 80008
rect 499294 79828 499350 79884
rect 499418 79828 499474 79884
rect 499294 79704 499350 79760
rect 499418 79704 499474 79760
rect 499294 79580 499350 79636
rect 499418 79580 499474 79636
rect 499294 79456 499350 79512
rect 499418 79456 499474 79512
rect 499294 79332 499350 79388
rect 499418 79332 499474 79388
rect 499294 79208 499350 79264
rect 499418 79208 499474 79264
rect 494294 78552 494350 78608
rect 494418 78552 494474 78608
rect 494294 78428 494350 78484
rect 494418 78428 494474 78484
rect 494294 78304 494350 78360
rect 494418 78304 494474 78360
rect 494294 78180 494350 78236
rect 494418 78180 494474 78236
rect 494294 78056 494350 78112
rect 494418 78056 494474 78112
rect 494294 77932 494350 77988
rect 494418 77932 494474 77988
rect 494294 77808 494350 77864
rect 494418 77808 494474 77864
rect 509294 79952 509350 80008
rect 509418 79952 509474 80008
rect 509294 79828 509350 79884
rect 509418 79828 509474 79884
rect 509294 79704 509350 79760
rect 509418 79704 509474 79760
rect 509294 79580 509350 79636
rect 509418 79580 509474 79636
rect 509294 79456 509350 79512
rect 509418 79456 509474 79512
rect 509294 79332 509350 79388
rect 509418 79332 509474 79388
rect 509294 79208 509350 79264
rect 509418 79208 509474 79264
rect 504294 78552 504350 78608
rect 504418 78552 504474 78608
rect 504294 78428 504350 78484
rect 504418 78428 504474 78484
rect 504294 78304 504350 78360
rect 504418 78304 504474 78360
rect 504294 78180 504350 78236
rect 504418 78180 504474 78236
rect 504294 78056 504350 78112
rect 504418 78056 504474 78112
rect 504294 77932 504350 77988
rect 504418 77932 504474 77988
rect 504294 77808 504350 77864
rect 504418 77808 504474 77864
rect 519294 79952 519350 80008
rect 519418 79952 519474 80008
rect 519294 79828 519350 79884
rect 519418 79828 519474 79884
rect 519294 79704 519350 79760
rect 519418 79704 519474 79760
rect 519294 79580 519350 79636
rect 519418 79580 519474 79636
rect 519294 79456 519350 79512
rect 519418 79456 519474 79512
rect 519294 79332 519350 79388
rect 519418 79332 519474 79388
rect 519294 79208 519350 79264
rect 519418 79208 519474 79264
rect 514294 78552 514350 78608
rect 514418 78552 514474 78608
rect 514294 78428 514350 78484
rect 514418 78428 514474 78484
rect 514294 78304 514350 78360
rect 514418 78304 514474 78360
rect 514294 78180 514350 78236
rect 514418 78180 514474 78236
rect 514294 78056 514350 78112
rect 514418 78056 514474 78112
rect 514294 77932 514350 77988
rect 514418 77932 514474 77988
rect 514294 77808 514350 77864
rect 514418 77808 514474 77864
rect 529294 79952 529350 80008
rect 529418 79952 529474 80008
rect 529294 79828 529350 79884
rect 529418 79828 529474 79884
rect 529294 79704 529350 79760
rect 529418 79704 529474 79760
rect 529294 79580 529350 79636
rect 529418 79580 529474 79636
rect 529294 79456 529350 79512
rect 529418 79456 529474 79512
rect 529294 79332 529350 79388
rect 529418 79332 529474 79388
rect 529294 79208 529350 79264
rect 529418 79208 529474 79264
rect 524294 78552 524350 78608
rect 524418 78552 524474 78608
rect 524294 78428 524350 78484
rect 524418 78428 524474 78484
rect 524294 78304 524350 78360
rect 524418 78304 524474 78360
rect 524294 78180 524350 78236
rect 524418 78180 524474 78236
rect 524294 78056 524350 78112
rect 524418 78056 524474 78112
rect 524294 77932 524350 77988
rect 524418 77932 524474 77988
rect 524294 77808 524350 77864
rect 524418 77808 524474 77864
rect 539294 79952 539350 80008
rect 539418 79952 539474 80008
rect 539294 79828 539350 79884
rect 539418 79828 539474 79884
rect 539294 79704 539350 79760
rect 539418 79704 539474 79760
rect 539294 79580 539350 79636
rect 539418 79580 539474 79636
rect 539294 79456 539350 79512
rect 539418 79456 539474 79512
rect 539294 79332 539350 79388
rect 539418 79332 539474 79388
rect 539294 79208 539350 79264
rect 539418 79208 539474 79264
rect 534294 78552 534350 78608
rect 534418 78552 534474 78608
rect 534294 78428 534350 78484
rect 534418 78428 534474 78484
rect 534294 78304 534350 78360
rect 534418 78304 534474 78360
rect 534294 78180 534350 78236
rect 534418 78180 534474 78236
rect 534294 78056 534350 78112
rect 534418 78056 534474 78112
rect 534294 77932 534350 77988
rect 534418 77932 534474 77988
rect 534294 77808 534350 77864
rect 534418 77808 534474 77864
rect 549294 79952 549350 80008
rect 549418 79952 549474 80008
rect 549294 79828 549350 79884
rect 549418 79828 549474 79884
rect 549294 79704 549350 79760
rect 549418 79704 549474 79760
rect 549294 79580 549350 79636
rect 549418 79580 549474 79636
rect 549294 79456 549350 79512
rect 549418 79456 549474 79512
rect 549294 79332 549350 79388
rect 549418 79332 549474 79388
rect 549294 79208 549350 79264
rect 549418 79208 549474 79264
rect 544294 78552 544350 78608
rect 544418 78552 544474 78608
rect 544294 78428 544350 78484
rect 544418 78428 544474 78484
rect 544294 78304 544350 78360
rect 544418 78304 544474 78360
rect 544294 78180 544350 78236
rect 544418 78180 544474 78236
rect 544294 78056 544350 78112
rect 544418 78056 544474 78112
rect 544294 77932 544350 77988
rect 544418 77932 544474 77988
rect 544294 77808 544350 77864
rect 544418 77808 544474 77864
rect 590970 79952 591026 80008
rect 591094 79952 591150 80008
rect 591218 79952 591274 80008
rect 591342 79952 591398 80008
rect 591466 79952 591522 80008
rect 591590 79952 591646 80008
rect 591714 79952 591770 80008
rect 590970 79828 591026 79884
rect 591094 79828 591150 79884
rect 591218 79828 591274 79884
rect 591342 79828 591398 79884
rect 591466 79828 591522 79884
rect 591590 79828 591646 79884
rect 591714 79828 591770 79884
rect 590970 79704 591026 79760
rect 591094 79704 591150 79760
rect 591218 79704 591274 79760
rect 591342 79704 591398 79760
rect 591466 79704 591522 79760
rect 591590 79704 591646 79760
rect 591714 79704 591770 79760
rect 590970 79580 591026 79636
rect 591094 79580 591150 79636
rect 591218 79580 591274 79636
rect 591342 79580 591398 79636
rect 591466 79580 591522 79636
rect 591590 79580 591646 79636
rect 591714 79580 591770 79636
rect 590970 79456 591026 79512
rect 591094 79456 591150 79512
rect 591218 79456 591274 79512
rect 591342 79456 591398 79512
rect 591466 79456 591522 79512
rect 591590 79456 591646 79512
rect 591714 79456 591770 79512
rect 590970 79332 591026 79388
rect 591094 79332 591150 79388
rect 591218 79332 591274 79388
rect 591342 79332 591398 79388
rect 591466 79332 591522 79388
rect 591590 79332 591646 79388
rect 591714 79332 591770 79388
rect 590970 79208 591026 79264
rect 591094 79208 591150 79264
rect 591218 79208 591274 79264
rect 591342 79208 591398 79264
rect 591466 79208 591522 79264
rect 591590 79208 591646 79264
rect 591714 79208 591770 79264
rect 592310 305670 592366 305726
rect 592434 305670 592490 305726
rect 592558 305670 592614 305726
rect 592682 305670 592738 305726
rect 592806 305670 592862 305726
rect 592930 305670 592986 305726
rect 593054 305670 593110 305726
rect 592310 305546 592366 305602
rect 592434 305546 592490 305602
rect 592558 305546 592614 305602
rect 592682 305546 592738 305602
rect 592806 305546 592862 305602
rect 592930 305546 592986 305602
rect 593054 305546 593110 305602
rect 592310 305422 592366 305478
rect 592434 305422 592490 305478
rect 592558 305422 592614 305478
rect 592682 305422 592738 305478
rect 592806 305422 592862 305478
rect 592930 305422 592986 305478
rect 593054 305422 593110 305478
rect 592310 305298 592366 305354
rect 592434 305298 592490 305354
rect 592558 305298 592614 305354
rect 592682 305298 592738 305354
rect 592806 305298 592862 305354
rect 592930 305298 592986 305354
rect 593054 305298 593110 305354
rect 592310 305174 592366 305230
rect 592434 305174 592490 305230
rect 592558 305174 592614 305230
rect 592682 305174 592738 305230
rect 592806 305174 592862 305230
rect 592930 305174 592986 305230
rect 593054 305174 593110 305230
rect 592310 305050 592366 305106
rect 592434 305050 592490 305106
rect 592558 305050 592614 305106
rect 592682 305050 592738 305106
rect 592806 305050 592862 305106
rect 592930 305050 592986 305106
rect 593054 305050 593110 305106
rect 592310 304926 592366 304982
rect 592434 304926 592490 304982
rect 592558 304926 592614 304982
rect 592682 304926 592738 304982
rect 592806 304926 592862 304982
rect 592930 304926 592986 304982
rect 593054 304926 593110 304982
rect 634860 307130 634916 307186
rect 634984 307130 635040 307186
rect 634860 307006 634916 307062
rect 634984 307006 635040 307062
rect 634860 306882 634916 306938
rect 634984 306882 635040 306938
rect 634860 306758 634916 306814
rect 634984 306758 635040 306814
rect 634860 306634 634916 306690
rect 634984 306634 635040 306690
rect 634860 306510 634916 306566
rect 634984 306510 635040 306566
rect 634860 306386 634916 306442
rect 634984 306386 635040 306442
rect 633265 305730 633321 305786
rect 633389 305730 633445 305786
rect 633265 305606 633321 305662
rect 633389 305606 633445 305662
rect 633265 305482 633321 305538
rect 633389 305482 633445 305538
rect 633265 305358 633321 305414
rect 633389 305358 633445 305414
rect 633265 305234 633321 305290
rect 633389 305234 633445 305290
rect 633265 305110 633321 305166
rect 633389 305110 633445 305166
rect 633265 304986 633321 305042
rect 633389 304986 633445 305042
rect 638050 307130 638106 307186
rect 638174 307130 638230 307186
rect 638050 307006 638106 307062
rect 638174 307006 638230 307062
rect 638050 306882 638106 306938
rect 638174 306882 638230 306938
rect 638050 306758 638106 306814
rect 638174 306758 638230 306814
rect 638050 306634 638106 306690
rect 638174 306634 638230 306690
rect 638050 306510 638106 306566
rect 638174 306510 638230 306566
rect 638050 306386 638106 306442
rect 638174 306386 638230 306442
rect 636455 305730 636511 305786
rect 636579 305730 636635 305786
rect 636455 305606 636511 305662
rect 636579 305606 636635 305662
rect 636455 305482 636511 305538
rect 636579 305482 636635 305538
rect 636455 305358 636511 305414
rect 636579 305358 636635 305414
rect 636455 305234 636511 305290
rect 636579 305234 636635 305290
rect 636455 305110 636511 305166
rect 636579 305110 636635 305166
rect 636455 304986 636511 305042
rect 636579 304986 636635 305042
rect 641240 307130 641296 307186
rect 641364 307130 641420 307186
rect 641240 307006 641296 307062
rect 641364 307006 641420 307062
rect 641240 306882 641296 306938
rect 641364 306882 641420 306938
rect 641240 306758 641296 306814
rect 641364 306758 641420 306814
rect 641240 306634 641296 306690
rect 641364 306634 641420 306690
rect 641240 306510 641296 306566
rect 641364 306510 641420 306566
rect 641240 306386 641296 306442
rect 641364 306386 641420 306442
rect 639645 305730 639701 305786
rect 639769 305730 639825 305786
rect 639645 305606 639701 305662
rect 639769 305606 639825 305662
rect 639645 305482 639701 305538
rect 639769 305482 639825 305538
rect 639645 305358 639701 305414
rect 639769 305358 639825 305414
rect 639645 305234 639701 305290
rect 639769 305234 639825 305290
rect 639645 305110 639701 305166
rect 639769 305110 639825 305166
rect 639645 304986 639701 305042
rect 639769 304986 639825 305042
rect 642835 305730 642891 305786
rect 642959 305730 643015 305786
rect 642835 305606 642891 305662
rect 642959 305606 643015 305662
rect 642835 305482 642891 305538
rect 642959 305482 643015 305538
rect 642835 305358 642891 305414
rect 642959 305358 643015 305414
rect 642835 305234 642891 305290
rect 642959 305234 643015 305290
rect 642835 305110 642891 305166
rect 642959 305110 643015 305166
rect 642835 304986 642891 305042
rect 642959 304986 643015 305042
rect 698044 313378 698100 313434
rect 698344 313378 698400 313434
rect 698644 313378 698700 313434
rect 698052 307130 698108 307186
rect 698176 307130 698232 307186
rect 698300 307130 698356 307186
rect 698424 307130 698480 307186
rect 698548 307130 698604 307186
rect 698672 307130 698728 307186
rect 698796 307130 698852 307186
rect 698052 307006 698108 307062
rect 698176 307006 698232 307062
rect 698300 307006 698356 307062
rect 698424 307006 698480 307062
rect 698548 307006 698604 307062
rect 698672 307006 698728 307062
rect 698796 307006 698852 307062
rect 698052 306882 698108 306938
rect 698176 306882 698232 306938
rect 698300 306882 698356 306938
rect 698424 306882 698480 306938
rect 698548 306882 698604 306938
rect 698672 306882 698728 306938
rect 698796 306882 698852 306938
rect 698052 306758 698108 306814
rect 698176 306758 698232 306814
rect 698300 306758 698356 306814
rect 698424 306758 698480 306814
rect 698548 306758 698604 306814
rect 698672 306758 698728 306814
rect 698796 306758 698852 306814
rect 698052 306634 698108 306690
rect 698176 306634 698232 306690
rect 698300 306634 698356 306690
rect 698424 306634 698480 306690
rect 698548 306634 698604 306690
rect 698672 306634 698728 306690
rect 698796 306634 698852 306690
rect 698052 306510 698108 306566
rect 698176 306510 698232 306566
rect 698300 306510 698356 306566
rect 698424 306510 698480 306566
rect 698548 306510 698604 306566
rect 698672 306510 698728 306566
rect 698796 306510 698852 306566
rect 698052 306386 698108 306442
rect 698176 306386 698232 306442
rect 698300 306386 698356 306442
rect 698424 306386 698480 306442
rect 698548 306386 698604 306442
rect 698672 306386 698728 306442
rect 698796 306386 698852 306442
rect 592370 281916 592426 281972
rect 592494 281916 592550 281972
rect 592618 281916 592674 281972
rect 592742 281916 592798 281972
rect 592866 281916 592922 281972
rect 592990 281916 593046 281972
rect 593114 281916 593170 281972
rect 592370 281792 592426 281848
rect 592494 281792 592550 281848
rect 592618 281792 592674 281848
rect 592742 281792 592798 281848
rect 592866 281792 592922 281848
rect 592990 281792 593046 281848
rect 593114 281792 593170 281848
rect 592370 281668 592426 281724
rect 592494 281668 592550 281724
rect 592618 281668 592674 281724
rect 592742 281668 592798 281724
rect 592866 281668 592922 281724
rect 592990 281668 593046 281724
rect 593114 281668 593170 281724
rect 592370 281544 592426 281600
rect 592494 281544 592550 281600
rect 592618 281544 592674 281600
rect 592742 281544 592798 281600
rect 592866 281544 592922 281600
rect 592990 281544 593046 281600
rect 593114 281544 593170 281600
rect 592370 281420 592426 281476
rect 592494 281420 592550 281476
rect 592618 281420 592674 281476
rect 592742 281420 592798 281476
rect 592866 281420 592922 281476
rect 592990 281420 593046 281476
rect 593114 281420 593170 281476
rect 592370 281296 592426 281352
rect 592494 281296 592550 281352
rect 592618 281296 592674 281352
rect 592742 281296 592798 281352
rect 592866 281296 592922 281352
rect 592990 281296 593046 281352
rect 593114 281296 593170 281352
rect 592370 281172 592426 281228
rect 592494 281172 592550 281228
rect 592618 281172 592674 281228
rect 592742 281172 592798 281228
rect 592866 281172 592922 281228
rect 592990 281172 593046 281228
rect 593114 281172 593170 281228
rect 592370 268316 592426 268372
rect 592494 268316 592550 268372
rect 592618 268316 592674 268372
rect 592742 268316 592798 268372
rect 592866 268316 592922 268372
rect 592990 268316 593046 268372
rect 593114 268316 593170 268372
rect 592370 268192 592426 268248
rect 592494 268192 592550 268248
rect 592618 268192 592674 268248
rect 592742 268192 592798 268248
rect 592866 268192 592922 268248
rect 592990 268192 593046 268248
rect 593114 268192 593170 268248
rect 592370 242316 592426 242372
rect 592494 242316 592550 242372
rect 592618 242316 592674 242372
rect 592742 242316 592798 242372
rect 592866 242316 592922 242372
rect 592990 242316 593046 242372
rect 593114 242316 593170 242372
rect 592370 242192 592426 242248
rect 592494 242192 592550 242248
rect 592618 242192 592674 242248
rect 592742 242192 592798 242248
rect 592866 242192 592922 242248
rect 592990 242192 593046 242248
rect 593114 242192 593170 242248
rect 592370 216316 592426 216372
rect 592494 216316 592550 216372
rect 592618 216316 592674 216372
rect 592742 216316 592798 216372
rect 592866 216316 592922 216372
rect 592990 216316 593046 216372
rect 593114 216316 593170 216372
rect 592370 216192 592426 216248
rect 592494 216192 592550 216248
rect 592618 216192 592674 216248
rect 592742 216192 592798 216248
rect 592866 216192 592922 216248
rect 592990 216192 593046 216248
rect 593114 216192 593170 216248
rect 592370 190316 592426 190372
rect 592494 190316 592550 190372
rect 592618 190316 592674 190372
rect 592742 190316 592798 190372
rect 592866 190316 592922 190372
rect 592990 190316 593046 190372
rect 593114 190316 593170 190372
rect 592370 190192 592426 190248
rect 592494 190192 592550 190248
rect 592618 190192 592674 190248
rect 592742 190192 592798 190248
rect 592866 190192 592922 190248
rect 592990 190192 593046 190248
rect 593114 190192 593170 190248
rect 592370 164316 592426 164372
rect 592494 164316 592550 164372
rect 592618 164316 592674 164372
rect 592742 164316 592798 164372
rect 592866 164316 592922 164372
rect 592990 164316 593046 164372
rect 593114 164316 593170 164372
rect 592370 164192 592426 164248
rect 592494 164192 592550 164248
rect 592618 164192 592674 164248
rect 592742 164192 592798 164248
rect 592866 164192 592922 164248
rect 592990 164192 593046 164248
rect 593114 164192 593170 164248
rect 592370 138316 592426 138372
rect 592494 138316 592550 138372
rect 592618 138316 592674 138372
rect 592742 138316 592798 138372
rect 592866 138316 592922 138372
rect 592990 138316 593046 138372
rect 593114 138316 593170 138372
rect 592370 138192 592426 138248
rect 592494 138192 592550 138248
rect 592618 138192 592674 138248
rect 592742 138192 592798 138248
rect 592866 138192 592922 138248
rect 592990 138192 593046 138248
rect 593114 138192 593170 138248
rect 592359 121635 592415 121691
rect 592659 121635 592715 121691
rect 592959 121635 593015 121691
rect 592359 118527 592415 118583
rect 592659 118527 592715 118583
rect 592959 118527 593015 118583
rect 592359 115419 592415 115475
rect 592659 115419 592715 115475
rect 592959 115419 593015 115475
rect 592370 112316 592426 112372
rect 592494 112316 592550 112372
rect 592618 112316 592674 112372
rect 592742 112316 592798 112372
rect 592866 112316 592922 112372
rect 592990 112316 593046 112372
rect 593114 112316 593170 112372
rect 592370 112192 592426 112248
rect 592494 112192 592550 112248
rect 592618 112192 592674 112248
rect 592742 112192 592798 112248
rect 592866 112192 592922 112248
rect 592990 112192 593046 112248
rect 593114 112192 593170 112248
rect 698060 289952 698116 290008
rect 698360 289952 698416 290008
rect 698660 289952 698716 290008
rect 698044 283869 698100 283925
rect 698344 283869 698400 283925
rect 698644 283869 698700 283925
rect 698044 277378 698100 277434
rect 698344 277378 698400 277434
rect 698644 277378 698700 277434
rect 698044 270378 698100 270434
rect 698344 270378 698400 270434
rect 698644 270378 698700 270434
rect 698044 263378 698100 263434
rect 698344 263378 698400 263434
rect 698644 263378 698700 263434
rect 698044 253233 698100 253289
rect 698344 253233 698400 253289
rect 698644 253233 698700 253289
rect 698060 246952 698116 247008
rect 698360 246952 698416 247008
rect 698660 246952 698716 247008
rect 698044 234378 698100 234434
rect 698344 234378 698400 234434
rect 698644 234378 698700 234434
rect 698044 227378 698100 227434
rect 698344 227378 698400 227434
rect 698644 227378 698700 227434
rect 698044 222597 698100 222653
rect 698344 222597 698400 222653
rect 698644 222597 698700 222653
rect 698044 220378 698100 220434
rect 698344 220378 698400 220434
rect 698644 220378 698700 220434
rect 698060 203952 698116 204008
rect 698360 203952 698416 204008
rect 698660 203952 698716 204008
rect 698044 191961 698100 192017
rect 698344 191961 698400 192017
rect 698644 191961 698700 192017
rect 698044 191378 698100 191434
rect 698344 191378 698400 191434
rect 698644 191378 698700 191434
rect 698044 184378 698100 184434
rect 698344 184378 698400 184434
rect 698644 184378 698700 184434
rect 698044 177378 698100 177434
rect 698344 177378 698400 177434
rect 698644 177378 698700 177434
rect 698044 161325 698100 161381
rect 698344 161325 698400 161381
rect 698644 161325 698700 161381
rect 698060 160952 698116 161008
rect 698360 160952 698416 161008
rect 698660 160952 698716 161008
rect 698044 148378 698100 148434
rect 698344 148378 698400 148434
rect 698644 148378 698700 148434
rect 698044 141378 698100 141434
rect 698344 141378 698400 141434
rect 698644 141378 698700 141434
rect 698044 134362 698100 134418
rect 698344 134362 698400 134418
rect 698644 134362 698700 134418
rect 698044 132947 698100 133003
rect 698344 132947 698400 133003
rect 698644 132947 698700 133003
rect 698060 117952 698116 118008
rect 698360 117952 698416 118008
rect 698660 117952 698716 118008
rect 698044 105378 698100 105434
rect 698344 105378 698400 105434
rect 698644 105378 698700 105434
rect 592370 86316 592426 86372
rect 592494 86316 592550 86372
rect 592618 86316 592674 86372
rect 592742 86316 592798 86372
rect 592866 86316 592922 86372
rect 592990 86316 593046 86372
rect 593114 86316 593170 86372
rect 592370 86192 592426 86248
rect 592494 86192 592550 86248
rect 592618 86192 592674 86248
rect 592742 86192 592798 86248
rect 592866 86192 592922 86248
rect 592990 86192 593046 86248
rect 593114 86192 593170 86248
rect 554294 78552 554350 78608
rect 554418 78552 554474 78608
rect 554294 78428 554350 78484
rect 554418 78428 554474 78484
rect 554294 78304 554350 78360
rect 554418 78304 554474 78360
rect 554294 78180 554350 78236
rect 554418 78180 554474 78236
rect 554294 78056 554350 78112
rect 554418 78056 554474 78112
rect 554294 77932 554350 77988
rect 554418 77932 554474 77988
rect 554294 77808 554350 77864
rect 554418 77808 554474 77864
rect 668060 99453 668116 99509
rect 668184 99453 668240 99509
rect 668308 99453 668364 99509
rect 668432 99453 668488 99509
rect 668556 99453 668612 99509
rect 668680 99453 668736 99509
rect 668060 99329 668116 99385
rect 668184 99329 668240 99385
rect 668308 99329 668364 99385
rect 668432 99329 668488 99385
rect 668556 99329 668612 99385
rect 668680 99329 668736 99385
rect 668060 99205 668116 99261
rect 668184 99205 668240 99261
rect 668308 99205 668364 99261
rect 668432 99205 668488 99261
rect 668556 99205 668612 99261
rect 668680 99205 668736 99261
rect 668060 99081 668116 99137
rect 668184 99081 668240 99137
rect 668308 99081 668364 99137
rect 668432 99081 668488 99137
rect 668556 99081 668612 99137
rect 668680 99081 668736 99137
rect 668060 98957 668116 99013
rect 668184 98957 668240 99013
rect 668308 98957 668364 99013
rect 668432 98957 668488 99013
rect 668556 98957 668612 99013
rect 668680 98957 668736 99013
rect 668060 98833 668116 98889
rect 668184 98833 668240 98889
rect 668308 98833 668364 98889
rect 668432 98833 668488 98889
rect 668556 98833 668612 98889
rect 668680 98833 668736 98889
rect 668060 98709 668116 98765
rect 668184 98709 668240 98765
rect 668308 98709 668364 98765
rect 668432 98709 668488 98765
rect 668556 98709 668612 98765
rect 668680 98709 668736 98765
rect 592370 78552 592426 78608
rect 592494 78552 592550 78608
rect 592618 78552 592674 78608
rect 592742 78552 592798 78608
rect 592866 78552 592922 78608
rect 592990 78552 593046 78608
rect 593114 78552 593170 78608
rect 592370 78428 592426 78484
rect 592494 78428 592550 78484
rect 592618 78428 592674 78484
rect 592742 78428 592798 78484
rect 592866 78428 592922 78484
rect 592990 78428 593046 78484
rect 593114 78428 593170 78484
rect 592370 78304 592426 78360
rect 592494 78304 592550 78360
rect 592618 78304 592674 78360
rect 592742 78304 592798 78360
rect 592866 78304 592922 78360
rect 592990 78304 593046 78360
rect 593114 78304 593170 78360
rect 592370 78180 592426 78236
rect 592494 78180 592550 78236
rect 592618 78180 592674 78236
rect 592742 78180 592798 78236
rect 592866 78180 592922 78236
rect 592990 78180 593046 78236
rect 593114 78180 593170 78236
rect 592370 78056 592426 78112
rect 592494 78056 592550 78112
rect 592618 78056 592674 78112
rect 592742 78056 592798 78112
rect 592866 78056 592922 78112
rect 592990 78056 593046 78112
rect 593114 78056 593170 78112
rect 592370 77932 592426 77988
rect 592494 77932 592550 77988
rect 592618 77932 592674 77988
rect 592742 77932 592798 77988
rect 592866 77932 592922 77988
rect 592990 77932 593046 77988
rect 593114 77932 593170 77988
rect 592370 77808 592426 77864
rect 592494 77808 592550 77864
rect 592618 77808 592674 77864
rect 592742 77808 592798 77864
rect 592866 77808 592922 77864
rect 592990 77808 593046 77864
rect 593114 77808 593170 77864
rect 602330 79952 602386 80008
rect 602454 79952 602510 80008
rect 602578 79952 602634 80008
rect 602702 79952 602758 80008
rect 602826 79952 602882 80008
rect 602950 79952 603006 80008
rect 603074 79952 603130 80008
rect 603198 79952 603254 80008
rect 603322 79952 603378 80008
rect 603446 79952 603502 80008
rect 603570 79952 603626 80008
rect 603694 79952 603750 80008
rect 603818 79952 603874 80008
rect 603942 79952 603998 80008
rect 604066 79952 604122 80008
rect 602330 79828 602386 79884
rect 602454 79828 602510 79884
rect 602578 79828 602634 79884
rect 602702 79828 602758 79884
rect 602826 79828 602882 79884
rect 602950 79828 603006 79884
rect 603074 79828 603130 79884
rect 603198 79828 603254 79884
rect 603322 79828 603378 79884
rect 603446 79828 603502 79884
rect 603570 79828 603626 79884
rect 603694 79828 603750 79884
rect 603818 79828 603874 79884
rect 603942 79828 603998 79884
rect 604066 79828 604122 79884
rect 602330 79704 602386 79760
rect 602454 79704 602510 79760
rect 602578 79704 602634 79760
rect 602702 79704 602758 79760
rect 602826 79704 602882 79760
rect 602950 79704 603006 79760
rect 603074 79704 603130 79760
rect 603198 79704 603254 79760
rect 603322 79704 603378 79760
rect 603446 79704 603502 79760
rect 603570 79704 603626 79760
rect 603694 79704 603750 79760
rect 603818 79704 603874 79760
rect 603942 79704 603998 79760
rect 604066 79704 604122 79760
rect 602330 79580 602386 79636
rect 602454 79580 602510 79636
rect 602578 79580 602634 79636
rect 602702 79580 602758 79636
rect 602826 79580 602882 79636
rect 602950 79580 603006 79636
rect 603074 79580 603130 79636
rect 603198 79580 603254 79636
rect 603322 79580 603378 79636
rect 603446 79580 603502 79636
rect 603570 79580 603626 79636
rect 603694 79580 603750 79636
rect 603818 79580 603874 79636
rect 603942 79580 603998 79636
rect 604066 79580 604122 79636
rect 602330 79456 602386 79512
rect 602454 79456 602510 79512
rect 602578 79456 602634 79512
rect 602702 79456 602758 79512
rect 602826 79456 602882 79512
rect 602950 79456 603006 79512
rect 603074 79456 603130 79512
rect 603198 79456 603254 79512
rect 603322 79456 603378 79512
rect 603446 79456 603502 79512
rect 603570 79456 603626 79512
rect 603694 79456 603750 79512
rect 603818 79456 603874 79512
rect 603942 79456 603998 79512
rect 604066 79456 604122 79512
rect 602330 79332 602386 79388
rect 602454 79332 602510 79388
rect 602578 79332 602634 79388
rect 602702 79332 602758 79388
rect 602826 79332 602882 79388
rect 602950 79332 603006 79388
rect 603074 79332 603130 79388
rect 603198 79332 603254 79388
rect 603322 79332 603378 79388
rect 603446 79332 603502 79388
rect 603570 79332 603626 79388
rect 603694 79332 603750 79388
rect 603818 79332 603874 79388
rect 603942 79332 603998 79388
rect 604066 79332 604122 79388
rect 602330 79208 602386 79264
rect 602454 79208 602510 79264
rect 602578 79208 602634 79264
rect 602702 79208 602758 79264
rect 602826 79208 602882 79264
rect 602950 79208 603006 79264
rect 603074 79208 603130 79264
rect 603198 79208 603254 79264
rect 603322 79208 603378 79264
rect 603446 79208 603502 79264
rect 603570 79208 603626 79264
rect 603694 79208 603750 79264
rect 603818 79208 603874 79264
rect 603942 79208 603998 79264
rect 604066 79208 604122 79264
rect 604810 79952 604866 80008
rect 604934 79952 604990 80008
rect 605058 79952 605114 80008
rect 605182 79952 605238 80008
rect 605306 79952 605362 80008
rect 605430 79952 605486 80008
rect 605554 79952 605610 80008
rect 605678 79952 605734 80008
rect 605802 79952 605858 80008
rect 605926 79952 605982 80008
rect 606050 79952 606106 80008
rect 606174 79952 606230 80008
rect 606298 79952 606354 80008
rect 606422 79952 606478 80008
rect 606546 79952 606602 80008
rect 606670 79952 606726 80008
rect 604810 79828 604866 79884
rect 604934 79828 604990 79884
rect 605058 79828 605114 79884
rect 605182 79828 605238 79884
rect 605306 79828 605362 79884
rect 605430 79828 605486 79884
rect 605554 79828 605610 79884
rect 605678 79828 605734 79884
rect 605802 79828 605858 79884
rect 605926 79828 605982 79884
rect 606050 79828 606106 79884
rect 606174 79828 606230 79884
rect 606298 79828 606354 79884
rect 606422 79828 606478 79884
rect 606546 79828 606602 79884
rect 606670 79828 606726 79884
rect 604810 79704 604866 79760
rect 604934 79704 604990 79760
rect 605058 79704 605114 79760
rect 605182 79704 605238 79760
rect 605306 79704 605362 79760
rect 605430 79704 605486 79760
rect 605554 79704 605610 79760
rect 605678 79704 605734 79760
rect 605802 79704 605858 79760
rect 605926 79704 605982 79760
rect 606050 79704 606106 79760
rect 606174 79704 606230 79760
rect 606298 79704 606354 79760
rect 606422 79704 606478 79760
rect 606546 79704 606602 79760
rect 606670 79704 606726 79760
rect 604810 79580 604866 79636
rect 604934 79580 604990 79636
rect 605058 79580 605114 79636
rect 605182 79580 605238 79636
rect 605306 79580 605362 79636
rect 605430 79580 605486 79636
rect 605554 79580 605610 79636
rect 605678 79580 605734 79636
rect 605802 79580 605858 79636
rect 605926 79580 605982 79636
rect 606050 79580 606106 79636
rect 606174 79580 606230 79636
rect 606298 79580 606354 79636
rect 606422 79580 606478 79636
rect 606546 79580 606602 79636
rect 606670 79580 606726 79636
rect 604810 79456 604866 79512
rect 604934 79456 604990 79512
rect 605058 79456 605114 79512
rect 605182 79456 605238 79512
rect 605306 79456 605362 79512
rect 605430 79456 605486 79512
rect 605554 79456 605610 79512
rect 605678 79456 605734 79512
rect 605802 79456 605858 79512
rect 605926 79456 605982 79512
rect 606050 79456 606106 79512
rect 606174 79456 606230 79512
rect 606298 79456 606354 79512
rect 606422 79456 606478 79512
rect 606546 79456 606602 79512
rect 606670 79456 606726 79512
rect 604810 79332 604866 79388
rect 604934 79332 604990 79388
rect 605058 79332 605114 79388
rect 605182 79332 605238 79388
rect 605306 79332 605362 79388
rect 605430 79332 605486 79388
rect 605554 79332 605610 79388
rect 605678 79332 605734 79388
rect 605802 79332 605858 79388
rect 605926 79332 605982 79388
rect 606050 79332 606106 79388
rect 606174 79332 606230 79388
rect 606298 79332 606354 79388
rect 606422 79332 606478 79388
rect 606546 79332 606602 79388
rect 606670 79332 606726 79388
rect 604810 79208 604866 79264
rect 604934 79208 604990 79264
rect 605058 79208 605114 79264
rect 605182 79208 605238 79264
rect 605306 79208 605362 79264
rect 605430 79208 605486 79264
rect 605554 79208 605610 79264
rect 605678 79208 605734 79264
rect 605802 79208 605858 79264
rect 605926 79208 605982 79264
rect 606050 79208 606106 79264
rect 606174 79208 606230 79264
rect 606298 79208 606354 79264
rect 606422 79208 606478 79264
rect 606546 79208 606602 79264
rect 606670 79208 606726 79264
rect 607180 79952 607236 80008
rect 607304 79952 607360 80008
rect 607428 79952 607484 80008
rect 607552 79952 607608 80008
rect 607676 79952 607732 80008
rect 607800 79952 607856 80008
rect 607924 79952 607980 80008
rect 608048 79952 608104 80008
rect 608172 79952 608228 80008
rect 608296 79952 608352 80008
rect 608420 79952 608476 80008
rect 608544 79952 608600 80008
rect 608668 79952 608724 80008
rect 608792 79952 608848 80008
rect 608916 79952 608972 80008
rect 609040 79952 609096 80008
rect 607180 79828 607236 79884
rect 607304 79828 607360 79884
rect 607428 79828 607484 79884
rect 607552 79828 607608 79884
rect 607676 79828 607732 79884
rect 607800 79828 607856 79884
rect 607924 79828 607980 79884
rect 608048 79828 608104 79884
rect 608172 79828 608228 79884
rect 608296 79828 608352 79884
rect 608420 79828 608476 79884
rect 608544 79828 608600 79884
rect 608668 79828 608724 79884
rect 608792 79828 608848 79884
rect 608916 79828 608972 79884
rect 609040 79828 609096 79884
rect 607180 79704 607236 79760
rect 607304 79704 607360 79760
rect 607428 79704 607484 79760
rect 607552 79704 607608 79760
rect 607676 79704 607732 79760
rect 607800 79704 607856 79760
rect 607924 79704 607980 79760
rect 608048 79704 608104 79760
rect 608172 79704 608228 79760
rect 608296 79704 608352 79760
rect 608420 79704 608476 79760
rect 608544 79704 608600 79760
rect 608668 79704 608724 79760
rect 608792 79704 608848 79760
rect 608916 79704 608972 79760
rect 609040 79704 609096 79760
rect 607180 79580 607236 79636
rect 607304 79580 607360 79636
rect 607428 79580 607484 79636
rect 607552 79580 607608 79636
rect 607676 79580 607732 79636
rect 607800 79580 607856 79636
rect 607924 79580 607980 79636
rect 608048 79580 608104 79636
rect 608172 79580 608228 79636
rect 608296 79580 608352 79636
rect 608420 79580 608476 79636
rect 608544 79580 608600 79636
rect 608668 79580 608724 79636
rect 608792 79580 608848 79636
rect 608916 79580 608972 79636
rect 609040 79580 609096 79636
rect 607180 79456 607236 79512
rect 607304 79456 607360 79512
rect 607428 79456 607484 79512
rect 607552 79456 607608 79512
rect 607676 79456 607732 79512
rect 607800 79456 607856 79512
rect 607924 79456 607980 79512
rect 608048 79456 608104 79512
rect 608172 79456 608228 79512
rect 608296 79456 608352 79512
rect 608420 79456 608476 79512
rect 608544 79456 608600 79512
rect 608668 79456 608724 79512
rect 608792 79456 608848 79512
rect 608916 79456 608972 79512
rect 609040 79456 609096 79512
rect 607180 79332 607236 79388
rect 607304 79332 607360 79388
rect 607428 79332 607484 79388
rect 607552 79332 607608 79388
rect 607676 79332 607732 79388
rect 607800 79332 607856 79388
rect 607924 79332 607980 79388
rect 608048 79332 608104 79388
rect 608172 79332 608228 79388
rect 608296 79332 608352 79388
rect 608420 79332 608476 79388
rect 608544 79332 608600 79388
rect 608668 79332 608724 79388
rect 608792 79332 608848 79388
rect 608916 79332 608972 79388
rect 609040 79332 609096 79388
rect 607180 79208 607236 79264
rect 607304 79208 607360 79264
rect 607428 79208 607484 79264
rect 607552 79208 607608 79264
rect 607676 79208 607732 79264
rect 607800 79208 607856 79264
rect 607924 79208 607980 79264
rect 608048 79208 608104 79264
rect 608172 79208 608228 79264
rect 608296 79208 608352 79264
rect 608420 79208 608476 79264
rect 608544 79208 608600 79264
rect 608668 79208 608724 79264
rect 608792 79208 608848 79264
rect 608916 79208 608972 79264
rect 609040 79208 609096 79264
rect 609886 79952 609942 80008
rect 610010 79952 610066 80008
rect 610134 79952 610190 80008
rect 610258 79952 610314 80008
rect 610382 79952 610438 80008
rect 610506 79952 610562 80008
rect 610630 79952 610686 80008
rect 610754 79952 610810 80008
rect 610878 79952 610934 80008
rect 611002 79952 611058 80008
rect 611126 79952 611182 80008
rect 611250 79952 611306 80008
rect 611374 79952 611430 80008
rect 611498 79952 611554 80008
rect 611622 79952 611678 80008
rect 611746 79952 611802 80008
rect 609886 79828 609942 79884
rect 610010 79828 610066 79884
rect 610134 79828 610190 79884
rect 610258 79828 610314 79884
rect 610382 79828 610438 79884
rect 610506 79828 610562 79884
rect 610630 79828 610686 79884
rect 610754 79828 610810 79884
rect 610878 79828 610934 79884
rect 611002 79828 611058 79884
rect 611126 79828 611182 79884
rect 611250 79828 611306 79884
rect 611374 79828 611430 79884
rect 611498 79828 611554 79884
rect 611622 79828 611678 79884
rect 611746 79828 611802 79884
rect 609886 79704 609942 79760
rect 610010 79704 610066 79760
rect 610134 79704 610190 79760
rect 610258 79704 610314 79760
rect 610382 79704 610438 79760
rect 610506 79704 610562 79760
rect 610630 79704 610686 79760
rect 610754 79704 610810 79760
rect 610878 79704 610934 79760
rect 611002 79704 611058 79760
rect 611126 79704 611182 79760
rect 611250 79704 611306 79760
rect 611374 79704 611430 79760
rect 611498 79704 611554 79760
rect 611622 79704 611678 79760
rect 611746 79704 611802 79760
rect 609886 79580 609942 79636
rect 610010 79580 610066 79636
rect 610134 79580 610190 79636
rect 610258 79580 610314 79636
rect 610382 79580 610438 79636
rect 610506 79580 610562 79636
rect 610630 79580 610686 79636
rect 610754 79580 610810 79636
rect 610878 79580 610934 79636
rect 611002 79580 611058 79636
rect 611126 79580 611182 79636
rect 611250 79580 611306 79636
rect 611374 79580 611430 79636
rect 611498 79580 611554 79636
rect 611622 79580 611678 79636
rect 611746 79580 611802 79636
rect 609886 79456 609942 79512
rect 610010 79456 610066 79512
rect 610134 79456 610190 79512
rect 610258 79456 610314 79512
rect 610382 79456 610438 79512
rect 610506 79456 610562 79512
rect 610630 79456 610686 79512
rect 610754 79456 610810 79512
rect 610878 79456 610934 79512
rect 611002 79456 611058 79512
rect 611126 79456 611182 79512
rect 611250 79456 611306 79512
rect 611374 79456 611430 79512
rect 611498 79456 611554 79512
rect 611622 79456 611678 79512
rect 611746 79456 611802 79512
rect 609886 79332 609942 79388
rect 610010 79332 610066 79388
rect 610134 79332 610190 79388
rect 610258 79332 610314 79388
rect 610382 79332 610438 79388
rect 610506 79332 610562 79388
rect 610630 79332 610686 79388
rect 610754 79332 610810 79388
rect 610878 79332 610934 79388
rect 611002 79332 611058 79388
rect 611126 79332 611182 79388
rect 611250 79332 611306 79388
rect 611374 79332 611430 79388
rect 611498 79332 611554 79388
rect 611622 79332 611678 79388
rect 611746 79332 611802 79388
rect 609886 79208 609942 79264
rect 610010 79208 610066 79264
rect 610134 79208 610190 79264
rect 610258 79208 610314 79264
rect 610382 79208 610438 79264
rect 610506 79208 610562 79264
rect 610630 79208 610686 79264
rect 610754 79208 610810 79264
rect 610878 79208 610934 79264
rect 611002 79208 611058 79264
rect 611126 79208 611182 79264
rect 611250 79208 611306 79264
rect 611374 79208 611430 79264
rect 611498 79208 611554 79264
rect 611622 79208 611678 79264
rect 611746 79208 611802 79264
rect 612256 79952 612312 80008
rect 612380 79952 612436 80008
rect 612504 79952 612560 80008
rect 612628 79952 612684 80008
rect 612752 79952 612808 80008
rect 612876 79952 612932 80008
rect 613000 79952 613056 80008
rect 613124 79952 613180 80008
rect 613248 79952 613304 80008
rect 613372 79952 613428 80008
rect 613496 79952 613552 80008
rect 613620 79952 613676 80008
rect 613744 79952 613800 80008
rect 613868 79952 613924 80008
rect 613992 79952 614048 80008
rect 614116 79952 614172 80008
rect 612256 79828 612312 79884
rect 612380 79828 612436 79884
rect 612504 79828 612560 79884
rect 612628 79828 612684 79884
rect 612752 79828 612808 79884
rect 612876 79828 612932 79884
rect 613000 79828 613056 79884
rect 613124 79828 613180 79884
rect 613248 79828 613304 79884
rect 613372 79828 613428 79884
rect 613496 79828 613552 79884
rect 613620 79828 613676 79884
rect 613744 79828 613800 79884
rect 613868 79828 613924 79884
rect 613992 79828 614048 79884
rect 614116 79828 614172 79884
rect 612256 79704 612312 79760
rect 612380 79704 612436 79760
rect 612504 79704 612560 79760
rect 612628 79704 612684 79760
rect 612752 79704 612808 79760
rect 612876 79704 612932 79760
rect 613000 79704 613056 79760
rect 613124 79704 613180 79760
rect 613248 79704 613304 79760
rect 613372 79704 613428 79760
rect 613496 79704 613552 79760
rect 613620 79704 613676 79760
rect 613744 79704 613800 79760
rect 613868 79704 613924 79760
rect 613992 79704 614048 79760
rect 614116 79704 614172 79760
rect 612256 79580 612312 79636
rect 612380 79580 612436 79636
rect 612504 79580 612560 79636
rect 612628 79580 612684 79636
rect 612752 79580 612808 79636
rect 612876 79580 612932 79636
rect 613000 79580 613056 79636
rect 613124 79580 613180 79636
rect 613248 79580 613304 79636
rect 613372 79580 613428 79636
rect 613496 79580 613552 79636
rect 613620 79580 613676 79636
rect 613744 79580 613800 79636
rect 613868 79580 613924 79636
rect 613992 79580 614048 79636
rect 614116 79580 614172 79636
rect 612256 79456 612312 79512
rect 612380 79456 612436 79512
rect 612504 79456 612560 79512
rect 612628 79456 612684 79512
rect 612752 79456 612808 79512
rect 612876 79456 612932 79512
rect 613000 79456 613056 79512
rect 613124 79456 613180 79512
rect 613248 79456 613304 79512
rect 613372 79456 613428 79512
rect 613496 79456 613552 79512
rect 613620 79456 613676 79512
rect 613744 79456 613800 79512
rect 613868 79456 613924 79512
rect 613992 79456 614048 79512
rect 614116 79456 614172 79512
rect 612256 79332 612312 79388
rect 612380 79332 612436 79388
rect 612504 79332 612560 79388
rect 612628 79332 612684 79388
rect 612752 79332 612808 79388
rect 612876 79332 612932 79388
rect 613000 79332 613056 79388
rect 613124 79332 613180 79388
rect 613248 79332 613304 79388
rect 613372 79332 613428 79388
rect 613496 79332 613552 79388
rect 613620 79332 613676 79388
rect 613744 79332 613800 79388
rect 613868 79332 613924 79388
rect 613992 79332 614048 79388
rect 614116 79332 614172 79388
rect 612256 79208 612312 79264
rect 612380 79208 612436 79264
rect 612504 79208 612560 79264
rect 612628 79208 612684 79264
rect 612752 79208 612808 79264
rect 612876 79208 612932 79264
rect 613000 79208 613056 79264
rect 613124 79208 613180 79264
rect 613248 79208 613304 79264
rect 613372 79208 613428 79264
rect 613496 79208 613552 79264
rect 613620 79208 613676 79264
rect 613744 79208 613800 79264
rect 613868 79208 613924 79264
rect 613992 79208 614048 79264
rect 614116 79208 614172 79264
rect 614860 79952 614916 80008
rect 614984 79952 615040 80008
rect 615108 79952 615164 80008
rect 615232 79952 615288 80008
rect 615356 79952 615412 80008
rect 615480 79952 615536 80008
rect 615604 79952 615660 80008
rect 615728 79952 615784 80008
rect 615852 79952 615908 80008
rect 615976 79952 616032 80008
rect 616100 79952 616156 80008
rect 616224 79952 616280 80008
rect 616348 79952 616404 80008
rect 616472 79952 616528 80008
rect 616596 79952 616652 80008
rect 614860 79828 614916 79884
rect 614984 79828 615040 79884
rect 615108 79828 615164 79884
rect 615232 79828 615288 79884
rect 615356 79828 615412 79884
rect 615480 79828 615536 79884
rect 615604 79828 615660 79884
rect 615728 79828 615784 79884
rect 615852 79828 615908 79884
rect 615976 79828 616032 79884
rect 616100 79828 616156 79884
rect 616224 79828 616280 79884
rect 616348 79828 616404 79884
rect 616472 79828 616528 79884
rect 616596 79828 616652 79884
rect 614860 79704 614916 79760
rect 614984 79704 615040 79760
rect 615108 79704 615164 79760
rect 615232 79704 615288 79760
rect 615356 79704 615412 79760
rect 615480 79704 615536 79760
rect 615604 79704 615660 79760
rect 615728 79704 615784 79760
rect 615852 79704 615908 79760
rect 615976 79704 616032 79760
rect 616100 79704 616156 79760
rect 616224 79704 616280 79760
rect 616348 79704 616404 79760
rect 616472 79704 616528 79760
rect 616596 79704 616652 79760
rect 614860 79580 614916 79636
rect 614984 79580 615040 79636
rect 615108 79580 615164 79636
rect 615232 79580 615288 79636
rect 615356 79580 615412 79636
rect 615480 79580 615536 79636
rect 615604 79580 615660 79636
rect 615728 79580 615784 79636
rect 615852 79580 615908 79636
rect 615976 79580 616032 79636
rect 616100 79580 616156 79636
rect 616224 79580 616280 79636
rect 616348 79580 616404 79636
rect 616472 79580 616528 79636
rect 616596 79580 616652 79636
rect 614860 79456 614916 79512
rect 614984 79456 615040 79512
rect 615108 79456 615164 79512
rect 615232 79456 615288 79512
rect 615356 79456 615412 79512
rect 615480 79456 615536 79512
rect 615604 79456 615660 79512
rect 615728 79456 615784 79512
rect 615852 79456 615908 79512
rect 615976 79456 616032 79512
rect 616100 79456 616156 79512
rect 616224 79456 616280 79512
rect 616348 79456 616404 79512
rect 616472 79456 616528 79512
rect 616596 79456 616652 79512
rect 614860 79332 614916 79388
rect 614984 79332 615040 79388
rect 615108 79332 615164 79388
rect 615232 79332 615288 79388
rect 615356 79332 615412 79388
rect 615480 79332 615536 79388
rect 615604 79332 615660 79388
rect 615728 79332 615784 79388
rect 615852 79332 615908 79388
rect 615976 79332 616032 79388
rect 616100 79332 616156 79388
rect 616224 79332 616280 79388
rect 616348 79332 616404 79388
rect 616472 79332 616528 79388
rect 616596 79332 616652 79388
rect 614860 79208 614916 79264
rect 614984 79208 615040 79264
rect 615108 79208 615164 79264
rect 615232 79208 615288 79264
rect 615356 79208 615412 79264
rect 615480 79208 615536 79264
rect 615604 79208 615660 79264
rect 615728 79208 615784 79264
rect 615852 79208 615908 79264
rect 615976 79208 616032 79264
rect 616100 79208 616156 79264
rect 616224 79208 616280 79264
rect 616348 79208 616404 79264
rect 616472 79208 616528 79264
rect 616596 79208 616652 79264
rect 628697 79952 628753 80008
rect 628821 79952 628877 80008
rect 628697 79828 628753 79884
rect 628821 79828 628877 79884
rect 628697 79704 628753 79760
rect 628821 79704 628877 79760
rect 628697 79580 628753 79636
rect 628821 79580 628877 79636
rect 628697 79456 628753 79512
rect 628821 79456 628877 79512
rect 628697 79332 628753 79388
rect 628821 79332 628877 79388
rect 628697 79208 628753 79264
rect 628821 79208 628877 79264
rect 624727 78552 624783 78608
rect 624851 78552 624907 78608
rect 624727 78428 624783 78484
rect 624851 78428 624907 78484
rect 624727 78304 624783 78360
rect 624851 78304 624907 78360
rect 624727 78180 624783 78236
rect 624851 78180 624907 78236
rect 624727 78056 624783 78112
rect 624851 78056 624907 78112
rect 624727 77932 624783 77988
rect 624851 77932 624907 77988
rect 624727 77808 624783 77864
rect 624851 77808 624907 77864
rect 636637 79952 636693 80008
rect 636761 79952 636817 80008
rect 636637 79828 636693 79884
rect 636761 79828 636817 79884
rect 636637 79704 636693 79760
rect 636761 79704 636817 79760
rect 636637 79580 636693 79636
rect 636761 79580 636817 79636
rect 636637 79456 636693 79512
rect 636761 79456 636817 79512
rect 636637 79332 636693 79388
rect 636761 79332 636817 79388
rect 636637 79208 636693 79264
rect 636761 79208 636817 79264
rect 632667 78552 632723 78608
rect 632791 78552 632847 78608
rect 632667 78428 632723 78484
rect 632791 78428 632847 78484
rect 632667 78304 632723 78360
rect 632791 78304 632847 78360
rect 632667 78180 632723 78236
rect 632791 78180 632847 78236
rect 632667 78056 632723 78112
rect 632791 78056 632847 78112
rect 632667 77932 632723 77988
rect 632791 77932 632847 77988
rect 632667 77808 632723 77864
rect 632791 77808 632847 77864
rect 644577 79952 644633 80008
rect 644701 79952 644757 80008
rect 644577 79828 644633 79884
rect 644701 79828 644757 79884
rect 644577 79704 644633 79760
rect 644701 79704 644757 79760
rect 644577 79580 644633 79636
rect 644701 79580 644757 79636
rect 644577 79456 644633 79512
rect 644701 79456 644757 79512
rect 644577 79332 644633 79388
rect 644701 79332 644757 79388
rect 644577 79208 644633 79264
rect 644701 79208 644757 79264
rect 640607 78552 640663 78608
rect 640731 78552 640787 78608
rect 640607 78428 640663 78484
rect 640731 78428 640787 78484
rect 640607 78304 640663 78360
rect 640731 78304 640787 78360
rect 640607 78180 640663 78236
rect 640731 78180 640787 78236
rect 640607 78056 640663 78112
rect 640731 78056 640787 78112
rect 640607 77932 640663 77988
rect 640731 77932 640787 77988
rect 640607 77808 640663 77864
rect 640731 77808 640787 77864
rect 670090 99453 670146 99509
rect 670214 99453 670270 99509
rect 670338 99453 670394 99509
rect 670462 99453 670518 99509
rect 670586 99453 670642 99509
rect 670710 99453 670766 99509
rect 670090 99329 670146 99385
rect 670214 99329 670270 99385
rect 670338 99329 670394 99385
rect 670462 99329 670518 99385
rect 670586 99329 670642 99385
rect 670710 99329 670766 99385
rect 670090 99205 670146 99261
rect 670214 99205 670270 99261
rect 670338 99205 670394 99261
rect 670462 99205 670518 99261
rect 670586 99205 670642 99261
rect 670710 99205 670766 99261
rect 670090 99081 670146 99137
rect 670214 99081 670270 99137
rect 670338 99081 670394 99137
rect 670462 99081 670518 99137
rect 670586 99081 670642 99137
rect 670710 99081 670766 99137
rect 670090 98957 670146 99013
rect 670214 98957 670270 99013
rect 670338 98957 670394 99013
rect 670462 98957 670518 99013
rect 670586 98957 670642 99013
rect 670710 98957 670766 99013
rect 670090 98833 670146 98889
rect 670214 98833 670270 98889
rect 670338 98833 670394 98889
rect 670462 98833 670518 98889
rect 670586 98833 670642 98889
rect 670710 98833 670766 98889
rect 670090 98709 670146 98765
rect 670214 98709 670270 98765
rect 670338 98709 670394 98765
rect 670462 98709 670518 98765
rect 670586 98709 670642 98765
rect 670710 98709 670766 98765
rect 670090 79952 670146 80008
rect 670214 79952 670270 80008
rect 670338 79952 670394 80008
rect 670462 79952 670518 80008
rect 670586 79952 670642 80008
rect 670710 79952 670766 80008
rect 670090 79828 670146 79884
rect 670214 79828 670270 79884
rect 670338 79828 670394 79884
rect 670462 79828 670518 79884
rect 670586 79828 670642 79884
rect 670710 79828 670766 79884
rect 670090 79704 670146 79760
rect 670214 79704 670270 79760
rect 670338 79704 670394 79760
rect 670462 79704 670518 79760
rect 670586 79704 670642 79760
rect 670710 79704 670766 79760
rect 670090 79580 670146 79636
rect 670214 79580 670270 79636
rect 670338 79580 670394 79636
rect 670462 79580 670518 79636
rect 670586 79580 670642 79636
rect 670710 79580 670766 79636
rect 670090 79456 670146 79512
rect 670214 79456 670270 79512
rect 670338 79456 670394 79512
rect 670462 79456 670518 79512
rect 670586 79456 670642 79512
rect 670710 79456 670766 79512
rect 670090 79332 670146 79388
rect 670214 79332 670270 79388
rect 670338 79332 670394 79388
rect 670462 79332 670518 79388
rect 670586 79332 670642 79388
rect 670710 79332 670766 79388
rect 670090 79208 670146 79264
rect 670214 79208 670270 79264
rect 670338 79208 670394 79264
rect 670462 79208 670518 79264
rect 670586 79208 670642 79264
rect 670710 79208 670766 79264
rect 698044 98378 698100 98434
rect 698344 98378 698400 98434
rect 698644 98378 698700 98434
rect 698044 91378 698100 91434
rect 698344 91378 698400 91434
rect 698644 91378 698700 91434
rect 698052 79952 698108 80008
rect 698176 79952 698232 80008
rect 698300 79952 698356 80008
rect 698424 79952 698480 80008
rect 698548 79952 698604 80008
rect 698672 79952 698728 80008
rect 698796 79952 698852 80008
rect 698052 79828 698108 79884
rect 698176 79828 698232 79884
rect 698300 79828 698356 79884
rect 698424 79828 698480 79884
rect 698548 79828 698604 79884
rect 698672 79828 698728 79884
rect 698796 79828 698852 79884
rect 698052 79704 698108 79760
rect 698176 79704 698232 79760
rect 698300 79704 698356 79760
rect 698424 79704 698480 79760
rect 698548 79704 698604 79760
rect 698672 79704 698728 79760
rect 698796 79704 698852 79760
rect 698052 79580 698108 79636
rect 698176 79580 698232 79636
rect 698300 79580 698356 79636
rect 698424 79580 698480 79636
rect 698548 79580 698604 79636
rect 698672 79580 698728 79636
rect 698796 79580 698852 79636
rect 698052 79456 698108 79512
rect 698176 79456 698232 79512
rect 698300 79456 698356 79512
rect 698424 79456 698480 79512
rect 698548 79456 698604 79512
rect 698672 79456 698728 79512
rect 698796 79456 698852 79512
rect 698052 79332 698108 79388
rect 698176 79332 698232 79388
rect 698300 79332 698356 79388
rect 698424 79332 698480 79388
rect 698548 79332 698604 79388
rect 698672 79332 698728 79388
rect 698796 79332 698852 79388
rect 698052 79208 698108 79264
rect 698176 79208 698232 79264
rect 698300 79208 698356 79264
rect 698424 79208 698480 79264
rect 698548 79208 698604 79264
rect 698672 79208 698728 79264
rect 698796 79208 698852 79264
rect 648547 78552 648603 78608
rect 648671 78552 648727 78608
rect 648547 78428 648603 78484
rect 648671 78428 648727 78484
rect 648547 78304 648603 78360
rect 648671 78304 648727 78360
rect 648547 78180 648603 78236
rect 648671 78180 648727 78236
rect 648547 78056 648603 78112
rect 648671 78056 648727 78112
rect 648547 77932 648603 77988
rect 648671 77932 648727 77988
rect 648547 77808 648603 77864
rect 648671 77808 648727 77864
rect 657330 78552 657386 78608
rect 657454 78552 657510 78608
rect 657578 78552 657634 78608
rect 657702 78552 657758 78608
rect 657826 78552 657882 78608
rect 657950 78552 658006 78608
rect 658074 78552 658130 78608
rect 658198 78552 658254 78608
rect 658322 78552 658378 78608
rect 658446 78552 658502 78608
rect 658570 78552 658626 78608
rect 658694 78552 658750 78608
rect 658818 78552 658874 78608
rect 658942 78552 658998 78608
rect 659066 78552 659122 78608
rect 657330 78428 657386 78484
rect 657454 78428 657510 78484
rect 657578 78428 657634 78484
rect 657702 78428 657758 78484
rect 657826 78428 657882 78484
rect 657950 78428 658006 78484
rect 658074 78428 658130 78484
rect 658198 78428 658254 78484
rect 658322 78428 658378 78484
rect 658446 78428 658502 78484
rect 658570 78428 658626 78484
rect 658694 78428 658750 78484
rect 658818 78428 658874 78484
rect 658942 78428 658998 78484
rect 659066 78428 659122 78484
rect 657330 78304 657386 78360
rect 657454 78304 657510 78360
rect 657578 78304 657634 78360
rect 657702 78304 657758 78360
rect 657826 78304 657882 78360
rect 657950 78304 658006 78360
rect 658074 78304 658130 78360
rect 658198 78304 658254 78360
rect 658322 78304 658378 78360
rect 658446 78304 658502 78360
rect 658570 78304 658626 78360
rect 658694 78304 658750 78360
rect 658818 78304 658874 78360
rect 658942 78304 658998 78360
rect 659066 78304 659122 78360
rect 657330 78180 657386 78236
rect 657454 78180 657510 78236
rect 657578 78180 657634 78236
rect 657702 78180 657758 78236
rect 657826 78180 657882 78236
rect 657950 78180 658006 78236
rect 658074 78180 658130 78236
rect 658198 78180 658254 78236
rect 658322 78180 658378 78236
rect 658446 78180 658502 78236
rect 658570 78180 658626 78236
rect 658694 78180 658750 78236
rect 658818 78180 658874 78236
rect 658942 78180 658998 78236
rect 659066 78180 659122 78236
rect 657330 78056 657386 78112
rect 657454 78056 657510 78112
rect 657578 78056 657634 78112
rect 657702 78056 657758 78112
rect 657826 78056 657882 78112
rect 657950 78056 658006 78112
rect 658074 78056 658130 78112
rect 658198 78056 658254 78112
rect 658322 78056 658378 78112
rect 658446 78056 658502 78112
rect 658570 78056 658626 78112
rect 658694 78056 658750 78112
rect 658818 78056 658874 78112
rect 658942 78056 658998 78112
rect 659066 78056 659122 78112
rect 657330 77932 657386 77988
rect 657454 77932 657510 77988
rect 657578 77932 657634 77988
rect 657702 77932 657758 77988
rect 657826 77932 657882 77988
rect 657950 77932 658006 77988
rect 658074 77932 658130 77988
rect 658198 77932 658254 77988
rect 658322 77932 658378 77988
rect 658446 77932 658502 77988
rect 658570 77932 658626 77988
rect 658694 77932 658750 77988
rect 658818 77932 658874 77988
rect 658942 77932 658998 77988
rect 659066 77932 659122 77988
rect 657330 77808 657386 77864
rect 657454 77808 657510 77864
rect 657578 77808 657634 77864
rect 657702 77808 657758 77864
rect 657826 77808 657882 77864
rect 657950 77808 658006 77864
rect 658074 77808 658130 77864
rect 658198 77808 658254 77864
rect 658322 77808 658378 77864
rect 658446 77808 658502 77864
rect 658570 77808 658626 77864
rect 658694 77808 658750 77864
rect 658818 77808 658874 77864
rect 658942 77808 658998 77864
rect 659066 77808 659122 77864
rect 659810 78552 659866 78608
rect 659934 78552 659990 78608
rect 660058 78552 660114 78608
rect 660182 78552 660238 78608
rect 660306 78552 660362 78608
rect 660430 78552 660486 78608
rect 660554 78552 660610 78608
rect 660678 78552 660734 78608
rect 660802 78552 660858 78608
rect 660926 78552 660982 78608
rect 661050 78552 661106 78608
rect 661174 78552 661230 78608
rect 661298 78552 661354 78608
rect 661422 78552 661478 78608
rect 661546 78552 661602 78608
rect 661670 78552 661726 78608
rect 659810 78428 659866 78484
rect 659934 78428 659990 78484
rect 660058 78428 660114 78484
rect 660182 78428 660238 78484
rect 660306 78428 660362 78484
rect 660430 78428 660486 78484
rect 660554 78428 660610 78484
rect 660678 78428 660734 78484
rect 660802 78428 660858 78484
rect 660926 78428 660982 78484
rect 661050 78428 661106 78484
rect 661174 78428 661230 78484
rect 661298 78428 661354 78484
rect 661422 78428 661478 78484
rect 661546 78428 661602 78484
rect 661670 78428 661726 78484
rect 659810 78304 659866 78360
rect 659934 78304 659990 78360
rect 660058 78304 660114 78360
rect 660182 78304 660238 78360
rect 660306 78304 660362 78360
rect 660430 78304 660486 78360
rect 660554 78304 660610 78360
rect 660678 78304 660734 78360
rect 660802 78304 660858 78360
rect 660926 78304 660982 78360
rect 661050 78304 661106 78360
rect 661174 78304 661230 78360
rect 661298 78304 661354 78360
rect 661422 78304 661478 78360
rect 661546 78304 661602 78360
rect 661670 78304 661726 78360
rect 659810 78180 659866 78236
rect 659934 78180 659990 78236
rect 660058 78180 660114 78236
rect 660182 78180 660238 78236
rect 660306 78180 660362 78236
rect 660430 78180 660486 78236
rect 660554 78180 660610 78236
rect 660678 78180 660734 78236
rect 660802 78180 660858 78236
rect 660926 78180 660982 78236
rect 661050 78180 661106 78236
rect 661174 78180 661230 78236
rect 661298 78180 661354 78236
rect 661422 78180 661478 78236
rect 661546 78180 661602 78236
rect 661670 78180 661726 78236
rect 659810 78056 659866 78112
rect 659934 78056 659990 78112
rect 660058 78056 660114 78112
rect 660182 78056 660238 78112
rect 660306 78056 660362 78112
rect 660430 78056 660486 78112
rect 660554 78056 660610 78112
rect 660678 78056 660734 78112
rect 660802 78056 660858 78112
rect 660926 78056 660982 78112
rect 661050 78056 661106 78112
rect 661174 78056 661230 78112
rect 661298 78056 661354 78112
rect 661422 78056 661478 78112
rect 661546 78056 661602 78112
rect 661670 78056 661726 78112
rect 659810 77932 659866 77988
rect 659934 77932 659990 77988
rect 660058 77932 660114 77988
rect 660182 77932 660238 77988
rect 660306 77932 660362 77988
rect 660430 77932 660486 77988
rect 660554 77932 660610 77988
rect 660678 77932 660734 77988
rect 660802 77932 660858 77988
rect 660926 77932 660982 77988
rect 661050 77932 661106 77988
rect 661174 77932 661230 77988
rect 661298 77932 661354 77988
rect 661422 77932 661478 77988
rect 661546 77932 661602 77988
rect 661670 77932 661726 77988
rect 659810 77808 659866 77864
rect 659934 77808 659990 77864
rect 660058 77808 660114 77864
rect 660182 77808 660238 77864
rect 660306 77808 660362 77864
rect 660430 77808 660486 77864
rect 660554 77808 660610 77864
rect 660678 77808 660734 77864
rect 660802 77808 660858 77864
rect 660926 77808 660982 77864
rect 661050 77808 661106 77864
rect 661174 77808 661230 77864
rect 661298 77808 661354 77864
rect 661422 77808 661478 77864
rect 661546 77808 661602 77864
rect 661670 77808 661726 77864
rect 662180 78552 662236 78608
rect 662304 78552 662360 78608
rect 662428 78552 662484 78608
rect 662552 78552 662608 78608
rect 662676 78552 662732 78608
rect 662800 78552 662856 78608
rect 662924 78552 662980 78608
rect 663048 78552 663104 78608
rect 663172 78552 663228 78608
rect 663296 78552 663352 78608
rect 663420 78552 663476 78608
rect 663544 78552 663600 78608
rect 663668 78552 663724 78608
rect 663792 78552 663848 78608
rect 663916 78552 663972 78608
rect 664040 78552 664096 78608
rect 662180 78428 662236 78484
rect 662304 78428 662360 78484
rect 662428 78428 662484 78484
rect 662552 78428 662608 78484
rect 662676 78428 662732 78484
rect 662800 78428 662856 78484
rect 662924 78428 662980 78484
rect 663048 78428 663104 78484
rect 663172 78428 663228 78484
rect 663296 78428 663352 78484
rect 663420 78428 663476 78484
rect 663544 78428 663600 78484
rect 663668 78428 663724 78484
rect 663792 78428 663848 78484
rect 663916 78428 663972 78484
rect 664040 78428 664096 78484
rect 662180 78304 662236 78360
rect 662304 78304 662360 78360
rect 662428 78304 662484 78360
rect 662552 78304 662608 78360
rect 662676 78304 662732 78360
rect 662800 78304 662856 78360
rect 662924 78304 662980 78360
rect 663048 78304 663104 78360
rect 663172 78304 663228 78360
rect 663296 78304 663352 78360
rect 663420 78304 663476 78360
rect 663544 78304 663600 78360
rect 663668 78304 663724 78360
rect 663792 78304 663848 78360
rect 663916 78304 663972 78360
rect 664040 78304 664096 78360
rect 662180 78180 662236 78236
rect 662304 78180 662360 78236
rect 662428 78180 662484 78236
rect 662552 78180 662608 78236
rect 662676 78180 662732 78236
rect 662800 78180 662856 78236
rect 662924 78180 662980 78236
rect 663048 78180 663104 78236
rect 663172 78180 663228 78236
rect 663296 78180 663352 78236
rect 663420 78180 663476 78236
rect 663544 78180 663600 78236
rect 663668 78180 663724 78236
rect 663792 78180 663848 78236
rect 663916 78180 663972 78236
rect 664040 78180 664096 78236
rect 662180 78056 662236 78112
rect 662304 78056 662360 78112
rect 662428 78056 662484 78112
rect 662552 78056 662608 78112
rect 662676 78056 662732 78112
rect 662800 78056 662856 78112
rect 662924 78056 662980 78112
rect 663048 78056 663104 78112
rect 663172 78056 663228 78112
rect 663296 78056 663352 78112
rect 663420 78056 663476 78112
rect 663544 78056 663600 78112
rect 663668 78056 663724 78112
rect 663792 78056 663848 78112
rect 663916 78056 663972 78112
rect 664040 78056 664096 78112
rect 662180 77932 662236 77988
rect 662304 77932 662360 77988
rect 662428 77932 662484 77988
rect 662552 77932 662608 77988
rect 662676 77932 662732 77988
rect 662800 77932 662856 77988
rect 662924 77932 662980 77988
rect 663048 77932 663104 77988
rect 663172 77932 663228 77988
rect 663296 77932 663352 77988
rect 663420 77932 663476 77988
rect 663544 77932 663600 77988
rect 663668 77932 663724 77988
rect 663792 77932 663848 77988
rect 663916 77932 663972 77988
rect 664040 77932 664096 77988
rect 662180 77808 662236 77864
rect 662304 77808 662360 77864
rect 662428 77808 662484 77864
rect 662552 77808 662608 77864
rect 662676 77808 662732 77864
rect 662800 77808 662856 77864
rect 662924 77808 662980 77864
rect 663048 77808 663104 77864
rect 663172 77808 663228 77864
rect 663296 77808 663352 77864
rect 663420 77808 663476 77864
rect 663544 77808 663600 77864
rect 663668 77808 663724 77864
rect 663792 77808 663848 77864
rect 663916 77808 663972 77864
rect 664040 77808 664096 77864
rect 664886 78552 664942 78608
rect 665010 78552 665066 78608
rect 665134 78552 665190 78608
rect 665258 78552 665314 78608
rect 665382 78552 665438 78608
rect 665506 78552 665562 78608
rect 665630 78552 665686 78608
rect 665754 78552 665810 78608
rect 665878 78552 665934 78608
rect 666002 78552 666058 78608
rect 666126 78552 666182 78608
rect 666250 78552 666306 78608
rect 666374 78552 666430 78608
rect 666498 78552 666554 78608
rect 666622 78552 666678 78608
rect 666746 78552 666802 78608
rect 664886 78428 664942 78484
rect 665010 78428 665066 78484
rect 665134 78428 665190 78484
rect 665258 78428 665314 78484
rect 665382 78428 665438 78484
rect 665506 78428 665562 78484
rect 665630 78428 665686 78484
rect 665754 78428 665810 78484
rect 665878 78428 665934 78484
rect 666002 78428 666058 78484
rect 666126 78428 666182 78484
rect 666250 78428 666306 78484
rect 666374 78428 666430 78484
rect 666498 78428 666554 78484
rect 666622 78428 666678 78484
rect 666746 78428 666802 78484
rect 664886 78304 664942 78360
rect 665010 78304 665066 78360
rect 665134 78304 665190 78360
rect 665258 78304 665314 78360
rect 665382 78304 665438 78360
rect 665506 78304 665562 78360
rect 665630 78304 665686 78360
rect 665754 78304 665810 78360
rect 665878 78304 665934 78360
rect 666002 78304 666058 78360
rect 666126 78304 666182 78360
rect 666250 78304 666306 78360
rect 666374 78304 666430 78360
rect 666498 78304 666554 78360
rect 666622 78304 666678 78360
rect 666746 78304 666802 78360
rect 664886 78180 664942 78236
rect 665010 78180 665066 78236
rect 665134 78180 665190 78236
rect 665258 78180 665314 78236
rect 665382 78180 665438 78236
rect 665506 78180 665562 78236
rect 665630 78180 665686 78236
rect 665754 78180 665810 78236
rect 665878 78180 665934 78236
rect 666002 78180 666058 78236
rect 666126 78180 666182 78236
rect 666250 78180 666306 78236
rect 666374 78180 666430 78236
rect 666498 78180 666554 78236
rect 666622 78180 666678 78236
rect 666746 78180 666802 78236
rect 664886 78056 664942 78112
rect 665010 78056 665066 78112
rect 665134 78056 665190 78112
rect 665258 78056 665314 78112
rect 665382 78056 665438 78112
rect 665506 78056 665562 78112
rect 665630 78056 665686 78112
rect 665754 78056 665810 78112
rect 665878 78056 665934 78112
rect 666002 78056 666058 78112
rect 666126 78056 666182 78112
rect 666250 78056 666306 78112
rect 666374 78056 666430 78112
rect 666498 78056 666554 78112
rect 666622 78056 666678 78112
rect 666746 78056 666802 78112
rect 664886 77932 664942 77988
rect 665010 77932 665066 77988
rect 665134 77932 665190 77988
rect 665258 77932 665314 77988
rect 665382 77932 665438 77988
rect 665506 77932 665562 77988
rect 665630 77932 665686 77988
rect 665754 77932 665810 77988
rect 665878 77932 665934 77988
rect 666002 77932 666058 77988
rect 666126 77932 666182 77988
rect 666250 77932 666306 77988
rect 666374 77932 666430 77988
rect 666498 77932 666554 77988
rect 666622 77932 666678 77988
rect 666746 77932 666802 77988
rect 664886 77808 664942 77864
rect 665010 77808 665066 77864
rect 665134 77808 665190 77864
rect 665258 77808 665314 77864
rect 665382 77808 665438 77864
rect 665506 77808 665562 77864
rect 665630 77808 665686 77864
rect 665754 77808 665810 77864
rect 665878 77808 665934 77864
rect 666002 77808 666058 77864
rect 666126 77808 666182 77864
rect 666250 77808 666306 77864
rect 666374 77808 666430 77864
rect 666498 77808 666554 77864
rect 666622 77808 666678 77864
rect 666746 77808 666802 77864
rect 667256 78552 667312 78608
rect 667380 78552 667436 78608
rect 667504 78552 667560 78608
rect 667628 78552 667684 78608
rect 667752 78552 667808 78608
rect 667876 78552 667932 78608
rect 668000 78552 668056 78608
rect 668124 78552 668180 78608
rect 668248 78552 668304 78608
rect 668372 78552 668428 78608
rect 668496 78552 668552 78608
rect 668620 78552 668676 78608
rect 668744 78552 668800 78608
rect 668868 78552 668924 78608
rect 668992 78552 669048 78608
rect 669116 78552 669172 78608
rect 667256 78428 667312 78484
rect 667380 78428 667436 78484
rect 667504 78428 667560 78484
rect 667628 78428 667684 78484
rect 667752 78428 667808 78484
rect 667876 78428 667932 78484
rect 668000 78428 668056 78484
rect 668124 78428 668180 78484
rect 668248 78428 668304 78484
rect 668372 78428 668428 78484
rect 668496 78428 668552 78484
rect 668620 78428 668676 78484
rect 668744 78428 668800 78484
rect 668868 78428 668924 78484
rect 668992 78428 669048 78484
rect 669116 78428 669172 78484
rect 667256 78304 667312 78360
rect 667380 78304 667436 78360
rect 667504 78304 667560 78360
rect 667628 78304 667684 78360
rect 667752 78304 667808 78360
rect 667876 78304 667932 78360
rect 668000 78304 668056 78360
rect 668124 78304 668180 78360
rect 668248 78304 668304 78360
rect 668372 78304 668428 78360
rect 668496 78304 668552 78360
rect 668620 78304 668676 78360
rect 668744 78304 668800 78360
rect 668868 78304 668924 78360
rect 668992 78304 669048 78360
rect 669116 78304 669172 78360
rect 667256 78180 667312 78236
rect 667380 78180 667436 78236
rect 667504 78180 667560 78236
rect 667628 78180 667684 78236
rect 667752 78180 667808 78236
rect 667876 78180 667932 78236
rect 668000 78180 668056 78236
rect 668124 78180 668180 78236
rect 668248 78180 668304 78236
rect 668372 78180 668428 78236
rect 668496 78180 668552 78236
rect 668620 78180 668676 78236
rect 668744 78180 668800 78236
rect 668868 78180 668924 78236
rect 668992 78180 669048 78236
rect 669116 78180 669172 78236
rect 667256 78056 667312 78112
rect 667380 78056 667436 78112
rect 667504 78056 667560 78112
rect 667628 78056 667684 78112
rect 667752 78056 667808 78112
rect 667876 78056 667932 78112
rect 668000 78056 668056 78112
rect 668124 78056 668180 78112
rect 668248 78056 668304 78112
rect 668372 78056 668428 78112
rect 668496 78056 668552 78112
rect 668620 78056 668676 78112
rect 668744 78056 668800 78112
rect 668868 78056 668924 78112
rect 668992 78056 669048 78112
rect 669116 78056 669172 78112
rect 667256 77932 667312 77988
rect 667380 77932 667436 77988
rect 667504 77932 667560 77988
rect 667628 77932 667684 77988
rect 667752 77932 667808 77988
rect 667876 77932 667932 77988
rect 668000 77932 668056 77988
rect 668124 77932 668180 77988
rect 668248 77932 668304 77988
rect 668372 77932 668428 77988
rect 668496 77932 668552 77988
rect 668620 77932 668676 77988
rect 668744 77932 668800 77988
rect 668868 77932 668924 77988
rect 668992 77932 669048 77988
rect 669116 77932 669172 77988
rect 667256 77808 667312 77864
rect 667380 77808 667436 77864
rect 667504 77808 667560 77864
rect 667628 77808 667684 77864
rect 667752 77808 667808 77864
rect 667876 77808 667932 77864
rect 668000 77808 668056 77864
rect 668124 77808 668180 77864
rect 668248 77808 668304 77864
rect 668372 77808 668428 77864
rect 668496 77808 668552 77864
rect 668620 77808 668676 77864
rect 668744 77808 668800 77864
rect 668868 77808 668924 77864
rect 668992 77808 669048 77864
rect 669116 77808 669172 77864
rect 669860 78552 669916 78608
rect 669984 78552 670040 78608
rect 670108 78552 670164 78608
rect 670232 78552 670288 78608
rect 670356 78552 670412 78608
rect 670480 78552 670536 78608
rect 670604 78552 670660 78608
rect 670728 78552 670784 78608
rect 670852 78552 670908 78608
rect 670976 78552 671032 78608
rect 671100 78552 671156 78608
rect 671224 78552 671280 78608
rect 671348 78552 671404 78608
rect 671472 78552 671528 78608
rect 671596 78552 671652 78608
rect 669860 78428 669916 78484
rect 669984 78428 670040 78484
rect 670108 78428 670164 78484
rect 670232 78428 670288 78484
rect 670356 78428 670412 78484
rect 670480 78428 670536 78484
rect 670604 78428 670660 78484
rect 670728 78428 670784 78484
rect 670852 78428 670908 78484
rect 670976 78428 671032 78484
rect 671100 78428 671156 78484
rect 671224 78428 671280 78484
rect 671348 78428 671404 78484
rect 671472 78428 671528 78484
rect 671596 78428 671652 78484
rect 669860 78304 669916 78360
rect 669984 78304 670040 78360
rect 670108 78304 670164 78360
rect 670232 78304 670288 78360
rect 670356 78304 670412 78360
rect 670480 78304 670536 78360
rect 670604 78304 670660 78360
rect 670728 78304 670784 78360
rect 670852 78304 670908 78360
rect 670976 78304 671032 78360
rect 671100 78304 671156 78360
rect 671224 78304 671280 78360
rect 671348 78304 671404 78360
rect 671472 78304 671528 78360
rect 671596 78304 671652 78360
rect 669860 78180 669916 78236
rect 669984 78180 670040 78236
rect 670108 78180 670164 78236
rect 670232 78180 670288 78236
rect 670356 78180 670412 78236
rect 670480 78180 670536 78236
rect 670604 78180 670660 78236
rect 670728 78180 670784 78236
rect 670852 78180 670908 78236
rect 670976 78180 671032 78236
rect 671100 78180 671156 78236
rect 671224 78180 671280 78236
rect 671348 78180 671404 78236
rect 671472 78180 671528 78236
rect 671596 78180 671652 78236
rect 669860 78056 669916 78112
rect 669984 78056 670040 78112
rect 670108 78056 670164 78112
rect 670232 78056 670288 78112
rect 670356 78056 670412 78112
rect 670480 78056 670536 78112
rect 670604 78056 670660 78112
rect 670728 78056 670784 78112
rect 670852 78056 670908 78112
rect 670976 78056 671032 78112
rect 671100 78056 671156 78112
rect 671224 78056 671280 78112
rect 671348 78056 671404 78112
rect 671472 78056 671528 78112
rect 671596 78056 671652 78112
rect 669860 77932 669916 77988
rect 669984 77932 670040 77988
rect 670108 77932 670164 77988
rect 670232 77932 670288 77988
rect 670356 77932 670412 77988
rect 670480 77932 670536 77988
rect 670604 77932 670660 77988
rect 670728 77932 670784 77988
rect 670852 77932 670908 77988
rect 670976 77932 671032 77988
rect 671100 77932 671156 77988
rect 671224 77932 671280 77988
rect 671348 77932 671404 77988
rect 671472 77932 671528 77988
rect 671596 77932 671652 77988
rect 669860 77808 669916 77864
rect 669984 77808 670040 77864
rect 670108 77808 670164 77864
rect 670232 77808 670288 77864
rect 670356 77808 670412 77864
rect 670480 77808 670536 77864
rect 670604 77808 670660 77864
rect 670728 77808 670784 77864
rect 670852 77808 670908 77864
rect 670976 77808 671032 77864
rect 671100 77808 671156 77864
rect 671224 77808 671280 77864
rect 671348 77808 671404 77864
rect 671472 77808 671528 77864
rect 671596 77808 671652 77864
rect 699444 925898 699500 925954
rect 699744 925898 699800 925954
rect 700044 925898 700100 925954
rect 699444 918898 699500 918954
rect 699744 918898 699800 918954
rect 700044 918898 700100 918954
rect 699544 914373 699600 914429
rect 699844 914373 699900 914429
rect 700144 914373 700200 914429
rect 699544 914173 699600 914229
rect 699844 914173 699900 914229
rect 700144 914173 700200 914229
rect 699444 911898 699500 911954
rect 699744 911898 699800 911954
rect 700044 911898 700100 911954
rect 699497 892367 699553 892423
rect 699797 892367 699853 892423
rect 700097 892367 700153 892423
rect 699392 883596 699448 883652
rect 699516 883596 699572 883652
rect 699640 883596 699696 883652
rect 699764 883596 699820 883652
rect 699888 883596 699944 883652
rect 700012 883596 700068 883652
rect 700136 883596 700192 883652
rect 699392 883472 699448 883528
rect 699516 883472 699572 883528
rect 699640 883472 699696 883528
rect 699764 883472 699820 883528
rect 699888 883472 699944 883528
rect 700012 883472 700068 883528
rect 700136 883472 700192 883528
rect 699392 883348 699448 883404
rect 699516 883348 699572 883404
rect 699640 883348 699696 883404
rect 699764 883348 699820 883404
rect 699888 883348 699944 883404
rect 700012 883348 700068 883404
rect 700136 883348 700192 883404
rect 699392 883224 699448 883280
rect 699516 883224 699572 883280
rect 699640 883224 699696 883280
rect 699764 883224 699820 883280
rect 699888 883224 699944 883280
rect 700012 883224 700068 883280
rect 700136 883224 700192 883280
rect 699392 883100 699448 883156
rect 699516 883100 699572 883156
rect 699640 883100 699696 883156
rect 699764 883100 699820 883156
rect 699888 883100 699944 883156
rect 700012 883100 700068 883156
rect 700136 883100 700192 883156
rect 699392 882976 699448 883032
rect 699516 882976 699572 883032
rect 699640 882976 699696 883032
rect 699764 882976 699820 883032
rect 699888 882976 699944 883032
rect 700012 882976 700068 883032
rect 700136 882976 700192 883032
rect 699392 882852 699448 882908
rect 699516 882852 699572 882908
rect 699640 882852 699696 882908
rect 699764 882852 699820 882908
rect 699888 882852 699944 882908
rect 700012 882852 700068 882908
rect 700136 882852 700192 882908
rect 699392 882728 699448 882784
rect 699516 882728 699572 882784
rect 699640 882728 699696 882784
rect 699764 882728 699820 882784
rect 699888 882728 699944 882784
rect 700012 882728 700068 882784
rect 700136 882728 700192 882784
rect 699392 882604 699448 882660
rect 699516 882604 699572 882660
rect 699640 882604 699696 882660
rect 699764 882604 699820 882660
rect 699888 882604 699944 882660
rect 700012 882604 700068 882660
rect 700136 882604 700192 882660
rect 699392 882480 699448 882536
rect 699516 882480 699572 882536
rect 699640 882480 699696 882536
rect 699764 882480 699820 882536
rect 699888 882480 699944 882536
rect 700012 882480 700068 882536
rect 700136 882480 700192 882536
rect 699392 882356 699448 882412
rect 699516 882356 699572 882412
rect 699640 882356 699696 882412
rect 699764 882356 699820 882412
rect 699888 882356 699944 882412
rect 700012 882356 700068 882412
rect 700136 882356 700192 882412
rect 699392 882232 699448 882288
rect 699516 882232 699572 882288
rect 699640 882232 699696 882288
rect 699764 882232 699820 882288
rect 699888 882232 699944 882288
rect 700012 882232 700068 882288
rect 700136 882232 700192 882288
rect 699392 882108 699448 882164
rect 699516 882108 699572 882164
rect 699640 882108 699696 882164
rect 699764 882108 699820 882164
rect 699888 882108 699944 882164
rect 700012 882108 700068 882164
rect 700136 882108 700192 882164
rect 699392 881984 699448 882040
rect 699516 881984 699572 882040
rect 699640 881984 699696 882040
rect 699764 881984 699820 882040
rect 699888 881984 699944 882040
rect 700012 881984 700068 882040
rect 700136 881984 700192 882040
rect 699392 881860 699448 881916
rect 699516 881860 699572 881916
rect 699640 881860 699696 881916
rect 699764 881860 699820 881916
rect 699888 881860 699944 881916
rect 700012 881860 700068 881916
rect 700136 881860 700192 881916
rect 707870 883602 707926 883658
rect 707870 883478 707926 883534
rect 707870 883354 707926 883410
rect 707870 883230 707926 883286
rect 707870 883106 707926 883162
rect 707870 882982 707926 883038
rect 707870 882858 707926 882914
rect 707870 882734 707926 882790
rect 707870 882610 707926 882666
rect 707870 882486 707926 882542
rect 707870 882362 707926 882418
rect 707870 882238 707926 882294
rect 707870 882114 707926 882170
rect 707870 881990 707926 882046
rect 707870 881866 707926 881922
rect 699392 881116 699448 881172
rect 699516 881116 699572 881172
rect 699640 881116 699696 881172
rect 699764 881116 699820 881172
rect 699888 881116 699944 881172
rect 700012 881116 700068 881172
rect 700136 881116 700192 881172
rect 699392 880992 699448 881048
rect 699516 880992 699572 881048
rect 699640 880992 699696 881048
rect 699764 880992 699820 881048
rect 699888 880992 699944 881048
rect 700012 880992 700068 881048
rect 700136 880992 700192 881048
rect 699392 880868 699448 880924
rect 699516 880868 699572 880924
rect 699640 880868 699696 880924
rect 699764 880868 699820 880924
rect 699888 880868 699944 880924
rect 700012 880868 700068 880924
rect 700136 880868 700192 880924
rect 699392 880744 699448 880800
rect 699516 880744 699572 880800
rect 699640 880744 699696 880800
rect 699764 880744 699820 880800
rect 699888 880744 699944 880800
rect 700012 880744 700068 880800
rect 700136 880744 700192 880800
rect 699392 880620 699448 880676
rect 699516 880620 699572 880676
rect 699640 880620 699696 880676
rect 699764 880620 699820 880676
rect 699888 880620 699944 880676
rect 700012 880620 700068 880676
rect 700136 880620 700192 880676
rect 699392 880496 699448 880552
rect 699516 880496 699572 880552
rect 699640 880496 699696 880552
rect 699764 880496 699820 880552
rect 699888 880496 699944 880552
rect 700012 880496 700068 880552
rect 700136 880496 700192 880552
rect 699392 880372 699448 880428
rect 699516 880372 699572 880428
rect 699640 880372 699696 880428
rect 699764 880372 699820 880428
rect 699888 880372 699944 880428
rect 700012 880372 700068 880428
rect 700136 880372 700192 880428
rect 699392 880248 699448 880304
rect 699516 880248 699572 880304
rect 699640 880248 699696 880304
rect 699764 880248 699820 880304
rect 699888 880248 699944 880304
rect 700012 880248 700068 880304
rect 700136 880248 700192 880304
rect 699392 880124 699448 880180
rect 699516 880124 699572 880180
rect 699640 880124 699696 880180
rect 699764 880124 699820 880180
rect 699888 880124 699944 880180
rect 700012 880124 700068 880180
rect 700136 880124 700192 880180
rect 699392 880000 699448 880056
rect 699516 880000 699572 880056
rect 699640 880000 699696 880056
rect 699764 880000 699820 880056
rect 699888 880000 699944 880056
rect 700012 880000 700068 880056
rect 700136 880000 700192 880056
rect 699392 879876 699448 879932
rect 699516 879876 699572 879932
rect 699640 879876 699696 879932
rect 699764 879876 699820 879932
rect 699888 879876 699944 879932
rect 700012 879876 700068 879932
rect 700136 879876 700192 879932
rect 699392 879752 699448 879808
rect 699516 879752 699572 879808
rect 699640 879752 699696 879808
rect 699764 879752 699820 879808
rect 699888 879752 699944 879808
rect 700012 879752 700068 879808
rect 700136 879752 700192 879808
rect 699392 879628 699448 879684
rect 699516 879628 699572 879684
rect 699640 879628 699696 879684
rect 699764 879628 699820 879684
rect 699888 879628 699944 879684
rect 700012 879628 700068 879684
rect 700136 879628 700192 879684
rect 699392 879504 699448 879560
rect 699516 879504 699572 879560
rect 699640 879504 699696 879560
rect 699764 879504 699820 879560
rect 699888 879504 699944 879560
rect 700012 879504 700068 879560
rect 700136 879504 700192 879560
rect 699392 879380 699448 879436
rect 699516 879380 699572 879436
rect 699640 879380 699696 879436
rect 699764 879380 699820 879436
rect 699888 879380 699944 879436
rect 700012 879380 700068 879436
rect 700136 879380 700192 879436
rect 699392 879256 699448 879312
rect 699516 879256 699572 879312
rect 699640 879256 699696 879312
rect 699764 879256 699820 879312
rect 699888 879256 699944 879312
rect 700012 879256 700068 879312
rect 700136 879256 700192 879312
rect 707870 881122 707926 881178
rect 707870 880998 707926 881054
rect 707870 880874 707926 880930
rect 707870 880750 707926 880806
rect 707870 880626 707926 880682
rect 707870 880502 707926 880558
rect 707870 880378 707926 880434
rect 707870 880254 707926 880310
rect 707870 880130 707926 880186
rect 707870 880006 707926 880062
rect 707870 879882 707926 879938
rect 707870 879758 707926 879814
rect 707870 879634 707926 879690
rect 707870 879510 707926 879566
rect 707870 879386 707926 879442
rect 707870 879262 707926 879318
rect 699392 878746 699448 878802
rect 699516 878746 699572 878802
rect 699640 878746 699696 878802
rect 699764 878746 699820 878802
rect 699888 878746 699944 878802
rect 700012 878746 700068 878802
rect 700136 878746 700192 878802
rect 699392 878622 699448 878678
rect 699516 878622 699572 878678
rect 699640 878622 699696 878678
rect 699764 878622 699820 878678
rect 699888 878622 699944 878678
rect 700012 878622 700068 878678
rect 700136 878622 700192 878678
rect 699392 878498 699448 878554
rect 699516 878498 699572 878554
rect 699640 878498 699696 878554
rect 699764 878498 699820 878554
rect 699888 878498 699944 878554
rect 700012 878498 700068 878554
rect 700136 878498 700192 878554
rect 699392 878374 699448 878430
rect 699516 878374 699572 878430
rect 699640 878374 699696 878430
rect 699764 878374 699820 878430
rect 699888 878374 699944 878430
rect 700012 878374 700068 878430
rect 700136 878374 700192 878430
rect 699392 878250 699448 878306
rect 699516 878250 699572 878306
rect 699640 878250 699696 878306
rect 699764 878250 699820 878306
rect 699888 878250 699944 878306
rect 700012 878250 700068 878306
rect 700136 878250 700192 878306
rect 699392 878126 699448 878182
rect 699516 878126 699572 878182
rect 699640 878126 699696 878182
rect 699764 878126 699820 878182
rect 699888 878126 699944 878182
rect 700012 878126 700068 878182
rect 700136 878126 700192 878182
rect 699392 878002 699448 878058
rect 699516 878002 699572 878058
rect 699640 878002 699696 878058
rect 699764 878002 699820 878058
rect 699888 878002 699944 878058
rect 700012 878002 700068 878058
rect 700136 878002 700192 878058
rect 699392 877878 699448 877934
rect 699516 877878 699572 877934
rect 699640 877878 699696 877934
rect 699764 877878 699820 877934
rect 699888 877878 699944 877934
rect 700012 877878 700068 877934
rect 700136 877878 700192 877934
rect 699392 877754 699448 877810
rect 699516 877754 699572 877810
rect 699640 877754 699696 877810
rect 699764 877754 699820 877810
rect 699888 877754 699944 877810
rect 700012 877754 700068 877810
rect 700136 877754 700192 877810
rect 699392 877630 699448 877686
rect 699516 877630 699572 877686
rect 699640 877630 699696 877686
rect 699764 877630 699820 877686
rect 699888 877630 699944 877686
rect 700012 877630 700068 877686
rect 700136 877630 700192 877686
rect 699392 877506 699448 877562
rect 699516 877506 699572 877562
rect 699640 877506 699696 877562
rect 699764 877506 699820 877562
rect 699888 877506 699944 877562
rect 700012 877506 700068 877562
rect 700136 877506 700192 877562
rect 699392 877382 699448 877438
rect 699516 877382 699572 877438
rect 699640 877382 699696 877438
rect 699764 877382 699820 877438
rect 699888 877382 699944 877438
rect 700012 877382 700068 877438
rect 700136 877382 700192 877438
rect 699392 877258 699448 877314
rect 699516 877258 699572 877314
rect 699640 877258 699696 877314
rect 699764 877258 699820 877314
rect 699888 877258 699944 877314
rect 700012 877258 700068 877314
rect 700136 877258 700192 877314
rect 699392 877134 699448 877190
rect 699516 877134 699572 877190
rect 699640 877134 699696 877190
rect 699764 877134 699820 877190
rect 699888 877134 699944 877190
rect 700012 877134 700068 877190
rect 700136 877134 700192 877190
rect 699392 877010 699448 877066
rect 699516 877010 699572 877066
rect 699640 877010 699696 877066
rect 699764 877010 699820 877066
rect 699888 877010 699944 877066
rect 700012 877010 700068 877066
rect 700136 877010 700192 877066
rect 699392 876886 699448 876942
rect 699516 876886 699572 876942
rect 699640 876886 699696 876942
rect 699764 876886 699820 876942
rect 699888 876886 699944 876942
rect 700012 876886 700068 876942
rect 700136 876886 700192 876942
rect 707870 878752 707926 878808
rect 707870 878628 707926 878684
rect 707870 878504 707926 878560
rect 707870 878380 707926 878436
rect 707870 878256 707926 878312
rect 707870 878132 707926 878188
rect 707870 878008 707926 878064
rect 707870 877884 707926 877940
rect 707870 877760 707926 877816
rect 707870 877636 707926 877692
rect 707870 877512 707926 877568
rect 707870 877388 707926 877444
rect 707870 877264 707926 877320
rect 707870 877140 707926 877196
rect 707870 877016 707926 877072
rect 707870 876892 707926 876948
rect 699392 876040 699448 876096
rect 699516 876040 699572 876096
rect 699640 876040 699696 876096
rect 699764 876040 699820 876096
rect 699888 876040 699944 876096
rect 700012 876040 700068 876096
rect 700136 876040 700192 876096
rect 699392 875916 699448 875972
rect 699516 875916 699572 875972
rect 699640 875916 699696 875972
rect 699764 875916 699820 875972
rect 699888 875916 699944 875972
rect 700012 875916 700068 875972
rect 700136 875916 700192 875972
rect 699392 875792 699448 875848
rect 699516 875792 699572 875848
rect 699640 875792 699696 875848
rect 699764 875792 699820 875848
rect 699888 875792 699944 875848
rect 700012 875792 700068 875848
rect 700136 875792 700192 875848
rect 699392 875668 699448 875724
rect 699516 875668 699572 875724
rect 699640 875668 699696 875724
rect 699764 875668 699820 875724
rect 699888 875668 699944 875724
rect 700012 875668 700068 875724
rect 700136 875668 700192 875724
rect 699392 875544 699448 875600
rect 699516 875544 699572 875600
rect 699640 875544 699696 875600
rect 699764 875544 699820 875600
rect 699888 875544 699944 875600
rect 700012 875544 700068 875600
rect 700136 875544 700192 875600
rect 699392 875420 699448 875476
rect 699516 875420 699572 875476
rect 699640 875420 699696 875476
rect 699764 875420 699820 875476
rect 699888 875420 699944 875476
rect 700012 875420 700068 875476
rect 700136 875420 700192 875476
rect 699392 875296 699448 875352
rect 699516 875296 699572 875352
rect 699640 875296 699696 875352
rect 699764 875296 699820 875352
rect 699888 875296 699944 875352
rect 700012 875296 700068 875352
rect 700136 875296 700192 875352
rect 699392 875172 699448 875228
rect 699516 875172 699572 875228
rect 699640 875172 699696 875228
rect 699764 875172 699820 875228
rect 699888 875172 699944 875228
rect 700012 875172 700068 875228
rect 700136 875172 700192 875228
rect 699392 875048 699448 875104
rect 699516 875048 699572 875104
rect 699640 875048 699696 875104
rect 699764 875048 699820 875104
rect 699888 875048 699944 875104
rect 700012 875048 700068 875104
rect 700136 875048 700192 875104
rect 699392 874924 699448 874980
rect 699516 874924 699572 874980
rect 699640 874924 699696 874980
rect 699764 874924 699820 874980
rect 699888 874924 699944 874980
rect 700012 874924 700068 874980
rect 700136 874924 700192 874980
rect 699392 874800 699448 874856
rect 699516 874800 699572 874856
rect 699640 874800 699696 874856
rect 699764 874800 699820 874856
rect 699888 874800 699944 874856
rect 700012 874800 700068 874856
rect 700136 874800 700192 874856
rect 699392 874676 699448 874732
rect 699516 874676 699572 874732
rect 699640 874676 699696 874732
rect 699764 874676 699820 874732
rect 699888 874676 699944 874732
rect 700012 874676 700068 874732
rect 700136 874676 700192 874732
rect 699392 874552 699448 874608
rect 699516 874552 699572 874608
rect 699640 874552 699696 874608
rect 699764 874552 699820 874608
rect 699888 874552 699944 874608
rect 700012 874552 700068 874608
rect 700136 874552 700192 874608
rect 699392 874428 699448 874484
rect 699516 874428 699572 874484
rect 699640 874428 699696 874484
rect 699764 874428 699820 874484
rect 699888 874428 699944 874484
rect 700012 874428 700068 874484
rect 700136 874428 700192 874484
rect 699392 874304 699448 874360
rect 699516 874304 699572 874360
rect 699640 874304 699696 874360
rect 699764 874304 699820 874360
rect 699888 874304 699944 874360
rect 700012 874304 700068 874360
rect 700136 874304 700192 874360
rect 699392 874180 699448 874236
rect 699516 874180 699572 874236
rect 699640 874180 699696 874236
rect 699764 874180 699820 874236
rect 699888 874180 699944 874236
rect 700012 874180 700068 874236
rect 700136 874180 700192 874236
rect 707870 876046 707926 876102
rect 707870 875922 707926 875978
rect 707870 875798 707926 875854
rect 707870 875674 707926 875730
rect 707870 875550 707926 875606
rect 707870 875426 707926 875482
rect 707870 875302 707926 875358
rect 707870 875178 707926 875234
rect 707870 875054 707926 875110
rect 707870 874930 707926 874986
rect 707870 874806 707926 874862
rect 707870 874682 707926 874738
rect 707870 874558 707926 874614
rect 707870 874434 707926 874490
rect 707870 874310 707926 874366
rect 707870 874186 707926 874242
rect 699392 873670 699448 873726
rect 699516 873670 699572 873726
rect 699640 873670 699696 873726
rect 699764 873670 699820 873726
rect 699888 873670 699944 873726
rect 700012 873670 700068 873726
rect 700136 873670 700192 873726
rect 699392 873546 699448 873602
rect 699516 873546 699572 873602
rect 699640 873546 699696 873602
rect 699764 873546 699820 873602
rect 699888 873546 699944 873602
rect 700012 873546 700068 873602
rect 700136 873546 700192 873602
rect 699392 873422 699448 873478
rect 699516 873422 699572 873478
rect 699640 873422 699696 873478
rect 699764 873422 699820 873478
rect 699888 873422 699944 873478
rect 700012 873422 700068 873478
rect 700136 873422 700192 873478
rect 699392 873298 699448 873354
rect 699516 873298 699572 873354
rect 699640 873298 699696 873354
rect 699764 873298 699820 873354
rect 699888 873298 699944 873354
rect 700012 873298 700068 873354
rect 700136 873298 700192 873354
rect 699392 873174 699448 873230
rect 699516 873174 699572 873230
rect 699640 873174 699696 873230
rect 699764 873174 699820 873230
rect 699888 873174 699944 873230
rect 700012 873174 700068 873230
rect 700136 873174 700192 873230
rect 699392 873050 699448 873106
rect 699516 873050 699572 873106
rect 699640 873050 699696 873106
rect 699764 873050 699820 873106
rect 699888 873050 699944 873106
rect 700012 873050 700068 873106
rect 700136 873050 700192 873106
rect 699392 872926 699448 872982
rect 699516 872926 699572 872982
rect 699640 872926 699696 872982
rect 699764 872926 699820 872982
rect 699888 872926 699944 872982
rect 700012 872926 700068 872982
rect 700136 872926 700192 872982
rect 699392 872802 699448 872858
rect 699516 872802 699572 872858
rect 699640 872802 699696 872858
rect 699764 872802 699820 872858
rect 699888 872802 699944 872858
rect 700012 872802 700068 872858
rect 700136 872802 700192 872858
rect 699392 872678 699448 872734
rect 699516 872678 699572 872734
rect 699640 872678 699696 872734
rect 699764 872678 699820 872734
rect 699888 872678 699944 872734
rect 700012 872678 700068 872734
rect 700136 872678 700192 872734
rect 699392 872554 699448 872610
rect 699516 872554 699572 872610
rect 699640 872554 699696 872610
rect 699764 872554 699820 872610
rect 699888 872554 699944 872610
rect 700012 872554 700068 872610
rect 700136 872554 700192 872610
rect 699392 872430 699448 872486
rect 699516 872430 699572 872486
rect 699640 872430 699696 872486
rect 699764 872430 699820 872486
rect 699888 872430 699944 872486
rect 700012 872430 700068 872486
rect 700136 872430 700192 872486
rect 699392 872306 699448 872362
rect 699516 872306 699572 872362
rect 699640 872306 699696 872362
rect 699764 872306 699820 872362
rect 699888 872306 699944 872362
rect 700012 872306 700068 872362
rect 700136 872306 700192 872362
rect 699392 872182 699448 872238
rect 699516 872182 699572 872238
rect 699640 872182 699696 872238
rect 699764 872182 699820 872238
rect 699888 872182 699944 872238
rect 700012 872182 700068 872238
rect 700136 872182 700192 872238
rect 699392 872058 699448 872114
rect 699516 872058 699572 872114
rect 699640 872058 699696 872114
rect 699764 872058 699820 872114
rect 699888 872058 699944 872114
rect 700012 872058 700068 872114
rect 700136 872058 700192 872114
rect 699392 871934 699448 871990
rect 699516 871934 699572 871990
rect 699640 871934 699696 871990
rect 699764 871934 699820 871990
rect 699888 871934 699944 871990
rect 700012 871934 700068 871990
rect 700136 871934 700192 871990
rect 699392 871810 699448 871866
rect 699516 871810 699572 871866
rect 699640 871810 699696 871866
rect 699764 871810 699820 871866
rect 699888 871810 699944 871866
rect 700012 871810 700068 871866
rect 700136 871810 700192 871866
rect 707870 873676 707926 873732
rect 707870 873552 707926 873608
rect 707870 873428 707926 873484
rect 707870 873304 707926 873360
rect 707870 873180 707926 873236
rect 707870 873056 707926 873112
rect 707870 872932 707926 872988
rect 707870 872808 707926 872864
rect 707870 872684 707926 872740
rect 707870 872560 707926 872616
rect 707870 872436 707926 872492
rect 707870 872312 707926 872368
rect 707870 872188 707926 872244
rect 707870 872064 707926 872120
rect 707870 871940 707926 871996
rect 707870 871816 707926 871872
rect 699392 871066 699448 871122
rect 699516 871066 699572 871122
rect 699640 871066 699696 871122
rect 699764 871066 699820 871122
rect 699888 871066 699944 871122
rect 700012 871066 700068 871122
rect 700136 871066 700192 871122
rect 699392 870942 699448 870998
rect 699516 870942 699572 870998
rect 699640 870942 699696 870998
rect 699764 870942 699820 870998
rect 699888 870942 699944 870998
rect 700012 870942 700068 870998
rect 700136 870942 700192 870998
rect 699392 870818 699448 870874
rect 699516 870818 699572 870874
rect 699640 870818 699696 870874
rect 699764 870818 699820 870874
rect 699888 870818 699944 870874
rect 700012 870818 700068 870874
rect 700136 870818 700192 870874
rect 699392 870694 699448 870750
rect 699516 870694 699572 870750
rect 699640 870694 699696 870750
rect 699764 870694 699820 870750
rect 699888 870694 699944 870750
rect 700012 870694 700068 870750
rect 700136 870694 700192 870750
rect 699392 870570 699448 870626
rect 699516 870570 699572 870626
rect 699640 870570 699696 870626
rect 699764 870570 699820 870626
rect 699888 870570 699944 870626
rect 700012 870570 700068 870626
rect 700136 870570 700192 870626
rect 699392 870446 699448 870502
rect 699516 870446 699572 870502
rect 699640 870446 699696 870502
rect 699764 870446 699820 870502
rect 699888 870446 699944 870502
rect 700012 870446 700068 870502
rect 700136 870446 700192 870502
rect 699392 870322 699448 870378
rect 699516 870322 699572 870378
rect 699640 870322 699696 870378
rect 699764 870322 699820 870378
rect 699888 870322 699944 870378
rect 700012 870322 700068 870378
rect 700136 870322 700192 870378
rect 699392 870198 699448 870254
rect 699516 870198 699572 870254
rect 699640 870198 699696 870254
rect 699764 870198 699820 870254
rect 699888 870198 699944 870254
rect 700012 870198 700068 870254
rect 700136 870198 700192 870254
rect 699392 870074 699448 870130
rect 699516 870074 699572 870130
rect 699640 870074 699696 870130
rect 699764 870074 699820 870130
rect 699888 870074 699944 870130
rect 700012 870074 700068 870130
rect 700136 870074 700192 870130
rect 699392 869950 699448 870006
rect 699516 869950 699572 870006
rect 699640 869950 699696 870006
rect 699764 869950 699820 870006
rect 699888 869950 699944 870006
rect 700012 869950 700068 870006
rect 700136 869950 700192 870006
rect 699392 869826 699448 869882
rect 699516 869826 699572 869882
rect 699640 869826 699696 869882
rect 699764 869826 699820 869882
rect 699888 869826 699944 869882
rect 700012 869826 700068 869882
rect 700136 869826 700192 869882
rect 699392 869702 699448 869758
rect 699516 869702 699572 869758
rect 699640 869702 699696 869758
rect 699764 869702 699820 869758
rect 699888 869702 699944 869758
rect 700012 869702 700068 869758
rect 700136 869702 700192 869758
rect 699392 869578 699448 869634
rect 699516 869578 699572 869634
rect 699640 869578 699696 869634
rect 699764 869578 699820 869634
rect 699888 869578 699944 869634
rect 700012 869578 700068 869634
rect 700136 869578 700192 869634
rect 699392 869454 699448 869510
rect 699516 869454 699572 869510
rect 699640 869454 699696 869510
rect 699764 869454 699820 869510
rect 699888 869454 699944 869510
rect 700012 869454 700068 869510
rect 700136 869454 700192 869510
rect 699392 869330 699448 869386
rect 699516 869330 699572 869386
rect 699640 869330 699696 869386
rect 699764 869330 699820 869386
rect 699888 869330 699944 869386
rect 700012 869330 700068 869386
rect 700136 869330 700192 869386
rect 707870 871078 707926 871134
rect 707870 870954 707926 871010
rect 707870 870830 707926 870886
rect 707870 870706 707926 870762
rect 707870 870582 707926 870638
rect 707870 870458 707926 870514
rect 707870 870334 707926 870390
rect 707870 870210 707926 870266
rect 707870 870086 707926 870142
rect 707870 869962 707926 870018
rect 707870 869838 707926 869894
rect 707870 869714 707926 869770
rect 707870 869590 707926 869646
rect 707870 869466 707926 869522
rect 707870 869342 707926 869398
rect 699544 842373 699600 842429
rect 699844 842373 699900 842429
rect 700144 842373 700200 842429
rect 699544 842173 699600 842229
rect 699844 842173 699900 842229
rect 700144 842173 700200 842229
rect 699444 839898 699500 839954
rect 699744 839898 699800 839954
rect 700044 839898 700100 839954
rect 699444 832898 699500 832954
rect 699744 832898 699800 832954
rect 700044 832898 700100 832954
rect 699444 825898 699500 825954
rect 699744 825898 699800 825954
rect 700044 825898 700100 825954
rect 699497 806367 699553 806423
rect 699797 806367 699853 806423
rect 700097 806367 700153 806423
rect 699392 797596 699448 797652
rect 699516 797596 699572 797652
rect 699640 797596 699696 797652
rect 699764 797596 699820 797652
rect 699888 797596 699944 797652
rect 700012 797596 700068 797652
rect 700136 797596 700192 797652
rect 699392 797472 699448 797528
rect 699516 797472 699572 797528
rect 699640 797472 699696 797528
rect 699764 797472 699820 797528
rect 699888 797472 699944 797528
rect 700012 797472 700068 797528
rect 700136 797472 700192 797528
rect 699392 797348 699448 797404
rect 699516 797348 699572 797404
rect 699640 797348 699696 797404
rect 699764 797348 699820 797404
rect 699888 797348 699944 797404
rect 700012 797348 700068 797404
rect 700136 797348 700192 797404
rect 699392 797224 699448 797280
rect 699516 797224 699572 797280
rect 699640 797224 699696 797280
rect 699764 797224 699820 797280
rect 699888 797224 699944 797280
rect 700012 797224 700068 797280
rect 700136 797224 700192 797280
rect 699392 797100 699448 797156
rect 699516 797100 699572 797156
rect 699640 797100 699696 797156
rect 699764 797100 699820 797156
rect 699888 797100 699944 797156
rect 700012 797100 700068 797156
rect 700136 797100 700192 797156
rect 699392 796976 699448 797032
rect 699516 796976 699572 797032
rect 699640 796976 699696 797032
rect 699764 796976 699820 797032
rect 699888 796976 699944 797032
rect 700012 796976 700068 797032
rect 700136 796976 700192 797032
rect 699392 796852 699448 796908
rect 699516 796852 699572 796908
rect 699640 796852 699696 796908
rect 699764 796852 699820 796908
rect 699888 796852 699944 796908
rect 700012 796852 700068 796908
rect 700136 796852 700192 796908
rect 699392 796728 699448 796784
rect 699516 796728 699572 796784
rect 699640 796728 699696 796784
rect 699764 796728 699820 796784
rect 699888 796728 699944 796784
rect 700012 796728 700068 796784
rect 700136 796728 700192 796784
rect 699392 796604 699448 796660
rect 699516 796604 699572 796660
rect 699640 796604 699696 796660
rect 699764 796604 699820 796660
rect 699888 796604 699944 796660
rect 700012 796604 700068 796660
rect 700136 796604 700192 796660
rect 699392 796480 699448 796536
rect 699516 796480 699572 796536
rect 699640 796480 699696 796536
rect 699764 796480 699820 796536
rect 699888 796480 699944 796536
rect 700012 796480 700068 796536
rect 700136 796480 700192 796536
rect 699392 796356 699448 796412
rect 699516 796356 699572 796412
rect 699640 796356 699696 796412
rect 699764 796356 699820 796412
rect 699888 796356 699944 796412
rect 700012 796356 700068 796412
rect 700136 796356 700192 796412
rect 699392 796232 699448 796288
rect 699516 796232 699572 796288
rect 699640 796232 699696 796288
rect 699764 796232 699820 796288
rect 699888 796232 699944 796288
rect 700012 796232 700068 796288
rect 700136 796232 700192 796288
rect 699392 796108 699448 796164
rect 699516 796108 699572 796164
rect 699640 796108 699696 796164
rect 699764 796108 699820 796164
rect 699888 796108 699944 796164
rect 700012 796108 700068 796164
rect 700136 796108 700192 796164
rect 699392 795984 699448 796040
rect 699516 795984 699572 796040
rect 699640 795984 699696 796040
rect 699764 795984 699820 796040
rect 699888 795984 699944 796040
rect 700012 795984 700068 796040
rect 700136 795984 700192 796040
rect 699392 795860 699448 795916
rect 699516 795860 699572 795916
rect 699640 795860 699696 795916
rect 699764 795860 699820 795916
rect 699888 795860 699944 795916
rect 700012 795860 700068 795916
rect 700136 795860 700192 795916
rect 707870 797602 707926 797658
rect 707870 797478 707926 797534
rect 707870 797354 707926 797410
rect 707870 797230 707926 797286
rect 707870 797106 707926 797162
rect 707870 796982 707926 797038
rect 707870 796858 707926 796914
rect 707870 796734 707926 796790
rect 707870 796610 707926 796666
rect 707870 796486 707926 796542
rect 707870 796362 707926 796418
rect 707870 796238 707926 796294
rect 707870 796114 707926 796170
rect 707870 795990 707926 796046
rect 707870 795866 707926 795922
rect 699392 795116 699448 795172
rect 699516 795116 699572 795172
rect 699640 795116 699696 795172
rect 699764 795116 699820 795172
rect 699888 795116 699944 795172
rect 700012 795116 700068 795172
rect 700136 795116 700192 795172
rect 699392 794992 699448 795048
rect 699516 794992 699572 795048
rect 699640 794992 699696 795048
rect 699764 794992 699820 795048
rect 699888 794992 699944 795048
rect 700012 794992 700068 795048
rect 700136 794992 700192 795048
rect 699392 794868 699448 794924
rect 699516 794868 699572 794924
rect 699640 794868 699696 794924
rect 699764 794868 699820 794924
rect 699888 794868 699944 794924
rect 700012 794868 700068 794924
rect 700136 794868 700192 794924
rect 699392 794744 699448 794800
rect 699516 794744 699572 794800
rect 699640 794744 699696 794800
rect 699764 794744 699820 794800
rect 699888 794744 699944 794800
rect 700012 794744 700068 794800
rect 700136 794744 700192 794800
rect 699392 794620 699448 794676
rect 699516 794620 699572 794676
rect 699640 794620 699696 794676
rect 699764 794620 699820 794676
rect 699888 794620 699944 794676
rect 700012 794620 700068 794676
rect 700136 794620 700192 794676
rect 699392 794496 699448 794552
rect 699516 794496 699572 794552
rect 699640 794496 699696 794552
rect 699764 794496 699820 794552
rect 699888 794496 699944 794552
rect 700012 794496 700068 794552
rect 700136 794496 700192 794552
rect 699392 794372 699448 794428
rect 699516 794372 699572 794428
rect 699640 794372 699696 794428
rect 699764 794372 699820 794428
rect 699888 794372 699944 794428
rect 700012 794372 700068 794428
rect 700136 794372 700192 794428
rect 699392 794248 699448 794304
rect 699516 794248 699572 794304
rect 699640 794248 699696 794304
rect 699764 794248 699820 794304
rect 699888 794248 699944 794304
rect 700012 794248 700068 794304
rect 700136 794248 700192 794304
rect 699392 794124 699448 794180
rect 699516 794124 699572 794180
rect 699640 794124 699696 794180
rect 699764 794124 699820 794180
rect 699888 794124 699944 794180
rect 700012 794124 700068 794180
rect 700136 794124 700192 794180
rect 699392 794000 699448 794056
rect 699516 794000 699572 794056
rect 699640 794000 699696 794056
rect 699764 794000 699820 794056
rect 699888 794000 699944 794056
rect 700012 794000 700068 794056
rect 700136 794000 700192 794056
rect 699392 793876 699448 793932
rect 699516 793876 699572 793932
rect 699640 793876 699696 793932
rect 699764 793876 699820 793932
rect 699888 793876 699944 793932
rect 700012 793876 700068 793932
rect 700136 793876 700192 793932
rect 699392 793752 699448 793808
rect 699516 793752 699572 793808
rect 699640 793752 699696 793808
rect 699764 793752 699820 793808
rect 699888 793752 699944 793808
rect 700012 793752 700068 793808
rect 700136 793752 700192 793808
rect 699392 793628 699448 793684
rect 699516 793628 699572 793684
rect 699640 793628 699696 793684
rect 699764 793628 699820 793684
rect 699888 793628 699944 793684
rect 700012 793628 700068 793684
rect 700136 793628 700192 793684
rect 699392 793504 699448 793560
rect 699516 793504 699572 793560
rect 699640 793504 699696 793560
rect 699764 793504 699820 793560
rect 699888 793504 699944 793560
rect 700012 793504 700068 793560
rect 700136 793504 700192 793560
rect 699392 793380 699448 793436
rect 699516 793380 699572 793436
rect 699640 793380 699696 793436
rect 699764 793380 699820 793436
rect 699888 793380 699944 793436
rect 700012 793380 700068 793436
rect 700136 793380 700192 793436
rect 699392 793256 699448 793312
rect 699516 793256 699572 793312
rect 699640 793256 699696 793312
rect 699764 793256 699820 793312
rect 699888 793256 699944 793312
rect 700012 793256 700068 793312
rect 700136 793256 700192 793312
rect 707870 795122 707926 795178
rect 707870 794998 707926 795054
rect 707870 794874 707926 794930
rect 707870 794750 707926 794806
rect 707870 794626 707926 794682
rect 707870 794502 707926 794558
rect 707870 794378 707926 794434
rect 707870 794254 707926 794310
rect 707870 794130 707926 794186
rect 707870 794006 707926 794062
rect 707870 793882 707926 793938
rect 707870 793758 707926 793814
rect 707870 793634 707926 793690
rect 707870 793510 707926 793566
rect 707870 793386 707926 793442
rect 707870 793262 707926 793318
rect 699392 792746 699448 792802
rect 699516 792746 699572 792802
rect 699640 792746 699696 792802
rect 699764 792746 699820 792802
rect 699888 792746 699944 792802
rect 700012 792746 700068 792802
rect 700136 792746 700192 792802
rect 699392 792622 699448 792678
rect 699516 792622 699572 792678
rect 699640 792622 699696 792678
rect 699764 792622 699820 792678
rect 699888 792622 699944 792678
rect 700012 792622 700068 792678
rect 700136 792622 700192 792678
rect 699392 792498 699448 792554
rect 699516 792498 699572 792554
rect 699640 792498 699696 792554
rect 699764 792498 699820 792554
rect 699888 792498 699944 792554
rect 700012 792498 700068 792554
rect 700136 792498 700192 792554
rect 699392 792374 699448 792430
rect 699516 792374 699572 792430
rect 699640 792374 699696 792430
rect 699764 792374 699820 792430
rect 699888 792374 699944 792430
rect 700012 792374 700068 792430
rect 700136 792374 700192 792430
rect 699392 792250 699448 792306
rect 699516 792250 699572 792306
rect 699640 792250 699696 792306
rect 699764 792250 699820 792306
rect 699888 792250 699944 792306
rect 700012 792250 700068 792306
rect 700136 792250 700192 792306
rect 699392 792126 699448 792182
rect 699516 792126 699572 792182
rect 699640 792126 699696 792182
rect 699764 792126 699820 792182
rect 699888 792126 699944 792182
rect 700012 792126 700068 792182
rect 700136 792126 700192 792182
rect 699392 792002 699448 792058
rect 699516 792002 699572 792058
rect 699640 792002 699696 792058
rect 699764 792002 699820 792058
rect 699888 792002 699944 792058
rect 700012 792002 700068 792058
rect 700136 792002 700192 792058
rect 699392 791878 699448 791934
rect 699516 791878 699572 791934
rect 699640 791878 699696 791934
rect 699764 791878 699820 791934
rect 699888 791878 699944 791934
rect 700012 791878 700068 791934
rect 700136 791878 700192 791934
rect 699392 791754 699448 791810
rect 699516 791754 699572 791810
rect 699640 791754 699696 791810
rect 699764 791754 699820 791810
rect 699888 791754 699944 791810
rect 700012 791754 700068 791810
rect 700136 791754 700192 791810
rect 699392 791630 699448 791686
rect 699516 791630 699572 791686
rect 699640 791630 699696 791686
rect 699764 791630 699820 791686
rect 699888 791630 699944 791686
rect 700012 791630 700068 791686
rect 700136 791630 700192 791686
rect 699392 791506 699448 791562
rect 699516 791506 699572 791562
rect 699640 791506 699696 791562
rect 699764 791506 699820 791562
rect 699888 791506 699944 791562
rect 700012 791506 700068 791562
rect 700136 791506 700192 791562
rect 699392 791382 699448 791438
rect 699516 791382 699572 791438
rect 699640 791382 699696 791438
rect 699764 791382 699820 791438
rect 699888 791382 699944 791438
rect 700012 791382 700068 791438
rect 700136 791382 700192 791438
rect 699392 791258 699448 791314
rect 699516 791258 699572 791314
rect 699640 791258 699696 791314
rect 699764 791258 699820 791314
rect 699888 791258 699944 791314
rect 700012 791258 700068 791314
rect 700136 791258 700192 791314
rect 699392 791134 699448 791190
rect 699516 791134 699572 791190
rect 699640 791134 699696 791190
rect 699764 791134 699820 791190
rect 699888 791134 699944 791190
rect 700012 791134 700068 791190
rect 700136 791134 700192 791190
rect 699392 791010 699448 791066
rect 699516 791010 699572 791066
rect 699640 791010 699696 791066
rect 699764 791010 699820 791066
rect 699888 791010 699944 791066
rect 700012 791010 700068 791066
rect 700136 791010 700192 791066
rect 699392 790886 699448 790942
rect 699516 790886 699572 790942
rect 699640 790886 699696 790942
rect 699764 790886 699820 790942
rect 699888 790886 699944 790942
rect 700012 790886 700068 790942
rect 700136 790886 700192 790942
rect 707870 792752 707926 792808
rect 707870 792628 707926 792684
rect 707870 792504 707926 792560
rect 707870 792380 707926 792436
rect 707870 792256 707926 792312
rect 707870 792132 707926 792188
rect 707870 792008 707926 792064
rect 707870 791884 707926 791940
rect 707870 791760 707926 791816
rect 707870 791636 707926 791692
rect 707870 791512 707926 791568
rect 707870 791388 707926 791444
rect 707870 791264 707926 791320
rect 707870 791140 707926 791196
rect 707870 791016 707926 791072
rect 707870 790892 707926 790948
rect 699392 790040 699448 790096
rect 699516 790040 699572 790096
rect 699640 790040 699696 790096
rect 699764 790040 699820 790096
rect 699888 790040 699944 790096
rect 700012 790040 700068 790096
rect 700136 790040 700192 790096
rect 699392 789916 699448 789972
rect 699516 789916 699572 789972
rect 699640 789916 699696 789972
rect 699764 789916 699820 789972
rect 699888 789916 699944 789972
rect 700012 789916 700068 789972
rect 700136 789916 700192 789972
rect 699392 789792 699448 789848
rect 699516 789792 699572 789848
rect 699640 789792 699696 789848
rect 699764 789792 699820 789848
rect 699888 789792 699944 789848
rect 700012 789792 700068 789848
rect 700136 789792 700192 789848
rect 699392 789668 699448 789724
rect 699516 789668 699572 789724
rect 699640 789668 699696 789724
rect 699764 789668 699820 789724
rect 699888 789668 699944 789724
rect 700012 789668 700068 789724
rect 700136 789668 700192 789724
rect 699392 789544 699448 789600
rect 699516 789544 699572 789600
rect 699640 789544 699696 789600
rect 699764 789544 699820 789600
rect 699888 789544 699944 789600
rect 700012 789544 700068 789600
rect 700136 789544 700192 789600
rect 699392 789420 699448 789476
rect 699516 789420 699572 789476
rect 699640 789420 699696 789476
rect 699764 789420 699820 789476
rect 699888 789420 699944 789476
rect 700012 789420 700068 789476
rect 700136 789420 700192 789476
rect 699392 789296 699448 789352
rect 699516 789296 699572 789352
rect 699640 789296 699696 789352
rect 699764 789296 699820 789352
rect 699888 789296 699944 789352
rect 700012 789296 700068 789352
rect 700136 789296 700192 789352
rect 699392 789172 699448 789228
rect 699516 789172 699572 789228
rect 699640 789172 699696 789228
rect 699764 789172 699820 789228
rect 699888 789172 699944 789228
rect 700012 789172 700068 789228
rect 700136 789172 700192 789228
rect 699392 789048 699448 789104
rect 699516 789048 699572 789104
rect 699640 789048 699696 789104
rect 699764 789048 699820 789104
rect 699888 789048 699944 789104
rect 700012 789048 700068 789104
rect 700136 789048 700192 789104
rect 699392 788924 699448 788980
rect 699516 788924 699572 788980
rect 699640 788924 699696 788980
rect 699764 788924 699820 788980
rect 699888 788924 699944 788980
rect 700012 788924 700068 788980
rect 700136 788924 700192 788980
rect 699392 788800 699448 788856
rect 699516 788800 699572 788856
rect 699640 788800 699696 788856
rect 699764 788800 699820 788856
rect 699888 788800 699944 788856
rect 700012 788800 700068 788856
rect 700136 788800 700192 788856
rect 699392 788676 699448 788732
rect 699516 788676 699572 788732
rect 699640 788676 699696 788732
rect 699764 788676 699820 788732
rect 699888 788676 699944 788732
rect 700012 788676 700068 788732
rect 700136 788676 700192 788732
rect 699392 788552 699448 788608
rect 699516 788552 699572 788608
rect 699640 788552 699696 788608
rect 699764 788552 699820 788608
rect 699888 788552 699944 788608
rect 700012 788552 700068 788608
rect 700136 788552 700192 788608
rect 699392 788428 699448 788484
rect 699516 788428 699572 788484
rect 699640 788428 699696 788484
rect 699764 788428 699820 788484
rect 699888 788428 699944 788484
rect 700012 788428 700068 788484
rect 700136 788428 700192 788484
rect 699392 788304 699448 788360
rect 699516 788304 699572 788360
rect 699640 788304 699696 788360
rect 699764 788304 699820 788360
rect 699888 788304 699944 788360
rect 700012 788304 700068 788360
rect 700136 788304 700192 788360
rect 699392 788180 699448 788236
rect 699516 788180 699572 788236
rect 699640 788180 699696 788236
rect 699764 788180 699820 788236
rect 699888 788180 699944 788236
rect 700012 788180 700068 788236
rect 700136 788180 700192 788236
rect 707870 790046 707926 790102
rect 707870 789922 707926 789978
rect 707870 789798 707926 789854
rect 707870 789674 707926 789730
rect 707870 789550 707926 789606
rect 707870 789426 707926 789482
rect 707870 789302 707926 789358
rect 707870 789178 707926 789234
rect 707870 789054 707926 789110
rect 707870 788930 707926 788986
rect 707870 788806 707926 788862
rect 707870 788682 707926 788738
rect 707870 788558 707926 788614
rect 707870 788434 707926 788490
rect 707870 788310 707926 788366
rect 707870 788186 707926 788242
rect 699392 787670 699448 787726
rect 699516 787670 699572 787726
rect 699640 787670 699696 787726
rect 699764 787670 699820 787726
rect 699888 787670 699944 787726
rect 700012 787670 700068 787726
rect 700136 787670 700192 787726
rect 699392 787546 699448 787602
rect 699516 787546 699572 787602
rect 699640 787546 699696 787602
rect 699764 787546 699820 787602
rect 699888 787546 699944 787602
rect 700012 787546 700068 787602
rect 700136 787546 700192 787602
rect 699392 787422 699448 787478
rect 699516 787422 699572 787478
rect 699640 787422 699696 787478
rect 699764 787422 699820 787478
rect 699888 787422 699944 787478
rect 700012 787422 700068 787478
rect 700136 787422 700192 787478
rect 699392 787298 699448 787354
rect 699516 787298 699572 787354
rect 699640 787298 699696 787354
rect 699764 787298 699820 787354
rect 699888 787298 699944 787354
rect 700012 787298 700068 787354
rect 700136 787298 700192 787354
rect 699392 787174 699448 787230
rect 699516 787174 699572 787230
rect 699640 787174 699696 787230
rect 699764 787174 699820 787230
rect 699888 787174 699944 787230
rect 700012 787174 700068 787230
rect 700136 787174 700192 787230
rect 699392 787050 699448 787106
rect 699516 787050 699572 787106
rect 699640 787050 699696 787106
rect 699764 787050 699820 787106
rect 699888 787050 699944 787106
rect 700012 787050 700068 787106
rect 700136 787050 700192 787106
rect 699392 786926 699448 786982
rect 699516 786926 699572 786982
rect 699640 786926 699696 786982
rect 699764 786926 699820 786982
rect 699888 786926 699944 786982
rect 700012 786926 700068 786982
rect 700136 786926 700192 786982
rect 699392 786802 699448 786858
rect 699516 786802 699572 786858
rect 699640 786802 699696 786858
rect 699764 786802 699820 786858
rect 699888 786802 699944 786858
rect 700012 786802 700068 786858
rect 700136 786802 700192 786858
rect 699392 786678 699448 786734
rect 699516 786678 699572 786734
rect 699640 786678 699696 786734
rect 699764 786678 699820 786734
rect 699888 786678 699944 786734
rect 700012 786678 700068 786734
rect 700136 786678 700192 786734
rect 699392 786554 699448 786610
rect 699516 786554 699572 786610
rect 699640 786554 699696 786610
rect 699764 786554 699820 786610
rect 699888 786554 699944 786610
rect 700012 786554 700068 786610
rect 700136 786554 700192 786610
rect 699392 786430 699448 786486
rect 699516 786430 699572 786486
rect 699640 786430 699696 786486
rect 699764 786430 699820 786486
rect 699888 786430 699944 786486
rect 700012 786430 700068 786486
rect 700136 786430 700192 786486
rect 699392 786306 699448 786362
rect 699516 786306 699572 786362
rect 699640 786306 699696 786362
rect 699764 786306 699820 786362
rect 699888 786306 699944 786362
rect 700012 786306 700068 786362
rect 700136 786306 700192 786362
rect 699392 786182 699448 786238
rect 699516 786182 699572 786238
rect 699640 786182 699696 786238
rect 699764 786182 699820 786238
rect 699888 786182 699944 786238
rect 700012 786182 700068 786238
rect 700136 786182 700192 786238
rect 699392 786058 699448 786114
rect 699516 786058 699572 786114
rect 699640 786058 699696 786114
rect 699764 786058 699820 786114
rect 699888 786058 699944 786114
rect 700012 786058 700068 786114
rect 700136 786058 700192 786114
rect 699392 785934 699448 785990
rect 699516 785934 699572 785990
rect 699640 785934 699696 785990
rect 699764 785934 699820 785990
rect 699888 785934 699944 785990
rect 700012 785934 700068 785990
rect 700136 785934 700192 785990
rect 699392 785810 699448 785866
rect 699516 785810 699572 785866
rect 699640 785810 699696 785866
rect 699764 785810 699820 785866
rect 699888 785810 699944 785866
rect 700012 785810 700068 785866
rect 700136 785810 700192 785866
rect 707870 787676 707926 787732
rect 707870 787552 707926 787608
rect 707870 787428 707926 787484
rect 707870 787304 707926 787360
rect 707870 787180 707926 787236
rect 707870 787056 707926 787112
rect 707870 786932 707926 786988
rect 707870 786808 707926 786864
rect 707870 786684 707926 786740
rect 707870 786560 707926 786616
rect 707870 786436 707926 786492
rect 707870 786312 707926 786368
rect 707870 786188 707926 786244
rect 707870 786064 707926 786120
rect 707870 785940 707926 785996
rect 707870 785816 707926 785872
rect 699392 785066 699448 785122
rect 699516 785066 699572 785122
rect 699640 785066 699696 785122
rect 699764 785066 699820 785122
rect 699888 785066 699944 785122
rect 700012 785066 700068 785122
rect 700136 785066 700192 785122
rect 699392 784942 699448 784998
rect 699516 784942 699572 784998
rect 699640 784942 699696 784998
rect 699764 784942 699820 784998
rect 699888 784942 699944 784998
rect 700012 784942 700068 784998
rect 700136 784942 700192 784998
rect 699392 784818 699448 784874
rect 699516 784818 699572 784874
rect 699640 784818 699696 784874
rect 699764 784818 699820 784874
rect 699888 784818 699944 784874
rect 700012 784818 700068 784874
rect 700136 784818 700192 784874
rect 699392 784694 699448 784750
rect 699516 784694 699572 784750
rect 699640 784694 699696 784750
rect 699764 784694 699820 784750
rect 699888 784694 699944 784750
rect 700012 784694 700068 784750
rect 700136 784694 700192 784750
rect 699392 784570 699448 784626
rect 699516 784570 699572 784626
rect 699640 784570 699696 784626
rect 699764 784570 699820 784626
rect 699888 784570 699944 784626
rect 700012 784570 700068 784626
rect 700136 784570 700192 784626
rect 699392 784446 699448 784502
rect 699516 784446 699572 784502
rect 699640 784446 699696 784502
rect 699764 784446 699820 784502
rect 699888 784446 699944 784502
rect 700012 784446 700068 784502
rect 700136 784446 700192 784502
rect 699392 784322 699448 784378
rect 699516 784322 699572 784378
rect 699640 784322 699696 784378
rect 699764 784322 699820 784378
rect 699888 784322 699944 784378
rect 700012 784322 700068 784378
rect 700136 784322 700192 784378
rect 699392 784198 699448 784254
rect 699516 784198 699572 784254
rect 699640 784198 699696 784254
rect 699764 784198 699820 784254
rect 699888 784198 699944 784254
rect 700012 784198 700068 784254
rect 700136 784198 700192 784254
rect 699392 784074 699448 784130
rect 699516 784074 699572 784130
rect 699640 784074 699696 784130
rect 699764 784074 699820 784130
rect 699888 784074 699944 784130
rect 700012 784074 700068 784130
rect 700136 784074 700192 784130
rect 699392 783950 699448 784006
rect 699516 783950 699572 784006
rect 699640 783950 699696 784006
rect 699764 783950 699820 784006
rect 699888 783950 699944 784006
rect 700012 783950 700068 784006
rect 700136 783950 700192 784006
rect 699392 783826 699448 783882
rect 699516 783826 699572 783882
rect 699640 783826 699696 783882
rect 699764 783826 699820 783882
rect 699888 783826 699944 783882
rect 700012 783826 700068 783882
rect 700136 783826 700192 783882
rect 699392 783702 699448 783758
rect 699516 783702 699572 783758
rect 699640 783702 699696 783758
rect 699764 783702 699820 783758
rect 699888 783702 699944 783758
rect 700012 783702 700068 783758
rect 700136 783702 700192 783758
rect 699392 783578 699448 783634
rect 699516 783578 699572 783634
rect 699640 783578 699696 783634
rect 699764 783578 699820 783634
rect 699888 783578 699944 783634
rect 700012 783578 700068 783634
rect 700136 783578 700192 783634
rect 699392 783454 699448 783510
rect 699516 783454 699572 783510
rect 699640 783454 699696 783510
rect 699764 783454 699820 783510
rect 699888 783454 699944 783510
rect 700012 783454 700068 783510
rect 700136 783454 700192 783510
rect 699392 783330 699448 783386
rect 699516 783330 699572 783386
rect 699640 783330 699696 783386
rect 699764 783330 699820 783386
rect 699888 783330 699944 783386
rect 700012 783330 700068 783386
rect 700136 783330 700192 783386
rect 707870 785078 707926 785134
rect 707870 784954 707926 785010
rect 707870 784830 707926 784886
rect 707870 784706 707926 784762
rect 707870 784582 707926 784638
rect 707870 784458 707926 784514
rect 707870 784334 707926 784390
rect 707870 784210 707926 784266
rect 707870 784086 707926 784142
rect 707870 783962 707926 784018
rect 707870 783838 707926 783894
rect 707870 783714 707926 783770
rect 707870 783590 707926 783646
rect 707870 783466 707926 783522
rect 707870 783342 707926 783398
rect 699544 770373 699600 770429
rect 699844 770373 699900 770429
rect 700144 770373 700200 770429
rect 699544 770173 699600 770229
rect 699844 770173 699900 770229
rect 700144 770173 700200 770229
rect 699444 753898 699500 753954
rect 699744 753898 699800 753954
rect 700044 753898 700100 753954
rect 699444 746898 699500 746954
rect 699744 746898 699800 746954
rect 700044 746898 700100 746954
rect 699444 739898 699500 739954
rect 699744 739898 699800 739954
rect 700044 739898 700100 739954
rect 699544 734373 699600 734429
rect 699844 734373 699900 734429
rect 700144 734373 700200 734429
rect 699544 734173 699600 734229
rect 699844 734173 699900 734229
rect 700144 734173 700200 734229
rect 699497 720367 699553 720423
rect 699797 720367 699853 720423
rect 700097 720367 700153 720423
rect 699444 710898 699500 710954
rect 699744 710898 699800 710954
rect 700044 710898 700100 710954
rect 699444 703898 699500 703954
rect 699744 703898 699800 703954
rect 700044 703898 700100 703954
rect 699544 698373 699600 698429
rect 699844 698373 699900 698429
rect 700144 698373 700200 698429
rect 699544 698173 699600 698229
rect 699844 698173 699900 698229
rect 700144 698173 700200 698229
rect 699444 696898 699500 696954
rect 699744 696898 699800 696954
rect 700044 696898 700100 696954
rect 699497 677367 699553 677423
rect 699797 677367 699853 677423
rect 700097 677367 700153 677423
rect 699444 667898 699500 667954
rect 699744 667898 699800 667954
rect 700044 667898 700100 667954
rect 699544 662373 699600 662429
rect 699844 662373 699900 662429
rect 700144 662373 700200 662429
rect 699544 662173 699600 662229
rect 699844 662173 699900 662229
rect 700144 662173 700200 662229
rect 699444 660898 699500 660954
rect 699744 660898 699800 660954
rect 700044 660898 700100 660954
rect 699444 653898 699500 653954
rect 699744 653898 699800 653954
rect 700044 653898 700100 653954
rect 699497 634367 699553 634423
rect 699797 634367 699853 634423
rect 700097 634367 700153 634423
rect 699544 626373 699600 626429
rect 699844 626373 699900 626429
rect 700144 626373 700200 626429
rect 699544 626173 699600 626229
rect 699844 626173 699900 626229
rect 700144 626173 700200 626229
rect 699444 624898 699500 624954
rect 699744 624898 699800 624954
rect 700044 624898 700100 624954
rect 699444 617898 699500 617954
rect 699744 617898 699800 617954
rect 700044 617898 700100 617954
rect 699444 610898 699500 610954
rect 699744 610898 699800 610954
rect 700044 610898 700100 610954
rect 699497 591367 699553 591423
rect 699797 591367 699853 591423
rect 700097 591367 700153 591423
rect 699544 590373 699600 590429
rect 699844 590373 699900 590429
rect 700144 590373 700200 590429
rect 699544 590173 699600 590229
rect 699844 590173 699900 590229
rect 700144 590173 700200 590229
rect 699444 581898 699500 581954
rect 699744 581898 699800 581954
rect 700044 581898 700100 581954
rect 699444 574898 699500 574954
rect 699744 574898 699800 574954
rect 700044 574898 700100 574954
rect 699444 567898 699500 567954
rect 699744 567898 699800 567954
rect 700044 567898 700100 567954
rect 699544 554373 699600 554429
rect 699844 554373 699900 554429
rect 700144 554373 700200 554429
rect 699544 554173 699600 554229
rect 699844 554173 699900 554229
rect 700144 554173 700200 554229
rect 699497 548367 699553 548423
rect 699797 548367 699853 548423
rect 700097 548367 700153 548423
rect 699444 538898 699500 538954
rect 699744 538898 699800 538954
rect 700044 538898 700100 538954
rect 699444 531898 699500 531954
rect 699744 531898 699800 531954
rect 700044 531898 700100 531954
rect 699444 524898 699500 524954
rect 699744 524898 699800 524954
rect 700044 524898 700100 524954
rect 699544 518373 699600 518429
rect 699844 518373 699900 518429
rect 700144 518373 700200 518429
rect 699544 518173 699600 518229
rect 699844 518173 699900 518229
rect 700144 518173 700200 518229
rect 699497 505367 699553 505423
rect 699797 505367 699853 505423
rect 700097 505367 700153 505423
rect 699392 496596 699448 496652
rect 699516 496596 699572 496652
rect 699640 496596 699696 496652
rect 699764 496596 699820 496652
rect 699888 496596 699944 496652
rect 700012 496596 700068 496652
rect 700136 496596 700192 496652
rect 699392 496472 699448 496528
rect 699516 496472 699572 496528
rect 699640 496472 699696 496528
rect 699764 496472 699820 496528
rect 699888 496472 699944 496528
rect 700012 496472 700068 496528
rect 700136 496472 700192 496528
rect 699392 496348 699448 496404
rect 699516 496348 699572 496404
rect 699640 496348 699696 496404
rect 699764 496348 699820 496404
rect 699888 496348 699944 496404
rect 700012 496348 700068 496404
rect 700136 496348 700192 496404
rect 699392 496224 699448 496280
rect 699516 496224 699572 496280
rect 699640 496224 699696 496280
rect 699764 496224 699820 496280
rect 699888 496224 699944 496280
rect 700012 496224 700068 496280
rect 700136 496224 700192 496280
rect 699392 496100 699448 496156
rect 699516 496100 699572 496156
rect 699640 496100 699696 496156
rect 699764 496100 699820 496156
rect 699888 496100 699944 496156
rect 700012 496100 700068 496156
rect 700136 496100 700192 496156
rect 699392 495976 699448 496032
rect 699516 495976 699572 496032
rect 699640 495976 699696 496032
rect 699764 495976 699820 496032
rect 699888 495976 699944 496032
rect 700012 495976 700068 496032
rect 700136 495976 700192 496032
rect 699392 495852 699448 495908
rect 699516 495852 699572 495908
rect 699640 495852 699696 495908
rect 699764 495852 699820 495908
rect 699888 495852 699944 495908
rect 700012 495852 700068 495908
rect 700136 495852 700192 495908
rect 699392 495728 699448 495784
rect 699516 495728 699572 495784
rect 699640 495728 699696 495784
rect 699764 495728 699820 495784
rect 699888 495728 699944 495784
rect 700012 495728 700068 495784
rect 700136 495728 700192 495784
rect 699392 495604 699448 495660
rect 699516 495604 699572 495660
rect 699640 495604 699696 495660
rect 699764 495604 699820 495660
rect 699888 495604 699944 495660
rect 700012 495604 700068 495660
rect 700136 495604 700192 495660
rect 699392 495480 699448 495536
rect 699516 495480 699572 495536
rect 699640 495480 699696 495536
rect 699764 495480 699820 495536
rect 699888 495480 699944 495536
rect 700012 495480 700068 495536
rect 700136 495480 700192 495536
rect 699392 495356 699448 495412
rect 699516 495356 699572 495412
rect 699640 495356 699696 495412
rect 699764 495356 699820 495412
rect 699888 495356 699944 495412
rect 700012 495356 700068 495412
rect 700136 495356 700192 495412
rect 699392 495232 699448 495288
rect 699516 495232 699572 495288
rect 699640 495232 699696 495288
rect 699764 495232 699820 495288
rect 699888 495232 699944 495288
rect 700012 495232 700068 495288
rect 700136 495232 700192 495288
rect 699392 495108 699448 495164
rect 699516 495108 699572 495164
rect 699640 495108 699696 495164
rect 699764 495108 699820 495164
rect 699888 495108 699944 495164
rect 700012 495108 700068 495164
rect 700136 495108 700192 495164
rect 699392 494984 699448 495040
rect 699516 494984 699572 495040
rect 699640 494984 699696 495040
rect 699764 494984 699820 495040
rect 699888 494984 699944 495040
rect 700012 494984 700068 495040
rect 700136 494984 700192 495040
rect 699392 494860 699448 494916
rect 699516 494860 699572 494916
rect 699640 494860 699696 494916
rect 699764 494860 699820 494916
rect 699888 494860 699944 494916
rect 700012 494860 700068 494916
rect 700136 494860 700192 494916
rect 707870 496602 707926 496658
rect 707870 496478 707926 496534
rect 707870 496354 707926 496410
rect 707870 496230 707926 496286
rect 707870 496106 707926 496162
rect 707870 495982 707926 496038
rect 707870 495858 707926 495914
rect 707870 495734 707926 495790
rect 707870 495610 707926 495666
rect 707870 495486 707926 495542
rect 707870 495362 707926 495418
rect 707870 495238 707926 495294
rect 707870 495114 707926 495170
rect 707870 494990 707926 495046
rect 707870 494866 707926 494922
rect 699392 494116 699448 494172
rect 699516 494116 699572 494172
rect 699640 494116 699696 494172
rect 699764 494116 699820 494172
rect 699888 494116 699944 494172
rect 700012 494116 700068 494172
rect 700136 494116 700192 494172
rect 699392 493992 699448 494048
rect 699516 493992 699572 494048
rect 699640 493992 699696 494048
rect 699764 493992 699820 494048
rect 699888 493992 699944 494048
rect 700012 493992 700068 494048
rect 700136 493992 700192 494048
rect 699392 493868 699448 493924
rect 699516 493868 699572 493924
rect 699640 493868 699696 493924
rect 699764 493868 699820 493924
rect 699888 493868 699944 493924
rect 700012 493868 700068 493924
rect 700136 493868 700192 493924
rect 699392 493744 699448 493800
rect 699516 493744 699572 493800
rect 699640 493744 699696 493800
rect 699764 493744 699820 493800
rect 699888 493744 699944 493800
rect 700012 493744 700068 493800
rect 700136 493744 700192 493800
rect 699392 493620 699448 493676
rect 699516 493620 699572 493676
rect 699640 493620 699696 493676
rect 699764 493620 699820 493676
rect 699888 493620 699944 493676
rect 700012 493620 700068 493676
rect 700136 493620 700192 493676
rect 699392 493496 699448 493552
rect 699516 493496 699572 493552
rect 699640 493496 699696 493552
rect 699764 493496 699820 493552
rect 699888 493496 699944 493552
rect 700012 493496 700068 493552
rect 700136 493496 700192 493552
rect 699392 493372 699448 493428
rect 699516 493372 699572 493428
rect 699640 493372 699696 493428
rect 699764 493372 699820 493428
rect 699888 493372 699944 493428
rect 700012 493372 700068 493428
rect 700136 493372 700192 493428
rect 699392 493248 699448 493304
rect 699516 493248 699572 493304
rect 699640 493248 699696 493304
rect 699764 493248 699820 493304
rect 699888 493248 699944 493304
rect 700012 493248 700068 493304
rect 700136 493248 700192 493304
rect 699392 493124 699448 493180
rect 699516 493124 699572 493180
rect 699640 493124 699696 493180
rect 699764 493124 699820 493180
rect 699888 493124 699944 493180
rect 700012 493124 700068 493180
rect 700136 493124 700192 493180
rect 699392 493000 699448 493056
rect 699516 493000 699572 493056
rect 699640 493000 699696 493056
rect 699764 493000 699820 493056
rect 699888 493000 699944 493056
rect 700012 493000 700068 493056
rect 700136 493000 700192 493056
rect 699392 492876 699448 492932
rect 699516 492876 699572 492932
rect 699640 492876 699696 492932
rect 699764 492876 699820 492932
rect 699888 492876 699944 492932
rect 700012 492876 700068 492932
rect 700136 492876 700192 492932
rect 699392 492752 699448 492808
rect 699516 492752 699572 492808
rect 699640 492752 699696 492808
rect 699764 492752 699820 492808
rect 699888 492752 699944 492808
rect 700012 492752 700068 492808
rect 700136 492752 700192 492808
rect 699392 492628 699448 492684
rect 699516 492628 699572 492684
rect 699640 492628 699696 492684
rect 699764 492628 699820 492684
rect 699888 492628 699944 492684
rect 700012 492628 700068 492684
rect 700136 492628 700192 492684
rect 699392 492504 699448 492560
rect 699516 492504 699572 492560
rect 699640 492504 699696 492560
rect 699764 492504 699820 492560
rect 699888 492504 699944 492560
rect 700012 492504 700068 492560
rect 700136 492504 700192 492560
rect 699392 492380 699448 492436
rect 699516 492380 699572 492436
rect 699640 492380 699696 492436
rect 699764 492380 699820 492436
rect 699888 492380 699944 492436
rect 700012 492380 700068 492436
rect 700136 492380 700192 492436
rect 699392 492256 699448 492312
rect 699516 492256 699572 492312
rect 699640 492256 699696 492312
rect 699764 492256 699820 492312
rect 699888 492256 699944 492312
rect 700012 492256 700068 492312
rect 700136 492256 700192 492312
rect 707870 494122 707926 494178
rect 707870 493998 707926 494054
rect 707870 493874 707926 493930
rect 707870 493750 707926 493806
rect 707870 493626 707926 493682
rect 707870 493502 707926 493558
rect 707870 493378 707926 493434
rect 707870 493254 707926 493310
rect 707870 493130 707926 493186
rect 707870 493006 707926 493062
rect 707870 492882 707926 492938
rect 707870 492758 707926 492814
rect 707870 492634 707926 492690
rect 707870 492510 707926 492566
rect 707870 492386 707926 492442
rect 707870 492262 707926 492318
rect 699392 491746 699448 491802
rect 699516 491746 699572 491802
rect 699640 491746 699696 491802
rect 699764 491746 699820 491802
rect 699888 491746 699944 491802
rect 700012 491746 700068 491802
rect 700136 491746 700192 491802
rect 699392 491622 699448 491678
rect 699516 491622 699572 491678
rect 699640 491622 699696 491678
rect 699764 491622 699820 491678
rect 699888 491622 699944 491678
rect 700012 491622 700068 491678
rect 700136 491622 700192 491678
rect 699392 491498 699448 491554
rect 699516 491498 699572 491554
rect 699640 491498 699696 491554
rect 699764 491498 699820 491554
rect 699888 491498 699944 491554
rect 700012 491498 700068 491554
rect 700136 491498 700192 491554
rect 699392 491374 699448 491430
rect 699516 491374 699572 491430
rect 699640 491374 699696 491430
rect 699764 491374 699820 491430
rect 699888 491374 699944 491430
rect 700012 491374 700068 491430
rect 700136 491374 700192 491430
rect 699392 491250 699448 491306
rect 699516 491250 699572 491306
rect 699640 491250 699696 491306
rect 699764 491250 699820 491306
rect 699888 491250 699944 491306
rect 700012 491250 700068 491306
rect 700136 491250 700192 491306
rect 699392 491126 699448 491182
rect 699516 491126 699572 491182
rect 699640 491126 699696 491182
rect 699764 491126 699820 491182
rect 699888 491126 699944 491182
rect 700012 491126 700068 491182
rect 700136 491126 700192 491182
rect 699392 491002 699448 491058
rect 699516 491002 699572 491058
rect 699640 491002 699696 491058
rect 699764 491002 699820 491058
rect 699888 491002 699944 491058
rect 700012 491002 700068 491058
rect 700136 491002 700192 491058
rect 699392 490878 699448 490934
rect 699516 490878 699572 490934
rect 699640 490878 699696 490934
rect 699764 490878 699820 490934
rect 699888 490878 699944 490934
rect 700012 490878 700068 490934
rect 700136 490878 700192 490934
rect 699392 490754 699448 490810
rect 699516 490754 699572 490810
rect 699640 490754 699696 490810
rect 699764 490754 699820 490810
rect 699888 490754 699944 490810
rect 700012 490754 700068 490810
rect 700136 490754 700192 490810
rect 699392 490630 699448 490686
rect 699516 490630 699572 490686
rect 699640 490630 699696 490686
rect 699764 490630 699820 490686
rect 699888 490630 699944 490686
rect 700012 490630 700068 490686
rect 700136 490630 700192 490686
rect 699392 490506 699448 490562
rect 699516 490506 699572 490562
rect 699640 490506 699696 490562
rect 699764 490506 699820 490562
rect 699888 490506 699944 490562
rect 700012 490506 700068 490562
rect 700136 490506 700192 490562
rect 699392 490382 699448 490438
rect 699516 490382 699572 490438
rect 699640 490382 699696 490438
rect 699764 490382 699820 490438
rect 699888 490382 699944 490438
rect 700012 490382 700068 490438
rect 700136 490382 700192 490438
rect 699392 490258 699448 490314
rect 699516 490258 699572 490314
rect 699640 490258 699696 490314
rect 699764 490258 699820 490314
rect 699888 490258 699944 490314
rect 700012 490258 700068 490314
rect 700136 490258 700192 490314
rect 699392 490134 699448 490190
rect 699516 490134 699572 490190
rect 699640 490134 699696 490190
rect 699764 490134 699820 490190
rect 699888 490134 699944 490190
rect 700012 490134 700068 490190
rect 700136 490134 700192 490190
rect 699392 490010 699448 490066
rect 699516 490010 699572 490066
rect 699640 490010 699696 490066
rect 699764 490010 699820 490066
rect 699888 490010 699944 490066
rect 700012 490010 700068 490066
rect 700136 490010 700192 490066
rect 699392 489886 699448 489942
rect 699516 489886 699572 489942
rect 699640 489886 699696 489942
rect 699764 489886 699820 489942
rect 699888 489886 699944 489942
rect 700012 489886 700068 489942
rect 700136 489886 700192 489942
rect 707870 491752 707926 491808
rect 707870 491628 707926 491684
rect 707870 491504 707926 491560
rect 707870 491380 707926 491436
rect 707870 491256 707926 491312
rect 707870 491132 707926 491188
rect 707870 491008 707926 491064
rect 707870 490884 707926 490940
rect 707870 490760 707926 490816
rect 707870 490636 707926 490692
rect 707870 490512 707926 490568
rect 707870 490388 707926 490444
rect 707870 490264 707926 490320
rect 707870 490140 707926 490196
rect 707870 490016 707926 490072
rect 707870 489892 707926 489948
rect 699392 489040 699448 489096
rect 699516 489040 699572 489096
rect 699640 489040 699696 489096
rect 699764 489040 699820 489096
rect 699888 489040 699944 489096
rect 700012 489040 700068 489096
rect 700136 489040 700192 489096
rect 699392 488916 699448 488972
rect 699516 488916 699572 488972
rect 699640 488916 699696 488972
rect 699764 488916 699820 488972
rect 699888 488916 699944 488972
rect 700012 488916 700068 488972
rect 700136 488916 700192 488972
rect 699392 488792 699448 488848
rect 699516 488792 699572 488848
rect 699640 488792 699696 488848
rect 699764 488792 699820 488848
rect 699888 488792 699944 488848
rect 700012 488792 700068 488848
rect 700136 488792 700192 488848
rect 699392 488668 699448 488724
rect 699516 488668 699572 488724
rect 699640 488668 699696 488724
rect 699764 488668 699820 488724
rect 699888 488668 699944 488724
rect 700012 488668 700068 488724
rect 700136 488668 700192 488724
rect 699392 488544 699448 488600
rect 699516 488544 699572 488600
rect 699640 488544 699696 488600
rect 699764 488544 699820 488600
rect 699888 488544 699944 488600
rect 700012 488544 700068 488600
rect 700136 488544 700192 488600
rect 699392 488420 699448 488476
rect 699516 488420 699572 488476
rect 699640 488420 699696 488476
rect 699764 488420 699820 488476
rect 699888 488420 699944 488476
rect 700012 488420 700068 488476
rect 700136 488420 700192 488476
rect 699392 488296 699448 488352
rect 699516 488296 699572 488352
rect 699640 488296 699696 488352
rect 699764 488296 699820 488352
rect 699888 488296 699944 488352
rect 700012 488296 700068 488352
rect 700136 488296 700192 488352
rect 699392 488172 699448 488228
rect 699516 488172 699572 488228
rect 699640 488172 699696 488228
rect 699764 488172 699820 488228
rect 699888 488172 699944 488228
rect 700012 488172 700068 488228
rect 700136 488172 700192 488228
rect 699392 488048 699448 488104
rect 699516 488048 699572 488104
rect 699640 488048 699696 488104
rect 699764 488048 699820 488104
rect 699888 488048 699944 488104
rect 700012 488048 700068 488104
rect 700136 488048 700192 488104
rect 699392 487924 699448 487980
rect 699516 487924 699572 487980
rect 699640 487924 699696 487980
rect 699764 487924 699820 487980
rect 699888 487924 699944 487980
rect 700012 487924 700068 487980
rect 700136 487924 700192 487980
rect 699392 487800 699448 487856
rect 699516 487800 699572 487856
rect 699640 487800 699696 487856
rect 699764 487800 699820 487856
rect 699888 487800 699944 487856
rect 700012 487800 700068 487856
rect 700136 487800 700192 487856
rect 699392 487676 699448 487732
rect 699516 487676 699572 487732
rect 699640 487676 699696 487732
rect 699764 487676 699820 487732
rect 699888 487676 699944 487732
rect 700012 487676 700068 487732
rect 700136 487676 700192 487732
rect 699392 487552 699448 487608
rect 699516 487552 699572 487608
rect 699640 487552 699696 487608
rect 699764 487552 699820 487608
rect 699888 487552 699944 487608
rect 700012 487552 700068 487608
rect 700136 487552 700192 487608
rect 699392 487428 699448 487484
rect 699516 487428 699572 487484
rect 699640 487428 699696 487484
rect 699764 487428 699820 487484
rect 699888 487428 699944 487484
rect 700012 487428 700068 487484
rect 700136 487428 700192 487484
rect 699392 487304 699448 487360
rect 699516 487304 699572 487360
rect 699640 487304 699696 487360
rect 699764 487304 699820 487360
rect 699888 487304 699944 487360
rect 700012 487304 700068 487360
rect 700136 487304 700192 487360
rect 699392 487180 699448 487236
rect 699516 487180 699572 487236
rect 699640 487180 699696 487236
rect 699764 487180 699820 487236
rect 699888 487180 699944 487236
rect 700012 487180 700068 487236
rect 700136 487180 700192 487236
rect 707870 489046 707926 489102
rect 707870 488922 707926 488978
rect 707870 488798 707926 488854
rect 707870 488674 707926 488730
rect 707870 488550 707926 488606
rect 707870 488426 707926 488482
rect 707870 488302 707926 488358
rect 707870 488178 707926 488234
rect 707870 488054 707926 488110
rect 707870 487930 707926 487986
rect 707870 487806 707926 487862
rect 707870 487682 707926 487738
rect 707870 487558 707926 487614
rect 707870 487434 707926 487490
rect 707870 487310 707926 487366
rect 707870 487186 707926 487242
rect 699392 486670 699448 486726
rect 699516 486670 699572 486726
rect 699640 486670 699696 486726
rect 699764 486670 699820 486726
rect 699888 486670 699944 486726
rect 700012 486670 700068 486726
rect 700136 486670 700192 486726
rect 699392 486546 699448 486602
rect 699516 486546 699572 486602
rect 699640 486546 699696 486602
rect 699764 486546 699820 486602
rect 699888 486546 699944 486602
rect 700012 486546 700068 486602
rect 700136 486546 700192 486602
rect 699392 486422 699448 486478
rect 699516 486422 699572 486478
rect 699640 486422 699696 486478
rect 699764 486422 699820 486478
rect 699888 486422 699944 486478
rect 700012 486422 700068 486478
rect 700136 486422 700192 486478
rect 699392 486298 699448 486354
rect 699516 486298 699572 486354
rect 699640 486298 699696 486354
rect 699764 486298 699820 486354
rect 699888 486298 699944 486354
rect 700012 486298 700068 486354
rect 700136 486298 700192 486354
rect 699392 486174 699448 486230
rect 699516 486174 699572 486230
rect 699640 486174 699696 486230
rect 699764 486174 699820 486230
rect 699888 486174 699944 486230
rect 700012 486174 700068 486230
rect 700136 486174 700192 486230
rect 699392 486050 699448 486106
rect 699516 486050 699572 486106
rect 699640 486050 699696 486106
rect 699764 486050 699820 486106
rect 699888 486050 699944 486106
rect 700012 486050 700068 486106
rect 700136 486050 700192 486106
rect 699392 485926 699448 485982
rect 699516 485926 699572 485982
rect 699640 485926 699696 485982
rect 699764 485926 699820 485982
rect 699888 485926 699944 485982
rect 700012 485926 700068 485982
rect 700136 485926 700192 485982
rect 699392 485802 699448 485858
rect 699516 485802 699572 485858
rect 699640 485802 699696 485858
rect 699764 485802 699820 485858
rect 699888 485802 699944 485858
rect 700012 485802 700068 485858
rect 700136 485802 700192 485858
rect 699392 485678 699448 485734
rect 699516 485678 699572 485734
rect 699640 485678 699696 485734
rect 699764 485678 699820 485734
rect 699888 485678 699944 485734
rect 700012 485678 700068 485734
rect 700136 485678 700192 485734
rect 699392 485554 699448 485610
rect 699516 485554 699572 485610
rect 699640 485554 699696 485610
rect 699764 485554 699820 485610
rect 699888 485554 699944 485610
rect 700012 485554 700068 485610
rect 700136 485554 700192 485610
rect 699392 485430 699448 485486
rect 699516 485430 699572 485486
rect 699640 485430 699696 485486
rect 699764 485430 699820 485486
rect 699888 485430 699944 485486
rect 700012 485430 700068 485486
rect 700136 485430 700192 485486
rect 699392 485306 699448 485362
rect 699516 485306 699572 485362
rect 699640 485306 699696 485362
rect 699764 485306 699820 485362
rect 699888 485306 699944 485362
rect 700012 485306 700068 485362
rect 700136 485306 700192 485362
rect 699392 485182 699448 485238
rect 699516 485182 699572 485238
rect 699640 485182 699696 485238
rect 699764 485182 699820 485238
rect 699888 485182 699944 485238
rect 700012 485182 700068 485238
rect 700136 485182 700192 485238
rect 699392 485058 699448 485114
rect 699516 485058 699572 485114
rect 699640 485058 699696 485114
rect 699764 485058 699820 485114
rect 699888 485058 699944 485114
rect 700012 485058 700068 485114
rect 700136 485058 700192 485114
rect 699392 484934 699448 484990
rect 699516 484934 699572 484990
rect 699640 484934 699696 484990
rect 699764 484934 699820 484990
rect 699888 484934 699944 484990
rect 700012 484934 700068 484990
rect 700136 484934 700192 484990
rect 699392 484810 699448 484866
rect 699516 484810 699572 484866
rect 699640 484810 699696 484866
rect 699764 484810 699820 484866
rect 699888 484810 699944 484866
rect 700012 484810 700068 484866
rect 700136 484810 700192 484866
rect 707870 486676 707926 486732
rect 707870 486552 707926 486608
rect 707870 486428 707926 486484
rect 707870 486304 707926 486360
rect 707870 486180 707926 486236
rect 707870 486056 707926 486112
rect 707870 485932 707926 485988
rect 707870 485808 707926 485864
rect 707870 485684 707926 485740
rect 707870 485560 707926 485616
rect 707870 485436 707926 485492
rect 707870 485312 707926 485368
rect 707870 485188 707926 485244
rect 707870 485064 707926 485120
rect 707870 484940 707926 484996
rect 707870 484816 707926 484872
rect 699392 484066 699448 484122
rect 699516 484066 699572 484122
rect 699640 484066 699696 484122
rect 699764 484066 699820 484122
rect 699888 484066 699944 484122
rect 700012 484066 700068 484122
rect 700136 484066 700192 484122
rect 699392 483942 699448 483998
rect 699516 483942 699572 483998
rect 699640 483942 699696 483998
rect 699764 483942 699820 483998
rect 699888 483942 699944 483998
rect 700012 483942 700068 483998
rect 700136 483942 700192 483998
rect 699392 483818 699448 483874
rect 699516 483818 699572 483874
rect 699640 483818 699696 483874
rect 699764 483818 699820 483874
rect 699888 483818 699944 483874
rect 700012 483818 700068 483874
rect 700136 483818 700192 483874
rect 699392 483694 699448 483750
rect 699516 483694 699572 483750
rect 699640 483694 699696 483750
rect 699764 483694 699820 483750
rect 699888 483694 699944 483750
rect 700012 483694 700068 483750
rect 700136 483694 700192 483750
rect 699392 483570 699448 483626
rect 699516 483570 699572 483626
rect 699640 483570 699696 483626
rect 699764 483570 699820 483626
rect 699888 483570 699944 483626
rect 700012 483570 700068 483626
rect 700136 483570 700192 483626
rect 699392 483446 699448 483502
rect 699516 483446 699572 483502
rect 699640 483446 699696 483502
rect 699764 483446 699820 483502
rect 699888 483446 699944 483502
rect 700012 483446 700068 483502
rect 700136 483446 700192 483502
rect 699392 483322 699448 483378
rect 699516 483322 699572 483378
rect 699640 483322 699696 483378
rect 699764 483322 699820 483378
rect 699888 483322 699944 483378
rect 700012 483322 700068 483378
rect 700136 483322 700192 483378
rect 699392 483198 699448 483254
rect 699516 483198 699572 483254
rect 699640 483198 699696 483254
rect 699764 483198 699820 483254
rect 699888 483198 699944 483254
rect 700012 483198 700068 483254
rect 700136 483198 700192 483254
rect 699392 483074 699448 483130
rect 699516 483074 699572 483130
rect 699640 483074 699696 483130
rect 699764 483074 699820 483130
rect 699888 483074 699944 483130
rect 700012 483074 700068 483130
rect 700136 483074 700192 483130
rect 699392 482950 699448 483006
rect 699516 482950 699572 483006
rect 699640 482950 699696 483006
rect 699764 482950 699820 483006
rect 699888 482950 699944 483006
rect 700012 482950 700068 483006
rect 700136 482950 700192 483006
rect 699392 482826 699448 482882
rect 699516 482826 699572 482882
rect 699640 482826 699696 482882
rect 699764 482826 699820 482882
rect 699888 482826 699944 482882
rect 700012 482826 700068 482882
rect 700136 482826 700192 482882
rect 699392 482702 699448 482758
rect 699516 482702 699572 482758
rect 699640 482702 699696 482758
rect 699764 482702 699820 482758
rect 699888 482702 699944 482758
rect 700012 482702 700068 482758
rect 700136 482702 700192 482758
rect 699392 482578 699448 482634
rect 699516 482578 699572 482634
rect 699640 482578 699696 482634
rect 699764 482578 699820 482634
rect 699888 482578 699944 482634
rect 700012 482578 700068 482634
rect 700136 482578 700192 482634
rect 699392 482454 699448 482510
rect 699516 482454 699572 482510
rect 699640 482454 699696 482510
rect 699764 482454 699820 482510
rect 699888 482454 699944 482510
rect 700012 482454 700068 482510
rect 700136 482454 700192 482510
rect 699392 482330 699448 482386
rect 699516 482330 699572 482386
rect 699640 482330 699696 482386
rect 699764 482330 699820 482386
rect 699888 482330 699944 482386
rect 700012 482330 700068 482386
rect 700136 482330 700192 482386
rect 707870 484078 707926 484134
rect 707870 483954 707926 484010
rect 707870 483830 707926 483886
rect 707870 483706 707926 483762
rect 707870 483582 707926 483638
rect 707870 483458 707926 483514
rect 707870 483334 707926 483390
rect 707870 483210 707926 483266
rect 707870 483086 707926 483142
rect 707870 482962 707926 483018
rect 707870 482838 707926 482894
rect 707870 482714 707926 482770
rect 707870 482590 707926 482646
rect 707870 482466 707926 482522
rect 707870 482342 707926 482398
rect 707870 453602 707926 453658
rect 707870 453478 707926 453534
rect 707870 453354 707926 453410
rect 707870 453230 707926 453286
rect 707870 453106 707926 453162
rect 707870 452982 707926 453038
rect 707870 452858 707926 452914
rect 707870 452734 707926 452790
rect 707870 452610 707926 452666
rect 707870 452486 707926 452542
rect 707870 452362 707926 452418
rect 707870 452238 707926 452294
rect 707870 452114 707926 452170
rect 707870 451990 707926 452046
rect 707870 451866 707926 451922
rect 707870 451122 707926 451178
rect 707870 450998 707926 451054
rect 707870 450874 707926 450930
rect 707870 450750 707926 450806
rect 707870 450626 707926 450682
rect 707870 450502 707926 450558
rect 707870 450378 707926 450434
rect 707870 450254 707926 450310
rect 707870 450130 707926 450186
rect 707870 450006 707926 450062
rect 707870 449882 707926 449938
rect 707870 449758 707926 449814
rect 707870 449634 707926 449690
rect 707870 449510 707926 449566
rect 707870 449386 707926 449442
rect 707870 449262 707926 449318
rect 707870 448752 707926 448808
rect 707870 448628 707926 448684
rect 707870 448504 707926 448560
rect 707870 448380 707926 448436
rect 707870 448256 707926 448312
rect 707870 448132 707926 448188
rect 707870 448008 707926 448064
rect 707870 447884 707926 447940
rect 707870 447760 707926 447816
rect 707870 447636 707926 447692
rect 707870 447512 707926 447568
rect 707870 447388 707926 447444
rect 707870 447264 707926 447320
rect 707870 447140 707926 447196
rect 707870 447016 707926 447072
rect 707870 446892 707926 446948
rect 707870 446046 707926 446102
rect 707870 445922 707926 445978
rect 707870 445798 707926 445854
rect 707870 445674 707926 445730
rect 707870 445550 707926 445606
rect 707870 445426 707926 445482
rect 707870 445302 707926 445358
rect 707870 445178 707926 445234
rect 707870 445054 707926 445110
rect 707870 444930 707926 444986
rect 707870 444806 707926 444862
rect 707870 444682 707926 444738
rect 707870 444558 707926 444614
rect 707870 444434 707926 444490
rect 707870 444310 707926 444366
rect 707870 444186 707926 444242
rect 707870 443676 707926 443732
rect 707870 443552 707926 443608
rect 707870 443428 707926 443484
rect 707870 443304 707926 443360
rect 707870 443180 707926 443236
rect 707870 443056 707926 443112
rect 707870 442932 707926 442988
rect 707870 442808 707926 442864
rect 707870 442684 707926 442740
rect 707870 442560 707926 442616
rect 707870 442436 707926 442492
rect 707870 442312 707926 442368
rect 707870 442188 707926 442244
rect 707870 442064 707926 442120
rect 707870 441940 707926 441996
rect 707870 441816 707926 441872
rect 707870 441078 707926 441134
rect 707870 440954 707926 441010
rect 707870 440830 707926 440886
rect 707870 440706 707926 440762
rect 707870 440582 707926 440638
rect 707870 440458 707926 440514
rect 707870 440334 707926 440390
rect 707870 440210 707926 440266
rect 707870 440086 707926 440142
rect 707870 439962 707926 440018
rect 707870 439838 707926 439894
rect 707870 439714 707926 439770
rect 707870 439590 707926 439646
rect 707870 439466 707926 439522
rect 707870 439342 707926 439398
rect 707870 410602 707926 410658
rect 707870 410478 707926 410534
rect 707870 410354 707926 410410
rect 707870 410230 707926 410286
rect 707870 410106 707926 410162
rect 707870 409982 707926 410038
rect 707870 409858 707926 409914
rect 707870 409734 707926 409790
rect 707870 409610 707926 409666
rect 707870 409486 707926 409542
rect 707870 409362 707926 409418
rect 707870 409238 707926 409294
rect 707870 409114 707926 409170
rect 707870 408990 707926 409046
rect 707870 408866 707926 408922
rect 707870 408122 707926 408178
rect 707870 407998 707926 408054
rect 707870 407874 707926 407930
rect 707870 407750 707926 407806
rect 707870 407626 707926 407682
rect 707870 407502 707926 407558
rect 707870 407378 707926 407434
rect 707870 407254 707926 407310
rect 707870 407130 707926 407186
rect 707870 407006 707926 407062
rect 707870 406882 707926 406938
rect 707870 406758 707926 406814
rect 707870 406634 707926 406690
rect 707870 406510 707926 406566
rect 707870 406386 707926 406442
rect 707870 406262 707926 406318
rect 707870 405752 707926 405808
rect 707870 405628 707926 405684
rect 707870 405504 707926 405560
rect 707870 405380 707926 405436
rect 707870 405256 707926 405312
rect 707870 405132 707926 405188
rect 707870 405008 707926 405064
rect 707870 404884 707926 404940
rect 707870 404760 707926 404816
rect 707870 404636 707926 404692
rect 707870 404512 707926 404568
rect 707870 404388 707926 404444
rect 707870 404264 707926 404320
rect 707870 404140 707926 404196
rect 707870 404016 707926 404072
rect 707870 403892 707926 403948
rect 707870 403046 707926 403102
rect 707870 402922 707926 402978
rect 707870 402798 707926 402854
rect 707870 402674 707926 402730
rect 707870 402550 707926 402606
rect 707870 402426 707926 402482
rect 707870 402302 707926 402358
rect 707870 402178 707926 402234
rect 707870 402054 707926 402110
rect 707870 401930 707926 401986
rect 707870 401806 707926 401862
rect 707870 401682 707926 401738
rect 707870 401558 707926 401614
rect 707870 401434 707926 401490
rect 707870 401310 707926 401366
rect 707870 401186 707926 401242
rect 707870 400676 707926 400732
rect 707870 400552 707926 400608
rect 707870 400428 707926 400484
rect 707870 400304 707926 400360
rect 707870 400180 707926 400236
rect 707870 400056 707926 400112
rect 707870 399932 707926 399988
rect 707870 399808 707926 399864
rect 707870 399684 707926 399740
rect 707870 399560 707926 399616
rect 707870 399436 707926 399492
rect 707870 399312 707926 399368
rect 707870 399188 707926 399244
rect 707870 399064 707926 399120
rect 707870 398940 707926 398996
rect 707870 398816 707926 398872
rect 707870 398078 707926 398134
rect 707870 397954 707926 398010
rect 707870 397830 707926 397886
rect 707870 397706 707926 397762
rect 707870 397582 707926 397638
rect 707870 397458 707926 397514
rect 707870 397334 707926 397390
rect 707870 397210 707926 397266
rect 707870 397086 707926 397142
rect 707870 396962 707926 397018
rect 707870 396838 707926 396894
rect 707870 396714 707926 396770
rect 707870 396590 707926 396646
rect 707870 396466 707926 396522
rect 707870 396342 707926 396398
rect 699544 374373 699600 374429
rect 699844 374373 699900 374429
rect 700144 374373 700200 374429
rect 699544 374173 699600 374229
rect 699844 374173 699900 374229
rect 700144 374173 700200 374229
rect 699444 366898 699500 366954
rect 699744 366898 699800 366954
rect 700044 366898 700100 366954
rect 699444 359898 699500 359954
rect 699744 359898 699800 359954
rect 700044 359898 700100 359954
rect 699444 352898 699500 352954
rect 699744 352898 699800 352954
rect 700044 352898 700100 352954
rect 699544 338373 699600 338429
rect 699844 338373 699900 338429
rect 700144 338373 700200 338429
rect 699544 338173 699600 338229
rect 699844 338173 699900 338229
rect 700144 338173 700200 338229
rect 699497 333367 699553 333423
rect 699797 333367 699853 333423
rect 700097 333367 700153 333423
rect 699452 329584 699508 329640
rect 699576 329584 699632 329640
rect 699700 329584 699756 329640
rect 699824 329584 699880 329640
rect 699948 329584 700004 329640
rect 700072 329584 700128 329640
rect 700196 329584 700252 329640
rect 699452 329460 699508 329516
rect 699576 329460 699632 329516
rect 699700 329460 699756 329516
rect 699824 329460 699880 329516
rect 699948 329460 700004 329516
rect 700072 329460 700128 329516
rect 700196 329460 700252 329516
rect 699452 329336 699508 329392
rect 699576 329336 699632 329392
rect 699700 329336 699756 329392
rect 699824 329336 699880 329392
rect 699948 329336 700004 329392
rect 700072 329336 700128 329392
rect 700196 329336 700252 329392
rect 699452 329212 699508 329268
rect 699576 329212 699632 329268
rect 699700 329212 699756 329268
rect 699824 329212 699880 329268
rect 699948 329212 700004 329268
rect 700072 329212 700128 329268
rect 700196 329212 700252 329268
rect 699452 329088 699508 329144
rect 699576 329088 699632 329144
rect 699700 329088 699756 329144
rect 699824 329088 699880 329144
rect 699948 329088 700004 329144
rect 700072 329088 700128 329144
rect 700196 329088 700252 329144
rect 699452 328964 699508 329020
rect 699576 328964 699632 329020
rect 699700 328964 699756 329020
rect 699824 328964 699880 329020
rect 699948 328964 700004 329020
rect 700072 328964 700128 329020
rect 700196 328964 700252 329020
rect 699452 328840 699508 328896
rect 699576 328840 699632 328896
rect 699700 328840 699756 328896
rect 699824 328840 699880 328896
rect 699948 328840 700004 328896
rect 700072 328840 700128 328896
rect 700196 328840 700252 328896
rect 699444 323898 699500 323954
rect 699744 323898 699800 323954
rect 700044 323898 700100 323954
rect 699444 316898 699500 316954
rect 699744 316898 699800 316954
rect 700044 316898 700100 316954
rect 699444 309898 699500 309954
rect 699744 309898 699800 309954
rect 700044 309898 700100 309954
rect 699452 305730 699508 305786
rect 699576 305730 699632 305786
rect 699700 305730 699756 305786
rect 699824 305730 699880 305786
rect 699948 305730 700004 305786
rect 700072 305730 700128 305786
rect 700196 305730 700252 305786
rect 699452 305606 699508 305662
rect 699576 305606 699632 305662
rect 699700 305606 699756 305662
rect 699824 305606 699880 305662
rect 699948 305606 700004 305662
rect 700072 305606 700128 305662
rect 700196 305606 700252 305662
rect 699452 305482 699508 305538
rect 699576 305482 699632 305538
rect 699700 305482 699756 305538
rect 699824 305482 699880 305538
rect 699948 305482 700004 305538
rect 700072 305482 700128 305538
rect 700196 305482 700252 305538
rect 699452 305358 699508 305414
rect 699576 305358 699632 305414
rect 699700 305358 699756 305414
rect 699824 305358 699880 305414
rect 699948 305358 700004 305414
rect 700072 305358 700128 305414
rect 700196 305358 700252 305414
rect 699452 305234 699508 305290
rect 699576 305234 699632 305290
rect 699700 305234 699756 305290
rect 699824 305234 699880 305290
rect 699948 305234 700004 305290
rect 700072 305234 700128 305290
rect 700196 305234 700252 305290
rect 699452 305110 699508 305166
rect 699576 305110 699632 305166
rect 699700 305110 699756 305166
rect 699824 305110 699880 305166
rect 699948 305110 700004 305166
rect 700072 305110 700128 305166
rect 700196 305110 700252 305166
rect 699452 304986 699508 305042
rect 699576 304986 699632 305042
rect 699700 304986 699756 305042
rect 699824 304986 699880 305042
rect 699948 304986 700004 305042
rect 700072 304986 700128 305042
rect 700196 304986 700252 305042
rect 699497 290367 699553 290423
rect 699797 290367 699853 290423
rect 700097 290367 700153 290423
rect 699444 280898 699500 280954
rect 699744 280898 699800 280954
rect 700044 280898 700100 280954
rect 699444 273898 699500 273954
rect 699744 273898 699800 273954
rect 700044 273898 700100 273954
rect 699444 268551 699500 268607
rect 699744 268551 699800 268607
rect 700044 268551 700100 268607
rect 699444 266898 699500 266954
rect 699744 266898 699800 266954
rect 700044 266898 700100 266954
rect 699497 247367 699553 247423
rect 699797 247367 699853 247423
rect 700097 247367 700153 247423
rect 699444 237915 699500 237971
rect 699744 237915 699800 237971
rect 700044 237915 700100 237971
rect 699444 230898 699500 230954
rect 699744 230898 699800 230954
rect 700044 230898 700100 230954
rect 699444 223898 699500 223954
rect 699744 223898 699800 223954
rect 700044 223898 700100 223954
rect 699444 207279 699500 207335
rect 699744 207279 699800 207335
rect 700044 207279 700100 207335
rect 699497 204367 699553 204423
rect 699797 204367 699853 204423
rect 700097 204367 700153 204423
rect 699444 194898 699500 194954
rect 699744 194898 699800 194954
rect 700044 194898 700100 194954
rect 699444 187898 699500 187954
rect 699744 187898 699800 187954
rect 700044 187898 700100 187954
rect 699444 180898 699500 180954
rect 699744 180898 699800 180954
rect 700044 180898 700100 180954
rect 699444 176643 699500 176699
rect 699744 176643 699800 176699
rect 700044 176643 700100 176699
rect 699497 161367 699553 161423
rect 699797 161367 699853 161423
rect 700097 161367 700153 161423
rect 699444 151898 699500 151954
rect 699744 151898 699800 151954
rect 700044 151898 700100 151954
rect 699444 146007 699500 146063
rect 699744 146007 699800 146063
rect 700044 146007 700100 146063
rect 699444 144898 699500 144954
rect 699744 144898 699800 144954
rect 700044 144898 700100 144954
rect 699444 137898 699500 137954
rect 699744 137898 699800 137954
rect 700044 137898 700100 137954
rect 699444 133747 699500 133803
rect 699744 133747 699800 133803
rect 700044 133747 700100 133803
rect 699497 118367 699553 118423
rect 699797 118367 699853 118423
rect 700097 118367 700153 118423
rect 699444 108898 699500 108954
rect 699744 108898 699800 108954
rect 700044 108898 700100 108954
rect 699444 101898 699500 101954
rect 699744 101898 699800 101954
rect 700044 101898 700100 101954
rect 699444 94898 699500 94954
rect 699744 94898 699800 94954
rect 700044 94898 700100 94954
rect 699452 78552 699508 78608
rect 699576 78552 699632 78608
rect 699700 78552 699756 78608
rect 699824 78552 699880 78608
rect 699948 78552 700004 78608
rect 700072 78552 700128 78608
rect 700196 78552 700252 78608
rect 699452 78428 699508 78484
rect 699576 78428 699632 78484
rect 699700 78428 699756 78484
rect 699824 78428 699880 78484
rect 699948 78428 700004 78484
rect 700072 78428 700128 78484
rect 700196 78428 700252 78484
rect 699452 78304 699508 78360
rect 699576 78304 699632 78360
rect 699700 78304 699756 78360
rect 699824 78304 699880 78360
rect 699948 78304 700004 78360
rect 700072 78304 700128 78360
rect 700196 78304 700252 78360
rect 699452 78180 699508 78236
rect 699576 78180 699632 78236
rect 699700 78180 699756 78236
rect 699824 78180 699880 78236
rect 699948 78180 700004 78236
rect 700072 78180 700128 78236
rect 700196 78180 700252 78236
rect 699452 78056 699508 78112
rect 699576 78056 699632 78112
rect 699700 78056 699756 78112
rect 699824 78056 699880 78112
rect 699948 78056 700004 78112
rect 700072 78056 700128 78112
rect 700196 78056 700252 78112
rect 699452 77932 699508 77988
rect 699576 77932 699632 77988
rect 699700 77932 699756 77988
rect 699824 77932 699880 77988
rect 699948 77932 700004 77988
rect 700072 77932 700128 77988
rect 700196 77932 700252 77988
rect 699452 77808 699508 77864
rect 699576 77808 699632 77864
rect 699700 77808 699756 77864
rect 699824 77808 699880 77864
rect 699948 77808 700004 77864
rect 700072 77808 700128 77864
rect 700196 77808 700252 77864
rect 699497 75367 699553 75423
rect 699797 75367 699853 75423
rect 700097 75367 700153 75423
rect 698060 74952 698116 75008
rect 698360 74952 698416 75008
rect 698660 74952 698716 75008
<< metal5 >>
rect 76115 946048 80078 946110
rect 76115 945992 79284 946048
rect 79340 945992 79584 946048
rect 79640 945992 79884 946048
rect 79940 945992 80078 946048
rect 76115 945910 80078 945992
rect 76115 945510 76435 945910
rect 76915 945633 78678 945710
rect 76915 945577 77847 945633
rect 77903 945577 78147 945633
rect 78203 945577 78447 945633
rect 78503 945577 78678 945633
rect 76915 945510 78678 945577
rect 106924 942322 107244 944688
rect 110424 943435 110744 944624
rect 110424 943379 110548 943435
rect 110604 943379 110744 943435
rect 110424 943304 110744 943379
rect 113924 942322 114244 944688
rect 117424 943435 117744 944624
rect 117424 943379 117548 943435
rect 117604 943379 117744 943435
rect 117424 943304 117744 943379
rect 120924 942322 121244 944688
rect 124424 943435 124744 944624
rect 124424 943379 124548 943435
rect 124604 943379 124744 943435
rect 124424 943304 124744 943379
rect 161924 942322 162244 944688
rect 165424 943435 165744 944624
rect 165424 943379 165548 943435
rect 165604 943379 165744 943435
rect 165424 943304 165744 943379
rect 168924 942322 169244 944688
rect 172424 943435 172744 944624
rect 172424 943379 172548 943435
rect 172604 943379 172744 943435
rect 172424 943304 172744 943379
rect 175924 942322 176244 944688
rect 179424 943435 179744 944624
rect 179424 943379 179548 943435
rect 179604 943379 179744 943435
rect 179424 943304 179744 943379
rect 216924 942322 217244 944688
rect 220424 943435 220744 944624
rect 220424 943379 220548 943435
rect 220604 943379 220744 943435
rect 220424 943304 220744 943379
rect 223924 942322 224244 944688
rect 227424 943435 227744 944624
rect 227424 943379 227548 943435
rect 227604 943379 227744 943435
rect 227424 943304 227744 943379
rect 230924 942322 231244 944688
rect 234424 943435 234744 944624
rect 234424 943379 234548 943435
rect 234604 943379 234744 943435
rect 234424 943304 234744 943379
rect 271924 942322 272244 944688
rect 275424 943435 275744 944624
rect 275424 943379 275548 943435
rect 275604 943379 275744 943435
rect 275424 943304 275744 943379
rect 278924 942322 279244 944688
rect 282424 943435 282744 944624
rect 282424 943379 282548 943435
rect 282604 943379 282744 943435
rect 282424 943304 282744 943379
rect 285924 942322 286244 944688
rect 289424 943435 289744 944624
rect 289424 943379 289548 943435
rect 289604 943379 289744 943435
rect 289424 943304 289744 943379
rect 326924 942322 327244 944688
rect 330424 943435 330744 944624
rect 330424 943379 330548 943435
rect 330604 943379 330744 943435
rect 330424 943304 330744 943379
rect 333924 942322 334244 944688
rect 337424 943435 337744 944624
rect 337424 943379 337548 943435
rect 337604 943379 337744 943435
rect 337424 943304 337744 943379
rect 340924 942322 341244 944688
rect 344424 943435 344744 944624
rect 344424 943379 344548 943435
rect 344604 943379 344744 943435
rect 344424 943304 344744 943379
rect 436924 942322 437244 944688
rect 440424 943435 440744 944624
rect 440424 943379 440548 943435
rect 440604 943379 440744 943435
rect 440424 943304 440744 943379
rect 443924 942322 444244 944688
rect 447424 943435 447744 944624
rect 447424 943379 447548 943435
rect 447604 943379 447744 943435
rect 447424 943304 447744 943379
rect 450924 942322 451244 944688
rect 454424 943435 454744 944624
rect 454424 943379 454548 943435
rect 454604 943379 454744 943435
rect 454424 943304 454744 943379
rect 491924 942322 492244 944688
rect 495424 943435 495744 944624
rect 495424 943379 495548 943435
rect 495604 943379 495744 943435
rect 495424 943304 495744 943379
rect 498924 942322 499244 944688
rect 502424 943435 502744 944624
rect 502424 943379 502548 943435
rect 502604 943379 502744 943435
rect 502424 943304 502744 943379
rect 505924 942322 506244 944688
rect 509424 943435 509744 944624
rect 509424 943379 509548 943435
rect 509604 943379 509744 943435
rect 509424 943304 509744 943379
rect 546924 942322 547244 944688
rect 550424 943435 550744 944624
rect 550424 943379 550548 943435
rect 550604 943379 550744 943435
rect 550424 943304 550744 943379
rect 553924 942322 554244 944688
rect 557424 943435 557744 944624
rect 557424 943379 557548 943435
rect 557604 943379 557744 943435
rect 557424 943304 557744 943379
rect 560924 942322 561244 944688
rect 564424 943435 564744 944624
rect 564424 943379 564548 943435
rect 564604 943379 564744 943435
rect 564424 943304 564744 943379
rect 656924 942322 657244 944688
rect 660424 943435 660744 944624
rect 660424 943379 660548 943435
rect 660604 943379 660744 943435
rect 660424 943304 660744 943379
rect 663924 942322 664244 944688
rect 667424 943435 667744 944624
rect 667424 943379 667548 943435
rect 667604 943379 667744 943435
rect 667424 943304 667744 943379
rect 670924 942322 671244 944688
rect 674424 943435 674744 944624
rect 674424 943379 674548 943435
rect 674604 943379 674744 943435
rect 674424 943304 674744 943379
rect 77678 942252 700322 942322
rect 77678 942196 77748 942252
rect 77804 942196 77872 942252
rect 77928 942196 77996 942252
rect 78052 942196 78120 942252
rect 78176 942196 78244 942252
rect 78300 942196 78368 942252
rect 78424 942196 78492 942252
rect 78548 942200 700322 942252
rect 78548 942196 88207 942200
rect 77678 942144 88207 942196
rect 88263 942144 88407 942200
rect 88463 942153 160207 942200
rect 88463 942144 140406 942153
rect 77678 942128 140406 942144
rect 77678 942072 77748 942128
rect 77804 942072 77872 942128
rect 77928 942072 77996 942128
rect 78052 942072 78120 942128
rect 78176 942072 78244 942128
rect 78300 942072 78368 942128
rect 78424 942072 78492 942128
rect 78548 942097 140406 942128
rect 140462 942144 160207 942153
rect 160263 942144 160407 942200
rect 160463 942153 232207 942200
rect 160463 942144 195406 942153
rect 140462 942097 195406 942144
rect 195462 942144 232207 942153
rect 232263 942144 232407 942200
rect 232463 942153 268207 942200
rect 232463 942144 250406 942153
rect 195462 942097 250406 942144
rect 250462 942144 268207 942153
rect 268263 942144 268407 942200
rect 268463 942144 304207 942200
rect 304263 942144 304407 942200
rect 304463 942153 340207 942200
rect 304463 942144 305406 942153
rect 250462 942097 305406 942144
rect 305462 942144 340207 942153
rect 340263 942144 340407 942200
rect 340463 942153 376207 942200
rect 340463 942144 360406 942153
rect 305462 942097 360406 942144
rect 360462 942144 376207 942153
rect 376263 942144 376407 942200
rect 376463 942144 412207 942200
rect 412263 942144 412407 942200
rect 412463 942144 448207 942200
rect 448263 942144 448407 942200
rect 448463 942153 484207 942200
rect 448463 942144 470406 942153
rect 360462 942097 470406 942144
rect 470462 942144 484207 942153
rect 484263 942144 484407 942200
rect 484463 942144 520207 942200
rect 520263 942144 520407 942200
rect 520463 942153 556207 942200
rect 520463 942144 525406 942153
rect 470462 942097 525406 942144
rect 525462 942144 556207 942153
rect 556263 942144 556407 942200
rect 556463 942153 592207 942200
rect 556463 942144 580406 942153
rect 525462 942097 580406 942144
rect 580462 942144 592207 942153
rect 592263 942144 592407 942200
rect 592463 942144 628207 942200
rect 628263 942144 628407 942200
rect 628463 942144 664207 942200
rect 664263 942144 664407 942200
rect 664463 942192 700322 942200
rect 664463 942153 699452 942192
rect 664463 942144 690406 942153
rect 580462 942097 690406 942144
rect 690462 942136 699452 942153
rect 699508 942136 699576 942192
rect 699632 942136 699700 942192
rect 699756 942136 699824 942192
rect 699880 942136 699948 942192
rect 700004 942136 700072 942192
rect 700128 942136 700196 942192
rect 700252 942136 700322 942192
rect 690462 942097 700322 942136
rect 78548 942072 700322 942097
rect 77678 942068 700322 942072
rect 77678 942012 699452 942068
rect 699508 942012 699576 942068
rect 699632 942012 699700 942068
rect 699756 942012 699824 942068
rect 699880 942012 699948 942068
rect 700004 942012 700072 942068
rect 700128 942012 700196 942068
rect 700252 942012 700322 942068
rect 77678 942004 700322 942012
rect 77678 941948 77748 942004
rect 77804 941948 77872 942004
rect 77928 941948 77996 942004
rect 78052 941948 78120 942004
rect 78176 941948 78244 942004
rect 78300 941948 78368 942004
rect 78424 941948 78492 942004
rect 78548 941948 700322 942004
rect 77678 941944 700322 941948
rect 77678 941900 699452 941944
rect 77678 941880 88207 941900
rect 77678 941824 77748 941880
rect 77804 941824 77872 941880
rect 77928 941824 77996 941880
rect 78052 941824 78120 941880
rect 78176 941824 78244 941880
rect 78300 941824 78368 941880
rect 78424 941824 78492 941880
rect 78548 941844 88207 941880
rect 88263 941844 88407 941900
rect 88463 941853 160207 941900
rect 88463 941844 140406 941853
rect 78548 941824 140406 941844
rect 77678 941797 140406 941824
rect 140462 941844 160207 941853
rect 160263 941844 160407 941900
rect 160463 941853 232207 941900
rect 160463 941844 195406 941853
rect 140462 941797 195406 941844
rect 195462 941844 232207 941853
rect 232263 941844 232407 941900
rect 232463 941853 268207 941900
rect 232463 941844 250406 941853
rect 195462 941797 250406 941844
rect 250462 941844 268207 941853
rect 268263 941844 268407 941900
rect 268463 941844 304207 941900
rect 304263 941844 304407 941900
rect 304463 941853 340207 941900
rect 304463 941844 305406 941853
rect 250462 941797 305406 941844
rect 305462 941844 340207 941853
rect 340263 941844 340407 941900
rect 340463 941853 376207 941900
rect 340463 941844 360406 941853
rect 305462 941797 360406 941844
rect 360462 941844 376207 941853
rect 376263 941844 376407 941900
rect 376463 941844 412207 941900
rect 412263 941844 412407 941900
rect 412463 941844 448207 941900
rect 448263 941844 448407 941900
rect 448463 941853 484207 941900
rect 448463 941844 470406 941853
rect 360462 941797 470406 941844
rect 470462 941844 484207 941853
rect 484263 941844 484407 941900
rect 484463 941844 520207 941900
rect 520263 941844 520407 941900
rect 520463 941853 556207 941900
rect 520463 941844 525406 941853
rect 470462 941797 525406 941844
rect 525462 941844 556207 941853
rect 556263 941844 556407 941900
rect 556463 941853 592207 941900
rect 556463 941844 580406 941853
rect 525462 941797 580406 941844
rect 580462 941844 592207 941853
rect 592263 941844 592407 941900
rect 592463 941844 628207 941900
rect 628263 941844 628407 941900
rect 628463 941844 664207 941900
rect 664263 941844 664407 941900
rect 664463 941888 699452 941900
rect 699508 941888 699576 941944
rect 699632 941888 699700 941944
rect 699756 941888 699824 941944
rect 699880 941888 699948 941944
rect 700004 941888 700072 941944
rect 700128 941888 700196 941944
rect 700252 941888 700322 941944
rect 664463 941853 700322 941888
rect 664463 941844 690406 941853
rect 580462 941797 690406 941844
rect 690462 941820 700322 941853
rect 690462 941797 699452 941820
rect 77678 941764 699452 941797
rect 699508 941764 699576 941820
rect 699632 941764 699700 941820
rect 699756 941764 699824 941820
rect 699880 941764 699948 941820
rect 700004 941764 700072 941820
rect 700128 941764 700196 941820
rect 700252 941764 700322 941820
rect 77678 941756 700322 941764
rect 77678 941700 77748 941756
rect 77804 941700 77872 941756
rect 77928 941700 77996 941756
rect 78052 941700 78120 941756
rect 78176 941700 78244 941756
rect 78300 941700 78368 941756
rect 78424 941700 78492 941756
rect 78548 941700 700322 941756
rect 77678 941696 700322 941700
rect 77678 941640 699452 941696
rect 699508 941640 699576 941696
rect 699632 941640 699700 941696
rect 699756 941640 699824 941696
rect 699880 941640 699948 941696
rect 700004 941640 700072 941696
rect 700128 941640 700196 941696
rect 700252 941640 700322 941696
rect 77678 941632 700322 941640
rect 77678 941576 77748 941632
rect 77804 941576 77872 941632
rect 77928 941576 77996 941632
rect 78052 941576 78120 941632
rect 78176 941576 78244 941632
rect 78300 941576 78368 941632
rect 78424 941576 78492 941632
rect 78548 941600 700322 941632
rect 78548 941576 88207 941600
rect 77678 941544 88207 941576
rect 88263 941544 88407 941600
rect 88463 941553 160207 941600
rect 88463 941544 140406 941553
rect 77678 941508 140406 941544
rect 77678 941452 77748 941508
rect 77804 941452 77872 941508
rect 77928 941452 77996 941508
rect 78052 941452 78120 941508
rect 78176 941452 78244 941508
rect 78300 941452 78368 941508
rect 78424 941452 78492 941508
rect 78548 941497 140406 941508
rect 140462 941544 160207 941553
rect 160263 941544 160407 941600
rect 160463 941553 232207 941600
rect 160463 941544 195406 941553
rect 140462 941497 195406 941544
rect 195462 941544 232207 941553
rect 232263 941544 232407 941600
rect 232463 941553 268207 941600
rect 232463 941544 250406 941553
rect 195462 941497 250406 941544
rect 250462 941544 268207 941553
rect 268263 941544 268407 941600
rect 268463 941544 304207 941600
rect 304263 941544 304407 941600
rect 304463 941553 340207 941600
rect 304463 941544 305406 941553
rect 250462 941497 305406 941544
rect 305462 941544 340207 941553
rect 340263 941544 340407 941600
rect 340463 941553 376207 941600
rect 340463 941544 360406 941553
rect 305462 941497 360406 941544
rect 360462 941544 376207 941553
rect 376263 941544 376407 941600
rect 376463 941544 412207 941600
rect 412263 941544 412407 941600
rect 412463 941544 448207 941600
rect 448263 941544 448407 941600
rect 448463 941553 484207 941600
rect 448463 941544 470406 941553
rect 360462 941497 470406 941544
rect 470462 941544 484207 941553
rect 484263 941544 484407 941600
rect 484463 941544 520207 941600
rect 520263 941544 520407 941600
rect 520463 941553 556207 941600
rect 520463 941544 525406 941553
rect 470462 941497 525406 941544
rect 525462 941544 556207 941553
rect 556263 941544 556407 941600
rect 556463 941553 592207 941600
rect 556463 941544 580406 941553
rect 525462 941497 580406 941544
rect 580462 941544 592207 941553
rect 592263 941544 592407 941600
rect 592463 941544 628207 941600
rect 628263 941544 628407 941600
rect 628463 941544 664207 941600
rect 664263 941544 664407 941600
rect 664463 941572 700322 941600
rect 664463 941553 699452 941572
rect 664463 941544 690406 941553
rect 580462 941497 690406 941544
rect 690462 941516 699452 941553
rect 699508 941516 699576 941572
rect 699632 941516 699700 941572
rect 699756 941516 699824 941572
rect 699880 941516 699948 941572
rect 700004 941516 700072 941572
rect 700128 941516 700196 941572
rect 700252 941516 700322 941572
rect 690462 941497 700322 941516
rect 78548 941452 700322 941497
rect 77678 941448 700322 941452
rect 77678 941392 699452 941448
rect 699508 941392 699576 941448
rect 699632 941392 699700 941448
rect 699756 941392 699824 941448
rect 699880 941392 699948 941448
rect 700004 941392 700072 941448
rect 700128 941392 700196 941448
rect 700252 941392 700322 941448
rect 77678 941322 700322 941392
rect 79078 940852 698922 940922
rect 79078 940796 79148 940852
rect 79204 940796 79272 940852
rect 79328 940796 79396 940852
rect 79452 940796 79520 940852
rect 79576 940796 79644 940852
rect 79700 940796 79768 940852
rect 79824 940796 79892 940852
rect 79948 940800 698922 940852
rect 79948 940796 106207 940800
rect 79078 940744 106207 940796
rect 106263 940744 106407 940800
rect 106463 940744 142207 940800
rect 142263 940744 142407 940800
rect 142463 940744 178207 940800
rect 178263 940744 178407 940800
rect 178463 940744 214207 940800
rect 214263 940744 214407 940800
rect 214463 940744 250207 940800
rect 250263 940744 250407 940800
rect 250463 940744 286207 940800
rect 286263 940744 286407 940800
rect 286463 940744 322207 940800
rect 322263 940744 322407 940800
rect 322463 940744 358207 940800
rect 358263 940744 358407 940800
rect 358463 940792 430207 940800
rect 358463 940744 381348 940792
rect 79078 940736 381348 940744
rect 381404 940736 381472 940792
rect 381528 940736 381596 940792
rect 381652 940736 381720 940792
rect 381776 940736 381844 940792
rect 381900 940736 381968 940792
rect 382024 940736 382092 940792
rect 382148 940736 382216 940792
rect 382272 940736 382340 940792
rect 382396 940736 382464 940792
rect 382520 940736 382588 940792
rect 382644 940736 382712 940792
rect 382768 940736 382836 940792
rect 382892 940736 382960 940792
rect 383016 940736 383084 940792
rect 383140 940736 383828 940792
rect 383884 940736 383952 940792
rect 384008 940736 384076 940792
rect 384132 940736 384200 940792
rect 384256 940736 384324 940792
rect 384380 940736 384448 940792
rect 384504 940736 384572 940792
rect 384628 940736 384696 940792
rect 384752 940736 384820 940792
rect 384876 940736 384944 940792
rect 385000 940736 385068 940792
rect 385124 940736 385192 940792
rect 385248 940736 385316 940792
rect 385372 940736 385440 940792
rect 385496 940736 385564 940792
rect 385620 940736 385688 940792
rect 385744 940736 386198 940792
rect 386254 940736 386322 940792
rect 386378 940736 386446 940792
rect 386502 940736 386570 940792
rect 386626 940736 386694 940792
rect 386750 940736 386818 940792
rect 386874 940736 386942 940792
rect 386998 940736 387066 940792
rect 387122 940736 387190 940792
rect 387246 940736 387314 940792
rect 387370 940736 387438 940792
rect 387494 940736 387562 940792
rect 387618 940736 387686 940792
rect 387742 940736 387810 940792
rect 387866 940736 387934 940792
rect 387990 940736 388058 940792
rect 388114 940736 388904 940792
rect 388960 940736 389028 940792
rect 389084 940736 389152 940792
rect 389208 940736 389276 940792
rect 389332 940736 389400 940792
rect 389456 940736 389524 940792
rect 389580 940736 389648 940792
rect 389704 940736 389772 940792
rect 389828 940736 389896 940792
rect 389952 940736 390020 940792
rect 390076 940736 390144 940792
rect 390200 940736 390268 940792
rect 390324 940736 390392 940792
rect 390448 940736 390516 940792
rect 390572 940736 390640 940792
rect 390696 940736 390764 940792
rect 390820 940736 391274 940792
rect 391330 940736 391398 940792
rect 391454 940736 391522 940792
rect 391578 940736 391646 940792
rect 391702 940736 391770 940792
rect 391826 940736 391894 940792
rect 391950 940736 392018 940792
rect 392074 940736 392142 940792
rect 392198 940736 392266 940792
rect 392322 940736 392390 940792
rect 392446 940736 392514 940792
rect 392570 940736 392638 940792
rect 392694 940736 392762 940792
rect 392818 940736 392886 940792
rect 392942 940736 393010 940792
rect 393066 940736 393134 940792
rect 393190 940736 393878 940792
rect 393934 940736 394002 940792
rect 394058 940736 394126 940792
rect 394182 940736 394250 940792
rect 394306 940736 394374 940792
rect 394430 940736 394498 940792
rect 394554 940736 394622 940792
rect 394678 940736 394746 940792
rect 394802 940736 394870 940792
rect 394926 940736 394994 940792
rect 395050 940736 395118 940792
rect 395174 940736 395242 940792
rect 395298 940736 395366 940792
rect 395422 940736 395490 940792
rect 395546 940736 395614 940792
rect 395670 940744 430207 940792
rect 430263 940744 430407 940800
rect 430463 940744 466207 940800
rect 466263 940744 466407 940800
rect 466463 940744 502207 940800
rect 502263 940744 502407 940800
rect 502463 940744 538207 940800
rect 538263 940744 538407 940800
rect 538463 940744 574207 940800
rect 574263 940744 574407 940800
rect 574463 940792 646207 940800
rect 574463 940744 601348 940792
rect 395670 940736 601348 940744
rect 601404 940736 601472 940792
rect 601528 940736 601596 940792
rect 601652 940736 601720 940792
rect 601776 940736 601844 940792
rect 601900 940736 601968 940792
rect 602024 940736 602092 940792
rect 602148 940736 602216 940792
rect 602272 940736 602340 940792
rect 602396 940736 602464 940792
rect 602520 940736 602588 940792
rect 602644 940736 602712 940792
rect 602768 940736 602836 940792
rect 602892 940736 602960 940792
rect 603016 940736 603084 940792
rect 603140 940736 603828 940792
rect 603884 940736 603952 940792
rect 604008 940736 604076 940792
rect 604132 940736 604200 940792
rect 604256 940736 604324 940792
rect 604380 940736 604448 940792
rect 604504 940736 604572 940792
rect 604628 940736 604696 940792
rect 604752 940736 604820 940792
rect 604876 940736 604944 940792
rect 605000 940736 605068 940792
rect 605124 940736 605192 940792
rect 605248 940736 605316 940792
rect 605372 940736 605440 940792
rect 605496 940736 605564 940792
rect 605620 940736 605688 940792
rect 605744 940736 606198 940792
rect 606254 940736 606322 940792
rect 606378 940736 606446 940792
rect 606502 940736 606570 940792
rect 606626 940736 606694 940792
rect 606750 940736 606818 940792
rect 606874 940736 606942 940792
rect 606998 940736 607066 940792
rect 607122 940736 607190 940792
rect 607246 940736 607314 940792
rect 607370 940736 607438 940792
rect 607494 940736 607562 940792
rect 607618 940736 607686 940792
rect 607742 940736 607810 940792
rect 607866 940736 607934 940792
rect 607990 940736 608058 940792
rect 608114 940736 608904 940792
rect 608960 940736 609028 940792
rect 609084 940736 609152 940792
rect 609208 940736 609276 940792
rect 609332 940736 609400 940792
rect 609456 940736 609524 940792
rect 609580 940736 609648 940792
rect 609704 940736 609772 940792
rect 609828 940736 609896 940792
rect 609952 940736 610020 940792
rect 610076 940736 610144 940792
rect 610200 940736 610268 940792
rect 610324 940736 610392 940792
rect 610448 940736 610516 940792
rect 610572 940736 610640 940792
rect 610696 940736 610764 940792
rect 610820 940736 611274 940792
rect 611330 940736 611398 940792
rect 611454 940736 611522 940792
rect 611578 940736 611646 940792
rect 611702 940736 611770 940792
rect 611826 940736 611894 940792
rect 611950 940736 612018 940792
rect 612074 940736 612142 940792
rect 612198 940736 612266 940792
rect 612322 940736 612390 940792
rect 612446 940736 612514 940792
rect 612570 940736 612638 940792
rect 612694 940736 612762 940792
rect 612818 940736 612886 940792
rect 612942 940736 613010 940792
rect 613066 940736 613134 940792
rect 613190 940736 613878 940792
rect 613934 940736 614002 940792
rect 614058 940736 614126 940792
rect 614182 940736 614250 940792
rect 614306 940736 614374 940792
rect 614430 940736 614498 940792
rect 614554 940736 614622 940792
rect 614678 940736 614746 940792
rect 614802 940736 614870 940792
rect 614926 940736 614994 940792
rect 615050 940736 615118 940792
rect 615174 940736 615242 940792
rect 615298 940736 615366 940792
rect 615422 940736 615490 940792
rect 615546 940736 615614 940792
rect 615670 940744 646207 940792
rect 646263 940744 646407 940800
rect 646463 940744 682207 940800
rect 682263 940744 682407 940800
rect 682463 940792 698922 940800
rect 682463 940744 698052 940792
rect 615670 940736 698052 940744
rect 698108 940736 698176 940792
rect 698232 940736 698300 940792
rect 698356 940736 698424 940792
rect 698480 940736 698548 940792
rect 698604 940736 698672 940792
rect 698728 940736 698796 940792
rect 698852 940736 698922 940792
rect 79078 940728 698922 940736
rect 79078 940672 79148 940728
rect 79204 940672 79272 940728
rect 79328 940672 79396 940728
rect 79452 940672 79520 940728
rect 79576 940672 79644 940728
rect 79700 940672 79768 940728
rect 79824 940672 79892 940728
rect 79948 940716 698922 940728
rect 79948 940710 140821 940716
rect 79948 940672 110546 940710
rect 79078 940654 110546 940672
rect 110602 940654 117546 940710
rect 117602 940654 124546 940710
rect 124602 940660 140821 940710
rect 140877 940710 195821 940716
rect 140877 940660 165546 940710
rect 124602 940654 165546 940660
rect 165602 940654 172546 940710
rect 172602 940654 179546 940710
rect 179602 940660 195821 940710
rect 195877 940710 250821 940716
rect 195877 940660 220546 940710
rect 179602 940654 220546 940660
rect 220602 940654 227546 940710
rect 227602 940654 234546 940710
rect 234602 940660 250821 940710
rect 250877 940710 305821 940716
rect 250877 940660 275546 940710
rect 234602 940654 275546 940660
rect 275602 940654 282546 940710
rect 282602 940654 289546 940710
rect 289602 940660 305821 940710
rect 305877 940710 360821 940716
rect 305877 940660 330546 940710
rect 289602 940654 330546 940660
rect 330602 940654 337546 940710
rect 337602 940654 344546 940710
rect 344602 940660 360821 940710
rect 360877 940710 470821 940716
rect 360877 940668 440546 940710
rect 360877 940660 381348 940668
rect 344602 940654 381348 940660
rect 79078 940612 381348 940654
rect 381404 940612 381472 940668
rect 381528 940612 381596 940668
rect 381652 940612 381720 940668
rect 381776 940612 381844 940668
rect 381900 940612 381968 940668
rect 382024 940612 382092 940668
rect 382148 940612 382216 940668
rect 382272 940612 382340 940668
rect 382396 940612 382464 940668
rect 382520 940612 382588 940668
rect 382644 940612 382712 940668
rect 382768 940612 382836 940668
rect 382892 940612 382960 940668
rect 383016 940612 383084 940668
rect 383140 940612 383828 940668
rect 383884 940612 383952 940668
rect 384008 940612 384076 940668
rect 384132 940612 384200 940668
rect 384256 940612 384324 940668
rect 384380 940612 384448 940668
rect 384504 940612 384572 940668
rect 384628 940612 384696 940668
rect 384752 940612 384820 940668
rect 384876 940612 384944 940668
rect 385000 940612 385068 940668
rect 385124 940612 385192 940668
rect 385248 940612 385316 940668
rect 385372 940612 385440 940668
rect 385496 940612 385564 940668
rect 385620 940612 385688 940668
rect 385744 940612 386198 940668
rect 386254 940612 386322 940668
rect 386378 940612 386446 940668
rect 386502 940612 386570 940668
rect 386626 940612 386694 940668
rect 386750 940612 386818 940668
rect 386874 940612 386942 940668
rect 386998 940612 387066 940668
rect 387122 940612 387190 940668
rect 387246 940612 387314 940668
rect 387370 940612 387438 940668
rect 387494 940612 387562 940668
rect 387618 940612 387686 940668
rect 387742 940612 387810 940668
rect 387866 940612 387934 940668
rect 387990 940612 388058 940668
rect 388114 940612 388904 940668
rect 388960 940612 389028 940668
rect 389084 940612 389152 940668
rect 389208 940612 389276 940668
rect 389332 940612 389400 940668
rect 389456 940612 389524 940668
rect 389580 940612 389648 940668
rect 389704 940612 389772 940668
rect 389828 940612 389896 940668
rect 389952 940612 390020 940668
rect 390076 940612 390144 940668
rect 390200 940612 390268 940668
rect 390324 940612 390392 940668
rect 390448 940612 390516 940668
rect 390572 940612 390640 940668
rect 390696 940612 390764 940668
rect 390820 940612 391274 940668
rect 391330 940612 391398 940668
rect 391454 940612 391522 940668
rect 391578 940612 391646 940668
rect 391702 940612 391770 940668
rect 391826 940612 391894 940668
rect 391950 940612 392018 940668
rect 392074 940612 392142 940668
rect 392198 940612 392266 940668
rect 392322 940612 392390 940668
rect 392446 940612 392514 940668
rect 392570 940612 392638 940668
rect 392694 940612 392762 940668
rect 392818 940612 392886 940668
rect 392942 940612 393010 940668
rect 393066 940612 393134 940668
rect 393190 940612 393878 940668
rect 393934 940612 394002 940668
rect 394058 940612 394126 940668
rect 394182 940612 394250 940668
rect 394306 940612 394374 940668
rect 394430 940612 394498 940668
rect 394554 940612 394622 940668
rect 394678 940612 394746 940668
rect 394802 940612 394870 940668
rect 394926 940612 394994 940668
rect 395050 940612 395118 940668
rect 395174 940612 395242 940668
rect 395298 940612 395366 940668
rect 395422 940612 395490 940668
rect 395546 940612 395614 940668
rect 395670 940654 440546 940668
rect 440602 940654 447546 940710
rect 447602 940654 454546 940710
rect 454602 940660 470821 940710
rect 470877 940710 525821 940716
rect 470877 940660 495546 940710
rect 454602 940654 495546 940660
rect 495602 940654 502546 940710
rect 502602 940654 509546 940710
rect 509602 940660 525821 940710
rect 525877 940710 580821 940716
rect 525877 940660 550546 940710
rect 509602 940654 550546 940660
rect 550602 940654 557546 940710
rect 557602 940654 564546 940710
rect 564602 940660 580821 940710
rect 580877 940710 690821 940716
rect 580877 940668 660546 940710
rect 580877 940660 601348 940668
rect 564602 940654 601348 940660
rect 395670 940612 601348 940654
rect 601404 940612 601472 940668
rect 601528 940612 601596 940668
rect 601652 940612 601720 940668
rect 601776 940612 601844 940668
rect 601900 940612 601968 940668
rect 602024 940612 602092 940668
rect 602148 940612 602216 940668
rect 602272 940612 602340 940668
rect 602396 940612 602464 940668
rect 602520 940612 602588 940668
rect 602644 940612 602712 940668
rect 602768 940612 602836 940668
rect 602892 940612 602960 940668
rect 603016 940612 603084 940668
rect 603140 940612 603828 940668
rect 603884 940612 603952 940668
rect 604008 940612 604076 940668
rect 604132 940612 604200 940668
rect 604256 940612 604324 940668
rect 604380 940612 604448 940668
rect 604504 940612 604572 940668
rect 604628 940612 604696 940668
rect 604752 940612 604820 940668
rect 604876 940612 604944 940668
rect 605000 940612 605068 940668
rect 605124 940612 605192 940668
rect 605248 940612 605316 940668
rect 605372 940612 605440 940668
rect 605496 940612 605564 940668
rect 605620 940612 605688 940668
rect 605744 940612 606198 940668
rect 606254 940612 606322 940668
rect 606378 940612 606446 940668
rect 606502 940612 606570 940668
rect 606626 940612 606694 940668
rect 606750 940612 606818 940668
rect 606874 940612 606942 940668
rect 606998 940612 607066 940668
rect 607122 940612 607190 940668
rect 607246 940612 607314 940668
rect 607370 940612 607438 940668
rect 607494 940612 607562 940668
rect 607618 940612 607686 940668
rect 607742 940612 607810 940668
rect 607866 940612 607934 940668
rect 607990 940612 608058 940668
rect 608114 940612 608904 940668
rect 608960 940612 609028 940668
rect 609084 940612 609152 940668
rect 609208 940612 609276 940668
rect 609332 940612 609400 940668
rect 609456 940612 609524 940668
rect 609580 940612 609648 940668
rect 609704 940612 609772 940668
rect 609828 940612 609896 940668
rect 609952 940612 610020 940668
rect 610076 940612 610144 940668
rect 610200 940612 610268 940668
rect 610324 940612 610392 940668
rect 610448 940612 610516 940668
rect 610572 940612 610640 940668
rect 610696 940612 610764 940668
rect 610820 940612 611274 940668
rect 611330 940612 611398 940668
rect 611454 940612 611522 940668
rect 611578 940612 611646 940668
rect 611702 940612 611770 940668
rect 611826 940612 611894 940668
rect 611950 940612 612018 940668
rect 612074 940612 612142 940668
rect 612198 940612 612266 940668
rect 612322 940612 612390 940668
rect 612446 940612 612514 940668
rect 612570 940612 612638 940668
rect 612694 940612 612762 940668
rect 612818 940612 612886 940668
rect 612942 940612 613010 940668
rect 613066 940612 613134 940668
rect 613190 940612 613878 940668
rect 613934 940612 614002 940668
rect 614058 940612 614126 940668
rect 614182 940612 614250 940668
rect 614306 940612 614374 940668
rect 614430 940612 614498 940668
rect 614554 940612 614622 940668
rect 614678 940612 614746 940668
rect 614802 940612 614870 940668
rect 614926 940612 614994 940668
rect 615050 940612 615118 940668
rect 615174 940612 615242 940668
rect 615298 940612 615366 940668
rect 615422 940612 615490 940668
rect 615546 940612 615614 940668
rect 615670 940654 660546 940668
rect 660602 940654 667546 940710
rect 667602 940654 674546 940710
rect 674602 940660 690821 940710
rect 690877 940668 698922 940716
rect 690877 940660 698052 940668
rect 674602 940654 698052 940660
rect 615670 940612 698052 940654
rect 698108 940612 698176 940668
rect 698232 940612 698300 940668
rect 698356 940612 698424 940668
rect 698480 940612 698548 940668
rect 698604 940612 698672 940668
rect 698728 940612 698796 940668
rect 698852 940612 698922 940668
rect 79078 940604 698922 940612
rect 79078 940548 79148 940604
rect 79204 940548 79272 940604
rect 79328 940548 79396 940604
rect 79452 940548 79520 940604
rect 79576 940548 79644 940604
rect 79700 940548 79768 940604
rect 79824 940548 79892 940604
rect 79948 940548 698922 940604
rect 79078 940544 698922 940548
rect 79078 940500 381348 940544
rect 79078 940480 106207 940500
rect 79078 940424 79148 940480
rect 79204 940424 79272 940480
rect 79328 940424 79396 940480
rect 79452 940424 79520 940480
rect 79576 940424 79644 940480
rect 79700 940424 79768 940480
rect 79824 940424 79892 940480
rect 79948 940444 106207 940480
rect 106263 940444 106407 940500
rect 106463 940444 142207 940500
rect 142263 940444 142407 940500
rect 142463 940444 178207 940500
rect 178263 940444 178407 940500
rect 178463 940444 214207 940500
rect 214263 940444 214407 940500
rect 214463 940444 250207 940500
rect 250263 940444 250407 940500
rect 250463 940444 286207 940500
rect 286263 940444 286407 940500
rect 286463 940444 322207 940500
rect 322263 940444 322407 940500
rect 322463 940444 358207 940500
rect 358263 940444 358407 940500
rect 358463 940488 381348 940500
rect 381404 940488 381472 940544
rect 381528 940488 381596 940544
rect 381652 940488 381720 940544
rect 381776 940488 381844 940544
rect 381900 940488 381968 940544
rect 382024 940488 382092 940544
rect 382148 940488 382216 940544
rect 382272 940488 382340 940544
rect 382396 940488 382464 940544
rect 382520 940488 382588 940544
rect 382644 940488 382712 940544
rect 382768 940488 382836 940544
rect 382892 940488 382960 940544
rect 383016 940488 383084 940544
rect 383140 940488 383828 940544
rect 383884 940488 383952 940544
rect 384008 940488 384076 940544
rect 384132 940488 384200 940544
rect 384256 940488 384324 940544
rect 384380 940488 384448 940544
rect 384504 940488 384572 940544
rect 384628 940488 384696 940544
rect 384752 940488 384820 940544
rect 384876 940488 384944 940544
rect 385000 940488 385068 940544
rect 385124 940488 385192 940544
rect 385248 940488 385316 940544
rect 385372 940488 385440 940544
rect 385496 940488 385564 940544
rect 385620 940488 385688 940544
rect 385744 940488 386198 940544
rect 386254 940488 386322 940544
rect 386378 940488 386446 940544
rect 386502 940488 386570 940544
rect 386626 940488 386694 940544
rect 386750 940488 386818 940544
rect 386874 940488 386942 940544
rect 386998 940488 387066 940544
rect 387122 940488 387190 940544
rect 387246 940488 387314 940544
rect 387370 940488 387438 940544
rect 387494 940488 387562 940544
rect 387618 940488 387686 940544
rect 387742 940488 387810 940544
rect 387866 940488 387934 940544
rect 387990 940488 388058 940544
rect 388114 940488 388904 940544
rect 388960 940488 389028 940544
rect 389084 940488 389152 940544
rect 389208 940488 389276 940544
rect 389332 940488 389400 940544
rect 389456 940488 389524 940544
rect 389580 940488 389648 940544
rect 389704 940488 389772 940544
rect 389828 940488 389896 940544
rect 389952 940488 390020 940544
rect 390076 940488 390144 940544
rect 390200 940488 390268 940544
rect 390324 940488 390392 940544
rect 390448 940488 390516 940544
rect 390572 940488 390640 940544
rect 390696 940488 390764 940544
rect 390820 940488 391274 940544
rect 391330 940488 391398 940544
rect 391454 940488 391522 940544
rect 391578 940488 391646 940544
rect 391702 940488 391770 940544
rect 391826 940488 391894 940544
rect 391950 940488 392018 940544
rect 392074 940488 392142 940544
rect 392198 940488 392266 940544
rect 392322 940488 392390 940544
rect 392446 940488 392514 940544
rect 392570 940488 392638 940544
rect 392694 940488 392762 940544
rect 392818 940488 392886 940544
rect 392942 940488 393010 940544
rect 393066 940488 393134 940544
rect 393190 940488 393878 940544
rect 393934 940488 394002 940544
rect 394058 940488 394126 940544
rect 394182 940488 394250 940544
rect 394306 940488 394374 940544
rect 394430 940488 394498 940544
rect 394554 940488 394622 940544
rect 394678 940488 394746 940544
rect 394802 940488 394870 940544
rect 394926 940488 394994 940544
rect 395050 940488 395118 940544
rect 395174 940488 395242 940544
rect 395298 940488 395366 940544
rect 395422 940488 395490 940544
rect 395546 940488 395614 940544
rect 395670 940500 601348 940544
rect 395670 940488 430207 940500
rect 358463 940444 430207 940488
rect 430263 940444 430407 940500
rect 430463 940444 466207 940500
rect 466263 940444 466407 940500
rect 466463 940444 502207 940500
rect 502263 940444 502407 940500
rect 502463 940444 538207 940500
rect 538263 940444 538407 940500
rect 538463 940444 574207 940500
rect 574263 940444 574407 940500
rect 574463 940488 601348 940500
rect 601404 940488 601472 940544
rect 601528 940488 601596 940544
rect 601652 940488 601720 940544
rect 601776 940488 601844 940544
rect 601900 940488 601968 940544
rect 602024 940488 602092 940544
rect 602148 940488 602216 940544
rect 602272 940488 602340 940544
rect 602396 940488 602464 940544
rect 602520 940488 602588 940544
rect 602644 940488 602712 940544
rect 602768 940488 602836 940544
rect 602892 940488 602960 940544
rect 603016 940488 603084 940544
rect 603140 940488 603828 940544
rect 603884 940488 603952 940544
rect 604008 940488 604076 940544
rect 604132 940488 604200 940544
rect 604256 940488 604324 940544
rect 604380 940488 604448 940544
rect 604504 940488 604572 940544
rect 604628 940488 604696 940544
rect 604752 940488 604820 940544
rect 604876 940488 604944 940544
rect 605000 940488 605068 940544
rect 605124 940488 605192 940544
rect 605248 940488 605316 940544
rect 605372 940488 605440 940544
rect 605496 940488 605564 940544
rect 605620 940488 605688 940544
rect 605744 940488 606198 940544
rect 606254 940488 606322 940544
rect 606378 940488 606446 940544
rect 606502 940488 606570 940544
rect 606626 940488 606694 940544
rect 606750 940488 606818 940544
rect 606874 940488 606942 940544
rect 606998 940488 607066 940544
rect 607122 940488 607190 940544
rect 607246 940488 607314 940544
rect 607370 940488 607438 940544
rect 607494 940488 607562 940544
rect 607618 940488 607686 940544
rect 607742 940488 607810 940544
rect 607866 940488 607934 940544
rect 607990 940488 608058 940544
rect 608114 940488 608904 940544
rect 608960 940488 609028 940544
rect 609084 940488 609152 940544
rect 609208 940488 609276 940544
rect 609332 940488 609400 940544
rect 609456 940488 609524 940544
rect 609580 940488 609648 940544
rect 609704 940488 609772 940544
rect 609828 940488 609896 940544
rect 609952 940488 610020 940544
rect 610076 940488 610144 940544
rect 610200 940488 610268 940544
rect 610324 940488 610392 940544
rect 610448 940488 610516 940544
rect 610572 940488 610640 940544
rect 610696 940488 610764 940544
rect 610820 940488 611274 940544
rect 611330 940488 611398 940544
rect 611454 940488 611522 940544
rect 611578 940488 611646 940544
rect 611702 940488 611770 940544
rect 611826 940488 611894 940544
rect 611950 940488 612018 940544
rect 612074 940488 612142 940544
rect 612198 940488 612266 940544
rect 612322 940488 612390 940544
rect 612446 940488 612514 940544
rect 612570 940488 612638 940544
rect 612694 940488 612762 940544
rect 612818 940488 612886 940544
rect 612942 940488 613010 940544
rect 613066 940488 613134 940544
rect 613190 940488 613878 940544
rect 613934 940488 614002 940544
rect 614058 940488 614126 940544
rect 614182 940488 614250 940544
rect 614306 940488 614374 940544
rect 614430 940488 614498 940544
rect 614554 940488 614622 940544
rect 614678 940488 614746 940544
rect 614802 940488 614870 940544
rect 614926 940488 614994 940544
rect 615050 940488 615118 940544
rect 615174 940488 615242 940544
rect 615298 940488 615366 940544
rect 615422 940488 615490 940544
rect 615546 940488 615614 940544
rect 615670 940500 698052 940544
rect 615670 940488 646207 940500
rect 574463 940444 646207 940488
rect 646263 940444 646407 940500
rect 646463 940444 682207 940500
rect 682263 940444 682407 940500
rect 682463 940488 698052 940500
rect 698108 940488 698176 940544
rect 698232 940488 698300 940544
rect 698356 940488 698424 940544
rect 698480 940488 698548 940544
rect 698604 940488 698672 940544
rect 698728 940488 698796 940544
rect 698852 940488 698922 940544
rect 682463 940444 698922 940488
rect 79948 940424 698922 940444
rect 79078 940420 698922 940424
rect 79078 940416 381348 940420
rect 79078 940410 140821 940416
rect 79078 940356 110546 940410
rect 79078 940300 79148 940356
rect 79204 940300 79272 940356
rect 79328 940300 79396 940356
rect 79452 940300 79520 940356
rect 79576 940300 79644 940356
rect 79700 940300 79768 940356
rect 79824 940300 79892 940356
rect 79948 940354 110546 940356
rect 110602 940354 117546 940410
rect 117602 940354 124546 940410
rect 124602 940360 140821 940410
rect 140877 940410 195821 940416
rect 140877 940360 165546 940410
rect 124602 940354 165546 940360
rect 165602 940354 172546 940410
rect 172602 940354 179546 940410
rect 179602 940360 195821 940410
rect 195877 940410 250821 940416
rect 195877 940360 220546 940410
rect 179602 940354 220546 940360
rect 220602 940354 227546 940410
rect 227602 940354 234546 940410
rect 234602 940360 250821 940410
rect 250877 940410 305821 940416
rect 250877 940360 275546 940410
rect 234602 940354 275546 940360
rect 275602 940354 282546 940410
rect 282602 940354 289546 940410
rect 289602 940360 305821 940410
rect 305877 940410 360821 940416
rect 305877 940360 330546 940410
rect 289602 940354 330546 940360
rect 330602 940354 337546 940410
rect 337602 940354 344546 940410
rect 344602 940360 360821 940410
rect 360877 940364 381348 940416
rect 381404 940364 381472 940420
rect 381528 940364 381596 940420
rect 381652 940364 381720 940420
rect 381776 940364 381844 940420
rect 381900 940364 381968 940420
rect 382024 940364 382092 940420
rect 382148 940364 382216 940420
rect 382272 940364 382340 940420
rect 382396 940364 382464 940420
rect 382520 940364 382588 940420
rect 382644 940364 382712 940420
rect 382768 940364 382836 940420
rect 382892 940364 382960 940420
rect 383016 940364 383084 940420
rect 383140 940364 383828 940420
rect 383884 940364 383952 940420
rect 384008 940364 384076 940420
rect 384132 940364 384200 940420
rect 384256 940364 384324 940420
rect 384380 940364 384448 940420
rect 384504 940364 384572 940420
rect 384628 940364 384696 940420
rect 384752 940364 384820 940420
rect 384876 940364 384944 940420
rect 385000 940364 385068 940420
rect 385124 940364 385192 940420
rect 385248 940364 385316 940420
rect 385372 940364 385440 940420
rect 385496 940364 385564 940420
rect 385620 940364 385688 940420
rect 385744 940364 386198 940420
rect 386254 940364 386322 940420
rect 386378 940364 386446 940420
rect 386502 940364 386570 940420
rect 386626 940364 386694 940420
rect 386750 940364 386818 940420
rect 386874 940364 386942 940420
rect 386998 940364 387066 940420
rect 387122 940364 387190 940420
rect 387246 940364 387314 940420
rect 387370 940364 387438 940420
rect 387494 940364 387562 940420
rect 387618 940364 387686 940420
rect 387742 940364 387810 940420
rect 387866 940364 387934 940420
rect 387990 940364 388058 940420
rect 388114 940364 388904 940420
rect 388960 940364 389028 940420
rect 389084 940364 389152 940420
rect 389208 940364 389276 940420
rect 389332 940364 389400 940420
rect 389456 940364 389524 940420
rect 389580 940364 389648 940420
rect 389704 940364 389772 940420
rect 389828 940364 389896 940420
rect 389952 940364 390020 940420
rect 390076 940364 390144 940420
rect 390200 940364 390268 940420
rect 390324 940364 390392 940420
rect 390448 940364 390516 940420
rect 390572 940364 390640 940420
rect 390696 940364 390764 940420
rect 390820 940364 391274 940420
rect 391330 940364 391398 940420
rect 391454 940364 391522 940420
rect 391578 940364 391646 940420
rect 391702 940364 391770 940420
rect 391826 940364 391894 940420
rect 391950 940364 392018 940420
rect 392074 940364 392142 940420
rect 392198 940364 392266 940420
rect 392322 940364 392390 940420
rect 392446 940364 392514 940420
rect 392570 940364 392638 940420
rect 392694 940364 392762 940420
rect 392818 940364 392886 940420
rect 392942 940364 393010 940420
rect 393066 940364 393134 940420
rect 393190 940364 393878 940420
rect 393934 940364 394002 940420
rect 394058 940364 394126 940420
rect 394182 940364 394250 940420
rect 394306 940364 394374 940420
rect 394430 940364 394498 940420
rect 394554 940364 394622 940420
rect 394678 940364 394746 940420
rect 394802 940364 394870 940420
rect 394926 940364 394994 940420
rect 395050 940364 395118 940420
rect 395174 940364 395242 940420
rect 395298 940364 395366 940420
rect 395422 940364 395490 940420
rect 395546 940364 395614 940420
rect 395670 940416 601348 940420
rect 395670 940410 470821 940416
rect 395670 940364 440546 940410
rect 360877 940360 440546 940364
rect 344602 940354 440546 940360
rect 440602 940354 447546 940410
rect 447602 940354 454546 940410
rect 454602 940360 470821 940410
rect 470877 940410 525821 940416
rect 470877 940360 495546 940410
rect 454602 940354 495546 940360
rect 495602 940354 502546 940410
rect 502602 940354 509546 940410
rect 509602 940360 525821 940410
rect 525877 940410 580821 940416
rect 525877 940360 550546 940410
rect 509602 940354 550546 940360
rect 550602 940354 557546 940410
rect 557602 940354 564546 940410
rect 564602 940360 580821 940410
rect 580877 940364 601348 940416
rect 601404 940364 601472 940420
rect 601528 940364 601596 940420
rect 601652 940364 601720 940420
rect 601776 940364 601844 940420
rect 601900 940364 601968 940420
rect 602024 940364 602092 940420
rect 602148 940364 602216 940420
rect 602272 940364 602340 940420
rect 602396 940364 602464 940420
rect 602520 940364 602588 940420
rect 602644 940364 602712 940420
rect 602768 940364 602836 940420
rect 602892 940364 602960 940420
rect 603016 940364 603084 940420
rect 603140 940364 603828 940420
rect 603884 940364 603952 940420
rect 604008 940364 604076 940420
rect 604132 940364 604200 940420
rect 604256 940364 604324 940420
rect 604380 940364 604448 940420
rect 604504 940364 604572 940420
rect 604628 940364 604696 940420
rect 604752 940364 604820 940420
rect 604876 940364 604944 940420
rect 605000 940364 605068 940420
rect 605124 940364 605192 940420
rect 605248 940364 605316 940420
rect 605372 940364 605440 940420
rect 605496 940364 605564 940420
rect 605620 940364 605688 940420
rect 605744 940364 606198 940420
rect 606254 940364 606322 940420
rect 606378 940364 606446 940420
rect 606502 940364 606570 940420
rect 606626 940364 606694 940420
rect 606750 940364 606818 940420
rect 606874 940364 606942 940420
rect 606998 940364 607066 940420
rect 607122 940364 607190 940420
rect 607246 940364 607314 940420
rect 607370 940364 607438 940420
rect 607494 940364 607562 940420
rect 607618 940364 607686 940420
rect 607742 940364 607810 940420
rect 607866 940364 607934 940420
rect 607990 940364 608058 940420
rect 608114 940364 608904 940420
rect 608960 940364 609028 940420
rect 609084 940364 609152 940420
rect 609208 940364 609276 940420
rect 609332 940364 609400 940420
rect 609456 940364 609524 940420
rect 609580 940364 609648 940420
rect 609704 940364 609772 940420
rect 609828 940364 609896 940420
rect 609952 940364 610020 940420
rect 610076 940364 610144 940420
rect 610200 940364 610268 940420
rect 610324 940364 610392 940420
rect 610448 940364 610516 940420
rect 610572 940364 610640 940420
rect 610696 940364 610764 940420
rect 610820 940364 611274 940420
rect 611330 940364 611398 940420
rect 611454 940364 611522 940420
rect 611578 940364 611646 940420
rect 611702 940364 611770 940420
rect 611826 940364 611894 940420
rect 611950 940364 612018 940420
rect 612074 940364 612142 940420
rect 612198 940364 612266 940420
rect 612322 940364 612390 940420
rect 612446 940364 612514 940420
rect 612570 940364 612638 940420
rect 612694 940364 612762 940420
rect 612818 940364 612886 940420
rect 612942 940364 613010 940420
rect 613066 940364 613134 940420
rect 613190 940364 613878 940420
rect 613934 940364 614002 940420
rect 614058 940364 614126 940420
rect 614182 940364 614250 940420
rect 614306 940364 614374 940420
rect 614430 940364 614498 940420
rect 614554 940364 614622 940420
rect 614678 940364 614746 940420
rect 614802 940364 614870 940420
rect 614926 940364 614994 940420
rect 615050 940364 615118 940420
rect 615174 940364 615242 940420
rect 615298 940364 615366 940420
rect 615422 940364 615490 940420
rect 615546 940364 615614 940420
rect 615670 940416 698052 940420
rect 615670 940410 690821 940416
rect 615670 940364 660546 940410
rect 580877 940360 660546 940364
rect 564602 940354 660546 940360
rect 660602 940354 667546 940410
rect 667602 940354 674546 940410
rect 674602 940360 690821 940410
rect 690877 940364 698052 940416
rect 698108 940364 698176 940420
rect 698232 940364 698300 940420
rect 698356 940364 698424 940420
rect 698480 940364 698548 940420
rect 698604 940364 698672 940420
rect 698728 940364 698796 940420
rect 698852 940364 698922 940420
rect 690877 940360 698922 940364
rect 674602 940354 698922 940360
rect 79948 940300 698922 940354
rect 79078 940296 698922 940300
rect 79078 940240 381348 940296
rect 381404 940240 381472 940296
rect 381528 940240 381596 940296
rect 381652 940240 381720 940296
rect 381776 940240 381844 940296
rect 381900 940240 381968 940296
rect 382024 940240 382092 940296
rect 382148 940240 382216 940296
rect 382272 940240 382340 940296
rect 382396 940240 382464 940296
rect 382520 940240 382588 940296
rect 382644 940240 382712 940296
rect 382768 940240 382836 940296
rect 382892 940240 382960 940296
rect 383016 940240 383084 940296
rect 383140 940240 383828 940296
rect 383884 940240 383952 940296
rect 384008 940240 384076 940296
rect 384132 940240 384200 940296
rect 384256 940240 384324 940296
rect 384380 940240 384448 940296
rect 384504 940240 384572 940296
rect 384628 940240 384696 940296
rect 384752 940240 384820 940296
rect 384876 940240 384944 940296
rect 385000 940240 385068 940296
rect 385124 940240 385192 940296
rect 385248 940240 385316 940296
rect 385372 940240 385440 940296
rect 385496 940240 385564 940296
rect 385620 940240 385688 940296
rect 385744 940240 386198 940296
rect 386254 940240 386322 940296
rect 386378 940240 386446 940296
rect 386502 940240 386570 940296
rect 386626 940240 386694 940296
rect 386750 940240 386818 940296
rect 386874 940240 386942 940296
rect 386998 940240 387066 940296
rect 387122 940240 387190 940296
rect 387246 940240 387314 940296
rect 387370 940240 387438 940296
rect 387494 940240 387562 940296
rect 387618 940240 387686 940296
rect 387742 940240 387810 940296
rect 387866 940240 387934 940296
rect 387990 940240 388058 940296
rect 388114 940240 388904 940296
rect 388960 940240 389028 940296
rect 389084 940240 389152 940296
rect 389208 940240 389276 940296
rect 389332 940240 389400 940296
rect 389456 940240 389524 940296
rect 389580 940240 389648 940296
rect 389704 940240 389772 940296
rect 389828 940240 389896 940296
rect 389952 940240 390020 940296
rect 390076 940240 390144 940296
rect 390200 940240 390268 940296
rect 390324 940240 390392 940296
rect 390448 940240 390516 940296
rect 390572 940240 390640 940296
rect 390696 940240 390764 940296
rect 390820 940240 391274 940296
rect 391330 940240 391398 940296
rect 391454 940240 391522 940296
rect 391578 940240 391646 940296
rect 391702 940240 391770 940296
rect 391826 940240 391894 940296
rect 391950 940240 392018 940296
rect 392074 940240 392142 940296
rect 392198 940240 392266 940296
rect 392322 940240 392390 940296
rect 392446 940240 392514 940296
rect 392570 940240 392638 940296
rect 392694 940240 392762 940296
rect 392818 940240 392886 940296
rect 392942 940240 393010 940296
rect 393066 940240 393134 940296
rect 393190 940240 393878 940296
rect 393934 940240 394002 940296
rect 394058 940240 394126 940296
rect 394182 940240 394250 940296
rect 394306 940240 394374 940296
rect 394430 940240 394498 940296
rect 394554 940240 394622 940296
rect 394678 940240 394746 940296
rect 394802 940240 394870 940296
rect 394926 940240 394994 940296
rect 395050 940240 395118 940296
rect 395174 940240 395242 940296
rect 395298 940240 395366 940296
rect 395422 940240 395490 940296
rect 395546 940240 395614 940296
rect 395670 940240 601348 940296
rect 601404 940240 601472 940296
rect 601528 940240 601596 940296
rect 601652 940240 601720 940296
rect 601776 940240 601844 940296
rect 601900 940240 601968 940296
rect 602024 940240 602092 940296
rect 602148 940240 602216 940296
rect 602272 940240 602340 940296
rect 602396 940240 602464 940296
rect 602520 940240 602588 940296
rect 602644 940240 602712 940296
rect 602768 940240 602836 940296
rect 602892 940240 602960 940296
rect 603016 940240 603084 940296
rect 603140 940240 603828 940296
rect 603884 940240 603952 940296
rect 604008 940240 604076 940296
rect 604132 940240 604200 940296
rect 604256 940240 604324 940296
rect 604380 940240 604448 940296
rect 604504 940240 604572 940296
rect 604628 940240 604696 940296
rect 604752 940240 604820 940296
rect 604876 940240 604944 940296
rect 605000 940240 605068 940296
rect 605124 940240 605192 940296
rect 605248 940240 605316 940296
rect 605372 940240 605440 940296
rect 605496 940240 605564 940296
rect 605620 940240 605688 940296
rect 605744 940240 606198 940296
rect 606254 940240 606322 940296
rect 606378 940240 606446 940296
rect 606502 940240 606570 940296
rect 606626 940240 606694 940296
rect 606750 940240 606818 940296
rect 606874 940240 606942 940296
rect 606998 940240 607066 940296
rect 607122 940240 607190 940296
rect 607246 940240 607314 940296
rect 607370 940240 607438 940296
rect 607494 940240 607562 940296
rect 607618 940240 607686 940296
rect 607742 940240 607810 940296
rect 607866 940240 607934 940296
rect 607990 940240 608058 940296
rect 608114 940240 608904 940296
rect 608960 940240 609028 940296
rect 609084 940240 609152 940296
rect 609208 940240 609276 940296
rect 609332 940240 609400 940296
rect 609456 940240 609524 940296
rect 609580 940240 609648 940296
rect 609704 940240 609772 940296
rect 609828 940240 609896 940296
rect 609952 940240 610020 940296
rect 610076 940240 610144 940296
rect 610200 940240 610268 940296
rect 610324 940240 610392 940296
rect 610448 940240 610516 940296
rect 610572 940240 610640 940296
rect 610696 940240 610764 940296
rect 610820 940240 611274 940296
rect 611330 940240 611398 940296
rect 611454 940240 611522 940296
rect 611578 940240 611646 940296
rect 611702 940240 611770 940296
rect 611826 940240 611894 940296
rect 611950 940240 612018 940296
rect 612074 940240 612142 940296
rect 612198 940240 612266 940296
rect 612322 940240 612390 940296
rect 612446 940240 612514 940296
rect 612570 940240 612638 940296
rect 612694 940240 612762 940296
rect 612818 940240 612886 940296
rect 612942 940240 613010 940296
rect 613066 940240 613134 940296
rect 613190 940240 613878 940296
rect 613934 940240 614002 940296
rect 614058 940240 614126 940296
rect 614182 940240 614250 940296
rect 614306 940240 614374 940296
rect 614430 940240 614498 940296
rect 614554 940240 614622 940296
rect 614678 940240 614746 940296
rect 614802 940240 614870 940296
rect 614926 940240 614994 940296
rect 615050 940240 615118 940296
rect 615174 940240 615242 940296
rect 615298 940240 615366 940296
rect 615422 940240 615490 940296
rect 615546 940240 615614 940296
rect 615670 940240 698052 940296
rect 698108 940240 698176 940296
rect 698232 940240 698300 940296
rect 698356 940240 698424 940296
rect 698480 940240 698548 940296
rect 698604 940240 698672 940296
rect 698728 940240 698796 940296
rect 698852 940240 698922 940296
rect 79078 940232 698922 940240
rect 79078 940176 79148 940232
rect 79204 940176 79272 940232
rect 79328 940176 79396 940232
rect 79452 940176 79520 940232
rect 79576 940176 79644 940232
rect 79700 940176 79768 940232
rect 79824 940176 79892 940232
rect 79948 940200 698922 940232
rect 79948 940176 106207 940200
rect 79078 940144 106207 940176
rect 106263 940144 106407 940200
rect 106463 940144 142207 940200
rect 142263 940144 142407 940200
rect 142463 940144 178207 940200
rect 178263 940144 178407 940200
rect 178463 940144 214207 940200
rect 214263 940144 214407 940200
rect 214463 940144 250207 940200
rect 250263 940144 250407 940200
rect 250463 940144 286207 940200
rect 286263 940144 286407 940200
rect 286463 940144 322207 940200
rect 322263 940144 322407 940200
rect 322463 940144 358207 940200
rect 358263 940144 358407 940200
rect 358463 940172 430207 940200
rect 358463 940144 381348 940172
rect 79078 940116 381348 940144
rect 381404 940116 381472 940172
rect 381528 940116 381596 940172
rect 381652 940116 381720 940172
rect 381776 940116 381844 940172
rect 381900 940116 381968 940172
rect 382024 940116 382092 940172
rect 382148 940116 382216 940172
rect 382272 940116 382340 940172
rect 382396 940116 382464 940172
rect 382520 940116 382588 940172
rect 382644 940116 382712 940172
rect 382768 940116 382836 940172
rect 382892 940116 382960 940172
rect 383016 940116 383084 940172
rect 383140 940116 383828 940172
rect 383884 940116 383952 940172
rect 384008 940116 384076 940172
rect 384132 940116 384200 940172
rect 384256 940116 384324 940172
rect 384380 940116 384448 940172
rect 384504 940116 384572 940172
rect 384628 940116 384696 940172
rect 384752 940116 384820 940172
rect 384876 940116 384944 940172
rect 385000 940116 385068 940172
rect 385124 940116 385192 940172
rect 385248 940116 385316 940172
rect 385372 940116 385440 940172
rect 385496 940116 385564 940172
rect 385620 940116 385688 940172
rect 385744 940116 386198 940172
rect 386254 940116 386322 940172
rect 386378 940116 386446 940172
rect 386502 940116 386570 940172
rect 386626 940116 386694 940172
rect 386750 940116 386818 940172
rect 386874 940116 386942 940172
rect 386998 940116 387066 940172
rect 387122 940116 387190 940172
rect 387246 940116 387314 940172
rect 387370 940116 387438 940172
rect 387494 940116 387562 940172
rect 387618 940116 387686 940172
rect 387742 940116 387810 940172
rect 387866 940116 387934 940172
rect 387990 940116 388058 940172
rect 388114 940116 388904 940172
rect 388960 940116 389028 940172
rect 389084 940116 389152 940172
rect 389208 940116 389276 940172
rect 389332 940116 389400 940172
rect 389456 940116 389524 940172
rect 389580 940116 389648 940172
rect 389704 940116 389772 940172
rect 389828 940116 389896 940172
rect 389952 940116 390020 940172
rect 390076 940116 390144 940172
rect 390200 940116 390268 940172
rect 390324 940116 390392 940172
rect 390448 940116 390516 940172
rect 390572 940116 390640 940172
rect 390696 940116 390764 940172
rect 390820 940116 391274 940172
rect 391330 940116 391398 940172
rect 391454 940116 391522 940172
rect 391578 940116 391646 940172
rect 391702 940116 391770 940172
rect 391826 940116 391894 940172
rect 391950 940116 392018 940172
rect 392074 940116 392142 940172
rect 392198 940116 392266 940172
rect 392322 940116 392390 940172
rect 392446 940116 392514 940172
rect 392570 940116 392638 940172
rect 392694 940116 392762 940172
rect 392818 940116 392886 940172
rect 392942 940116 393010 940172
rect 393066 940116 393134 940172
rect 393190 940116 393878 940172
rect 393934 940116 394002 940172
rect 394058 940116 394126 940172
rect 394182 940116 394250 940172
rect 394306 940116 394374 940172
rect 394430 940116 394498 940172
rect 394554 940116 394622 940172
rect 394678 940116 394746 940172
rect 394802 940116 394870 940172
rect 394926 940116 394994 940172
rect 395050 940116 395118 940172
rect 395174 940116 395242 940172
rect 395298 940116 395366 940172
rect 395422 940116 395490 940172
rect 395546 940116 395614 940172
rect 395670 940144 430207 940172
rect 430263 940144 430407 940200
rect 430463 940144 466207 940200
rect 466263 940144 466407 940200
rect 466463 940144 502207 940200
rect 502263 940144 502407 940200
rect 502463 940144 538207 940200
rect 538263 940144 538407 940200
rect 538463 940144 574207 940200
rect 574263 940144 574407 940200
rect 574463 940172 646207 940200
rect 574463 940144 601348 940172
rect 395670 940116 601348 940144
rect 601404 940116 601472 940172
rect 601528 940116 601596 940172
rect 601652 940116 601720 940172
rect 601776 940116 601844 940172
rect 601900 940116 601968 940172
rect 602024 940116 602092 940172
rect 602148 940116 602216 940172
rect 602272 940116 602340 940172
rect 602396 940116 602464 940172
rect 602520 940116 602588 940172
rect 602644 940116 602712 940172
rect 602768 940116 602836 940172
rect 602892 940116 602960 940172
rect 603016 940116 603084 940172
rect 603140 940116 603828 940172
rect 603884 940116 603952 940172
rect 604008 940116 604076 940172
rect 604132 940116 604200 940172
rect 604256 940116 604324 940172
rect 604380 940116 604448 940172
rect 604504 940116 604572 940172
rect 604628 940116 604696 940172
rect 604752 940116 604820 940172
rect 604876 940116 604944 940172
rect 605000 940116 605068 940172
rect 605124 940116 605192 940172
rect 605248 940116 605316 940172
rect 605372 940116 605440 940172
rect 605496 940116 605564 940172
rect 605620 940116 605688 940172
rect 605744 940116 606198 940172
rect 606254 940116 606322 940172
rect 606378 940116 606446 940172
rect 606502 940116 606570 940172
rect 606626 940116 606694 940172
rect 606750 940116 606818 940172
rect 606874 940116 606942 940172
rect 606998 940116 607066 940172
rect 607122 940116 607190 940172
rect 607246 940116 607314 940172
rect 607370 940116 607438 940172
rect 607494 940116 607562 940172
rect 607618 940116 607686 940172
rect 607742 940116 607810 940172
rect 607866 940116 607934 940172
rect 607990 940116 608058 940172
rect 608114 940116 608904 940172
rect 608960 940116 609028 940172
rect 609084 940116 609152 940172
rect 609208 940116 609276 940172
rect 609332 940116 609400 940172
rect 609456 940116 609524 940172
rect 609580 940116 609648 940172
rect 609704 940116 609772 940172
rect 609828 940116 609896 940172
rect 609952 940116 610020 940172
rect 610076 940116 610144 940172
rect 610200 940116 610268 940172
rect 610324 940116 610392 940172
rect 610448 940116 610516 940172
rect 610572 940116 610640 940172
rect 610696 940116 610764 940172
rect 610820 940116 611274 940172
rect 611330 940116 611398 940172
rect 611454 940116 611522 940172
rect 611578 940116 611646 940172
rect 611702 940116 611770 940172
rect 611826 940116 611894 940172
rect 611950 940116 612018 940172
rect 612074 940116 612142 940172
rect 612198 940116 612266 940172
rect 612322 940116 612390 940172
rect 612446 940116 612514 940172
rect 612570 940116 612638 940172
rect 612694 940116 612762 940172
rect 612818 940116 612886 940172
rect 612942 940116 613010 940172
rect 613066 940116 613134 940172
rect 613190 940116 613878 940172
rect 613934 940116 614002 940172
rect 614058 940116 614126 940172
rect 614182 940116 614250 940172
rect 614306 940116 614374 940172
rect 614430 940116 614498 940172
rect 614554 940116 614622 940172
rect 614678 940116 614746 940172
rect 614802 940116 614870 940172
rect 614926 940116 614994 940172
rect 615050 940116 615118 940172
rect 615174 940116 615242 940172
rect 615298 940116 615366 940172
rect 615422 940116 615490 940172
rect 615546 940116 615614 940172
rect 615670 940144 646207 940172
rect 646263 940144 646407 940200
rect 646463 940144 682207 940200
rect 682263 940144 682407 940200
rect 682463 940172 698922 940200
rect 682463 940144 698052 940172
rect 615670 940116 698052 940144
rect 698108 940116 698176 940172
rect 698232 940116 698300 940172
rect 698356 940116 698424 940172
rect 698480 940116 698548 940172
rect 698604 940116 698672 940172
rect 698728 940116 698796 940172
rect 698852 940116 698922 940172
rect 79078 940110 140821 940116
rect 79078 940108 110546 940110
rect 79078 940052 79148 940108
rect 79204 940052 79272 940108
rect 79328 940052 79396 940108
rect 79452 940052 79520 940108
rect 79576 940052 79644 940108
rect 79700 940052 79768 940108
rect 79824 940052 79892 940108
rect 79948 940054 110546 940108
rect 110602 940054 117546 940110
rect 117602 940054 124546 940110
rect 124602 940060 140821 940110
rect 140877 940110 195821 940116
rect 140877 940060 165546 940110
rect 124602 940054 165546 940060
rect 165602 940054 172546 940110
rect 172602 940054 179546 940110
rect 179602 940060 195821 940110
rect 195877 940110 250821 940116
rect 195877 940060 220546 940110
rect 179602 940054 220546 940060
rect 220602 940054 227546 940110
rect 227602 940054 234546 940110
rect 234602 940060 250821 940110
rect 250877 940110 305821 940116
rect 250877 940060 275546 940110
rect 234602 940054 275546 940060
rect 275602 940054 282546 940110
rect 282602 940054 289546 940110
rect 289602 940060 305821 940110
rect 305877 940110 360821 940116
rect 305877 940060 330546 940110
rect 289602 940054 330546 940060
rect 330602 940054 337546 940110
rect 337602 940054 344546 940110
rect 344602 940060 360821 940110
rect 360877 940110 470821 940116
rect 360877 940060 440546 940110
rect 344602 940054 440546 940060
rect 440602 940054 447546 940110
rect 447602 940054 454546 940110
rect 454602 940060 470821 940110
rect 470877 940110 525821 940116
rect 470877 940060 495546 940110
rect 454602 940054 495546 940060
rect 495602 940054 502546 940110
rect 502602 940054 509546 940110
rect 509602 940060 525821 940110
rect 525877 940110 580821 940116
rect 525877 940060 550546 940110
rect 509602 940054 550546 940060
rect 550602 940054 557546 940110
rect 557602 940054 564546 940110
rect 564602 940060 580821 940110
rect 580877 940110 690821 940116
rect 580877 940060 660546 940110
rect 564602 940054 660546 940060
rect 660602 940054 667546 940110
rect 667602 940054 674546 940110
rect 674602 940060 690821 940110
rect 690877 940060 698922 940116
rect 674602 940054 698922 940060
rect 79948 940052 698922 940054
rect 79078 940048 698922 940052
rect 79078 939992 381348 940048
rect 381404 939992 381472 940048
rect 381528 939992 381596 940048
rect 381652 939992 381720 940048
rect 381776 939992 381844 940048
rect 381900 939992 381968 940048
rect 382024 939992 382092 940048
rect 382148 939992 382216 940048
rect 382272 939992 382340 940048
rect 382396 939992 382464 940048
rect 382520 939992 382588 940048
rect 382644 939992 382712 940048
rect 382768 939992 382836 940048
rect 382892 939992 382960 940048
rect 383016 939992 383084 940048
rect 383140 939992 383828 940048
rect 383884 939992 383952 940048
rect 384008 939992 384076 940048
rect 384132 939992 384200 940048
rect 384256 939992 384324 940048
rect 384380 939992 384448 940048
rect 384504 939992 384572 940048
rect 384628 939992 384696 940048
rect 384752 939992 384820 940048
rect 384876 939992 384944 940048
rect 385000 939992 385068 940048
rect 385124 939992 385192 940048
rect 385248 939992 385316 940048
rect 385372 939992 385440 940048
rect 385496 939992 385564 940048
rect 385620 939992 385688 940048
rect 385744 939992 386198 940048
rect 386254 939992 386322 940048
rect 386378 939992 386446 940048
rect 386502 939992 386570 940048
rect 386626 939992 386694 940048
rect 386750 939992 386818 940048
rect 386874 939992 386942 940048
rect 386998 939992 387066 940048
rect 387122 939992 387190 940048
rect 387246 939992 387314 940048
rect 387370 939992 387438 940048
rect 387494 939992 387562 940048
rect 387618 939992 387686 940048
rect 387742 939992 387810 940048
rect 387866 939992 387934 940048
rect 387990 939992 388058 940048
rect 388114 939992 388904 940048
rect 388960 939992 389028 940048
rect 389084 939992 389152 940048
rect 389208 939992 389276 940048
rect 389332 939992 389400 940048
rect 389456 939992 389524 940048
rect 389580 939992 389648 940048
rect 389704 939992 389772 940048
rect 389828 939992 389896 940048
rect 389952 939992 390020 940048
rect 390076 939992 390144 940048
rect 390200 939992 390268 940048
rect 390324 939992 390392 940048
rect 390448 939992 390516 940048
rect 390572 939992 390640 940048
rect 390696 939992 390764 940048
rect 390820 939992 391274 940048
rect 391330 939992 391398 940048
rect 391454 939992 391522 940048
rect 391578 939992 391646 940048
rect 391702 939992 391770 940048
rect 391826 939992 391894 940048
rect 391950 939992 392018 940048
rect 392074 939992 392142 940048
rect 392198 939992 392266 940048
rect 392322 939992 392390 940048
rect 392446 939992 392514 940048
rect 392570 939992 392638 940048
rect 392694 939992 392762 940048
rect 392818 939992 392886 940048
rect 392942 939992 393010 940048
rect 393066 939992 393134 940048
rect 393190 939992 393878 940048
rect 393934 939992 394002 940048
rect 394058 939992 394126 940048
rect 394182 939992 394250 940048
rect 394306 939992 394374 940048
rect 394430 939992 394498 940048
rect 394554 939992 394622 940048
rect 394678 939992 394746 940048
rect 394802 939992 394870 940048
rect 394926 939992 394994 940048
rect 395050 939992 395118 940048
rect 395174 939992 395242 940048
rect 395298 939992 395366 940048
rect 395422 939992 395490 940048
rect 395546 939992 395614 940048
rect 395670 939992 601348 940048
rect 601404 939992 601472 940048
rect 601528 939992 601596 940048
rect 601652 939992 601720 940048
rect 601776 939992 601844 940048
rect 601900 939992 601968 940048
rect 602024 939992 602092 940048
rect 602148 939992 602216 940048
rect 602272 939992 602340 940048
rect 602396 939992 602464 940048
rect 602520 939992 602588 940048
rect 602644 939992 602712 940048
rect 602768 939992 602836 940048
rect 602892 939992 602960 940048
rect 603016 939992 603084 940048
rect 603140 939992 603828 940048
rect 603884 939992 603952 940048
rect 604008 939992 604076 940048
rect 604132 939992 604200 940048
rect 604256 939992 604324 940048
rect 604380 939992 604448 940048
rect 604504 939992 604572 940048
rect 604628 939992 604696 940048
rect 604752 939992 604820 940048
rect 604876 939992 604944 940048
rect 605000 939992 605068 940048
rect 605124 939992 605192 940048
rect 605248 939992 605316 940048
rect 605372 939992 605440 940048
rect 605496 939992 605564 940048
rect 605620 939992 605688 940048
rect 605744 939992 606198 940048
rect 606254 939992 606322 940048
rect 606378 939992 606446 940048
rect 606502 939992 606570 940048
rect 606626 939992 606694 940048
rect 606750 939992 606818 940048
rect 606874 939992 606942 940048
rect 606998 939992 607066 940048
rect 607122 939992 607190 940048
rect 607246 939992 607314 940048
rect 607370 939992 607438 940048
rect 607494 939992 607562 940048
rect 607618 939992 607686 940048
rect 607742 939992 607810 940048
rect 607866 939992 607934 940048
rect 607990 939992 608058 940048
rect 608114 939992 608904 940048
rect 608960 939992 609028 940048
rect 609084 939992 609152 940048
rect 609208 939992 609276 940048
rect 609332 939992 609400 940048
rect 609456 939992 609524 940048
rect 609580 939992 609648 940048
rect 609704 939992 609772 940048
rect 609828 939992 609896 940048
rect 609952 939992 610020 940048
rect 610076 939992 610144 940048
rect 610200 939992 610268 940048
rect 610324 939992 610392 940048
rect 610448 939992 610516 940048
rect 610572 939992 610640 940048
rect 610696 939992 610764 940048
rect 610820 939992 611274 940048
rect 611330 939992 611398 940048
rect 611454 939992 611522 940048
rect 611578 939992 611646 940048
rect 611702 939992 611770 940048
rect 611826 939992 611894 940048
rect 611950 939992 612018 940048
rect 612074 939992 612142 940048
rect 612198 939992 612266 940048
rect 612322 939992 612390 940048
rect 612446 939992 612514 940048
rect 612570 939992 612638 940048
rect 612694 939992 612762 940048
rect 612818 939992 612886 940048
rect 612942 939992 613010 940048
rect 613066 939992 613134 940048
rect 613190 939992 613878 940048
rect 613934 939992 614002 940048
rect 614058 939992 614126 940048
rect 614182 939992 614250 940048
rect 614306 939992 614374 940048
rect 614430 939992 614498 940048
rect 614554 939992 614622 940048
rect 614678 939992 614746 940048
rect 614802 939992 614870 940048
rect 614926 939992 614994 940048
rect 615050 939992 615118 940048
rect 615174 939992 615242 940048
rect 615298 939992 615366 940048
rect 615422 939992 615490 940048
rect 615546 939992 615614 940048
rect 615670 939992 698052 940048
rect 698108 939992 698176 940048
rect 698232 939992 698300 940048
rect 698356 939992 698424 940048
rect 698480 939992 698548 940048
rect 698604 939992 698672 940048
rect 698728 939992 698796 940048
rect 698852 939992 698922 940048
rect 79078 939922 698922 939992
rect 75376 929622 80078 929744
rect 75376 929566 79300 929622
rect 79356 929566 79600 929622
rect 79656 929566 79900 929622
rect 79956 929566 80078 929622
rect 75376 929424 80078 929566
rect 75312 926102 78678 926244
rect 75312 926046 77900 926102
rect 77956 926046 78200 926102
rect 78256 926046 78500 926102
rect 78556 926046 78678 926102
rect 75312 925924 78678 926046
rect 699322 925954 702688 926076
rect 699322 925898 699444 925954
rect 699500 925898 699744 925954
rect 699800 925898 700044 925954
rect 700100 925898 702688 925954
rect 699322 925756 702688 925898
rect 75376 922622 80078 922744
rect 75376 922566 79300 922622
rect 79356 922566 79600 922622
rect 79656 922566 79900 922622
rect 79956 922566 80078 922622
rect 75376 922424 80078 922566
rect 697922 922434 702624 922576
rect 697922 922378 698044 922434
rect 698100 922378 698344 922434
rect 698400 922378 698644 922434
rect 698700 922378 702624 922434
rect 697922 922256 702624 922378
rect 75312 919102 78678 919244
rect 75312 919046 77900 919102
rect 77956 919046 78200 919102
rect 78256 919046 78500 919102
rect 78556 919046 78678 919102
rect 75312 918924 78678 919046
rect 699322 918954 702688 919076
rect 699322 918898 699444 918954
rect 699500 918898 699744 918954
rect 699800 918898 700044 918954
rect 700100 918898 702688 918954
rect 699322 918756 702688 918898
rect 75376 915622 80078 915744
rect 75376 915566 79300 915622
rect 79356 915566 79600 915622
rect 79656 915566 79900 915622
rect 79956 915566 80078 915622
rect 75376 915424 80078 915566
rect 697922 915434 702624 915576
rect 697922 915378 698044 915434
rect 698100 915378 698344 915434
rect 698400 915378 698644 915434
rect 698700 915378 702624 915434
rect 697922 915256 702624 915378
rect 77678 914429 84516 914630
rect 77678 914373 77800 914429
rect 77856 914373 78100 914429
rect 78156 914373 78400 914429
rect 78456 914373 84516 914429
rect 77678 914229 84516 914373
rect 77678 914173 77800 914229
rect 77856 914173 78100 914229
rect 78156 914173 78400 914229
rect 78456 914173 84516 914229
rect 77678 914010 84516 914173
rect 687412 914429 700322 914630
rect 687412 914373 699544 914429
rect 699600 914373 699844 914429
rect 699900 914373 700144 914429
rect 700200 914373 700322 914429
rect 687412 914229 700322 914373
rect 687412 914173 699544 914229
rect 699600 914173 699844 914229
rect 699900 914173 700144 914229
rect 700200 914173 700322 914229
rect 687412 914010 700322 914173
rect 75312 912102 78678 912244
rect 75312 912046 77900 912102
rect 77956 912046 78200 912102
rect 78256 912046 78500 912102
rect 78556 912046 78678 912102
rect 75312 911924 78678 912046
rect 699322 911954 702688 912076
rect 699322 911898 699444 911954
rect 699500 911898 699744 911954
rect 699800 911898 700044 911954
rect 700100 911898 702688 911954
rect 699322 911756 702688 911898
rect 697922 908434 702624 908576
rect 697922 908378 698044 908434
rect 698100 908378 698344 908434
rect 698400 908378 698644 908434
rect 698700 908378 702624 908434
rect 697922 908256 702624 908378
rect 79078 896429 83556 896630
rect 79078 896373 79200 896429
rect 79256 896373 79500 896429
rect 79556 896373 79800 896429
rect 79856 896373 83556 896429
rect 79078 896229 83556 896373
rect 79078 896173 79200 896229
rect 79256 896173 79500 896229
rect 79556 896173 79800 896229
rect 79856 896173 83556 896229
rect 79078 896010 83556 896173
rect 688372 896429 698922 896630
rect 688372 896373 698144 896429
rect 698200 896373 698444 896429
rect 698500 896373 698744 896429
rect 698800 896373 698922 896429
rect 688372 896229 698922 896373
rect 688372 896173 698144 896229
rect 698200 896173 698444 896229
rect 698500 896173 698744 896229
rect 698800 896173 698922 896229
rect 688372 896010 698922 896173
rect 699322 892423 701085 892490
rect 699322 892367 699497 892423
rect 699553 892367 699797 892423
rect 699853 892367 700097 892423
rect 700153 892367 701085 892423
rect 699322 892290 701085 892367
rect 701565 892090 701885 892490
rect 697922 892008 701885 892090
rect 697922 891952 698060 892008
rect 698116 891952 698360 892008
rect 698416 891952 698660 892008
rect 698716 891952 701885 892008
rect 697922 891890 701885 891952
rect 70000 884670 78678 884728
rect 70000 884658 77808 884670
rect 70000 884602 70074 884658
rect 70130 884614 77808 884658
rect 77864 884614 77932 884670
rect 77988 884614 78056 884670
rect 78112 884614 78180 884670
rect 78236 884614 78304 884670
rect 78360 884614 78428 884670
rect 78484 884614 78552 884670
rect 78608 884614 78678 884670
rect 70130 884602 78678 884614
rect 70000 884546 78678 884602
rect 70000 884534 77808 884546
rect 70000 884478 70074 884534
rect 70130 884490 77808 884534
rect 77864 884490 77932 884546
rect 77988 884490 78056 884546
rect 78112 884490 78180 884546
rect 78236 884490 78304 884546
rect 78360 884490 78428 884546
rect 78484 884490 78552 884546
rect 78608 884490 78678 884546
rect 70130 884478 78678 884490
rect 70000 884422 78678 884478
rect 70000 884410 77808 884422
rect 70000 884354 70074 884410
rect 70130 884366 77808 884410
rect 77864 884366 77932 884422
rect 77988 884366 78056 884422
rect 78112 884366 78180 884422
rect 78236 884366 78304 884422
rect 78360 884366 78428 884422
rect 78484 884366 78552 884422
rect 78608 884366 78678 884422
rect 70130 884354 78678 884366
rect 70000 884298 78678 884354
rect 70000 884286 77808 884298
rect 70000 884230 70074 884286
rect 70130 884242 77808 884286
rect 77864 884242 77932 884298
rect 77988 884242 78056 884298
rect 78112 884242 78180 884298
rect 78236 884242 78304 884298
rect 78360 884242 78428 884298
rect 78484 884242 78552 884298
rect 78608 884242 78678 884298
rect 70130 884230 78678 884242
rect 70000 884174 78678 884230
rect 70000 884162 77808 884174
rect 70000 884106 70074 884162
rect 70130 884118 77808 884162
rect 77864 884118 77932 884174
rect 77988 884118 78056 884174
rect 78112 884118 78180 884174
rect 78236 884118 78304 884174
rect 78360 884118 78428 884174
rect 78484 884118 78552 884174
rect 78608 884118 78678 884174
rect 70130 884106 78678 884118
rect 70000 884050 78678 884106
rect 70000 884038 77808 884050
rect 70000 883982 70074 884038
rect 70130 883994 77808 884038
rect 77864 883994 77932 884050
rect 77988 883994 78056 884050
rect 78112 883994 78180 884050
rect 78236 883994 78304 884050
rect 78360 883994 78428 884050
rect 78484 883994 78552 884050
rect 78608 883994 78678 884050
rect 70130 883982 78678 883994
rect 70000 883926 78678 883982
rect 70000 883914 77808 883926
rect 70000 883858 70074 883914
rect 70130 883870 77808 883914
rect 77864 883870 77932 883926
rect 77988 883870 78056 883926
rect 78112 883870 78180 883926
rect 78236 883870 78304 883926
rect 78360 883870 78428 883926
rect 78484 883870 78552 883926
rect 78608 883870 78678 883926
rect 70130 883858 78678 883870
rect 70000 883802 78678 883858
rect 70000 883790 77808 883802
rect 70000 883734 70074 883790
rect 70130 883746 77808 883790
rect 77864 883746 77932 883802
rect 77988 883746 78056 883802
rect 78112 883746 78180 883802
rect 78236 883746 78304 883802
rect 78360 883746 78428 883802
rect 78484 883746 78552 883802
rect 78608 883746 78678 883802
rect 70130 883734 78678 883746
rect 70000 883678 78678 883734
rect 70000 883666 77808 883678
rect 70000 883610 70074 883666
rect 70130 883622 77808 883666
rect 77864 883622 77932 883678
rect 77988 883622 78056 883678
rect 78112 883622 78180 883678
rect 78236 883622 78304 883678
rect 78360 883622 78428 883678
rect 78484 883622 78552 883678
rect 78608 883622 78678 883678
rect 70130 883610 78678 883622
rect 70000 883554 78678 883610
rect 70000 883542 77808 883554
rect 70000 883486 70074 883542
rect 70130 883498 77808 883542
rect 77864 883498 77932 883554
rect 77988 883498 78056 883554
rect 78112 883498 78180 883554
rect 78236 883498 78304 883554
rect 78360 883498 78428 883554
rect 78484 883498 78552 883554
rect 78608 883498 78678 883554
rect 70130 883486 78678 883498
rect 70000 883430 78678 883486
rect 70000 883418 77808 883430
rect 70000 883362 70074 883418
rect 70130 883374 77808 883418
rect 77864 883374 77932 883430
rect 77988 883374 78056 883430
rect 78112 883374 78180 883430
rect 78236 883374 78304 883430
rect 78360 883374 78428 883430
rect 78484 883374 78552 883430
rect 78608 883374 78678 883430
rect 70130 883362 78678 883374
rect 70000 883306 78678 883362
rect 70000 883294 77808 883306
rect 70000 883238 70074 883294
rect 70130 883250 77808 883294
rect 77864 883250 77932 883306
rect 77988 883250 78056 883306
rect 78112 883250 78180 883306
rect 78236 883250 78304 883306
rect 78360 883250 78428 883306
rect 78484 883250 78552 883306
rect 78608 883250 78678 883306
rect 70130 883238 78678 883250
rect 70000 883182 78678 883238
rect 70000 883170 77808 883182
rect 70000 883114 70074 883170
rect 70130 883126 77808 883170
rect 77864 883126 77932 883182
rect 77988 883126 78056 883182
rect 78112 883126 78180 883182
rect 78236 883126 78304 883182
rect 78360 883126 78428 883182
rect 78484 883126 78552 883182
rect 78608 883126 78678 883182
rect 70130 883114 78678 883126
rect 70000 883058 78678 883114
rect 70000 883046 77808 883058
rect 70000 882990 70074 883046
rect 70130 883002 77808 883046
rect 77864 883002 77932 883058
rect 77988 883002 78056 883058
rect 78112 883002 78180 883058
rect 78236 883002 78304 883058
rect 78360 883002 78428 883058
rect 78484 883002 78552 883058
rect 78608 883002 78678 883058
rect 70130 882990 78678 883002
rect 70000 882934 78678 882990
rect 70000 882922 77808 882934
rect 70000 882866 70074 882922
rect 70130 882878 77808 882922
rect 77864 882878 77932 882934
rect 77988 882878 78056 882934
rect 78112 882878 78180 882934
rect 78236 882878 78304 882934
rect 78360 882878 78428 882934
rect 78484 882878 78552 882934
rect 78608 882878 78678 882934
rect 70130 882866 78678 882878
rect 70000 882828 78678 882866
rect 699322 883658 708000 883728
rect 699322 883652 707870 883658
rect 699322 883596 699392 883652
rect 699448 883596 699516 883652
rect 699572 883596 699640 883652
rect 699696 883596 699764 883652
rect 699820 883596 699888 883652
rect 699944 883596 700012 883652
rect 700068 883596 700136 883652
rect 700192 883602 707870 883652
rect 707926 883602 708000 883658
rect 700192 883596 708000 883602
rect 699322 883534 708000 883596
rect 699322 883528 707870 883534
rect 699322 883472 699392 883528
rect 699448 883472 699516 883528
rect 699572 883472 699640 883528
rect 699696 883472 699764 883528
rect 699820 883472 699888 883528
rect 699944 883472 700012 883528
rect 700068 883472 700136 883528
rect 700192 883478 707870 883528
rect 707926 883478 708000 883534
rect 700192 883472 708000 883478
rect 699322 883410 708000 883472
rect 699322 883404 707870 883410
rect 699322 883348 699392 883404
rect 699448 883348 699516 883404
rect 699572 883348 699640 883404
rect 699696 883348 699764 883404
rect 699820 883348 699888 883404
rect 699944 883348 700012 883404
rect 700068 883348 700136 883404
rect 700192 883354 707870 883404
rect 707926 883354 708000 883410
rect 700192 883348 708000 883354
rect 699322 883286 708000 883348
rect 699322 883280 707870 883286
rect 699322 883224 699392 883280
rect 699448 883224 699516 883280
rect 699572 883224 699640 883280
rect 699696 883224 699764 883280
rect 699820 883224 699888 883280
rect 699944 883224 700012 883280
rect 700068 883224 700136 883280
rect 700192 883230 707870 883280
rect 707926 883230 708000 883286
rect 700192 883224 708000 883230
rect 699322 883162 708000 883224
rect 699322 883156 707870 883162
rect 699322 883100 699392 883156
rect 699448 883100 699516 883156
rect 699572 883100 699640 883156
rect 699696 883100 699764 883156
rect 699820 883100 699888 883156
rect 699944 883100 700012 883156
rect 700068 883100 700136 883156
rect 700192 883106 707870 883156
rect 707926 883106 708000 883162
rect 700192 883100 708000 883106
rect 699322 883038 708000 883100
rect 699322 883032 707870 883038
rect 699322 882976 699392 883032
rect 699448 882976 699516 883032
rect 699572 882976 699640 883032
rect 699696 882976 699764 883032
rect 699820 882976 699888 883032
rect 699944 882976 700012 883032
rect 700068 882976 700136 883032
rect 700192 882982 707870 883032
rect 707926 882982 708000 883038
rect 700192 882976 708000 882982
rect 699322 882914 708000 882976
rect 699322 882908 707870 882914
rect 699322 882852 699392 882908
rect 699448 882852 699516 882908
rect 699572 882852 699640 882908
rect 699696 882852 699764 882908
rect 699820 882852 699888 882908
rect 699944 882852 700012 882908
rect 700068 882852 700136 882908
rect 700192 882858 707870 882908
rect 707926 882858 708000 882914
rect 700192 882852 708000 882858
rect 699322 882790 708000 882852
rect 699322 882784 707870 882790
rect 699322 882728 699392 882784
rect 699448 882728 699516 882784
rect 699572 882728 699640 882784
rect 699696 882728 699764 882784
rect 699820 882728 699888 882784
rect 699944 882728 700012 882784
rect 700068 882728 700136 882784
rect 700192 882734 707870 882784
rect 707926 882734 708000 882790
rect 700192 882728 708000 882734
rect 699322 882666 708000 882728
rect 699322 882660 707870 882666
rect 699322 882604 699392 882660
rect 699448 882604 699516 882660
rect 699572 882604 699640 882660
rect 699696 882604 699764 882660
rect 699820 882604 699888 882660
rect 699944 882604 700012 882660
rect 700068 882604 700136 882660
rect 700192 882610 707870 882660
rect 707926 882610 708000 882666
rect 700192 882604 708000 882610
rect 699322 882542 708000 882604
rect 699322 882536 707870 882542
rect 699322 882480 699392 882536
rect 699448 882480 699516 882536
rect 699572 882480 699640 882536
rect 699696 882480 699764 882536
rect 699820 882480 699888 882536
rect 699944 882480 700012 882536
rect 700068 882480 700136 882536
rect 700192 882486 707870 882536
rect 707926 882486 708000 882542
rect 700192 882480 708000 882486
rect 699322 882418 708000 882480
rect 699322 882412 707870 882418
rect 699322 882356 699392 882412
rect 699448 882356 699516 882412
rect 699572 882356 699640 882412
rect 699696 882356 699764 882412
rect 699820 882356 699888 882412
rect 699944 882356 700012 882412
rect 700068 882356 700136 882412
rect 700192 882362 707870 882412
rect 707926 882362 708000 882418
rect 700192 882356 708000 882362
rect 699322 882294 708000 882356
rect 699322 882288 707870 882294
rect 70000 882190 78678 882248
rect 70000 882184 77808 882190
rect 70000 882128 70074 882184
rect 70130 882134 77808 882184
rect 77864 882134 77932 882190
rect 77988 882134 78056 882190
rect 78112 882134 78180 882190
rect 78236 882134 78304 882190
rect 78360 882134 78428 882190
rect 78484 882134 78552 882190
rect 78608 882134 78678 882190
rect 70130 882128 78678 882134
rect 70000 882066 78678 882128
rect 70000 882060 77808 882066
rect 70000 882004 70074 882060
rect 70130 882010 77808 882060
rect 77864 882010 77932 882066
rect 77988 882010 78056 882066
rect 78112 882010 78180 882066
rect 78236 882010 78304 882066
rect 78360 882010 78428 882066
rect 78484 882010 78552 882066
rect 78608 882010 78678 882066
rect 70130 882004 78678 882010
rect 70000 881942 78678 882004
rect 70000 881936 77808 881942
rect 70000 881880 70074 881936
rect 70130 881886 77808 881936
rect 77864 881886 77932 881942
rect 77988 881886 78056 881942
rect 78112 881886 78180 881942
rect 78236 881886 78304 881942
rect 78360 881886 78428 881942
rect 78484 881886 78552 881942
rect 78608 881886 78678 881942
rect 70130 881880 78678 881886
rect 70000 881818 78678 881880
rect 699322 882232 699392 882288
rect 699448 882232 699516 882288
rect 699572 882232 699640 882288
rect 699696 882232 699764 882288
rect 699820 882232 699888 882288
rect 699944 882232 700012 882288
rect 700068 882232 700136 882288
rect 700192 882238 707870 882288
rect 707926 882238 708000 882294
rect 700192 882232 708000 882238
rect 699322 882170 708000 882232
rect 699322 882164 707870 882170
rect 699322 882108 699392 882164
rect 699448 882108 699516 882164
rect 699572 882108 699640 882164
rect 699696 882108 699764 882164
rect 699820 882108 699888 882164
rect 699944 882108 700012 882164
rect 700068 882108 700136 882164
rect 700192 882114 707870 882164
rect 707926 882114 708000 882170
rect 700192 882108 708000 882114
rect 699322 882046 708000 882108
rect 699322 882040 707870 882046
rect 699322 881984 699392 882040
rect 699448 881984 699516 882040
rect 699572 881984 699640 882040
rect 699696 881984 699764 882040
rect 699820 881984 699888 882040
rect 699944 881984 700012 882040
rect 700068 881984 700136 882040
rect 700192 881990 707870 882040
rect 707926 881990 708000 882046
rect 700192 881984 708000 881990
rect 699322 881922 708000 881984
rect 699322 881916 707870 881922
rect 699322 881860 699392 881916
rect 699448 881860 699516 881916
rect 699572 881860 699640 881916
rect 699696 881860 699764 881916
rect 699820 881860 699888 881916
rect 699944 881860 700012 881916
rect 700068 881860 700136 881916
rect 700192 881866 707870 881916
rect 707926 881866 708000 881922
rect 700192 881860 708000 881866
rect 699322 881828 708000 881860
rect 70000 881812 77808 881818
rect 70000 881756 70074 881812
rect 70130 881762 77808 881812
rect 77864 881762 77932 881818
rect 77988 881762 78056 881818
rect 78112 881762 78180 881818
rect 78236 881762 78304 881818
rect 78360 881762 78428 881818
rect 78484 881762 78552 881818
rect 78608 881762 78678 881818
rect 70130 881756 78678 881762
rect 70000 881694 78678 881756
rect 70000 881688 77808 881694
rect 70000 881632 70074 881688
rect 70130 881638 77808 881688
rect 77864 881638 77932 881694
rect 77988 881638 78056 881694
rect 78112 881638 78180 881694
rect 78236 881638 78304 881694
rect 78360 881638 78428 881694
rect 78484 881638 78552 881694
rect 78608 881638 78678 881694
rect 70130 881632 78678 881638
rect 70000 881570 78678 881632
rect 70000 881564 77808 881570
rect 70000 881508 70074 881564
rect 70130 881514 77808 881564
rect 77864 881514 77932 881570
rect 77988 881514 78056 881570
rect 78112 881514 78180 881570
rect 78236 881514 78304 881570
rect 78360 881514 78428 881570
rect 78484 881514 78552 881570
rect 78608 881514 78678 881570
rect 70130 881508 78678 881514
rect 70000 881446 78678 881508
rect 70000 881440 77808 881446
rect 70000 881384 70074 881440
rect 70130 881390 77808 881440
rect 77864 881390 77932 881446
rect 77988 881390 78056 881446
rect 78112 881390 78180 881446
rect 78236 881390 78304 881446
rect 78360 881390 78428 881446
rect 78484 881390 78552 881446
rect 78608 881390 78678 881446
rect 70130 881384 78678 881390
rect 70000 881322 78678 881384
rect 70000 881316 77808 881322
rect 70000 881260 70074 881316
rect 70130 881266 77808 881316
rect 77864 881266 77932 881322
rect 77988 881266 78056 881322
rect 78112 881266 78180 881322
rect 78236 881266 78304 881322
rect 78360 881266 78428 881322
rect 78484 881266 78552 881322
rect 78608 881266 78678 881322
rect 70130 881260 78678 881266
rect 70000 881198 78678 881260
rect 70000 881192 77808 881198
rect 70000 881136 70074 881192
rect 70130 881142 77808 881192
rect 77864 881142 77932 881198
rect 77988 881142 78056 881198
rect 78112 881142 78180 881198
rect 78236 881142 78304 881198
rect 78360 881142 78428 881198
rect 78484 881142 78552 881198
rect 78608 881142 78678 881198
rect 70130 881136 78678 881142
rect 70000 881074 78678 881136
rect 70000 881068 77808 881074
rect 70000 881012 70074 881068
rect 70130 881018 77808 881068
rect 77864 881018 77932 881074
rect 77988 881018 78056 881074
rect 78112 881018 78180 881074
rect 78236 881018 78304 881074
rect 78360 881018 78428 881074
rect 78484 881018 78552 881074
rect 78608 881018 78678 881074
rect 70130 881012 78678 881018
rect 70000 880950 78678 881012
rect 70000 880944 77808 880950
rect 70000 880888 70074 880944
rect 70130 880894 77808 880944
rect 77864 880894 77932 880950
rect 77988 880894 78056 880950
rect 78112 880894 78180 880950
rect 78236 880894 78304 880950
rect 78360 880894 78428 880950
rect 78484 880894 78552 880950
rect 78608 880894 78678 880950
rect 70130 880888 78678 880894
rect 70000 880826 78678 880888
rect 70000 880820 77808 880826
rect 70000 880764 70074 880820
rect 70130 880770 77808 880820
rect 77864 880770 77932 880826
rect 77988 880770 78056 880826
rect 78112 880770 78180 880826
rect 78236 880770 78304 880826
rect 78360 880770 78428 880826
rect 78484 880770 78552 880826
rect 78608 880770 78678 880826
rect 70130 880764 78678 880770
rect 70000 880702 78678 880764
rect 70000 880696 77808 880702
rect 70000 880640 70074 880696
rect 70130 880646 77808 880696
rect 77864 880646 77932 880702
rect 77988 880646 78056 880702
rect 78112 880646 78180 880702
rect 78236 880646 78304 880702
rect 78360 880646 78428 880702
rect 78484 880646 78552 880702
rect 78608 880646 78678 880702
rect 70130 880640 78678 880646
rect 70000 880578 78678 880640
rect 70000 880572 77808 880578
rect 70000 880516 70074 880572
rect 70130 880522 77808 880572
rect 77864 880522 77932 880578
rect 77988 880522 78056 880578
rect 78112 880522 78180 880578
rect 78236 880522 78304 880578
rect 78360 880522 78428 880578
rect 78484 880522 78552 880578
rect 78608 880522 78678 880578
rect 70130 880516 78678 880522
rect 70000 880454 78678 880516
rect 70000 880448 77808 880454
rect 70000 880392 70074 880448
rect 70130 880398 77808 880448
rect 77864 880398 77932 880454
rect 77988 880398 78056 880454
rect 78112 880398 78180 880454
rect 78236 880398 78304 880454
rect 78360 880398 78428 880454
rect 78484 880398 78552 880454
rect 78608 880398 78678 880454
rect 70130 880392 78678 880398
rect 70000 880330 78678 880392
rect 70000 880324 77808 880330
rect 70000 880268 70074 880324
rect 70130 880274 77808 880324
rect 77864 880274 77932 880330
rect 77988 880274 78056 880330
rect 78112 880274 78180 880330
rect 78236 880274 78304 880330
rect 78360 880274 78428 880330
rect 78484 880274 78552 880330
rect 78608 880274 78678 880330
rect 70130 880268 78678 880274
rect 70000 880198 78678 880268
rect 699322 881178 708000 881248
rect 699322 881172 707870 881178
rect 699322 881116 699392 881172
rect 699448 881116 699516 881172
rect 699572 881116 699640 881172
rect 699696 881116 699764 881172
rect 699820 881116 699888 881172
rect 699944 881116 700012 881172
rect 700068 881116 700136 881172
rect 700192 881122 707870 881172
rect 707926 881122 708000 881178
rect 700192 881116 708000 881122
rect 699322 881054 708000 881116
rect 699322 881048 707870 881054
rect 699322 880992 699392 881048
rect 699448 880992 699516 881048
rect 699572 880992 699640 881048
rect 699696 880992 699764 881048
rect 699820 880992 699888 881048
rect 699944 880992 700012 881048
rect 700068 880992 700136 881048
rect 700192 880998 707870 881048
rect 707926 880998 708000 881054
rect 700192 880992 708000 880998
rect 699322 880930 708000 880992
rect 699322 880924 707870 880930
rect 699322 880868 699392 880924
rect 699448 880868 699516 880924
rect 699572 880868 699640 880924
rect 699696 880868 699764 880924
rect 699820 880868 699888 880924
rect 699944 880868 700012 880924
rect 700068 880868 700136 880924
rect 700192 880874 707870 880924
rect 707926 880874 708000 880930
rect 700192 880868 708000 880874
rect 699322 880806 708000 880868
rect 699322 880800 707870 880806
rect 699322 880744 699392 880800
rect 699448 880744 699516 880800
rect 699572 880744 699640 880800
rect 699696 880744 699764 880800
rect 699820 880744 699888 880800
rect 699944 880744 700012 880800
rect 700068 880744 700136 880800
rect 700192 880750 707870 880800
rect 707926 880750 708000 880806
rect 700192 880744 708000 880750
rect 699322 880682 708000 880744
rect 699322 880676 707870 880682
rect 699322 880620 699392 880676
rect 699448 880620 699516 880676
rect 699572 880620 699640 880676
rect 699696 880620 699764 880676
rect 699820 880620 699888 880676
rect 699944 880620 700012 880676
rect 700068 880620 700136 880676
rect 700192 880626 707870 880676
rect 707926 880626 708000 880682
rect 700192 880620 708000 880626
rect 699322 880558 708000 880620
rect 699322 880552 707870 880558
rect 699322 880496 699392 880552
rect 699448 880496 699516 880552
rect 699572 880496 699640 880552
rect 699696 880496 699764 880552
rect 699820 880496 699888 880552
rect 699944 880496 700012 880552
rect 700068 880496 700136 880552
rect 700192 880502 707870 880552
rect 707926 880502 708000 880558
rect 700192 880496 708000 880502
rect 699322 880434 708000 880496
rect 699322 880428 707870 880434
rect 699322 880372 699392 880428
rect 699448 880372 699516 880428
rect 699572 880372 699640 880428
rect 699696 880372 699764 880428
rect 699820 880372 699888 880428
rect 699944 880372 700012 880428
rect 700068 880372 700136 880428
rect 700192 880378 707870 880428
rect 707926 880378 708000 880434
rect 700192 880372 708000 880378
rect 699322 880310 708000 880372
rect 699322 880304 707870 880310
rect 699322 880248 699392 880304
rect 699448 880248 699516 880304
rect 699572 880248 699640 880304
rect 699696 880248 699764 880304
rect 699820 880248 699888 880304
rect 699944 880248 700012 880304
rect 700068 880248 700136 880304
rect 700192 880254 707870 880304
rect 707926 880254 708000 880310
rect 700192 880248 708000 880254
rect 699322 880186 708000 880248
rect 699322 880180 707870 880186
rect 699322 880124 699392 880180
rect 699448 880124 699516 880180
rect 699572 880124 699640 880180
rect 699696 880124 699764 880180
rect 699820 880124 699888 880180
rect 699944 880124 700012 880180
rect 700068 880124 700136 880180
rect 700192 880130 707870 880180
rect 707926 880130 708000 880186
rect 700192 880124 708000 880130
rect 699322 880062 708000 880124
rect 699322 880056 707870 880062
rect 699322 880000 699392 880056
rect 699448 880000 699516 880056
rect 699572 880000 699640 880056
rect 699696 880000 699764 880056
rect 699820 880000 699888 880056
rect 699944 880000 700012 880056
rect 700068 880000 700136 880056
rect 700192 880006 707870 880056
rect 707926 880006 708000 880062
rect 700192 880000 708000 880006
rect 699322 879938 708000 880000
rect 699322 879932 707870 879938
rect 70000 879820 78678 879878
rect 70000 879814 77808 879820
rect 70000 879758 70074 879814
rect 70130 879764 77808 879814
rect 77864 879764 77932 879820
rect 77988 879764 78056 879820
rect 78112 879764 78180 879820
rect 78236 879764 78304 879820
rect 78360 879764 78428 879820
rect 78484 879764 78552 879820
rect 78608 879764 78678 879820
rect 70130 879758 78678 879764
rect 70000 879696 78678 879758
rect 70000 879690 77808 879696
rect 70000 879634 70074 879690
rect 70130 879640 77808 879690
rect 77864 879640 77932 879696
rect 77988 879640 78056 879696
rect 78112 879640 78180 879696
rect 78236 879640 78304 879696
rect 78360 879640 78428 879696
rect 78484 879640 78552 879696
rect 78608 879640 78678 879696
rect 70130 879634 78678 879640
rect 70000 879572 78678 879634
rect 70000 879566 77808 879572
rect 70000 879510 70074 879566
rect 70130 879516 77808 879566
rect 77864 879516 77932 879572
rect 77988 879516 78056 879572
rect 78112 879516 78180 879572
rect 78236 879516 78304 879572
rect 78360 879516 78428 879572
rect 78484 879516 78552 879572
rect 78608 879516 78678 879572
rect 70130 879510 78678 879516
rect 70000 879448 78678 879510
rect 70000 879442 77808 879448
rect 70000 879386 70074 879442
rect 70130 879392 77808 879442
rect 77864 879392 77932 879448
rect 77988 879392 78056 879448
rect 78112 879392 78180 879448
rect 78236 879392 78304 879448
rect 78360 879392 78428 879448
rect 78484 879392 78552 879448
rect 78608 879392 78678 879448
rect 70130 879386 78678 879392
rect 70000 879324 78678 879386
rect 70000 879318 77808 879324
rect 70000 879262 70074 879318
rect 70130 879268 77808 879318
rect 77864 879268 77932 879324
rect 77988 879268 78056 879324
rect 78112 879268 78180 879324
rect 78236 879268 78304 879324
rect 78360 879268 78428 879324
rect 78484 879268 78552 879324
rect 78608 879268 78678 879324
rect 70130 879262 78678 879268
rect 70000 879200 78678 879262
rect 70000 879194 77808 879200
rect 70000 879138 70074 879194
rect 70130 879144 77808 879194
rect 77864 879144 77932 879200
rect 77988 879144 78056 879200
rect 78112 879144 78180 879200
rect 78236 879144 78304 879200
rect 78360 879144 78428 879200
rect 78484 879144 78552 879200
rect 78608 879144 78678 879200
rect 699322 879876 699392 879932
rect 699448 879876 699516 879932
rect 699572 879876 699640 879932
rect 699696 879876 699764 879932
rect 699820 879876 699888 879932
rect 699944 879876 700012 879932
rect 700068 879876 700136 879932
rect 700192 879882 707870 879932
rect 707926 879882 708000 879938
rect 700192 879876 708000 879882
rect 699322 879814 708000 879876
rect 699322 879808 707870 879814
rect 699322 879752 699392 879808
rect 699448 879752 699516 879808
rect 699572 879752 699640 879808
rect 699696 879752 699764 879808
rect 699820 879752 699888 879808
rect 699944 879752 700012 879808
rect 700068 879752 700136 879808
rect 700192 879758 707870 879808
rect 707926 879758 708000 879814
rect 700192 879752 708000 879758
rect 699322 879690 708000 879752
rect 699322 879684 707870 879690
rect 699322 879628 699392 879684
rect 699448 879628 699516 879684
rect 699572 879628 699640 879684
rect 699696 879628 699764 879684
rect 699820 879628 699888 879684
rect 699944 879628 700012 879684
rect 700068 879628 700136 879684
rect 700192 879634 707870 879684
rect 707926 879634 708000 879690
rect 700192 879628 708000 879634
rect 699322 879566 708000 879628
rect 699322 879560 707870 879566
rect 699322 879504 699392 879560
rect 699448 879504 699516 879560
rect 699572 879504 699640 879560
rect 699696 879504 699764 879560
rect 699820 879504 699888 879560
rect 699944 879504 700012 879560
rect 700068 879504 700136 879560
rect 700192 879510 707870 879560
rect 707926 879510 708000 879566
rect 700192 879504 708000 879510
rect 699322 879442 708000 879504
rect 699322 879436 707870 879442
rect 699322 879380 699392 879436
rect 699448 879380 699516 879436
rect 699572 879380 699640 879436
rect 699696 879380 699764 879436
rect 699820 879380 699888 879436
rect 699944 879380 700012 879436
rect 700068 879380 700136 879436
rect 700192 879386 707870 879436
rect 707926 879386 708000 879442
rect 700192 879380 708000 879386
rect 699322 879318 708000 879380
rect 699322 879312 707870 879318
rect 699322 879256 699392 879312
rect 699448 879256 699516 879312
rect 699572 879256 699640 879312
rect 699696 879256 699764 879312
rect 699820 879256 699888 879312
rect 699944 879256 700012 879312
rect 700068 879256 700136 879312
rect 700192 879262 707870 879312
rect 707926 879262 708000 879318
rect 700192 879256 708000 879262
rect 699322 879198 708000 879256
rect 70130 879138 78678 879144
rect 70000 879076 78678 879138
rect 70000 879070 77808 879076
rect 70000 879014 70074 879070
rect 70130 879020 77808 879070
rect 77864 879020 77932 879076
rect 77988 879020 78056 879076
rect 78112 879020 78180 879076
rect 78236 879020 78304 879076
rect 78360 879020 78428 879076
rect 78484 879020 78552 879076
rect 78608 879020 78678 879076
rect 70130 879014 78678 879020
rect 70000 878952 78678 879014
rect 70000 878946 77808 878952
rect 70000 878890 70074 878946
rect 70130 878896 77808 878946
rect 77864 878896 77932 878952
rect 77988 878896 78056 878952
rect 78112 878896 78180 878952
rect 78236 878896 78304 878952
rect 78360 878896 78428 878952
rect 78484 878896 78552 878952
rect 78608 878896 78678 878952
rect 70130 878890 78678 878896
rect 70000 878828 78678 878890
rect 70000 878822 77808 878828
rect 70000 878766 70074 878822
rect 70130 878772 77808 878822
rect 77864 878772 77932 878828
rect 77988 878772 78056 878828
rect 78112 878772 78180 878828
rect 78236 878772 78304 878828
rect 78360 878772 78428 878828
rect 78484 878772 78552 878828
rect 78608 878772 78678 878828
rect 70130 878766 78678 878772
rect 70000 878704 78678 878766
rect 70000 878698 77808 878704
rect 70000 878642 70074 878698
rect 70130 878648 77808 878698
rect 77864 878648 77932 878704
rect 77988 878648 78056 878704
rect 78112 878648 78180 878704
rect 78236 878648 78304 878704
rect 78360 878648 78428 878704
rect 78484 878648 78552 878704
rect 78608 878648 78678 878704
rect 70130 878642 78678 878648
rect 70000 878580 78678 878642
rect 70000 878574 77808 878580
rect 70000 878518 70074 878574
rect 70130 878524 77808 878574
rect 77864 878524 77932 878580
rect 77988 878524 78056 878580
rect 78112 878524 78180 878580
rect 78236 878524 78304 878580
rect 78360 878524 78428 878580
rect 78484 878524 78552 878580
rect 78608 878524 78678 878580
rect 70130 878518 78678 878524
rect 70000 878456 78678 878518
rect 70000 878450 77808 878456
rect 70000 878394 70074 878450
rect 70130 878400 77808 878450
rect 77864 878400 77932 878456
rect 77988 878400 78056 878456
rect 78112 878400 78180 878456
rect 78236 878400 78304 878456
rect 78360 878400 78428 878456
rect 78484 878400 78552 878456
rect 78608 878400 78678 878456
rect 70130 878394 78678 878400
rect 70000 878332 78678 878394
rect 70000 878326 77808 878332
rect 70000 878270 70074 878326
rect 70130 878276 77808 878326
rect 77864 878276 77932 878332
rect 77988 878276 78056 878332
rect 78112 878276 78180 878332
rect 78236 878276 78304 878332
rect 78360 878276 78428 878332
rect 78484 878276 78552 878332
rect 78608 878276 78678 878332
rect 70130 878270 78678 878276
rect 70000 878208 78678 878270
rect 70000 878202 77808 878208
rect 70000 878146 70074 878202
rect 70130 878152 77808 878202
rect 77864 878152 77932 878208
rect 77988 878152 78056 878208
rect 78112 878152 78180 878208
rect 78236 878152 78304 878208
rect 78360 878152 78428 878208
rect 78484 878152 78552 878208
rect 78608 878152 78678 878208
rect 70130 878146 78678 878152
rect 70000 878084 78678 878146
rect 70000 878078 77808 878084
rect 70000 878022 70074 878078
rect 70130 878028 77808 878078
rect 77864 878028 77932 878084
rect 77988 878028 78056 878084
rect 78112 878028 78180 878084
rect 78236 878028 78304 878084
rect 78360 878028 78428 878084
rect 78484 878028 78552 878084
rect 78608 878028 78678 878084
rect 70130 878022 78678 878028
rect 70000 877960 78678 878022
rect 70000 877954 77808 877960
rect 70000 877898 70074 877954
rect 70130 877904 77808 877954
rect 77864 877904 77932 877960
rect 77988 877904 78056 877960
rect 78112 877904 78180 877960
rect 78236 877904 78304 877960
rect 78360 877904 78428 877960
rect 78484 877904 78552 877960
rect 78608 877904 78678 877960
rect 70130 877898 78678 877904
rect 70000 877828 78678 877898
rect 699322 878808 708000 878878
rect 699322 878802 707870 878808
rect 699322 878746 699392 878802
rect 699448 878746 699516 878802
rect 699572 878746 699640 878802
rect 699696 878746 699764 878802
rect 699820 878746 699888 878802
rect 699944 878746 700012 878802
rect 700068 878746 700136 878802
rect 700192 878752 707870 878802
rect 707926 878752 708000 878808
rect 700192 878746 708000 878752
rect 699322 878684 708000 878746
rect 699322 878678 707870 878684
rect 699322 878622 699392 878678
rect 699448 878622 699516 878678
rect 699572 878622 699640 878678
rect 699696 878622 699764 878678
rect 699820 878622 699888 878678
rect 699944 878622 700012 878678
rect 700068 878622 700136 878678
rect 700192 878628 707870 878678
rect 707926 878628 708000 878684
rect 700192 878622 708000 878628
rect 699322 878560 708000 878622
rect 699322 878554 707870 878560
rect 699322 878498 699392 878554
rect 699448 878498 699516 878554
rect 699572 878498 699640 878554
rect 699696 878498 699764 878554
rect 699820 878498 699888 878554
rect 699944 878498 700012 878554
rect 700068 878498 700136 878554
rect 700192 878504 707870 878554
rect 707926 878504 708000 878560
rect 700192 878498 708000 878504
rect 699322 878436 708000 878498
rect 699322 878430 707870 878436
rect 699322 878374 699392 878430
rect 699448 878374 699516 878430
rect 699572 878374 699640 878430
rect 699696 878374 699764 878430
rect 699820 878374 699888 878430
rect 699944 878374 700012 878430
rect 700068 878374 700136 878430
rect 700192 878380 707870 878430
rect 707926 878380 708000 878436
rect 700192 878374 708000 878380
rect 699322 878312 708000 878374
rect 699322 878306 707870 878312
rect 699322 878250 699392 878306
rect 699448 878250 699516 878306
rect 699572 878250 699640 878306
rect 699696 878250 699764 878306
rect 699820 878250 699888 878306
rect 699944 878250 700012 878306
rect 700068 878250 700136 878306
rect 700192 878256 707870 878306
rect 707926 878256 708000 878312
rect 700192 878250 708000 878256
rect 699322 878188 708000 878250
rect 699322 878182 707870 878188
rect 699322 878126 699392 878182
rect 699448 878126 699516 878182
rect 699572 878126 699640 878182
rect 699696 878126 699764 878182
rect 699820 878126 699888 878182
rect 699944 878126 700012 878182
rect 700068 878126 700136 878182
rect 700192 878132 707870 878182
rect 707926 878132 708000 878188
rect 700192 878126 708000 878132
rect 699322 878064 708000 878126
rect 699322 878058 707870 878064
rect 699322 878002 699392 878058
rect 699448 878002 699516 878058
rect 699572 878002 699640 878058
rect 699696 878002 699764 878058
rect 699820 878002 699888 878058
rect 699944 878002 700012 878058
rect 700068 878002 700136 878058
rect 700192 878008 707870 878058
rect 707926 878008 708000 878064
rect 700192 878002 708000 878008
rect 699322 877940 708000 878002
rect 699322 877934 707870 877940
rect 699322 877878 699392 877934
rect 699448 877878 699516 877934
rect 699572 877878 699640 877934
rect 699696 877878 699764 877934
rect 699820 877878 699888 877934
rect 699944 877878 700012 877934
rect 700068 877878 700136 877934
rect 700192 877884 707870 877934
rect 707926 877884 708000 877940
rect 700192 877878 708000 877884
rect 699322 877816 708000 877878
rect 699322 877810 707870 877816
rect 699322 877754 699392 877810
rect 699448 877754 699516 877810
rect 699572 877754 699640 877810
rect 699696 877754 699764 877810
rect 699820 877754 699888 877810
rect 699944 877754 700012 877810
rect 700068 877754 700136 877810
rect 700192 877760 707870 877810
rect 707926 877760 708000 877816
rect 700192 877754 708000 877760
rect 699322 877692 708000 877754
rect 699322 877686 707870 877692
rect 699322 877630 699392 877686
rect 699448 877630 699516 877686
rect 699572 877630 699640 877686
rect 699696 877630 699764 877686
rect 699820 877630 699888 877686
rect 699944 877630 700012 877686
rect 700068 877630 700136 877686
rect 700192 877636 707870 877686
rect 707926 877636 708000 877692
rect 700192 877630 708000 877636
rect 699322 877568 708000 877630
rect 699322 877562 707870 877568
rect 699322 877506 699392 877562
rect 699448 877506 699516 877562
rect 699572 877506 699640 877562
rect 699696 877506 699764 877562
rect 699820 877506 699888 877562
rect 699944 877506 700012 877562
rect 700068 877506 700136 877562
rect 700192 877512 707870 877562
rect 707926 877512 708000 877568
rect 700192 877506 708000 877512
rect 699322 877444 708000 877506
rect 699322 877438 707870 877444
rect 699322 877382 699392 877438
rect 699448 877382 699516 877438
rect 699572 877382 699640 877438
rect 699696 877382 699764 877438
rect 699820 877382 699888 877438
rect 699944 877382 700012 877438
rect 700068 877382 700136 877438
rect 700192 877388 707870 877438
rect 707926 877388 708000 877444
rect 700192 877382 708000 877388
rect 699322 877320 708000 877382
rect 699322 877314 707870 877320
rect 699322 877258 699392 877314
rect 699448 877258 699516 877314
rect 699572 877258 699640 877314
rect 699696 877258 699764 877314
rect 699820 877258 699888 877314
rect 699944 877258 700012 877314
rect 700068 877258 700136 877314
rect 700192 877264 707870 877314
rect 707926 877264 708000 877320
rect 700192 877258 708000 877264
rect 699322 877196 708000 877258
rect 699322 877190 707870 877196
rect 70000 877114 78678 877172
rect 70000 877108 77808 877114
rect 70000 877052 70074 877108
rect 70130 877058 77808 877108
rect 77864 877058 77932 877114
rect 77988 877058 78056 877114
rect 78112 877058 78180 877114
rect 78236 877058 78304 877114
rect 78360 877058 78428 877114
rect 78484 877058 78552 877114
rect 78608 877058 78678 877114
rect 70130 877052 78678 877058
rect 70000 876990 78678 877052
rect 70000 876984 77808 876990
rect 70000 876928 70074 876984
rect 70130 876934 77808 876984
rect 77864 876934 77932 876990
rect 77988 876934 78056 876990
rect 78112 876934 78180 876990
rect 78236 876934 78304 876990
rect 78360 876934 78428 876990
rect 78484 876934 78552 876990
rect 78608 876934 78678 876990
rect 70130 876928 78678 876934
rect 70000 876866 78678 876928
rect 70000 876860 77808 876866
rect 70000 876804 70074 876860
rect 70130 876810 77808 876860
rect 77864 876810 77932 876866
rect 77988 876810 78056 876866
rect 78112 876810 78180 876866
rect 78236 876810 78304 876866
rect 78360 876810 78428 876866
rect 78484 876810 78552 876866
rect 78608 876810 78678 876866
rect 699322 877134 699392 877190
rect 699448 877134 699516 877190
rect 699572 877134 699640 877190
rect 699696 877134 699764 877190
rect 699820 877134 699888 877190
rect 699944 877134 700012 877190
rect 700068 877134 700136 877190
rect 700192 877140 707870 877190
rect 707926 877140 708000 877196
rect 700192 877134 708000 877140
rect 699322 877072 708000 877134
rect 699322 877066 707870 877072
rect 699322 877010 699392 877066
rect 699448 877010 699516 877066
rect 699572 877010 699640 877066
rect 699696 877010 699764 877066
rect 699820 877010 699888 877066
rect 699944 877010 700012 877066
rect 700068 877010 700136 877066
rect 700192 877016 707870 877066
rect 707926 877016 708000 877072
rect 700192 877010 708000 877016
rect 699322 876948 708000 877010
rect 699322 876942 707870 876948
rect 699322 876886 699392 876942
rect 699448 876886 699516 876942
rect 699572 876886 699640 876942
rect 699696 876886 699764 876942
rect 699820 876886 699888 876942
rect 699944 876886 700012 876942
rect 700068 876886 700136 876942
rect 700192 876892 707870 876942
rect 707926 876892 708000 876948
rect 700192 876886 708000 876892
rect 699322 876828 708000 876886
rect 70130 876804 78678 876810
rect 70000 876742 78678 876804
rect 70000 876736 77808 876742
rect 70000 876680 70074 876736
rect 70130 876686 77808 876736
rect 77864 876686 77932 876742
rect 77988 876686 78056 876742
rect 78112 876686 78180 876742
rect 78236 876686 78304 876742
rect 78360 876686 78428 876742
rect 78484 876686 78552 876742
rect 78608 876686 78678 876742
rect 70130 876680 78678 876686
rect 70000 876618 78678 876680
rect 70000 876612 77808 876618
rect 70000 876556 70074 876612
rect 70130 876562 77808 876612
rect 77864 876562 77932 876618
rect 77988 876562 78056 876618
rect 78112 876562 78180 876618
rect 78236 876562 78304 876618
rect 78360 876562 78428 876618
rect 78484 876562 78552 876618
rect 78608 876562 78678 876618
rect 70130 876556 78678 876562
rect 70000 876494 78678 876556
rect 70000 876488 77808 876494
rect 70000 876432 70074 876488
rect 70130 876438 77808 876488
rect 77864 876438 77932 876494
rect 77988 876438 78056 876494
rect 78112 876438 78180 876494
rect 78236 876438 78304 876494
rect 78360 876438 78428 876494
rect 78484 876438 78552 876494
rect 78608 876438 78678 876494
rect 70130 876432 78678 876438
rect 70000 876370 78678 876432
rect 70000 876364 77808 876370
rect 70000 876308 70074 876364
rect 70130 876314 77808 876364
rect 77864 876314 77932 876370
rect 77988 876314 78056 876370
rect 78112 876314 78180 876370
rect 78236 876314 78304 876370
rect 78360 876314 78428 876370
rect 78484 876314 78552 876370
rect 78608 876314 78678 876370
rect 70130 876308 78678 876314
rect 70000 876246 78678 876308
rect 70000 876240 77808 876246
rect 70000 876184 70074 876240
rect 70130 876190 77808 876240
rect 77864 876190 77932 876246
rect 77988 876190 78056 876246
rect 78112 876190 78180 876246
rect 78236 876190 78304 876246
rect 78360 876190 78428 876246
rect 78484 876190 78552 876246
rect 78608 876190 78678 876246
rect 70130 876184 78678 876190
rect 70000 876122 78678 876184
rect 70000 876116 77808 876122
rect 70000 876060 70074 876116
rect 70130 876066 77808 876116
rect 77864 876066 77932 876122
rect 77988 876066 78056 876122
rect 78112 876066 78180 876122
rect 78236 876066 78304 876122
rect 78360 876066 78428 876122
rect 78484 876066 78552 876122
rect 78608 876066 78678 876122
rect 70130 876060 78678 876066
rect 70000 875998 78678 876060
rect 70000 875992 77808 875998
rect 70000 875936 70074 875992
rect 70130 875942 77808 875992
rect 77864 875942 77932 875998
rect 77988 875942 78056 875998
rect 78112 875942 78180 875998
rect 78236 875942 78304 875998
rect 78360 875942 78428 875998
rect 78484 875942 78552 875998
rect 78608 875942 78678 875998
rect 70130 875936 78678 875942
rect 70000 875874 78678 875936
rect 70000 875868 77808 875874
rect 70000 875812 70074 875868
rect 70130 875818 77808 875868
rect 77864 875818 77932 875874
rect 77988 875818 78056 875874
rect 78112 875818 78180 875874
rect 78236 875818 78304 875874
rect 78360 875818 78428 875874
rect 78484 875818 78552 875874
rect 78608 875818 78678 875874
rect 70130 875812 78678 875818
rect 70000 875750 78678 875812
rect 70000 875744 77808 875750
rect 70000 875688 70074 875744
rect 70130 875694 77808 875744
rect 77864 875694 77932 875750
rect 77988 875694 78056 875750
rect 78112 875694 78180 875750
rect 78236 875694 78304 875750
rect 78360 875694 78428 875750
rect 78484 875694 78552 875750
rect 78608 875694 78678 875750
rect 70130 875688 78678 875694
rect 70000 875626 78678 875688
rect 70000 875620 77808 875626
rect 70000 875564 70074 875620
rect 70130 875570 77808 875620
rect 77864 875570 77932 875626
rect 77988 875570 78056 875626
rect 78112 875570 78180 875626
rect 78236 875570 78304 875626
rect 78360 875570 78428 875626
rect 78484 875570 78552 875626
rect 78608 875570 78678 875626
rect 70130 875564 78678 875570
rect 70000 875502 78678 875564
rect 70000 875496 77808 875502
rect 70000 875440 70074 875496
rect 70130 875446 77808 875496
rect 77864 875446 77932 875502
rect 77988 875446 78056 875502
rect 78112 875446 78180 875502
rect 78236 875446 78304 875502
rect 78360 875446 78428 875502
rect 78484 875446 78552 875502
rect 78608 875446 78678 875502
rect 70130 875440 78678 875446
rect 70000 875378 78678 875440
rect 70000 875372 77808 875378
rect 70000 875316 70074 875372
rect 70130 875322 77808 875372
rect 77864 875322 77932 875378
rect 77988 875322 78056 875378
rect 78112 875322 78180 875378
rect 78236 875322 78304 875378
rect 78360 875322 78428 875378
rect 78484 875322 78552 875378
rect 78608 875322 78678 875378
rect 70130 875316 78678 875322
rect 70000 875254 78678 875316
rect 70000 875248 77808 875254
rect 70000 875192 70074 875248
rect 70130 875198 77808 875248
rect 77864 875198 77932 875254
rect 77988 875198 78056 875254
rect 78112 875198 78180 875254
rect 78236 875198 78304 875254
rect 78360 875198 78428 875254
rect 78484 875198 78552 875254
rect 78608 875198 78678 875254
rect 70130 875192 78678 875198
rect 70000 875122 78678 875192
rect 699322 876102 708000 876172
rect 699322 876096 707870 876102
rect 699322 876040 699392 876096
rect 699448 876040 699516 876096
rect 699572 876040 699640 876096
rect 699696 876040 699764 876096
rect 699820 876040 699888 876096
rect 699944 876040 700012 876096
rect 700068 876040 700136 876096
rect 700192 876046 707870 876096
rect 707926 876046 708000 876102
rect 700192 876040 708000 876046
rect 699322 875978 708000 876040
rect 699322 875972 707870 875978
rect 699322 875916 699392 875972
rect 699448 875916 699516 875972
rect 699572 875916 699640 875972
rect 699696 875916 699764 875972
rect 699820 875916 699888 875972
rect 699944 875916 700012 875972
rect 700068 875916 700136 875972
rect 700192 875922 707870 875972
rect 707926 875922 708000 875978
rect 700192 875916 708000 875922
rect 699322 875854 708000 875916
rect 699322 875848 707870 875854
rect 699322 875792 699392 875848
rect 699448 875792 699516 875848
rect 699572 875792 699640 875848
rect 699696 875792 699764 875848
rect 699820 875792 699888 875848
rect 699944 875792 700012 875848
rect 700068 875792 700136 875848
rect 700192 875798 707870 875848
rect 707926 875798 708000 875854
rect 700192 875792 708000 875798
rect 699322 875730 708000 875792
rect 699322 875724 707870 875730
rect 699322 875668 699392 875724
rect 699448 875668 699516 875724
rect 699572 875668 699640 875724
rect 699696 875668 699764 875724
rect 699820 875668 699888 875724
rect 699944 875668 700012 875724
rect 700068 875668 700136 875724
rect 700192 875674 707870 875724
rect 707926 875674 708000 875730
rect 700192 875668 708000 875674
rect 699322 875606 708000 875668
rect 699322 875600 707870 875606
rect 699322 875544 699392 875600
rect 699448 875544 699516 875600
rect 699572 875544 699640 875600
rect 699696 875544 699764 875600
rect 699820 875544 699888 875600
rect 699944 875544 700012 875600
rect 700068 875544 700136 875600
rect 700192 875550 707870 875600
rect 707926 875550 708000 875606
rect 700192 875544 708000 875550
rect 699322 875482 708000 875544
rect 699322 875476 707870 875482
rect 699322 875420 699392 875476
rect 699448 875420 699516 875476
rect 699572 875420 699640 875476
rect 699696 875420 699764 875476
rect 699820 875420 699888 875476
rect 699944 875420 700012 875476
rect 700068 875420 700136 875476
rect 700192 875426 707870 875476
rect 707926 875426 708000 875482
rect 700192 875420 708000 875426
rect 699322 875358 708000 875420
rect 699322 875352 707870 875358
rect 699322 875296 699392 875352
rect 699448 875296 699516 875352
rect 699572 875296 699640 875352
rect 699696 875296 699764 875352
rect 699820 875296 699888 875352
rect 699944 875296 700012 875352
rect 700068 875296 700136 875352
rect 700192 875302 707870 875352
rect 707926 875302 708000 875358
rect 700192 875296 708000 875302
rect 699322 875234 708000 875296
rect 699322 875228 707870 875234
rect 699322 875172 699392 875228
rect 699448 875172 699516 875228
rect 699572 875172 699640 875228
rect 699696 875172 699764 875228
rect 699820 875172 699888 875228
rect 699944 875172 700012 875228
rect 700068 875172 700136 875228
rect 700192 875178 707870 875228
rect 707926 875178 708000 875234
rect 700192 875172 708000 875178
rect 699322 875110 708000 875172
rect 699322 875104 707870 875110
rect 699322 875048 699392 875104
rect 699448 875048 699516 875104
rect 699572 875048 699640 875104
rect 699696 875048 699764 875104
rect 699820 875048 699888 875104
rect 699944 875048 700012 875104
rect 700068 875048 700136 875104
rect 700192 875054 707870 875104
rect 707926 875054 708000 875110
rect 700192 875048 708000 875054
rect 699322 874986 708000 875048
rect 699322 874980 707870 874986
rect 699322 874924 699392 874980
rect 699448 874924 699516 874980
rect 699572 874924 699640 874980
rect 699696 874924 699764 874980
rect 699820 874924 699888 874980
rect 699944 874924 700012 874980
rect 700068 874924 700136 874980
rect 700192 874930 707870 874980
rect 707926 874930 708000 874986
rect 700192 874924 708000 874930
rect 699322 874862 708000 874924
rect 699322 874856 707870 874862
rect 70000 874744 78678 874802
rect 70000 874738 77808 874744
rect 70000 874682 70074 874738
rect 70130 874688 77808 874738
rect 77864 874688 77932 874744
rect 77988 874688 78056 874744
rect 78112 874688 78180 874744
rect 78236 874688 78304 874744
rect 78360 874688 78428 874744
rect 78484 874688 78552 874744
rect 78608 874688 78678 874744
rect 70130 874682 78678 874688
rect 70000 874620 78678 874682
rect 70000 874614 77808 874620
rect 70000 874558 70074 874614
rect 70130 874564 77808 874614
rect 77864 874564 77932 874620
rect 77988 874564 78056 874620
rect 78112 874564 78180 874620
rect 78236 874564 78304 874620
rect 78360 874564 78428 874620
rect 78484 874564 78552 874620
rect 78608 874564 78678 874620
rect 70130 874558 78678 874564
rect 70000 874496 78678 874558
rect 70000 874490 77808 874496
rect 70000 874434 70074 874490
rect 70130 874440 77808 874490
rect 77864 874440 77932 874496
rect 77988 874440 78056 874496
rect 78112 874440 78180 874496
rect 78236 874440 78304 874496
rect 78360 874440 78428 874496
rect 78484 874440 78552 874496
rect 78608 874440 78678 874496
rect 70130 874434 78678 874440
rect 70000 874372 78678 874434
rect 70000 874366 77808 874372
rect 70000 874310 70074 874366
rect 70130 874316 77808 874366
rect 77864 874316 77932 874372
rect 77988 874316 78056 874372
rect 78112 874316 78180 874372
rect 78236 874316 78304 874372
rect 78360 874316 78428 874372
rect 78484 874316 78552 874372
rect 78608 874316 78678 874372
rect 70130 874310 78678 874316
rect 70000 874248 78678 874310
rect 70000 874242 77808 874248
rect 70000 874186 70074 874242
rect 70130 874192 77808 874242
rect 77864 874192 77932 874248
rect 77988 874192 78056 874248
rect 78112 874192 78180 874248
rect 78236 874192 78304 874248
rect 78360 874192 78428 874248
rect 78484 874192 78552 874248
rect 78608 874192 78678 874248
rect 70130 874186 78678 874192
rect 70000 874124 78678 874186
rect 70000 874118 77808 874124
rect 70000 874062 70074 874118
rect 70130 874068 77808 874118
rect 77864 874068 77932 874124
rect 77988 874068 78056 874124
rect 78112 874068 78180 874124
rect 78236 874068 78304 874124
rect 78360 874068 78428 874124
rect 78484 874068 78552 874124
rect 78608 874068 78678 874124
rect 699322 874800 699392 874856
rect 699448 874800 699516 874856
rect 699572 874800 699640 874856
rect 699696 874800 699764 874856
rect 699820 874800 699888 874856
rect 699944 874800 700012 874856
rect 700068 874800 700136 874856
rect 700192 874806 707870 874856
rect 707926 874806 708000 874862
rect 700192 874800 708000 874806
rect 699322 874738 708000 874800
rect 699322 874732 707870 874738
rect 699322 874676 699392 874732
rect 699448 874676 699516 874732
rect 699572 874676 699640 874732
rect 699696 874676 699764 874732
rect 699820 874676 699888 874732
rect 699944 874676 700012 874732
rect 700068 874676 700136 874732
rect 700192 874682 707870 874732
rect 707926 874682 708000 874738
rect 700192 874676 708000 874682
rect 699322 874614 708000 874676
rect 699322 874608 707870 874614
rect 699322 874552 699392 874608
rect 699448 874552 699516 874608
rect 699572 874552 699640 874608
rect 699696 874552 699764 874608
rect 699820 874552 699888 874608
rect 699944 874552 700012 874608
rect 700068 874552 700136 874608
rect 700192 874558 707870 874608
rect 707926 874558 708000 874614
rect 700192 874552 708000 874558
rect 699322 874490 708000 874552
rect 699322 874484 707870 874490
rect 699322 874428 699392 874484
rect 699448 874428 699516 874484
rect 699572 874428 699640 874484
rect 699696 874428 699764 874484
rect 699820 874428 699888 874484
rect 699944 874428 700012 874484
rect 700068 874428 700136 874484
rect 700192 874434 707870 874484
rect 707926 874434 708000 874490
rect 700192 874428 708000 874434
rect 699322 874366 708000 874428
rect 699322 874360 707870 874366
rect 699322 874304 699392 874360
rect 699448 874304 699516 874360
rect 699572 874304 699640 874360
rect 699696 874304 699764 874360
rect 699820 874304 699888 874360
rect 699944 874304 700012 874360
rect 700068 874304 700136 874360
rect 700192 874310 707870 874360
rect 707926 874310 708000 874366
rect 700192 874304 708000 874310
rect 699322 874242 708000 874304
rect 699322 874236 707870 874242
rect 699322 874180 699392 874236
rect 699448 874180 699516 874236
rect 699572 874180 699640 874236
rect 699696 874180 699764 874236
rect 699820 874180 699888 874236
rect 699944 874180 700012 874236
rect 700068 874180 700136 874236
rect 700192 874186 707870 874236
rect 707926 874186 708000 874242
rect 700192 874180 708000 874186
rect 699322 874122 708000 874180
rect 70130 874062 78678 874068
rect 70000 874000 78678 874062
rect 70000 873994 77808 874000
rect 70000 873938 70074 873994
rect 70130 873944 77808 873994
rect 77864 873944 77932 874000
rect 77988 873944 78056 874000
rect 78112 873944 78180 874000
rect 78236 873944 78304 874000
rect 78360 873944 78428 874000
rect 78484 873944 78552 874000
rect 78608 873944 78678 874000
rect 70130 873938 78678 873944
rect 70000 873876 78678 873938
rect 70000 873870 77808 873876
rect 70000 873814 70074 873870
rect 70130 873820 77808 873870
rect 77864 873820 77932 873876
rect 77988 873820 78056 873876
rect 78112 873820 78180 873876
rect 78236 873820 78304 873876
rect 78360 873820 78428 873876
rect 78484 873820 78552 873876
rect 78608 873820 78678 873876
rect 70130 873814 78678 873820
rect 70000 873752 78678 873814
rect 70000 873746 77808 873752
rect 70000 873690 70074 873746
rect 70130 873696 77808 873746
rect 77864 873696 77932 873752
rect 77988 873696 78056 873752
rect 78112 873696 78180 873752
rect 78236 873696 78304 873752
rect 78360 873696 78428 873752
rect 78484 873696 78552 873752
rect 78608 873696 78678 873752
rect 70130 873690 78678 873696
rect 70000 873628 78678 873690
rect 70000 873622 77808 873628
rect 70000 873566 70074 873622
rect 70130 873572 77808 873622
rect 77864 873572 77932 873628
rect 77988 873572 78056 873628
rect 78112 873572 78180 873628
rect 78236 873572 78304 873628
rect 78360 873572 78428 873628
rect 78484 873572 78552 873628
rect 78608 873572 78678 873628
rect 70130 873566 78678 873572
rect 70000 873504 78678 873566
rect 70000 873498 77808 873504
rect 70000 873442 70074 873498
rect 70130 873448 77808 873498
rect 77864 873448 77932 873504
rect 77988 873448 78056 873504
rect 78112 873448 78180 873504
rect 78236 873448 78304 873504
rect 78360 873448 78428 873504
rect 78484 873448 78552 873504
rect 78608 873448 78678 873504
rect 70130 873442 78678 873448
rect 70000 873380 78678 873442
rect 70000 873374 77808 873380
rect 70000 873318 70074 873374
rect 70130 873324 77808 873374
rect 77864 873324 77932 873380
rect 77988 873324 78056 873380
rect 78112 873324 78180 873380
rect 78236 873324 78304 873380
rect 78360 873324 78428 873380
rect 78484 873324 78552 873380
rect 78608 873324 78678 873380
rect 70130 873318 78678 873324
rect 70000 873256 78678 873318
rect 70000 873250 77808 873256
rect 70000 873194 70074 873250
rect 70130 873200 77808 873250
rect 77864 873200 77932 873256
rect 77988 873200 78056 873256
rect 78112 873200 78180 873256
rect 78236 873200 78304 873256
rect 78360 873200 78428 873256
rect 78484 873200 78552 873256
rect 78608 873200 78678 873256
rect 70130 873194 78678 873200
rect 70000 873132 78678 873194
rect 70000 873126 77808 873132
rect 70000 873070 70074 873126
rect 70130 873076 77808 873126
rect 77864 873076 77932 873132
rect 77988 873076 78056 873132
rect 78112 873076 78180 873132
rect 78236 873076 78304 873132
rect 78360 873076 78428 873132
rect 78484 873076 78552 873132
rect 78608 873076 78678 873132
rect 70130 873070 78678 873076
rect 70000 873008 78678 873070
rect 70000 873002 77808 873008
rect 70000 872946 70074 873002
rect 70130 872952 77808 873002
rect 77864 872952 77932 873008
rect 77988 872952 78056 873008
rect 78112 872952 78180 873008
rect 78236 872952 78304 873008
rect 78360 872952 78428 873008
rect 78484 872952 78552 873008
rect 78608 872952 78678 873008
rect 70130 872946 78678 872952
rect 70000 872884 78678 872946
rect 70000 872878 77808 872884
rect 70000 872822 70074 872878
rect 70130 872828 77808 872878
rect 77864 872828 77932 872884
rect 77988 872828 78056 872884
rect 78112 872828 78180 872884
rect 78236 872828 78304 872884
rect 78360 872828 78428 872884
rect 78484 872828 78552 872884
rect 78608 872828 78678 872884
rect 70130 872822 78678 872828
rect 70000 872752 78678 872822
rect 699322 873732 708000 873802
rect 699322 873726 707870 873732
rect 699322 873670 699392 873726
rect 699448 873670 699516 873726
rect 699572 873670 699640 873726
rect 699696 873670 699764 873726
rect 699820 873670 699888 873726
rect 699944 873670 700012 873726
rect 700068 873670 700136 873726
rect 700192 873676 707870 873726
rect 707926 873676 708000 873732
rect 700192 873670 708000 873676
rect 699322 873608 708000 873670
rect 699322 873602 707870 873608
rect 699322 873546 699392 873602
rect 699448 873546 699516 873602
rect 699572 873546 699640 873602
rect 699696 873546 699764 873602
rect 699820 873546 699888 873602
rect 699944 873546 700012 873602
rect 700068 873546 700136 873602
rect 700192 873552 707870 873602
rect 707926 873552 708000 873608
rect 700192 873546 708000 873552
rect 699322 873484 708000 873546
rect 699322 873478 707870 873484
rect 699322 873422 699392 873478
rect 699448 873422 699516 873478
rect 699572 873422 699640 873478
rect 699696 873422 699764 873478
rect 699820 873422 699888 873478
rect 699944 873422 700012 873478
rect 700068 873422 700136 873478
rect 700192 873428 707870 873478
rect 707926 873428 708000 873484
rect 700192 873422 708000 873428
rect 699322 873360 708000 873422
rect 699322 873354 707870 873360
rect 699322 873298 699392 873354
rect 699448 873298 699516 873354
rect 699572 873298 699640 873354
rect 699696 873298 699764 873354
rect 699820 873298 699888 873354
rect 699944 873298 700012 873354
rect 700068 873298 700136 873354
rect 700192 873304 707870 873354
rect 707926 873304 708000 873360
rect 700192 873298 708000 873304
rect 699322 873236 708000 873298
rect 699322 873230 707870 873236
rect 699322 873174 699392 873230
rect 699448 873174 699516 873230
rect 699572 873174 699640 873230
rect 699696 873174 699764 873230
rect 699820 873174 699888 873230
rect 699944 873174 700012 873230
rect 700068 873174 700136 873230
rect 700192 873180 707870 873230
rect 707926 873180 708000 873236
rect 700192 873174 708000 873180
rect 699322 873112 708000 873174
rect 699322 873106 707870 873112
rect 699322 873050 699392 873106
rect 699448 873050 699516 873106
rect 699572 873050 699640 873106
rect 699696 873050 699764 873106
rect 699820 873050 699888 873106
rect 699944 873050 700012 873106
rect 700068 873050 700136 873106
rect 700192 873056 707870 873106
rect 707926 873056 708000 873112
rect 700192 873050 708000 873056
rect 699322 872988 708000 873050
rect 699322 872982 707870 872988
rect 699322 872926 699392 872982
rect 699448 872926 699516 872982
rect 699572 872926 699640 872982
rect 699696 872926 699764 872982
rect 699820 872926 699888 872982
rect 699944 872926 700012 872982
rect 700068 872926 700136 872982
rect 700192 872932 707870 872982
rect 707926 872932 708000 872988
rect 700192 872926 708000 872932
rect 699322 872864 708000 872926
rect 699322 872858 707870 872864
rect 699322 872802 699392 872858
rect 699448 872802 699516 872858
rect 699572 872802 699640 872858
rect 699696 872802 699764 872858
rect 699820 872802 699888 872858
rect 699944 872802 700012 872858
rect 700068 872802 700136 872858
rect 700192 872808 707870 872858
rect 707926 872808 708000 872864
rect 700192 872802 708000 872808
rect 699322 872740 708000 872802
rect 699322 872734 707870 872740
rect 699322 872678 699392 872734
rect 699448 872678 699516 872734
rect 699572 872678 699640 872734
rect 699696 872678 699764 872734
rect 699820 872678 699888 872734
rect 699944 872678 700012 872734
rect 700068 872678 700136 872734
rect 700192 872684 707870 872734
rect 707926 872684 708000 872740
rect 700192 872678 708000 872684
rect 699322 872616 708000 872678
rect 699322 872610 707870 872616
rect 699322 872554 699392 872610
rect 699448 872554 699516 872610
rect 699572 872554 699640 872610
rect 699696 872554 699764 872610
rect 699820 872554 699888 872610
rect 699944 872554 700012 872610
rect 700068 872554 700136 872610
rect 700192 872560 707870 872610
rect 707926 872560 708000 872616
rect 700192 872554 708000 872560
rect 699322 872492 708000 872554
rect 699322 872486 707870 872492
rect 699322 872430 699392 872486
rect 699448 872430 699516 872486
rect 699572 872430 699640 872486
rect 699696 872430 699764 872486
rect 699820 872430 699888 872486
rect 699944 872430 700012 872486
rect 700068 872430 700136 872486
rect 700192 872436 707870 872486
rect 707926 872436 708000 872492
rect 700192 872430 708000 872436
rect 699322 872368 708000 872430
rect 699322 872362 707870 872368
rect 699322 872306 699392 872362
rect 699448 872306 699516 872362
rect 699572 872306 699640 872362
rect 699696 872306 699764 872362
rect 699820 872306 699888 872362
rect 699944 872306 700012 872362
rect 700068 872306 700136 872362
rect 700192 872312 707870 872362
rect 707926 872312 708000 872368
rect 700192 872306 708000 872312
rect 699322 872244 708000 872306
rect 699322 872238 707870 872244
rect 699322 872182 699392 872238
rect 699448 872182 699516 872238
rect 699572 872182 699640 872238
rect 699696 872182 699764 872238
rect 699820 872182 699888 872238
rect 699944 872182 700012 872238
rect 700068 872182 700136 872238
rect 700192 872188 707870 872238
rect 707926 872188 708000 872244
rect 700192 872182 708000 872188
rect 70000 872140 78678 872172
rect 70000 872134 77808 872140
rect 70000 872078 70074 872134
rect 70130 872084 77808 872134
rect 77864 872084 77932 872140
rect 77988 872084 78056 872140
rect 78112 872084 78180 872140
rect 78236 872084 78304 872140
rect 78360 872084 78428 872140
rect 78484 872084 78552 872140
rect 78608 872084 78678 872140
rect 70130 872078 78678 872084
rect 70000 872016 78678 872078
rect 70000 872010 77808 872016
rect 70000 871954 70074 872010
rect 70130 871960 77808 872010
rect 77864 871960 77932 872016
rect 77988 871960 78056 872016
rect 78112 871960 78180 872016
rect 78236 871960 78304 872016
rect 78360 871960 78428 872016
rect 78484 871960 78552 872016
rect 78608 871960 78678 872016
rect 70130 871954 78678 871960
rect 70000 871892 78678 871954
rect 70000 871886 77808 871892
rect 70000 871830 70074 871886
rect 70130 871836 77808 871886
rect 77864 871836 77932 871892
rect 77988 871836 78056 871892
rect 78112 871836 78180 871892
rect 78236 871836 78304 871892
rect 78360 871836 78428 871892
rect 78484 871836 78552 871892
rect 78608 871836 78678 871892
rect 70130 871830 78678 871836
rect 70000 871768 78678 871830
rect 70000 871762 77808 871768
rect 70000 871706 70074 871762
rect 70130 871712 77808 871762
rect 77864 871712 77932 871768
rect 77988 871712 78056 871768
rect 78112 871712 78180 871768
rect 78236 871712 78304 871768
rect 78360 871712 78428 871768
rect 78484 871712 78552 871768
rect 78608 871712 78678 871768
rect 699322 872120 708000 872182
rect 699322 872114 707870 872120
rect 699322 872058 699392 872114
rect 699448 872058 699516 872114
rect 699572 872058 699640 872114
rect 699696 872058 699764 872114
rect 699820 872058 699888 872114
rect 699944 872058 700012 872114
rect 700068 872058 700136 872114
rect 700192 872064 707870 872114
rect 707926 872064 708000 872120
rect 700192 872058 708000 872064
rect 699322 871996 708000 872058
rect 699322 871990 707870 871996
rect 699322 871934 699392 871990
rect 699448 871934 699516 871990
rect 699572 871934 699640 871990
rect 699696 871934 699764 871990
rect 699820 871934 699888 871990
rect 699944 871934 700012 871990
rect 700068 871934 700136 871990
rect 700192 871940 707870 871990
rect 707926 871940 708000 871996
rect 700192 871934 708000 871940
rect 699322 871872 708000 871934
rect 699322 871866 707870 871872
rect 699322 871810 699392 871866
rect 699448 871810 699516 871866
rect 699572 871810 699640 871866
rect 699696 871810 699764 871866
rect 699820 871810 699888 871866
rect 699944 871810 700012 871866
rect 700068 871810 700136 871866
rect 700192 871816 707870 871866
rect 707926 871816 708000 871872
rect 700192 871810 708000 871816
rect 699322 871752 708000 871810
rect 70130 871706 78678 871712
rect 70000 871644 78678 871706
rect 70000 871638 77808 871644
rect 70000 871582 70074 871638
rect 70130 871588 77808 871638
rect 77864 871588 77932 871644
rect 77988 871588 78056 871644
rect 78112 871588 78180 871644
rect 78236 871588 78304 871644
rect 78360 871588 78428 871644
rect 78484 871588 78552 871644
rect 78608 871588 78678 871644
rect 70130 871582 78678 871588
rect 70000 871520 78678 871582
rect 70000 871514 77808 871520
rect 70000 871458 70074 871514
rect 70130 871464 77808 871514
rect 77864 871464 77932 871520
rect 77988 871464 78056 871520
rect 78112 871464 78180 871520
rect 78236 871464 78304 871520
rect 78360 871464 78428 871520
rect 78484 871464 78552 871520
rect 78608 871464 78678 871520
rect 70130 871458 78678 871464
rect 70000 871396 78678 871458
rect 70000 871390 77808 871396
rect 70000 871334 70074 871390
rect 70130 871340 77808 871390
rect 77864 871340 77932 871396
rect 77988 871340 78056 871396
rect 78112 871340 78180 871396
rect 78236 871340 78304 871396
rect 78360 871340 78428 871396
rect 78484 871340 78552 871396
rect 78608 871340 78678 871396
rect 70130 871334 78678 871340
rect 70000 871272 78678 871334
rect 70000 871266 77808 871272
rect 70000 871210 70074 871266
rect 70130 871216 77808 871266
rect 77864 871216 77932 871272
rect 77988 871216 78056 871272
rect 78112 871216 78180 871272
rect 78236 871216 78304 871272
rect 78360 871216 78428 871272
rect 78484 871216 78552 871272
rect 78608 871216 78678 871272
rect 70130 871210 78678 871216
rect 70000 871148 78678 871210
rect 70000 871142 77808 871148
rect 70000 871086 70074 871142
rect 70130 871092 77808 871142
rect 77864 871092 77932 871148
rect 77988 871092 78056 871148
rect 78112 871092 78180 871148
rect 78236 871092 78304 871148
rect 78360 871092 78428 871148
rect 78484 871092 78552 871148
rect 78608 871092 78678 871148
rect 70130 871086 78678 871092
rect 70000 871024 78678 871086
rect 70000 871018 77808 871024
rect 70000 870962 70074 871018
rect 70130 870968 77808 871018
rect 77864 870968 77932 871024
rect 77988 870968 78056 871024
rect 78112 870968 78180 871024
rect 78236 870968 78304 871024
rect 78360 870968 78428 871024
rect 78484 870968 78552 871024
rect 78608 870968 78678 871024
rect 70130 870962 78678 870968
rect 70000 870900 78678 870962
rect 70000 870894 77808 870900
rect 70000 870838 70074 870894
rect 70130 870844 77808 870894
rect 77864 870844 77932 870900
rect 77988 870844 78056 870900
rect 78112 870844 78180 870900
rect 78236 870844 78304 870900
rect 78360 870844 78428 870900
rect 78484 870844 78552 870900
rect 78608 870844 78678 870900
rect 70130 870838 78678 870844
rect 70000 870776 78678 870838
rect 70000 870770 77808 870776
rect 70000 870714 70074 870770
rect 70130 870720 77808 870770
rect 77864 870720 77932 870776
rect 77988 870720 78056 870776
rect 78112 870720 78180 870776
rect 78236 870720 78304 870776
rect 78360 870720 78428 870776
rect 78484 870720 78552 870776
rect 78608 870720 78678 870776
rect 70130 870714 78678 870720
rect 70000 870652 78678 870714
rect 70000 870646 77808 870652
rect 70000 870590 70074 870646
rect 70130 870596 77808 870646
rect 77864 870596 77932 870652
rect 77988 870596 78056 870652
rect 78112 870596 78180 870652
rect 78236 870596 78304 870652
rect 78360 870596 78428 870652
rect 78484 870596 78552 870652
rect 78608 870596 78678 870652
rect 70130 870590 78678 870596
rect 70000 870528 78678 870590
rect 70000 870522 77808 870528
rect 70000 870466 70074 870522
rect 70130 870472 77808 870522
rect 77864 870472 77932 870528
rect 77988 870472 78056 870528
rect 78112 870472 78180 870528
rect 78236 870472 78304 870528
rect 78360 870472 78428 870528
rect 78484 870472 78552 870528
rect 78608 870472 78678 870528
rect 70130 870466 78678 870472
rect 70000 870404 78678 870466
rect 70000 870398 77808 870404
rect 70000 870342 70074 870398
rect 70130 870348 77808 870398
rect 77864 870348 77932 870404
rect 77988 870348 78056 870404
rect 78112 870348 78180 870404
rect 78236 870348 78304 870404
rect 78360 870348 78428 870404
rect 78484 870348 78552 870404
rect 78608 870348 78678 870404
rect 70130 870342 78678 870348
rect 70000 870272 78678 870342
rect 699322 871134 708000 871172
rect 699322 871122 707870 871134
rect 699322 871066 699392 871122
rect 699448 871066 699516 871122
rect 699572 871066 699640 871122
rect 699696 871066 699764 871122
rect 699820 871066 699888 871122
rect 699944 871066 700012 871122
rect 700068 871066 700136 871122
rect 700192 871078 707870 871122
rect 707926 871078 708000 871134
rect 700192 871066 708000 871078
rect 699322 871010 708000 871066
rect 699322 870998 707870 871010
rect 699322 870942 699392 870998
rect 699448 870942 699516 870998
rect 699572 870942 699640 870998
rect 699696 870942 699764 870998
rect 699820 870942 699888 870998
rect 699944 870942 700012 870998
rect 700068 870942 700136 870998
rect 700192 870954 707870 870998
rect 707926 870954 708000 871010
rect 700192 870942 708000 870954
rect 699322 870886 708000 870942
rect 699322 870874 707870 870886
rect 699322 870818 699392 870874
rect 699448 870818 699516 870874
rect 699572 870818 699640 870874
rect 699696 870818 699764 870874
rect 699820 870818 699888 870874
rect 699944 870818 700012 870874
rect 700068 870818 700136 870874
rect 700192 870830 707870 870874
rect 707926 870830 708000 870886
rect 700192 870818 708000 870830
rect 699322 870762 708000 870818
rect 699322 870750 707870 870762
rect 699322 870694 699392 870750
rect 699448 870694 699516 870750
rect 699572 870694 699640 870750
rect 699696 870694 699764 870750
rect 699820 870694 699888 870750
rect 699944 870694 700012 870750
rect 700068 870694 700136 870750
rect 700192 870706 707870 870750
rect 707926 870706 708000 870762
rect 700192 870694 708000 870706
rect 699322 870638 708000 870694
rect 699322 870626 707870 870638
rect 699322 870570 699392 870626
rect 699448 870570 699516 870626
rect 699572 870570 699640 870626
rect 699696 870570 699764 870626
rect 699820 870570 699888 870626
rect 699944 870570 700012 870626
rect 700068 870570 700136 870626
rect 700192 870582 707870 870626
rect 707926 870582 708000 870638
rect 700192 870570 708000 870582
rect 699322 870514 708000 870570
rect 699322 870502 707870 870514
rect 699322 870446 699392 870502
rect 699448 870446 699516 870502
rect 699572 870446 699640 870502
rect 699696 870446 699764 870502
rect 699820 870446 699888 870502
rect 699944 870446 700012 870502
rect 700068 870446 700136 870502
rect 700192 870458 707870 870502
rect 707926 870458 708000 870514
rect 700192 870446 708000 870458
rect 699322 870390 708000 870446
rect 699322 870378 707870 870390
rect 699322 870322 699392 870378
rect 699448 870322 699516 870378
rect 699572 870322 699640 870378
rect 699696 870322 699764 870378
rect 699820 870322 699888 870378
rect 699944 870322 700012 870378
rect 700068 870322 700136 870378
rect 700192 870334 707870 870378
rect 707926 870334 708000 870390
rect 700192 870322 708000 870334
rect 699322 870266 708000 870322
rect 699322 870254 707870 870266
rect 699322 870198 699392 870254
rect 699448 870198 699516 870254
rect 699572 870198 699640 870254
rect 699696 870198 699764 870254
rect 699820 870198 699888 870254
rect 699944 870198 700012 870254
rect 700068 870198 700136 870254
rect 700192 870210 707870 870254
rect 707926 870210 708000 870266
rect 700192 870198 708000 870210
rect 699322 870142 708000 870198
rect 699322 870130 707870 870142
rect 699322 870074 699392 870130
rect 699448 870074 699516 870130
rect 699572 870074 699640 870130
rect 699696 870074 699764 870130
rect 699820 870074 699888 870130
rect 699944 870074 700012 870130
rect 700068 870074 700136 870130
rect 700192 870086 707870 870130
rect 707926 870086 708000 870142
rect 700192 870074 708000 870086
rect 699322 870018 708000 870074
rect 699322 870006 707870 870018
rect 699322 869950 699392 870006
rect 699448 869950 699516 870006
rect 699572 869950 699640 870006
rect 699696 869950 699764 870006
rect 699820 869950 699888 870006
rect 699944 869950 700012 870006
rect 700068 869950 700136 870006
rect 700192 869962 707870 870006
rect 707926 869962 708000 870018
rect 700192 869950 708000 869962
rect 699322 869894 708000 869950
rect 699322 869882 707870 869894
rect 699322 869826 699392 869882
rect 699448 869826 699516 869882
rect 699572 869826 699640 869882
rect 699696 869826 699764 869882
rect 699820 869826 699888 869882
rect 699944 869826 700012 869882
rect 700068 869826 700136 869882
rect 700192 869838 707870 869882
rect 707926 869838 708000 869894
rect 700192 869826 708000 869838
rect 699322 869770 708000 869826
rect 699322 869758 707870 869770
rect 699322 869702 699392 869758
rect 699448 869702 699516 869758
rect 699572 869702 699640 869758
rect 699696 869702 699764 869758
rect 699820 869702 699888 869758
rect 699944 869702 700012 869758
rect 700068 869702 700136 869758
rect 700192 869714 707870 869758
rect 707926 869714 708000 869770
rect 700192 869702 708000 869714
rect 699322 869646 708000 869702
rect 699322 869634 707870 869646
rect 699322 869578 699392 869634
rect 699448 869578 699516 869634
rect 699572 869578 699640 869634
rect 699696 869578 699764 869634
rect 699820 869578 699888 869634
rect 699944 869578 700012 869634
rect 700068 869578 700136 869634
rect 700192 869590 707870 869634
rect 707926 869590 708000 869646
rect 700192 869578 708000 869590
rect 699322 869522 708000 869578
rect 699322 869510 707870 869522
rect 699322 869454 699392 869510
rect 699448 869454 699516 869510
rect 699572 869454 699640 869510
rect 699696 869454 699764 869510
rect 699820 869454 699888 869510
rect 699944 869454 700012 869510
rect 700068 869454 700136 869510
rect 700192 869466 707870 869510
rect 707926 869466 708000 869522
rect 700192 869454 708000 869466
rect 699322 869398 708000 869454
rect 699322 869386 707870 869398
rect 699322 869330 699392 869386
rect 699448 869330 699516 869386
rect 699572 869330 699640 869386
rect 699696 869330 699764 869386
rect 699820 869330 699888 869386
rect 699944 869330 700012 869386
rect 700068 869330 700136 869386
rect 700192 869342 707870 869386
rect 707926 869342 708000 869398
rect 700192 869330 708000 869342
rect 699322 869272 708000 869330
rect 79078 860429 83556 860630
rect 79078 860373 79200 860429
rect 79256 860373 79500 860429
rect 79556 860373 79800 860429
rect 79856 860373 83556 860429
rect 79078 860229 83556 860373
rect 79078 860173 79200 860229
rect 79256 860173 79500 860229
rect 79556 860173 79800 860229
rect 79856 860173 83556 860229
rect 79078 860010 83556 860173
rect 688372 860429 698922 860630
rect 688372 860373 698144 860429
rect 698200 860373 698444 860429
rect 698500 860373 698744 860429
rect 698800 860373 698922 860429
rect 688372 860229 698922 860373
rect 688372 860173 698144 860229
rect 698200 860173 698444 860229
rect 698500 860173 698744 860229
rect 698800 860173 698922 860229
rect 688372 860010 698922 860173
rect 70000 843670 78678 843728
rect 70000 843658 77808 843670
rect 70000 843602 70074 843658
rect 70130 843614 77808 843658
rect 77864 843614 77932 843670
rect 77988 843614 78056 843670
rect 78112 843614 78180 843670
rect 78236 843614 78304 843670
rect 78360 843614 78428 843670
rect 78484 843614 78552 843670
rect 78608 843614 78678 843670
rect 70130 843602 78678 843614
rect 70000 843546 78678 843602
rect 70000 843534 77808 843546
rect 70000 843478 70074 843534
rect 70130 843490 77808 843534
rect 77864 843490 77932 843546
rect 77988 843490 78056 843546
rect 78112 843490 78180 843546
rect 78236 843490 78304 843546
rect 78360 843490 78428 843546
rect 78484 843490 78552 843546
rect 78608 843490 78678 843546
rect 70130 843478 78678 843490
rect 70000 843422 78678 843478
rect 70000 843410 77808 843422
rect 70000 843354 70074 843410
rect 70130 843366 77808 843410
rect 77864 843366 77932 843422
rect 77988 843366 78056 843422
rect 78112 843366 78180 843422
rect 78236 843366 78304 843422
rect 78360 843366 78428 843422
rect 78484 843366 78552 843422
rect 78608 843366 78678 843422
rect 70130 843354 78678 843366
rect 70000 843298 78678 843354
rect 70000 843286 77808 843298
rect 70000 843230 70074 843286
rect 70130 843242 77808 843286
rect 77864 843242 77932 843298
rect 77988 843242 78056 843298
rect 78112 843242 78180 843298
rect 78236 843242 78304 843298
rect 78360 843242 78428 843298
rect 78484 843242 78552 843298
rect 78608 843242 78678 843298
rect 70130 843230 78678 843242
rect 70000 843174 78678 843230
rect 70000 843162 77808 843174
rect 70000 843106 70074 843162
rect 70130 843118 77808 843162
rect 77864 843118 77932 843174
rect 77988 843118 78056 843174
rect 78112 843118 78180 843174
rect 78236 843118 78304 843174
rect 78360 843118 78428 843174
rect 78484 843118 78552 843174
rect 78608 843118 78678 843174
rect 70130 843106 78678 843118
rect 70000 843050 78678 843106
rect 70000 843038 77808 843050
rect 70000 842982 70074 843038
rect 70130 842994 77808 843038
rect 77864 842994 77932 843050
rect 77988 842994 78056 843050
rect 78112 842994 78180 843050
rect 78236 842994 78304 843050
rect 78360 842994 78428 843050
rect 78484 842994 78552 843050
rect 78608 842994 78678 843050
rect 70130 842982 78678 842994
rect 70000 842926 78678 842982
rect 70000 842914 77808 842926
rect 70000 842858 70074 842914
rect 70130 842870 77808 842914
rect 77864 842870 77932 842926
rect 77988 842870 78056 842926
rect 78112 842870 78180 842926
rect 78236 842870 78304 842926
rect 78360 842870 78428 842926
rect 78484 842870 78552 842926
rect 78608 842870 78678 842926
rect 70130 842858 78678 842870
rect 70000 842802 78678 842858
rect 70000 842790 77808 842802
rect 70000 842734 70074 842790
rect 70130 842746 77808 842790
rect 77864 842746 77932 842802
rect 77988 842746 78056 842802
rect 78112 842746 78180 842802
rect 78236 842746 78304 842802
rect 78360 842746 78428 842802
rect 78484 842746 78552 842802
rect 78608 842746 78678 842802
rect 70130 842734 78678 842746
rect 70000 842678 78678 842734
rect 70000 842666 77808 842678
rect 70000 842610 70074 842666
rect 70130 842622 77808 842666
rect 77864 842622 77932 842678
rect 77988 842622 78056 842678
rect 78112 842622 78180 842678
rect 78236 842622 78304 842678
rect 78360 842622 78428 842678
rect 78484 842622 78552 842678
rect 78608 842630 78678 842678
rect 78608 842622 84516 842630
rect 70130 842610 84516 842622
rect 70000 842554 84516 842610
rect 70000 842542 77808 842554
rect 70000 842486 70074 842542
rect 70130 842498 77808 842542
rect 77864 842498 77932 842554
rect 77988 842498 78056 842554
rect 78112 842498 78180 842554
rect 78236 842498 78304 842554
rect 78360 842498 78428 842554
rect 78484 842498 78552 842554
rect 78608 842498 84516 842554
rect 70130 842486 84516 842498
rect 70000 842430 84516 842486
rect 70000 842418 77808 842430
rect 70000 842362 70074 842418
rect 70130 842374 77808 842418
rect 77864 842374 77932 842430
rect 77988 842374 78056 842430
rect 78112 842374 78180 842430
rect 78236 842374 78304 842430
rect 78360 842374 78428 842430
rect 78484 842374 78552 842430
rect 78608 842374 84516 842430
rect 70130 842362 84516 842374
rect 70000 842306 84516 842362
rect 70000 842294 77808 842306
rect 70000 842238 70074 842294
rect 70130 842250 77808 842294
rect 77864 842250 77932 842306
rect 77988 842250 78056 842306
rect 78112 842250 78180 842306
rect 78236 842250 78304 842306
rect 78360 842250 78428 842306
rect 78484 842250 78552 842306
rect 78608 842250 84516 842306
rect 70130 842238 84516 842250
rect 70000 842182 84516 842238
rect 70000 842170 77808 842182
rect 70000 842114 70074 842170
rect 70130 842126 77808 842170
rect 77864 842126 77932 842182
rect 77988 842126 78056 842182
rect 78112 842126 78180 842182
rect 78236 842126 78304 842182
rect 78360 842126 78428 842182
rect 78484 842126 78552 842182
rect 78608 842126 84516 842182
rect 70130 842114 84516 842126
rect 70000 842058 84516 842114
rect 70000 842046 77808 842058
rect 70000 841990 70074 842046
rect 70130 842002 77808 842046
rect 77864 842002 77932 842058
rect 77988 842002 78056 842058
rect 78112 842002 78180 842058
rect 78236 842002 78304 842058
rect 78360 842002 78428 842058
rect 78484 842002 78552 842058
rect 78608 842010 84516 842058
rect 687412 842429 700322 842630
rect 687412 842373 699544 842429
rect 699600 842373 699844 842429
rect 699900 842373 700144 842429
rect 700200 842373 700322 842429
rect 687412 842229 700322 842373
rect 687412 842173 699544 842229
rect 699600 842173 699844 842229
rect 699900 842173 700144 842229
rect 700200 842173 700322 842229
rect 687412 842010 700322 842173
rect 78608 842002 78678 842010
rect 70130 841990 78678 842002
rect 70000 841934 78678 841990
rect 70000 841922 77808 841934
rect 70000 841866 70074 841922
rect 70130 841878 77808 841922
rect 77864 841878 77932 841934
rect 77988 841878 78056 841934
rect 78112 841878 78180 841934
rect 78236 841878 78304 841934
rect 78360 841878 78428 841934
rect 78484 841878 78552 841934
rect 78608 841878 78678 841934
rect 70130 841866 78678 841878
rect 70000 841828 78678 841866
rect 70000 841190 78678 841248
rect 70000 841184 77808 841190
rect 70000 841128 70074 841184
rect 70130 841134 77808 841184
rect 77864 841134 77932 841190
rect 77988 841134 78056 841190
rect 78112 841134 78180 841190
rect 78236 841134 78304 841190
rect 78360 841134 78428 841190
rect 78484 841134 78552 841190
rect 78608 841134 78678 841190
rect 70130 841128 78678 841134
rect 70000 841066 78678 841128
rect 70000 841060 77808 841066
rect 70000 841004 70074 841060
rect 70130 841010 77808 841060
rect 77864 841010 77932 841066
rect 77988 841010 78056 841066
rect 78112 841010 78180 841066
rect 78236 841010 78304 841066
rect 78360 841010 78428 841066
rect 78484 841010 78552 841066
rect 78608 841010 78678 841066
rect 70130 841004 78678 841010
rect 70000 840942 78678 841004
rect 70000 840936 77808 840942
rect 70000 840880 70074 840936
rect 70130 840886 77808 840936
rect 77864 840886 77932 840942
rect 77988 840886 78056 840942
rect 78112 840886 78180 840942
rect 78236 840886 78304 840942
rect 78360 840886 78428 840942
rect 78484 840886 78552 840942
rect 78608 840886 78678 840942
rect 70130 840880 78678 840886
rect 70000 840818 78678 840880
rect 70000 840812 77808 840818
rect 70000 840756 70074 840812
rect 70130 840762 77808 840812
rect 77864 840762 77932 840818
rect 77988 840762 78056 840818
rect 78112 840762 78180 840818
rect 78236 840762 78304 840818
rect 78360 840762 78428 840818
rect 78484 840762 78552 840818
rect 78608 840762 78678 840818
rect 70130 840756 78678 840762
rect 70000 840694 78678 840756
rect 70000 840688 77808 840694
rect 70000 840632 70074 840688
rect 70130 840638 77808 840688
rect 77864 840638 77932 840694
rect 77988 840638 78056 840694
rect 78112 840638 78180 840694
rect 78236 840638 78304 840694
rect 78360 840638 78428 840694
rect 78484 840638 78552 840694
rect 78608 840638 78678 840694
rect 70130 840632 78678 840638
rect 70000 840570 78678 840632
rect 70000 840564 77808 840570
rect 70000 840508 70074 840564
rect 70130 840514 77808 840564
rect 77864 840514 77932 840570
rect 77988 840514 78056 840570
rect 78112 840514 78180 840570
rect 78236 840514 78304 840570
rect 78360 840514 78428 840570
rect 78484 840514 78552 840570
rect 78608 840514 78678 840570
rect 70130 840508 78678 840514
rect 70000 840446 78678 840508
rect 70000 840440 77808 840446
rect 70000 840384 70074 840440
rect 70130 840390 77808 840440
rect 77864 840390 77932 840446
rect 77988 840390 78056 840446
rect 78112 840390 78180 840446
rect 78236 840390 78304 840446
rect 78360 840390 78428 840446
rect 78484 840390 78552 840446
rect 78608 840390 78678 840446
rect 70130 840384 78678 840390
rect 70000 840322 78678 840384
rect 70000 840316 77808 840322
rect 70000 840260 70074 840316
rect 70130 840266 77808 840316
rect 77864 840266 77932 840322
rect 77988 840266 78056 840322
rect 78112 840266 78180 840322
rect 78236 840266 78304 840322
rect 78360 840266 78428 840322
rect 78484 840266 78552 840322
rect 78608 840266 78678 840322
rect 70130 840260 78678 840266
rect 70000 840198 78678 840260
rect 70000 840192 77808 840198
rect 70000 840136 70074 840192
rect 70130 840142 77808 840192
rect 77864 840142 77932 840198
rect 77988 840142 78056 840198
rect 78112 840142 78180 840198
rect 78236 840142 78304 840198
rect 78360 840142 78428 840198
rect 78484 840142 78552 840198
rect 78608 840142 78678 840198
rect 70130 840136 78678 840142
rect 70000 840074 78678 840136
rect 70000 840068 77808 840074
rect 70000 840012 70074 840068
rect 70130 840018 77808 840068
rect 77864 840018 77932 840074
rect 77988 840018 78056 840074
rect 78112 840018 78180 840074
rect 78236 840018 78304 840074
rect 78360 840018 78428 840074
rect 78484 840018 78552 840074
rect 78608 840018 78678 840074
rect 70130 840012 78678 840018
rect 70000 839950 78678 840012
rect 70000 839944 77808 839950
rect 70000 839888 70074 839944
rect 70130 839894 77808 839944
rect 77864 839894 77932 839950
rect 77988 839894 78056 839950
rect 78112 839894 78180 839950
rect 78236 839894 78304 839950
rect 78360 839894 78428 839950
rect 78484 839894 78552 839950
rect 78608 839894 78678 839950
rect 70130 839888 78678 839894
rect 70000 839826 78678 839888
rect 70000 839820 77808 839826
rect 70000 839764 70074 839820
rect 70130 839770 77808 839820
rect 77864 839770 77932 839826
rect 77988 839770 78056 839826
rect 78112 839770 78180 839826
rect 78236 839770 78304 839826
rect 78360 839770 78428 839826
rect 78484 839770 78552 839826
rect 78608 839770 78678 839826
rect 70130 839764 78678 839770
rect 70000 839702 78678 839764
rect 699322 839954 702688 840076
rect 699322 839898 699444 839954
rect 699500 839898 699744 839954
rect 699800 839898 700044 839954
rect 700100 839898 702688 839954
rect 699322 839756 702688 839898
rect 70000 839696 77808 839702
rect 70000 839640 70074 839696
rect 70130 839646 77808 839696
rect 77864 839646 77932 839702
rect 77988 839646 78056 839702
rect 78112 839646 78180 839702
rect 78236 839646 78304 839702
rect 78360 839646 78428 839702
rect 78484 839646 78552 839702
rect 78608 839646 78678 839702
rect 70130 839640 78678 839646
rect 70000 839578 78678 839640
rect 70000 839572 77808 839578
rect 70000 839516 70074 839572
rect 70130 839522 77808 839572
rect 77864 839522 77932 839578
rect 77988 839522 78056 839578
rect 78112 839522 78180 839578
rect 78236 839522 78304 839578
rect 78360 839522 78428 839578
rect 78484 839522 78552 839578
rect 78608 839522 78678 839578
rect 70130 839516 78678 839522
rect 70000 839454 78678 839516
rect 70000 839448 77808 839454
rect 70000 839392 70074 839448
rect 70130 839398 77808 839448
rect 77864 839398 77932 839454
rect 77988 839398 78056 839454
rect 78112 839398 78180 839454
rect 78236 839398 78304 839454
rect 78360 839398 78428 839454
rect 78484 839398 78552 839454
rect 78608 839398 78678 839454
rect 70130 839392 78678 839398
rect 70000 839330 78678 839392
rect 70000 839324 77808 839330
rect 70000 839268 70074 839324
rect 70130 839274 77808 839324
rect 77864 839274 77932 839330
rect 77988 839274 78056 839330
rect 78112 839274 78180 839330
rect 78236 839274 78304 839330
rect 78360 839274 78428 839330
rect 78484 839274 78552 839330
rect 78608 839274 78678 839330
rect 70130 839268 78678 839274
rect 70000 839198 78678 839268
rect 70000 838820 78678 838878
rect 70000 838814 77808 838820
rect 70000 838758 70074 838814
rect 70130 838764 77808 838814
rect 77864 838764 77932 838820
rect 77988 838764 78056 838820
rect 78112 838764 78180 838820
rect 78236 838764 78304 838820
rect 78360 838764 78428 838820
rect 78484 838764 78552 838820
rect 78608 838764 78678 838820
rect 70130 838758 78678 838764
rect 70000 838696 78678 838758
rect 70000 838690 77808 838696
rect 70000 838634 70074 838690
rect 70130 838640 77808 838690
rect 77864 838640 77932 838696
rect 77988 838640 78056 838696
rect 78112 838640 78180 838696
rect 78236 838640 78304 838696
rect 78360 838640 78428 838696
rect 78484 838640 78552 838696
rect 78608 838640 78678 838696
rect 70130 838634 78678 838640
rect 70000 838572 78678 838634
rect 70000 838566 77808 838572
rect 70000 838510 70074 838566
rect 70130 838516 77808 838566
rect 77864 838516 77932 838572
rect 77988 838516 78056 838572
rect 78112 838516 78180 838572
rect 78236 838516 78304 838572
rect 78360 838516 78428 838572
rect 78484 838516 78552 838572
rect 78608 838516 78678 838572
rect 70130 838510 78678 838516
rect 70000 838448 78678 838510
rect 70000 838442 77808 838448
rect 70000 838386 70074 838442
rect 70130 838392 77808 838442
rect 77864 838392 77932 838448
rect 77988 838392 78056 838448
rect 78112 838392 78180 838448
rect 78236 838392 78304 838448
rect 78360 838392 78428 838448
rect 78484 838392 78552 838448
rect 78608 838392 78678 838448
rect 70130 838386 78678 838392
rect 70000 838324 78678 838386
rect 70000 838318 77808 838324
rect 70000 838262 70074 838318
rect 70130 838268 77808 838318
rect 77864 838268 77932 838324
rect 77988 838268 78056 838324
rect 78112 838268 78180 838324
rect 78236 838268 78304 838324
rect 78360 838268 78428 838324
rect 78484 838268 78552 838324
rect 78608 838268 78678 838324
rect 70130 838262 78678 838268
rect 70000 838200 78678 838262
rect 70000 838194 77808 838200
rect 70000 838138 70074 838194
rect 70130 838144 77808 838194
rect 77864 838144 77932 838200
rect 77988 838144 78056 838200
rect 78112 838144 78180 838200
rect 78236 838144 78304 838200
rect 78360 838144 78428 838200
rect 78484 838144 78552 838200
rect 78608 838144 78678 838200
rect 70130 838138 78678 838144
rect 70000 838076 78678 838138
rect 70000 838070 77808 838076
rect 70000 838014 70074 838070
rect 70130 838020 77808 838070
rect 77864 838020 77932 838076
rect 77988 838020 78056 838076
rect 78112 838020 78180 838076
rect 78236 838020 78304 838076
rect 78360 838020 78428 838076
rect 78484 838020 78552 838076
rect 78608 838020 78678 838076
rect 70130 838014 78678 838020
rect 70000 837952 78678 838014
rect 70000 837946 77808 837952
rect 70000 837890 70074 837946
rect 70130 837896 77808 837946
rect 77864 837896 77932 837952
rect 77988 837896 78056 837952
rect 78112 837896 78180 837952
rect 78236 837896 78304 837952
rect 78360 837896 78428 837952
rect 78484 837896 78552 837952
rect 78608 837896 78678 837952
rect 70130 837890 78678 837896
rect 70000 837828 78678 837890
rect 70000 837822 77808 837828
rect 70000 837766 70074 837822
rect 70130 837772 77808 837822
rect 77864 837772 77932 837828
rect 77988 837772 78056 837828
rect 78112 837772 78180 837828
rect 78236 837772 78304 837828
rect 78360 837772 78428 837828
rect 78484 837772 78552 837828
rect 78608 837772 78678 837828
rect 70130 837766 78678 837772
rect 70000 837704 78678 837766
rect 70000 837698 77808 837704
rect 70000 837642 70074 837698
rect 70130 837648 77808 837698
rect 77864 837648 77932 837704
rect 77988 837648 78056 837704
rect 78112 837648 78180 837704
rect 78236 837648 78304 837704
rect 78360 837648 78428 837704
rect 78484 837648 78552 837704
rect 78608 837648 78678 837704
rect 70130 837642 78678 837648
rect 70000 837580 78678 837642
rect 70000 837574 77808 837580
rect 70000 837518 70074 837574
rect 70130 837524 77808 837574
rect 77864 837524 77932 837580
rect 77988 837524 78056 837580
rect 78112 837524 78180 837580
rect 78236 837524 78304 837580
rect 78360 837524 78428 837580
rect 78484 837524 78552 837580
rect 78608 837524 78678 837580
rect 70130 837518 78678 837524
rect 70000 837456 78678 837518
rect 70000 837450 77808 837456
rect 70000 837394 70074 837450
rect 70130 837400 77808 837450
rect 77864 837400 77932 837456
rect 77988 837400 78056 837456
rect 78112 837400 78180 837456
rect 78236 837400 78304 837456
rect 78360 837400 78428 837456
rect 78484 837400 78552 837456
rect 78608 837400 78678 837456
rect 70130 837394 78678 837400
rect 70000 837332 78678 837394
rect 70000 837326 77808 837332
rect 70000 837270 70074 837326
rect 70130 837276 77808 837326
rect 77864 837276 77932 837332
rect 77988 837276 78056 837332
rect 78112 837276 78180 837332
rect 78236 837276 78304 837332
rect 78360 837276 78428 837332
rect 78484 837276 78552 837332
rect 78608 837276 78678 837332
rect 70130 837270 78678 837276
rect 70000 837208 78678 837270
rect 70000 837202 77808 837208
rect 70000 837146 70074 837202
rect 70130 837152 77808 837202
rect 77864 837152 77932 837208
rect 77988 837152 78056 837208
rect 78112 837152 78180 837208
rect 78236 837152 78304 837208
rect 78360 837152 78428 837208
rect 78484 837152 78552 837208
rect 78608 837152 78678 837208
rect 70130 837146 78678 837152
rect 70000 837084 78678 837146
rect 70000 837078 77808 837084
rect 70000 837022 70074 837078
rect 70130 837028 77808 837078
rect 77864 837028 77932 837084
rect 77988 837028 78056 837084
rect 78112 837028 78180 837084
rect 78236 837028 78304 837084
rect 78360 837028 78428 837084
rect 78484 837028 78552 837084
rect 78608 837028 78678 837084
rect 70130 837022 78678 837028
rect 70000 836960 78678 837022
rect 70000 836954 77808 836960
rect 70000 836898 70074 836954
rect 70130 836904 77808 836954
rect 77864 836904 77932 836960
rect 77988 836904 78056 836960
rect 78112 836904 78180 836960
rect 78236 836904 78304 836960
rect 78360 836904 78428 836960
rect 78484 836904 78552 836960
rect 78608 836904 78678 836960
rect 70130 836898 78678 836904
rect 70000 836828 78678 836898
rect 697922 836434 702624 836576
rect 697922 836378 698044 836434
rect 698100 836378 698344 836434
rect 698400 836378 698644 836434
rect 698700 836378 702624 836434
rect 697922 836256 702624 836378
rect 70000 836114 78678 836172
rect 70000 836108 77808 836114
rect 70000 836052 70074 836108
rect 70130 836058 77808 836108
rect 77864 836058 77932 836114
rect 77988 836058 78056 836114
rect 78112 836058 78180 836114
rect 78236 836058 78304 836114
rect 78360 836058 78428 836114
rect 78484 836058 78552 836114
rect 78608 836058 78678 836114
rect 70130 836052 78678 836058
rect 70000 835990 78678 836052
rect 70000 835984 77808 835990
rect 70000 835928 70074 835984
rect 70130 835934 77808 835984
rect 77864 835934 77932 835990
rect 77988 835934 78056 835990
rect 78112 835934 78180 835990
rect 78236 835934 78304 835990
rect 78360 835934 78428 835990
rect 78484 835934 78552 835990
rect 78608 835934 78678 835990
rect 70130 835928 78678 835934
rect 70000 835866 78678 835928
rect 70000 835860 77808 835866
rect 70000 835804 70074 835860
rect 70130 835810 77808 835860
rect 77864 835810 77932 835866
rect 77988 835810 78056 835866
rect 78112 835810 78180 835866
rect 78236 835810 78304 835866
rect 78360 835810 78428 835866
rect 78484 835810 78552 835866
rect 78608 835810 78678 835866
rect 70130 835804 78678 835810
rect 70000 835742 78678 835804
rect 70000 835736 77808 835742
rect 70000 835680 70074 835736
rect 70130 835686 77808 835736
rect 77864 835686 77932 835742
rect 77988 835686 78056 835742
rect 78112 835686 78180 835742
rect 78236 835686 78304 835742
rect 78360 835686 78428 835742
rect 78484 835686 78552 835742
rect 78608 835686 78678 835742
rect 70130 835680 78678 835686
rect 70000 835618 78678 835680
rect 70000 835612 77808 835618
rect 70000 835556 70074 835612
rect 70130 835562 77808 835612
rect 77864 835562 77932 835618
rect 77988 835562 78056 835618
rect 78112 835562 78180 835618
rect 78236 835562 78304 835618
rect 78360 835562 78428 835618
rect 78484 835562 78552 835618
rect 78608 835562 78678 835618
rect 70130 835556 78678 835562
rect 70000 835494 78678 835556
rect 70000 835488 77808 835494
rect 70000 835432 70074 835488
rect 70130 835438 77808 835488
rect 77864 835438 77932 835494
rect 77988 835438 78056 835494
rect 78112 835438 78180 835494
rect 78236 835438 78304 835494
rect 78360 835438 78428 835494
rect 78484 835438 78552 835494
rect 78608 835438 78678 835494
rect 70130 835432 78678 835438
rect 70000 835370 78678 835432
rect 70000 835364 77808 835370
rect 70000 835308 70074 835364
rect 70130 835314 77808 835364
rect 77864 835314 77932 835370
rect 77988 835314 78056 835370
rect 78112 835314 78180 835370
rect 78236 835314 78304 835370
rect 78360 835314 78428 835370
rect 78484 835314 78552 835370
rect 78608 835314 78678 835370
rect 70130 835308 78678 835314
rect 70000 835246 78678 835308
rect 70000 835240 77808 835246
rect 70000 835184 70074 835240
rect 70130 835190 77808 835240
rect 77864 835190 77932 835246
rect 77988 835190 78056 835246
rect 78112 835190 78180 835246
rect 78236 835190 78304 835246
rect 78360 835190 78428 835246
rect 78484 835190 78552 835246
rect 78608 835190 78678 835246
rect 70130 835184 78678 835190
rect 70000 835122 78678 835184
rect 70000 835116 77808 835122
rect 70000 835060 70074 835116
rect 70130 835066 77808 835116
rect 77864 835066 77932 835122
rect 77988 835066 78056 835122
rect 78112 835066 78180 835122
rect 78236 835066 78304 835122
rect 78360 835066 78428 835122
rect 78484 835066 78552 835122
rect 78608 835066 78678 835122
rect 70130 835060 78678 835066
rect 70000 834998 78678 835060
rect 70000 834992 77808 834998
rect 70000 834936 70074 834992
rect 70130 834942 77808 834992
rect 77864 834942 77932 834998
rect 77988 834942 78056 834998
rect 78112 834942 78180 834998
rect 78236 834942 78304 834998
rect 78360 834942 78428 834998
rect 78484 834942 78552 834998
rect 78608 834942 78678 834998
rect 70130 834936 78678 834942
rect 70000 834874 78678 834936
rect 70000 834868 77808 834874
rect 70000 834812 70074 834868
rect 70130 834818 77808 834868
rect 77864 834818 77932 834874
rect 77988 834818 78056 834874
rect 78112 834818 78180 834874
rect 78236 834818 78304 834874
rect 78360 834818 78428 834874
rect 78484 834818 78552 834874
rect 78608 834818 78678 834874
rect 70130 834812 78678 834818
rect 70000 834750 78678 834812
rect 70000 834744 77808 834750
rect 70000 834688 70074 834744
rect 70130 834694 77808 834744
rect 77864 834694 77932 834750
rect 77988 834694 78056 834750
rect 78112 834694 78180 834750
rect 78236 834694 78304 834750
rect 78360 834694 78428 834750
rect 78484 834694 78552 834750
rect 78608 834694 78678 834750
rect 70130 834688 78678 834694
rect 70000 834626 78678 834688
rect 70000 834620 77808 834626
rect 70000 834564 70074 834620
rect 70130 834570 77808 834620
rect 77864 834570 77932 834626
rect 77988 834570 78056 834626
rect 78112 834570 78180 834626
rect 78236 834570 78304 834626
rect 78360 834570 78428 834626
rect 78484 834570 78552 834626
rect 78608 834570 78678 834626
rect 70130 834564 78678 834570
rect 70000 834502 78678 834564
rect 70000 834496 77808 834502
rect 70000 834440 70074 834496
rect 70130 834446 77808 834496
rect 77864 834446 77932 834502
rect 77988 834446 78056 834502
rect 78112 834446 78180 834502
rect 78236 834446 78304 834502
rect 78360 834446 78428 834502
rect 78484 834446 78552 834502
rect 78608 834446 78678 834502
rect 70130 834440 78678 834446
rect 70000 834378 78678 834440
rect 70000 834372 77808 834378
rect 70000 834316 70074 834372
rect 70130 834322 77808 834372
rect 77864 834322 77932 834378
rect 77988 834322 78056 834378
rect 78112 834322 78180 834378
rect 78236 834322 78304 834378
rect 78360 834322 78428 834378
rect 78484 834322 78552 834378
rect 78608 834322 78678 834378
rect 70130 834316 78678 834322
rect 70000 834254 78678 834316
rect 70000 834248 77808 834254
rect 70000 834192 70074 834248
rect 70130 834198 77808 834248
rect 77864 834198 77932 834254
rect 77988 834198 78056 834254
rect 78112 834198 78180 834254
rect 78236 834198 78304 834254
rect 78360 834198 78428 834254
rect 78484 834198 78552 834254
rect 78608 834198 78678 834254
rect 70130 834192 78678 834198
rect 70000 834122 78678 834192
rect 70000 833744 78678 833802
rect 70000 833738 77808 833744
rect 70000 833682 70074 833738
rect 70130 833688 77808 833738
rect 77864 833688 77932 833744
rect 77988 833688 78056 833744
rect 78112 833688 78180 833744
rect 78236 833688 78304 833744
rect 78360 833688 78428 833744
rect 78484 833688 78552 833744
rect 78608 833688 78678 833744
rect 70130 833682 78678 833688
rect 70000 833620 78678 833682
rect 70000 833614 77808 833620
rect 70000 833558 70074 833614
rect 70130 833564 77808 833614
rect 77864 833564 77932 833620
rect 77988 833564 78056 833620
rect 78112 833564 78180 833620
rect 78236 833564 78304 833620
rect 78360 833564 78428 833620
rect 78484 833564 78552 833620
rect 78608 833564 78678 833620
rect 70130 833558 78678 833564
rect 70000 833496 78678 833558
rect 70000 833490 77808 833496
rect 70000 833434 70074 833490
rect 70130 833440 77808 833490
rect 77864 833440 77932 833496
rect 77988 833440 78056 833496
rect 78112 833440 78180 833496
rect 78236 833440 78304 833496
rect 78360 833440 78428 833496
rect 78484 833440 78552 833496
rect 78608 833440 78678 833496
rect 70130 833434 78678 833440
rect 70000 833372 78678 833434
rect 70000 833366 77808 833372
rect 70000 833310 70074 833366
rect 70130 833316 77808 833366
rect 77864 833316 77932 833372
rect 77988 833316 78056 833372
rect 78112 833316 78180 833372
rect 78236 833316 78304 833372
rect 78360 833316 78428 833372
rect 78484 833316 78552 833372
rect 78608 833316 78678 833372
rect 70130 833310 78678 833316
rect 70000 833248 78678 833310
rect 70000 833242 77808 833248
rect 70000 833186 70074 833242
rect 70130 833192 77808 833242
rect 77864 833192 77932 833248
rect 77988 833192 78056 833248
rect 78112 833192 78180 833248
rect 78236 833192 78304 833248
rect 78360 833192 78428 833248
rect 78484 833192 78552 833248
rect 78608 833192 78678 833248
rect 70130 833186 78678 833192
rect 70000 833124 78678 833186
rect 70000 833118 77808 833124
rect 70000 833062 70074 833118
rect 70130 833068 77808 833118
rect 77864 833068 77932 833124
rect 77988 833068 78056 833124
rect 78112 833068 78180 833124
rect 78236 833068 78304 833124
rect 78360 833068 78428 833124
rect 78484 833068 78552 833124
rect 78608 833068 78678 833124
rect 70130 833062 78678 833068
rect 70000 833000 78678 833062
rect 70000 832994 77808 833000
rect 70000 832938 70074 832994
rect 70130 832944 77808 832994
rect 77864 832944 77932 833000
rect 77988 832944 78056 833000
rect 78112 832944 78180 833000
rect 78236 832944 78304 833000
rect 78360 832944 78428 833000
rect 78484 832944 78552 833000
rect 78608 832944 78678 833000
rect 70130 832938 78678 832944
rect 70000 832876 78678 832938
rect 70000 832870 77808 832876
rect 70000 832814 70074 832870
rect 70130 832820 77808 832870
rect 77864 832820 77932 832876
rect 77988 832820 78056 832876
rect 78112 832820 78180 832876
rect 78236 832820 78304 832876
rect 78360 832820 78428 832876
rect 78484 832820 78552 832876
rect 78608 832820 78678 832876
rect 70130 832814 78678 832820
rect 70000 832752 78678 832814
rect 699322 832954 702688 833076
rect 699322 832898 699444 832954
rect 699500 832898 699744 832954
rect 699800 832898 700044 832954
rect 700100 832898 702688 832954
rect 699322 832756 702688 832898
rect 70000 832746 77808 832752
rect 70000 832690 70074 832746
rect 70130 832696 77808 832746
rect 77864 832696 77932 832752
rect 77988 832696 78056 832752
rect 78112 832696 78180 832752
rect 78236 832696 78304 832752
rect 78360 832696 78428 832752
rect 78484 832696 78552 832752
rect 78608 832696 78678 832752
rect 70130 832690 78678 832696
rect 70000 832628 78678 832690
rect 70000 832622 77808 832628
rect 70000 832566 70074 832622
rect 70130 832572 77808 832622
rect 77864 832572 77932 832628
rect 77988 832572 78056 832628
rect 78112 832572 78180 832628
rect 78236 832572 78304 832628
rect 78360 832572 78428 832628
rect 78484 832572 78552 832628
rect 78608 832572 78678 832628
rect 70130 832566 78678 832572
rect 70000 832504 78678 832566
rect 70000 832498 77808 832504
rect 70000 832442 70074 832498
rect 70130 832448 77808 832498
rect 77864 832448 77932 832504
rect 77988 832448 78056 832504
rect 78112 832448 78180 832504
rect 78236 832448 78304 832504
rect 78360 832448 78428 832504
rect 78484 832448 78552 832504
rect 78608 832448 78678 832504
rect 70130 832442 78678 832448
rect 70000 832380 78678 832442
rect 70000 832374 77808 832380
rect 70000 832318 70074 832374
rect 70130 832324 77808 832374
rect 77864 832324 77932 832380
rect 77988 832324 78056 832380
rect 78112 832324 78180 832380
rect 78236 832324 78304 832380
rect 78360 832324 78428 832380
rect 78484 832324 78552 832380
rect 78608 832324 78678 832380
rect 70130 832318 78678 832324
rect 70000 832256 78678 832318
rect 70000 832250 77808 832256
rect 70000 832194 70074 832250
rect 70130 832200 77808 832250
rect 77864 832200 77932 832256
rect 77988 832200 78056 832256
rect 78112 832200 78180 832256
rect 78236 832200 78304 832256
rect 78360 832200 78428 832256
rect 78484 832200 78552 832256
rect 78608 832200 78678 832256
rect 70130 832194 78678 832200
rect 70000 832132 78678 832194
rect 70000 832126 77808 832132
rect 70000 832070 70074 832126
rect 70130 832076 77808 832126
rect 77864 832076 77932 832132
rect 77988 832076 78056 832132
rect 78112 832076 78180 832132
rect 78236 832076 78304 832132
rect 78360 832076 78428 832132
rect 78484 832076 78552 832132
rect 78608 832076 78678 832132
rect 70130 832070 78678 832076
rect 70000 832008 78678 832070
rect 70000 832002 77808 832008
rect 70000 831946 70074 832002
rect 70130 831952 77808 832002
rect 77864 831952 77932 832008
rect 77988 831952 78056 832008
rect 78112 831952 78180 832008
rect 78236 831952 78304 832008
rect 78360 831952 78428 832008
rect 78484 831952 78552 832008
rect 78608 831952 78678 832008
rect 70130 831946 78678 831952
rect 70000 831884 78678 831946
rect 70000 831878 77808 831884
rect 70000 831822 70074 831878
rect 70130 831828 77808 831878
rect 77864 831828 77932 831884
rect 77988 831828 78056 831884
rect 78112 831828 78180 831884
rect 78236 831828 78304 831884
rect 78360 831828 78428 831884
rect 78484 831828 78552 831884
rect 78608 831828 78678 831884
rect 70130 831822 78678 831828
rect 70000 831752 78678 831822
rect 70000 831140 78678 831172
rect 70000 831134 77808 831140
rect 70000 831078 70074 831134
rect 70130 831084 77808 831134
rect 77864 831084 77932 831140
rect 77988 831084 78056 831140
rect 78112 831084 78180 831140
rect 78236 831084 78304 831140
rect 78360 831084 78428 831140
rect 78484 831084 78552 831140
rect 78608 831084 78678 831140
rect 70130 831078 78678 831084
rect 70000 831016 78678 831078
rect 70000 831010 77808 831016
rect 70000 830954 70074 831010
rect 70130 830960 77808 831010
rect 77864 830960 77932 831016
rect 77988 830960 78056 831016
rect 78112 830960 78180 831016
rect 78236 830960 78304 831016
rect 78360 830960 78428 831016
rect 78484 830960 78552 831016
rect 78608 830960 78678 831016
rect 70130 830954 78678 830960
rect 70000 830892 78678 830954
rect 70000 830886 77808 830892
rect 70000 830830 70074 830886
rect 70130 830836 77808 830886
rect 77864 830836 77932 830892
rect 77988 830836 78056 830892
rect 78112 830836 78180 830892
rect 78236 830836 78304 830892
rect 78360 830836 78428 830892
rect 78484 830836 78552 830892
rect 78608 830836 78678 830892
rect 70130 830830 78678 830836
rect 70000 830768 78678 830830
rect 70000 830762 77808 830768
rect 70000 830706 70074 830762
rect 70130 830712 77808 830762
rect 77864 830712 77932 830768
rect 77988 830712 78056 830768
rect 78112 830712 78180 830768
rect 78236 830712 78304 830768
rect 78360 830712 78428 830768
rect 78484 830712 78552 830768
rect 78608 830712 78678 830768
rect 70130 830706 78678 830712
rect 70000 830644 78678 830706
rect 70000 830638 77808 830644
rect 70000 830582 70074 830638
rect 70130 830588 77808 830638
rect 77864 830588 77932 830644
rect 77988 830588 78056 830644
rect 78112 830588 78180 830644
rect 78236 830588 78304 830644
rect 78360 830588 78428 830644
rect 78484 830588 78552 830644
rect 78608 830588 78678 830644
rect 70130 830582 78678 830588
rect 70000 830520 78678 830582
rect 70000 830514 77808 830520
rect 70000 830458 70074 830514
rect 70130 830464 77808 830514
rect 77864 830464 77932 830520
rect 77988 830464 78056 830520
rect 78112 830464 78180 830520
rect 78236 830464 78304 830520
rect 78360 830464 78428 830520
rect 78484 830464 78552 830520
rect 78608 830464 78678 830520
rect 70130 830458 78678 830464
rect 70000 830396 78678 830458
rect 70000 830390 77808 830396
rect 70000 830334 70074 830390
rect 70130 830340 77808 830390
rect 77864 830340 77932 830396
rect 77988 830340 78056 830396
rect 78112 830340 78180 830396
rect 78236 830340 78304 830396
rect 78360 830340 78428 830396
rect 78484 830340 78552 830396
rect 78608 830340 78678 830396
rect 70130 830334 78678 830340
rect 70000 830272 78678 830334
rect 70000 830266 77808 830272
rect 70000 830210 70074 830266
rect 70130 830216 77808 830266
rect 77864 830216 77932 830272
rect 77988 830216 78056 830272
rect 78112 830216 78180 830272
rect 78236 830216 78304 830272
rect 78360 830216 78428 830272
rect 78484 830216 78552 830272
rect 78608 830216 78678 830272
rect 70130 830210 78678 830216
rect 70000 830148 78678 830210
rect 70000 830142 77808 830148
rect 70000 830086 70074 830142
rect 70130 830092 77808 830142
rect 77864 830092 77932 830148
rect 77988 830092 78056 830148
rect 78112 830092 78180 830148
rect 78236 830092 78304 830148
rect 78360 830092 78428 830148
rect 78484 830092 78552 830148
rect 78608 830092 78678 830148
rect 70130 830086 78678 830092
rect 70000 830024 78678 830086
rect 70000 830018 77808 830024
rect 70000 829962 70074 830018
rect 70130 829968 77808 830018
rect 77864 829968 77932 830024
rect 77988 829968 78056 830024
rect 78112 829968 78180 830024
rect 78236 829968 78304 830024
rect 78360 829968 78428 830024
rect 78484 829968 78552 830024
rect 78608 829968 78678 830024
rect 70130 829962 78678 829968
rect 70000 829900 78678 829962
rect 70000 829894 77808 829900
rect 70000 829838 70074 829894
rect 70130 829844 77808 829894
rect 77864 829844 77932 829900
rect 77988 829844 78056 829900
rect 78112 829844 78180 829900
rect 78236 829844 78304 829900
rect 78360 829844 78428 829900
rect 78484 829844 78552 829900
rect 78608 829844 78678 829900
rect 70130 829838 78678 829844
rect 70000 829776 78678 829838
rect 70000 829770 77808 829776
rect 70000 829714 70074 829770
rect 70130 829720 77808 829770
rect 77864 829720 77932 829776
rect 77988 829720 78056 829776
rect 78112 829720 78180 829776
rect 78236 829720 78304 829776
rect 78360 829720 78428 829776
rect 78484 829720 78552 829776
rect 78608 829720 78678 829776
rect 70130 829714 78678 829720
rect 70000 829652 78678 829714
rect 70000 829646 77808 829652
rect 70000 829590 70074 829646
rect 70130 829596 77808 829646
rect 77864 829596 77932 829652
rect 77988 829596 78056 829652
rect 78112 829596 78180 829652
rect 78236 829596 78304 829652
rect 78360 829596 78428 829652
rect 78484 829596 78552 829652
rect 78608 829596 78678 829652
rect 70130 829590 78678 829596
rect 70000 829528 78678 829590
rect 70000 829522 77808 829528
rect 70000 829466 70074 829522
rect 70130 829472 77808 829522
rect 77864 829472 77932 829528
rect 77988 829472 78056 829528
rect 78112 829472 78180 829528
rect 78236 829472 78304 829528
rect 78360 829472 78428 829528
rect 78484 829472 78552 829528
rect 78608 829472 78678 829528
rect 70130 829466 78678 829472
rect 70000 829404 78678 829466
rect 70000 829398 77808 829404
rect 70000 829342 70074 829398
rect 70130 829348 77808 829398
rect 77864 829348 77932 829404
rect 77988 829348 78056 829404
rect 78112 829348 78180 829404
rect 78236 829348 78304 829404
rect 78360 829348 78428 829404
rect 78484 829348 78552 829404
rect 78608 829348 78678 829404
rect 70130 829342 78678 829348
rect 70000 829272 78678 829342
rect 697922 829434 702624 829576
rect 697922 829378 698044 829434
rect 698100 829378 698344 829434
rect 698400 829378 698644 829434
rect 698700 829378 702624 829434
rect 697922 829256 702624 829378
rect 699322 825954 702688 826076
rect 699322 825898 699444 825954
rect 699500 825898 699744 825954
rect 699800 825898 700044 825954
rect 700100 825898 702688 825954
rect 699322 825756 702688 825898
rect 79078 824429 83556 824630
rect 79078 824373 79200 824429
rect 79256 824373 79500 824429
rect 79556 824373 79800 824429
rect 79856 824373 83556 824429
rect 79078 824229 83556 824373
rect 79078 824173 79200 824229
rect 79256 824173 79500 824229
rect 79556 824173 79800 824229
rect 79856 824173 83556 824229
rect 79078 824010 83556 824173
rect 688372 824429 698922 824630
rect 688372 824373 698144 824429
rect 698200 824373 698444 824429
rect 698500 824373 698744 824429
rect 698800 824373 698922 824429
rect 688372 824229 698922 824373
rect 688372 824173 698144 824229
rect 698200 824173 698444 824229
rect 698500 824173 698744 824229
rect 698800 824173 698922 824229
rect 688372 824010 698922 824173
rect 697922 822434 702624 822576
rect 697922 822378 698044 822434
rect 698100 822378 698344 822434
rect 698400 822378 698644 822434
rect 698700 822378 702624 822434
rect 697922 822256 702624 822378
rect 77678 806429 84516 806630
rect 77678 806373 77800 806429
rect 77856 806373 78100 806429
rect 78156 806373 78400 806429
rect 78456 806373 84516 806429
rect 77678 806229 84516 806373
rect 699322 806423 701085 806490
rect 699322 806367 699497 806423
rect 699553 806367 699797 806423
rect 699853 806367 700097 806423
rect 700153 806367 701085 806423
rect 699322 806290 701085 806367
rect 77678 806173 77800 806229
rect 77856 806173 78100 806229
rect 78156 806173 78400 806229
rect 78456 806173 84516 806229
rect 77678 806010 84516 806173
rect 701565 806090 701885 806490
rect 697922 806008 701885 806090
rect 697922 805952 698060 806008
rect 698116 805952 698360 806008
rect 698416 805952 698660 806008
rect 698716 805952 701885 806008
rect 697922 805890 701885 805952
rect 70000 802670 80078 802728
rect 70000 802658 79208 802670
rect 70000 802602 70074 802658
rect 70130 802614 79208 802658
rect 79264 802614 79332 802670
rect 79388 802614 79456 802670
rect 79512 802614 79580 802670
rect 79636 802614 79704 802670
rect 79760 802614 79828 802670
rect 79884 802614 79952 802670
rect 80008 802614 80078 802670
rect 70130 802602 80078 802614
rect 70000 802546 80078 802602
rect 70000 802534 79208 802546
rect 70000 802478 70074 802534
rect 70130 802490 79208 802534
rect 79264 802490 79332 802546
rect 79388 802490 79456 802546
rect 79512 802490 79580 802546
rect 79636 802490 79704 802546
rect 79760 802490 79828 802546
rect 79884 802490 79952 802546
rect 80008 802490 80078 802546
rect 70130 802478 80078 802490
rect 70000 802422 80078 802478
rect 70000 802410 79208 802422
rect 70000 802354 70074 802410
rect 70130 802366 79208 802410
rect 79264 802366 79332 802422
rect 79388 802366 79456 802422
rect 79512 802366 79580 802422
rect 79636 802366 79704 802422
rect 79760 802366 79828 802422
rect 79884 802366 79952 802422
rect 80008 802366 80078 802422
rect 70130 802354 80078 802366
rect 70000 802298 80078 802354
rect 70000 802286 79208 802298
rect 70000 802230 70074 802286
rect 70130 802242 79208 802286
rect 79264 802242 79332 802298
rect 79388 802242 79456 802298
rect 79512 802242 79580 802298
rect 79636 802242 79704 802298
rect 79760 802242 79828 802298
rect 79884 802242 79952 802298
rect 80008 802242 80078 802298
rect 70130 802230 80078 802242
rect 70000 802174 80078 802230
rect 70000 802162 79208 802174
rect 70000 802106 70074 802162
rect 70130 802118 79208 802162
rect 79264 802118 79332 802174
rect 79388 802118 79456 802174
rect 79512 802118 79580 802174
rect 79636 802118 79704 802174
rect 79760 802118 79828 802174
rect 79884 802118 79952 802174
rect 80008 802118 80078 802174
rect 70130 802106 80078 802118
rect 70000 802050 80078 802106
rect 70000 802038 79208 802050
rect 70000 801982 70074 802038
rect 70130 801994 79208 802038
rect 79264 801994 79332 802050
rect 79388 801994 79456 802050
rect 79512 801994 79580 802050
rect 79636 801994 79704 802050
rect 79760 801994 79828 802050
rect 79884 801994 79952 802050
rect 80008 801994 80078 802050
rect 70130 801982 80078 801994
rect 70000 801926 80078 801982
rect 70000 801914 79208 801926
rect 70000 801858 70074 801914
rect 70130 801870 79208 801914
rect 79264 801870 79332 801926
rect 79388 801870 79456 801926
rect 79512 801870 79580 801926
rect 79636 801870 79704 801926
rect 79760 801870 79828 801926
rect 79884 801870 79952 801926
rect 80008 801870 80078 801926
rect 70130 801858 80078 801870
rect 70000 801802 80078 801858
rect 70000 801790 79208 801802
rect 70000 801734 70074 801790
rect 70130 801746 79208 801790
rect 79264 801746 79332 801802
rect 79388 801746 79456 801802
rect 79512 801746 79580 801802
rect 79636 801746 79704 801802
rect 79760 801746 79828 801802
rect 79884 801746 79952 801802
rect 80008 801746 80078 801802
rect 70130 801734 80078 801746
rect 70000 801678 80078 801734
rect 70000 801666 79208 801678
rect 70000 801610 70074 801666
rect 70130 801622 79208 801666
rect 79264 801622 79332 801678
rect 79388 801622 79456 801678
rect 79512 801622 79580 801678
rect 79636 801622 79704 801678
rect 79760 801622 79828 801678
rect 79884 801622 79952 801678
rect 80008 801622 80078 801678
rect 70130 801610 80078 801622
rect 70000 801554 80078 801610
rect 70000 801542 79208 801554
rect 70000 801486 70074 801542
rect 70130 801498 79208 801542
rect 79264 801498 79332 801554
rect 79388 801498 79456 801554
rect 79512 801498 79580 801554
rect 79636 801498 79704 801554
rect 79760 801498 79828 801554
rect 79884 801498 79952 801554
rect 80008 801498 80078 801554
rect 70130 801486 80078 801498
rect 70000 801430 80078 801486
rect 70000 801418 79208 801430
rect 70000 801362 70074 801418
rect 70130 801374 79208 801418
rect 79264 801374 79332 801430
rect 79388 801374 79456 801430
rect 79512 801374 79580 801430
rect 79636 801374 79704 801430
rect 79760 801374 79828 801430
rect 79884 801374 79952 801430
rect 80008 801374 80078 801430
rect 70130 801362 80078 801374
rect 70000 801306 80078 801362
rect 70000 801294 79208 801306
rect 70000 801238 70074 801294
rect 70130 801250 79208 801294
rect 79264 801250 79332 801306
rect 79388 801250 79456 801306
rect 79512 801250 79580 801306
rect 79636 801250 79704 801306
rect 79760 801250 79828 801306
rect 79884 801250 79952 801306
rect 80008 801250 80078 801306
rect 70130 801238 80078 801250
rect 70000 801182 80078 801238
rect 70000 801170 79208 801182
rect 70000 801114 70074 801170
rect 70130 801126 79208 801170
rect 79264 801126 79332 801182
rect 79388 801126 79456 801182
rect 79512 801126 79580 801182
rect 79636 801126 79704 801182
rect 79760 801126 79828 801182
rect 79884 801126 79952 801182
rect 80008 801126 80078 801182
rect 70130 801114 80078 801126
rect 70000 801058 80078 801114
rect 70000 801046 79208 801058
rect 70000 800990 70074 801046
rect 70130 801002 79208 801046
rect 79264 801002 79332 801058
rect 79388 801002 79456 801058
rect 79512 801002 79580 801058
rect 79636 801002 79704 801058
rect 79760 801002 79828 801058
rect 79884 801002 79952 801058
rect 80008 801002 80078 801058
rect 70130 800990 80078 801002
rect 70000 800934 80078 800990
rect 70000 800922 79208 800934
rect 70000 800866 70074 800922
rect 70130 800878 79208 800922
rect 79264 800878 79332 800934
rect 79388 800878 79456 800934
rect 79512 800878 79580 800934
rect 79636 800878 79704 800934
rect 79760 800878 79828 800934
rect 79884 800878 79952 800934
rect 80008 800878 80078 800934
rect 70130 800866 80078 800878
rect 70000 800828 80078 800866
rect 70000 800190 80078 800248
rect 70000 800184 79208 800190
rect 70000 800128 70074 800184
rect 70130 800134 79208 800184
rect 79264 800134 79332 800190
rect 79388 800134 79456 800190
rect 79512 800134 79580 800190
rect 79636 800134 79704 800190
rect 79760 800134 79828 800190
rect 79884 800134 79952 800190
rect 80008 800134 80078 800190
rect 70130 800128 80078 800134
rect 70000 800066 80078 800128
rect 70000 800060 79208 800066
rect 70000 800004 70074 800060
rect 70130 800010 79208 800060
rect 79264 800010 79332 800066
rect 79388 800010 79456 800066
rect 79512 800010 79580 800066
rect 79636 800010 79704 800066
rect 79760 800010 79828 800066
rect 79884 800010 79952 800066
rect 80008 800010 80078 800066
rect 70130 800004 80078 800010
rect 70000 799942 80078 800004
rect 70000 799936 79208 799942
rect 70000 799880 70074 799936
rect 70130 799886 79208 799936
rect 79264 799886 79332 799942
rect 79388 799886 79456 799942
rect 79512 799886 79580 799942
rect 79636 799886 79704 799942
rect 79760 799886 79828 799942
rect 79884 799886 79952 799942
rect 80008 799886 80078 799942
rect 70130 799880 80078 799886
rect 70000 799818 80078 799880
rect 70000 799812 79208 799818
rect 70000 799756 70074 799812
rect 70130 799762 79208 799812
rect 79264 799762 79332 799818
rect 79388 799762 79456 799818
rect 79512 799762 79580 799818
rect 79636 799762 79704 799818
rect 79760 799762 79828 799818
rect 79884 799762 79952 799818
rect 80008 799762 80078 799818
rect 70130 799756 80078 799762
rect 70000 799694 80078 799756
rect 70000 799688 79208 799694
rect 70000 799632 70074 799688
rect 70130 799638 79208 799688
rect 79264 799638 79332 799694
rect 79388 799638 79456 799694
rect 79512 799638 79580 799694
rect 79636 799638 79704 799694
rect 79760 799638 79828 799694
rect 79884 799638 79952 799694
rect 80008 799638 80078 799694
rect 70130 799632 80078 799638
rect 70000 799570 80078 799632
rect 70000 799564 79208 799570
rect 70000 799508 70074 799564
rect 70130 799514 79208 799564
rect 79264 799514 79332 799570
rect 79388 799514 79456 799570
rect 79512 799514 79580 799570
rect 79636 799514 79704 799570
rect 79760 799514 79828 799570
rect 79884 799514 79952 799570
rect 80008 799514 80078 799570
rect 70130 799508 80078 799514
rect 70000 799446 80078 799508
rect 70000 799440 79208 799446
rect 70000 799384 70074 799440
rect 70130 799390 79208 799440
rect 79264 799390 79332 799446
rect 79388 799390 79456 799446
rect 79512 799390 79580 799446
rect 79636 799390 79704 799446
rect 79760 799390 79828 799446
rect 79884 799390 79952 799446
rect 80008 799390 80078 799446
rect 70130 799384 80078 799390
rect 70000 799322 80078 799384
rect 70000 799316 79208 799322
rect 70000 799260 70074 799316
rect 70130 799266 79208 799316
rect 79264 799266 79332 799322
rect 79388 799266 79456 799322
rect 79512 799266 79580 799322
rect 79636 799266 79704 799322
rect 79760 799266 79828 799322
rect 79884 799266 79952 799322
rect 80008 799266 80078 799322
rect 70130 799260 80078 799266
rect 70000 799198 80078 799260
rect 70000 799192 79208 799198
rect 70000 799136 70074 799192
rect 70130 799142 79208 799192
rect 79264 799142 79332 799198
rect 79388 799142 79456 799198
rect 79512 799142 79580 799198
rect 79636 799142 79704 799198
rect 79760 799142 79828 799198
rect 79884 799142 79952 799198
rect 80008 799142 80078 799198
rect 70130 799136 80078 799142
rect 70000 799074 80078 799136
rect 70000 799068 79208 799074
rect 70000 799012 70074 799068
rect 70130 799018 79208 799068
rect 79264 799018 79332 799074
rect 79388 799018 79456 799074
rect 79512 799018 79580 799074
rect 79636 799018 79704 799074
rect 79760 799018 79828 799074
rect 79884 799018 79952 799074
rect 80008 799018 80078 799074
rect 70130 799012 80078 799018
rect 70000 798950 80078 799012
rect 70000 798944 79208 798950
rect 70000 798888 70074 798944
rect 70130 798894 79208 798944
rect 79264 798894 79332 798950
rect 79388 798894 79456 798950
rect 79512 798894 79580 798950
rect 79636 798894 79704 798950
rect 79760 798894 79828 798950
rect 79884 798894 79952 798950
rect 80008 798894 80078 798950
rect 70130 798888 80078 798894
rect 70000 798826 80078 798888
rect 70000 798820 79208 798826
rect 70000 798764 70074 798820
rect 70130 798770 79208 798820
rect 79264 798770 79332 798826
rect 79388 798770 79456 798826
rect 79512 798770 79580 798826
rect 79636 798770 79704 798826
rect 79760 798770 79828 798826
rect 79884 798770 79952 798826
rect 80008 798770 80078 798826
rect 70130 798764 80078 798770
rect 70000 798702 80078 798764
rect 70000 798696 79208 798702
rect 70000 798640 70074 798696
rect 70130 798646 79208 798696
rect 79264 798646 79332 798702
rect 79388 798646 79456 798702
rect 79512 798646 79580 798702
rect 79636 798646 79704 798702
rect 79760 798646 79828 798702
rect 79884 798646 79952 798702
rect 80008 798646 80078 798702
rect 70130 798640 80078 798646
rect 70000 798578 80078 798640
rect 70000 798572 79208 798578
rect 70000 798516 70074 798572
rect 70130 798522 79208 798572
rect 79264 798522 79332 798578
rect 79388 798522 79456 798578
rect 79512 798522 79580 798578
rect 79636 798522 79704 798578
rect 79760 798522 79828 798578
rect 79884 798522 79952 798578
rect 80008 798522 80078 798578
rect 70130 798516 80078 798522
rect 70000 798454 80078 798516
rect 70000 798448 79208 798454
rect 70000 798392 70074 798448
rect 70130 798398 79208 798448
rect 79264 798398 79332 798454
rect 79388 798398 79456 798454
rect 79512 798398 79580 798454
rect 79636 798398 79704 798454
rect 79760 798398 79828 798454
rect 79884 798398 79952 798454
rect 80008 798398 80078 798454
rect 70130 798392 80078 798398
rect 70000 798330 80078 798392
rect 70000 798324 79208 798330
rect 70000 798268 70074 798324
rect 70130 798274 79208 798324
rect 79264 798274 79332 798330
rect 79388 798274 79456 798330
rect 79512 798274 79580 798330
rect 79636 798274 79704 798330
rect 79760 798274 79828 798330
rect 79884 798274 79952 798330
rect 80008 798274 80078 798330
rect 70130 798268 80078 798274
rect 70000 798198 80078 798268
rect 70000 797820 80078 797878
rect 70000 797814 79208 797820
rect 70000 797758 70074 797814
rect 70130 797764 79208 797814
rect 79264 797764 79332 797820
rect 79388 797764 79456 797820
rect 79512 797764 79580 797820
rect 79636 797764 79704 797820
rect 79760 797764 79828 797820
rect 79884 797764 79952 797820
rect 80008 797764 80078 797820
rect 70130 797758 80078 797764
rect 70000 797696 80078 797758
rect 70000 797690 79208 797696
rect 70000 797634 70074 797690
rect 70130 797640 79208 797690
rect 79264 797640 79332 797696
rect 79388 797640 79456 797696
rect 79512 797640 79580 797696
rect 79636 797640 79704 797696
rect 79760 797640 79828 797696
rect 79884 797640 79952 797696
rect 80008 797640 80078 797696
rect 70130 797634 80078 797640
rect 70000 797572 80078 797634
rect 70000 797566 79208 797572
rect 70000 797510 70074 797566
rect 70130 797516 79208 797566
rect 79264 797516 79332 797572
rect 79388 797516 79456 797572
rect 79512 797516 79580 797572
rect 79636 797516 79704 797572
rect 79760 797516 79828 797572
rect 79884 797516 79952 797572
rect 80008 797516 80078 797572
rect 70130 797510 80078 797516
rect 70000 797448 80078 797510
rect 70000 797442 79208 797448
rect 70000 797386 70074 797442
rect 70130 797392 79208 797442
rect 79264 797392 79332 797448
rect 79388 797392 79456 797448
rect 79512 797392 79580 797448
rect 79636 797392 79704 797448
rect 79760 797392 79828 797448
rect 79884 797392 79952 797448
rect 80008 797392 80078 797448
rect 70130 797386 80078 797392
rect 70000 797324 80078 797386
rect 70000 797318 79208 797324
rect 70000 797262 70074 797318
rect 70130 797268 79208 797318
rect 79264 797268 79332 797324
rect 79388 797268 79456 797324
rect 79512 797268 79580 797324
rect 79636 797268 79704 797324
rect 79760 797268 79828 797324
rect 79884 797268 79952 797324
rect 80008 797268 80078 797324
rect 70130 797262 80078 797268
rect 70000 797200 80078 797262
rect 70000 797194 79208 797200
rect 70000 797138 70074 797194
rect 70130 797144 79208 797194
rect 79264 797144 79332 797200
rect 79388 797144 79456 797200
rect 79512 797144 79580 797200
rect 79636 797144 79704 797200
rect 79760 797144 79828 797200
rect 79884 797144 79952 797200
rect 80008 797144 80078 797200
rect 70130 797138 80078 797144
rect 70000 797076 80078 797138
rect 70000 797070 79208 797076
rect 70000 797014 70074 797070
rect 70130 797020 79208 797070
rect 79264 797020 79332 797076
rect 79388 797020 79456 797076
rect 79512 797020 79580 797076
rect 79636 797020 79704 797076
rect 79760 797020 79828 797076
rect 79884 797020 79952 797076
rect 80008 797020 80078 797076
rect 70130 797014 80078 797020
rect 70000 796952 80078 797014
rect 70000 796946 79208 796952
rect 70000 796890 70074 796946
rect 70130 796896 79208 796946
rect 79264 796896 79332 796952
rect 79388 796896 79456 796952
rect 79512 796896 79580 796952
rect 79636 796896 79704 796952
rect 79760 796896 79828 796952
rect 79884 796896 79952 796952
rect 80008 796896 80078 796952
rect 70130 796890 80078 796896
rect 70000 796828 80078 796890
rect 70000 796822 79208 796828
rect 70000 796766 70074 796822
rect 70130 796772 79208 796822
rect 79264 796772 79332 796828
rect 79388 796772 79456 796828
rect 79512 796772 79580 796828
rect 79636 796772 79704 796828
rect 79760 796772 79828 796828
rect 79884 796772 79952 796828
rect 80008 796772 80078 796828
rect 70130 796766 80078 796772
rect 70000 796704 80078 796766
rect 70000 796698 79208 796704
rect 70000 796642 70074 796698
rect 70130 796648 79208 796698
rect 79264 796648 79332 796704
rect 79388 796648 79456 796704
rect 79512 796648 79580 796704
rect 79636 796648 79704 796704
rect 79760 796648 79828 796704
rect 79884 796648 79952 796704
rect 80008 796648 80078 796704
rect 70130 796642 80078 796648
rect 70000 796580 80078 796642
rect 70000 796574 79208 796580
rect 70000 796518 70074 796574
rect 70130 796524 79208 796574
rect 79264 796524 79332 796580
rect 79388 796524 79456 796580
rect 79512 796524 79580 796580
rect 79636 796524 79704 796580
rect 79760 796524 79828 796580
rect 79884 796524 79952 796580
rect 80008 796524 80078 796580
rect 70130 796518 80078 796524
rect 70000 796456 80078 796518
rect 70000 796450 79208 796456
rect 70000 796394 70074 796450
rect 70130 796400 79208 796450
rect 79264 796400 79332 796456
rect 79388 796400 79456 796456
rect 79512 796400 79580 796456
rect 79636 796400 79704 796456
rect 79760 796400 79828 796456
rect 79884 796400 79952 796456
rect 80008 796400 80078 796456
rect 70130 796394 80078 796400
rect 70000 796332 80078 796394
rect 70000 796326 79208 796332
rect 70000 796270 70074 796326
rect 70130 796276 79208 796326
rect 79264 796276 79332 796332
rect 79388 796276 79456 796332
rect 79512 796276 79580 796332
rect 79636 796276 79704 796332
rect 79760 796276 79828 796332
rect 79884 796276 79952 796332
rect 80008 796276 80078 796332
rect 70130 796270 80078 796276
rect 70000 796208 80078 796270
rect 70000 796202 79208 796208
rect 70000 796146 70074 796202
rect 70130 796152 79208 796202
rect 79264 796152 79332 796208
rect 79388 796152 79456 796208
rect 79512 796152 79580 796208
rect 79636 796152 79704 796208
rect 79760 796152 79828 796208
rect 79884 796152 79952 796208
rect 80008 796152 80078 796208
rect 70130 796146 80078 796152
rect 70000 796084 80078 796146
rect 70000 796078 79208 796084
rect 70000 796022 70074 796078
rect 70130 796028 79208 796078
rect 79264 796028 79332 796084
rect 79388 796028 79456 796084
rect 79512 796028 79580 796084
rect 79636 796028 79704 796084
rect 79760 796028 79828 796084
rect 79884 796028 79952 796084
rect 80008 796028 80078 796084
rect 70130 796022 80078 796028
rect 70000 795960 80078 796022
rect 70000 795954 79208 795960
rect 70000 795898 70074 795954
rect 70130 795904 79208 795954
rect 79264 795904 79332 795960
rect 79388 795904 79456 795960
rect 79512 795904 79580 795960
rect 79636 795904 79704 795960
rect 79760 795904 79828 795960
rect 79884 795904 79952 795960
rect 80008 795904 80078 795960
rect 70130 795898 80078 795904
rect 70000 795828 80078 795898
rect 699322 797658 708000 797728
rect 699322 797652 707870 797658
rect 699322 797596 699392 797652
rect 699448 797596 699516 797652
rect 699572 797596 699640 797652
rect 699696 797596 699764 797652
rect 699820 797596 699888 797652
rect 699944 797596 700012 797652
rect 700068 797596 700136 797652
rect 700192 797602 707870 797652
rect 707926 797602 708000 797658
rect 700192 797596 708000 797602
rect 699322 797534 708000 797596
rect 699322 797528 707870 797534
rect 699322 797472 699392 797528
rect 699448 797472 699516 797528
rect 699572 797472 699640 797528
rect 699696 797472 699764 797528
rect 699820 797472 699888 797528
rect 699944 797472 700012 797528
rect 700068 797472 700136 797528
rect 700192 797478 707870 797528
rect 707926 797478 708000 797534
rect 700192 797472 708000 797478
rect 699322 797410 708000 797472
rect 699322 797404 707870 797410
rect 699322 797348 699392 797404
rect 699448 797348 699516 797404
rect 699572 797348 699640 797404
rect 699696 797348 699764 797404
rect 699820 797348 699888 797404
rect 699944 797348 700012 797404
rect 700068 797348 700136 797404
rect 700192 797354 707870 797404
rect 707926 797354 708000 797410
rect 700192 797348 708000 797354
rect 699322 797286 708000 797348
rect 699322 797280 707870 797286
rect 699322 797224 699392 797280
rect 699448 797224 699516 797280
rect 699572 797224 699640 797280
rect 699696 797224 699764 797280
rect 699820 797224 699888 797280
rect 699944 797224 700012 797280
rect 700068 797224 700136 797280
rect 700192 797230 707870 797280
rect 707926 797230 708000 797286
rect 700192 797224 708000 797230
rect 699322 797162 708000 797224
rect 699322 797156 707870 797162
rect 699322 797100 699392 797156
rect 699448 797100 699516 797156
rect 699572 797100 699640 797156
rect 699696 797100 699764 797156
rect 699820 797100 699888 797156
rect 699944 797100 700012 797156
rect 700068 797100 700136 797156
rect 700192 797106 707870 797156
rect 707926 797106 708000 797162
rect 700192 797100 708000 797106
rect 699322 797038 708000 797100
rect 699322 797032 707870 797038
rect 699322 796976 699392 797032
rect 699448 796976 699516 797032
rect 699572 796976 699640 797032
rect 699696 796976 699764 797032
rect 699820 796976 699888 797032
rect 699944 796976 700012 797032
rect 700068 796976 700136 797032
rect 700192 796982 707870 797032
rect 707926 796982 708000 797038
rect 700192 796976 708000 796982
rect 699322 796914 708000 796976
rect 699322 796908 707870 796914
rect 699322 796852 699392 796908
rect 699448 796852 699516 796908
rect 699572 796852 699640 796908
rect 699696 796852 699764 796908
rect 699820 796852 699888 796908
rect 699944 796852 700012 796908
rect 700068 796852 700136 796908
rect 700192 796858 707870 796908
rect 707926 796858 708000 796914
rect 700192 796852 708000 796858
rect 699322 796790 708000 796852
rect 699322 796784 707870 796790
rect 699322 796728 699392 796784
rect 699448 796728 699516 796784
rect 699572 796728 699640 796784
rect 699696 796728 699764 796784
rect 699820 796728 699888 796784
rect 699944 796728 700012 796784
rect 700068 796728 700136 796784
rect 700192 796734 707870 796784
rect 707926 796734 708000 796790
rect 700192 796728 708000 796734
rect 699322 796666 708000 796728
rect 699322 796660 707870 796666
rect 699322 796604 699392 796660
rect 699448 796604 699516 796660
rect 699572 796604 699640 796660
rect 699696 796604 699764 796660
rect 699820 796604 699888 796660
rect 699944 796604 700012 796660
rect 700068 796604 700136 796660
rect 700192 796610 707870 796660
rect 707926 796610 708000 796666
rect 700192 796604 708000 796610
rect 699322 796542 708000 796604
rect 699322 796536 707870 796542
rect 699322 796480 699392 796536
rect 699448 796480 699516 796536
rect 699572 796480 699640 796536
rect 699696 796480 699764 796536
rect 699820 796480 699888 796536
rect 699944 796480 700012 796536
rect 700068 796480 700136 796536
rect 700192 796486 707870 796536
rect 707926 796486 708000 796542
rect 700192 796480 708000 796486
rect 699322 796418 708000 796480
rect 699322 796412 707870 796418
rect 699322 796356 699392 796412
rect 699448 796356 699516 796412
rect 699572 796356 699640 796412
rect 699696 796356 699764 796412
rect 699820 796356 699888 796412
rect 699944 796356 700012 796412
rect 700068 796356 700136 796412
rect 700192 796362 707870 796412
rect 707926 796362 708000 796418
rect 700192 796356 708000 796362
rect 699322 796294 708000 796356
rect 699322 796288 707870 796294
rect 699322 796232 699392 796288
rect 699448 796232 699516 796288
rect 699572 796232 699640 796288
rect 699696 796232 699764 796288
rect 699820 796232 699888 796288
rect 699944 796232 700012 796288
rect 700068 796232 700136 796288
rect 700192 796238 707870 796288
rect 707926 796238 708000 796294
rect 700192 796232 708000 796238
rect 699322 796170 708000 796232
rect 699322 796164 707870 796170
rect 699322 796108 699392 796164
rect 699448 796108 699516 796164
rect 699572 796108 699640 796164
rect 699696 796108 699764 796164
rect 699820 796108 699888 796164
rect 699944 796108 700012 796164
rect 700068 796108 700136 796164
rect 700192 796114 707870 796164
rect 707926 796114 708000 796170
rect 700192 796108 708000 796114
rect 699322 796046 708000 796108
rect 699322 796040 707870 796046
rect 699322 795984 699392 796040
rect 699448 795984 699516 796040
rect 699572 795984 699640 796040
rect 699696 795984 699764 796040
rect 699820 795984 699888 796040
rect 699944 795984 700012 796040
rect 700068 795984 700136 796040
rect 700192 795990 707870 796040
rect 707926 795990 708000 796046
rect 700192 795984 708000 795990
rect 699322 795922 708000 795984
rect 699322 795916 707870 795922
rect 699322 795860 699392 795916
rect 699448 795860 699516 795916
rect 699572 795860 699640 795916
rect 699696 795860 699764 795916
rect 699820 795860 699888 795916
rect 699944 795860 700012 795916
rect 700068 795860 700136 795916
rect 700192 795866 707870 795916
rect 707926 795866 708000 795922
rect 700192 795860 708000 795866
rect 699322 795828 708000 795860
rect 699322 795178 708000 795248
rect 699322 795172 707870 795178
rect 70000 795114 80078 795172
rect 70000 795108 79208 795114
rect 70000 795052 70074 795108
rect 70130 795058 79208 795108
rect 79264 795058 79332 795114
rect 79388 795058 79456 795114
rect 79512 795058 79580 795114
rect 79636 795058 79704 795114
rect 79760 795058 79828 795114
rect 79884 795058 79952 795114
rect 80008 795058 80078 795114
rect 70130 795052 80078 795058
rect 70000 794990 80078 795052
rect 70000 794984 79208 794990
rect 70000 794928 70074 794984
rect 70130 794934 79208 794984
rect 79264 794934 79332 794990
rect 79388 794934 79456 794990
rect 79512 794934 79580 794990
rect 79636 794934 79704 794990
rect 79760 794934 79828 794990
rect 79884 794934 79952 794990
rect 80008 794934 80078 794990
rect 70130 794928 80078 794934
rect 70000 794866 80078 794928
rect 70000 794860 79208 794866
rect 70000 794804 70074 794860
rect 70130 794810 79208 794860
rect 79264 794810 79332 794866
rect 79388 794810 79456 794866
rect 79512 794810 79580 794866
rect 79636 794810 79704 794866
rect 79760 794810 79828 794866
rect 79884 794810 79952 794866
rect 80008 794810 80078 794866
rect 70130 794804 80078 794810
rect 70000 794742 80078 794804
rect 70000 794736 79208 794742
rect 70000 794680 70074 794736
rect 70130 794686 79208 794736
rect 79264 794686 79332 794742
rect 79388 794686 79456 794742
rect 79512 794686 79580 794742
rect 79636 794686 79704 794742
rect 79760 794686 79828 794742
rect 79884 794686 79952 794742
rect 80008 794686 80078 794742
rect 70130 794680 80078 794686
rect 70000 794618 80078 794680
rect 70000 794612 79208 794618
rect 70000 794556 70074 794612
rect 70130 794562 79208 794612
rect 79264 794562 79332 794618
rect 79388 794562 79456 794618
rect 79512 794562 79580 794618
rect 79636 794562 79704 794618
rect 79760 794562 79828 794618
rect 79884 794562 79952 794618
rect 80008 794562 80078 794618
rect 70130 794556 80078 794562
rect 70000 794494 80078 794556
rect 70000 794488 79208 794494
rect 70000 794432 70074 794488
rect 70130 794438 79208 794488
rect 79264 794438 79332 794494
rect 79388 794438 79456 794494
rect 79512 794438 79580 794494
rect 79636 794438 79704 794494
rect 79760 794438 79828 794494
rect 79884 794438 79952 794494
rect 80008 794438 80078 794494
rect 70130 794432 80078 794438
rect 70000 794370 80078 794432
rect 70000 794364 79208 794370
rect 70000 794308 70074 794364
rect 70130 794314 79208 794364
rect 79264 794314 79332 794370
rect 79388 794314 79456 794370
rect 79512 794314 79580 794370
rect 79636 794314 79704 794370
rect 79760 794314 79828 794370
rect 79884 794314 79952 794370
rect 80008 794314 80078 794370
rect 70130 794308 80078 794314
rect 70000 794246 80078 794308
rect 70000 794240 79208 794246
rect 70000 794184 70074 794240
rect 70130 794190 79208 794240
rect 79264 794190 79332 794246
rect 79388 794190 79456 794246
rect 79512 794190 79580 794246
rect 79636 794190 79704 794246
rect 79760 794190 79828 794246
rect 79884 794190 79952 794246
rect 80008 794190 80078 794246
rect 70130 794184 80078 794190
rect 70000 794122 80078 794184
rect 70000 794116 79208 794122
rect 70000 794060 70074 794116
rect 70130 794066 79208 794116
rect 79264 794066 79332 794122
rect 79388 794066 79456 794122
rect 79512 794066 79580 794122
rect 79636 794066 79704 794122
rect 79760 794066 79828 794122
rect 79884 794066 79952 794122
rect 80008 794066 80078 794122
rect 70130 794060 80078 794066
rect 70000 793998 80078 794060
rect 70000 793992 79208 793998
rect 70000 793936 70074 793992
rect 70130 793942 79208 793992
rect 79264 793942 79332 793998
rect 79388 793942 79456 793998
rect 79512 793942 79580 793998
rect 79636 793942 79704 793998
rect 79760 793942 79828 793998
rect 79884 793942 79952 793998
rect 80008 793942 80078 793998
rect 70130 793936 80078 793942
rect 70000 793874 80078 793936
rect 70000 793868 79208 793874
rect 70000 793812 70074 793868
rect 70130 793818 79208 793868
rect 79264 793818 79332 793874
rect 79388 793818 79456 793874
rect 79512 793818 79580 793874
rect 79636 793818 79704 793874
rect 79760 793818 79828 793874
rect 79884 793818 79952 793874
rect 80008 793818 80078 793874
rect 70130 793812 80078 793818
rect 70000 793750 80078 793812
rect 70000 793744 79208 793750
rect 70000 793688 70074 793744
rect 70130 793694 79208 793744
rect 79264 793694 79332 793750
rect 79388 793694 79456 793750
rect 79512 793694 79580 793750
rect 79636 793694 79704 793750
rect 79760 793694 79828 793750
rect 79884 793694 79952 793750
rect 80008 793694 80078 793750
rect 70130 793688 80078 793694
rect 70000 793626 80078 793688
rect 70000 793620 79208 793626
rect 70000 793564 70074 793620
rect 70130 793570 79208 793620
rect 79264 793570 79332 793626
rect 79388 793570 79456 793626
rect 79512 793570 79580 793626
rect 79636 793570 79704 793626
rect 79760 793570 79828 793626
rect 79884 793570 79952 793626
rect 80008 793570 80078 793626
rect 70130 793564 80078 793570
rect 70000 793502 80078 793564
rect 70000 793496 79208 793502
rect 70000 793440 70074 793496
rect 70130 793446 79208 793496
rect 79264 793446 79332 793502
rect 79388 793446 79456 793502
rect 79512 793446 79580 793502
rect 79636 793446 79704 793502
rect 79760 793446 79828 793502
rect 79884 793446 79952 793502
rect 80008 793446 80078 793502
rect 70130 793440 80078 793446
rect 70000 793378 80078 793440
rect 70000 793372 79208 793378
rect 70000 793316 70074 793372
rect 70130 793322 79208 793372
rect 79264 793322 79332 793378
rect 79388 793322 79456 793378
rect 79512 793322 79580 793378
rect 79636 793322 79704 793378
rect 79760 793322 79828 793378
rect 79884 793322 79952 793378
rect 80008 793322 80078 793378
rect 70130 793316 80078 793322
rect 70000 793254 80078 793316
rect 70000 793248 79208 793254
rect 70000 793192 70074 793248
rect 70130 793198 79208 793248
rect 79264 793198 79332 793254
rect 79388 793198 79456 793254
rect 79512 793198 79580 793254
rect 79636 793198 79704 793254
rect 79760 793198 79828 793254
rect 79884 793198 79952 793254
rect 80008 793198 80078 793254
rect 699322 795116 699392 795172
rect 699448 795116 699516 795172
rect 699572 795116 699640 795172
rect 699696 795116 699764 795172
rect 699820 795116 699888 795172
rect 699944 795116 700012 795172
rect 700068 795116 700136 795172
rect 700192 795122 707870 795172
rect 707926 795122 708000 795178
rect 700192 795116 708000 795122
rect 699322 795054 708000 795116
rect 699322 795048 707870 795054
rect 699322 794992 699392 795048
rect 699448 794992 699516 795048
rect 699572 794992 699640 795048
rect 699696 794992 699764 795048
rect 699820 794992 699888 795048
rect 699944 794992 700012 795048
rect 700068 794992 700136 795048
rect 700192 794998 707870 795048
rect 707926 794998 708000 795054
rect 700192 794992 708000 794998
rect 699322 794930 708000 794992
rect 699322 794924 707870 794930
rect 699322 794868 699392 794924
rect 699448 794868 699516 794924
rect 699572 794868 699640 794924
rect 699696 794868 699764 794924
rect 699820 794868 699888 794924
rect 699944 794868 700012 794924
rect 700068 794868 700136 794924
rect 700192 794874 707870 794924
rect 707926 794874 708000 794930
rect 700192 794868 708000 794874
rect 699322 794806 708000 794868
rect 699322 794800 707870 794806
rect 699322 794744 699392 794800
rect 699448 794744 699516 794800
rect 699572 794744 699640 794800
rect 699696 794744 699764 794800
rect 699820 794744 699888 794800
rect 699944 794744 700012 794800
rect 700068 794744 700136 794800
rect 700192 794750 707870 794800
rect 707926 794750 708000 794806
rect 700192 794744 708000 794750
rect 699322 794682 708000 794744
rect 699322 794676 707870 794682
rect 699322 794620 699392 794676
rect 699448 794620 699516 794676
rect 699572 794620 699640 794676
rect 699696 794620 699764 794676
rect 699820 794620 699888 794676
rect 699944 794620 700012 794676
rect 700068 794620 700136 794676
rect 700192 794626 707870 794676
rect 707926 794626 708000 794682
rect 700192 794620 708000 794626
rect 699322 794558 708000 794620
rect 699322 794552 707870 794558
rect 699322 794496 699392 794552
rect 699448 794496 699516 794552
rect 699572 794496 699640 794552
rect 699696 794496 699764 794552
rect 699820 794496 699888 794552
rect 699944 794496 700012 794552
rect 700068 794496 700136 794552
rect 700192 794502 707870 794552
rect 707926 794502 708000 794558
rect 700192 794496 708000 794502
rect 699322 794434 708000 794496
rect 699322 794428 707870 794434
rect 699322 794372 699392 794428
rect 699448 794372 699516 794428
rect 699572 794372 699640 794428
rect 699696 794372 699764 794428
rect 699820 794372 699888 794428
rect 699944 794372 700012 794428
rect 700068 794372 700136 794428
rect 700192 794378 707870 794428
rect 707926 794378 708000 794434
rect 700192 794372 708000 794378
rect 699322 794310 708000 794372
rect 699322 794304 707870 794310
rect 699322 794248 699392 794304
rect 699448 794248 699516 794304
rect 699572 794248 699640 794304
rect 699696 794248 699764 794304
rect 699820 794248 699888 794304
rect 699944 794248 700012 794304
rect 700068 794248 700136 794304
rect 700192 794254 707870 794304
rect 707926 794254 708000 794310
rect 700192 794248 708000 794254
rect 699322 794186 708000 794248
rect 699322 794180 707870 794186
rect 699322 794124 699392 794180
rect 699448 794124 699516 794180
rect 699572 794124 699640 794180
rect 699696 794124 699764 794180
rect 699820 794124 699888 794180
rect 699944 794124 700012 794180
rect 700068 794124 700136 794180
rect 700192 794130 707870 794180
rect 707926 794130 708000 794186
rect 700192 794124 708000 794130
rect 699322 794062 708000 794124
rect 699322 794056 707870 794062
rect 699322 794000 699392 794056
rect 699448 794000 699516 794056
rect 699572 794000 699640 794056
rect 699696 794000 699764 794056
rect 699820 794000 699888 794056
rect 699944 794000 700012 794056
rect 700068 794000 700136 794056
rect 700192 794006 707870 794056
rect 707926 794006 708000 794062
rect 700192 794000 708000 794006
rect 699322 793938 708000 794000
rect 699322 793932 707870 793938
rect 699322 793876 699392 793932
rect 699448 793876 699516 793932
rect 699572 793876 699640 793932
rect 699696 793876 699764 793932
rect 699820 793876 699888 793932
rect 699944 793876 700012 793932
rect 700068 793876 700136 793932
rect 700192 793882 707870 793932
rect 707926 793882 708000 793938
rect 700192 793876 708000 793882
rect 699322 793814 708000 793876
rect 699322 793808 707870 793814
rect 699322 793752 699392 793808
rect 699448 793752 699516 793808
rect 699572 793752 699640 793808
rect 699696 793752 699764 793808
rect 699820 793752 699888 793808
rect 699944 793752 700012 793808
rect 700068 793752 700136 793808
rect 700192 793758 707870 793808
rect 707926 793758 708000 793814
rect 700192 793752 708000 793758
rect 699322 793690 708000 793752
rect 699322 793684 707870 793690
rect 699322 793628 699392 793684
rect 699448 793628 699516 793684
rect 699572 793628 699640 793684
rect 699696 793628 699764 793684
rect 699820 793628 699888 793684
rect 699944 793628 700012 793684
rect 700068 793628 700136 793684
rect 700192 793634 707870 793684
rect 707926 793634 708000 793690
rect 700192 793628 708000 793634
rect 699322 793566 708000 793628
rect 699322 793560 707870 793566
rect 699322 793504 699392 793560
rect 699448 793504 699516 793560
rect 699572 793504 699640 793560
rect 699696 793504 699764 793560
rect 699820 793504 699888 793560
rect 699944 793504 700012 793560
rect 700068 793504 700136 793560
rect 700192 793510 707870 793560
rect 707926 793510 708000 793566
rect 700192 793504 708000 793510
rect 699322 793442 708000 793504
rect 699322 793436 707870 793442
rect 699322 793380 699392 793436
rect 699448 793380 699516 793436
rect 699572 793380 699640 793436
rect 699696 793380 699764 793436
rect 699820 793380 699888 793436
rect 699944 793380 700012 793436
rect 700068 793380 700136 793436
rect 700192 793386 707870 793436
rect 707926 793386 708000 793442
rect 700192 793380 708000 793386
rect 699322 793318 708000 793380
rect 699322 793312 707870 793318
rect 699322 793256 699392 793312
rect 699448 793256 699516 793312
rect 699572 793256 699640 793312
rect 699696 793256 699764 793312
rect 699820 793256 699888 793312
rect 699944 793256 700012 793312
rect 700068 793256 700136 793312
rect 700192 793262 707870 793312
rect 707926 793262 708000 793318
rect 700192 793256 708000 793262
rect 699322 793198 708000 793256
rect 70130 793192 80078 793198
rect 70000 793122 80078 793192
rect 699322 792808 708000 792878
rect 699322 792802 707870 792808
rect 70000 792744 80078 792802
rect 70000 792738 79208 792744
rect 70000 792682 70074 792738
rect 70130 792688 79208 792738
rect 79264 792688 79332 792744
rect 79388 792688 79456 792744
rect 79512 792688 79580 792744
rect 79636 792688 79704 792744
rect 79760 792688 79828 792744
rect 79884 792688 79952 792744
rect 80008 792688 80078 792744
rect 70130 792682 80078 792688
rect 70000 792620 80078 792682
rect 70000 792614 79208 792620
rect 70000 792558 70074 792614
rect 70130 792564 79208 792614
rect 79264 792564 79332 792620
rect 79388 792564 79456 792620
rect 79512 792564 79580 792620
rect 79636 792564 79704 792620
rect 79760 792564 79828 792620
rect 79884 792564 79952 792620
rect 80008 792564 80078 792620
rect 70130 792558 80078 792564
rect 70000 792496 80078 792558
rect 70000 792490 79208 792496
rect 70000 792434 70074 792490
rect 70130 792440 79208 792490
rect 79264 792440 79332 792496
rect 79388 792440 79456 792496
rect 79512 792440 79580 792496
rect 79636 792440 79704 792496
rect 79760 792440 79828 792496
rect 79884 792440 79952 792496
rect 80008 792440 80078 792496
rect 70130 792434 80078 792440
rect 70000 792372 80078 792434
rect 70000 792366 79208 792372
rect 70000 792310 70074 792366
rect 70130 792316 79208 792366
rect 79264 792316 79332 792372
rect 79388 792316 79456 792372
rect 79512 792316 79580 792372
rect 79636 792316 79704 792372
rect 79760 792316 79828 792372
rect 79884 792316 79952 792372
rect 80008 792316 80078 792372
rect 70130 792310 80078 792316
rect 70000 792248 80078 792310
rect 70000 792242 79208 792248
rect 70000 792186 70074 792242
rect 70130 792192 79208 792242
rect 79264 792192 79332 792248
rect 79388 792192 79456 792248
rect 79512 792192 79580 792248
rect 79636 792192 79704 792248
rect 79760 792192 79828 792248
rect 79884 792192 79952 792248
rect 80008 792192 80078 792248
rect 70130 792186 80078 792192
rect 70000 792124 80078 792186
rect 70000 792118 79208 792124
rect 70000 792062 70074 792118
rect 70130 792068 79208 792118
rect 79264 792068 79332 792124
rect 79388 792068 79456 792124
rect 79512 792068 79580 792124
rect 79636 792068 79704 792124
rect 79760 792068 79828 792124
rect 79884 792068 79952 792124
rect 80008 792068 80078 792124
rect 70130 792062 80078 792068
rect 70000 792000 80078 792062
rect 70000 791994 79208 792000
rect 70000 791938 70074 791994
rect 70130 791944 79208 791994
rect 79264 791944 79332 792000
rect 79388 791944 79456 792000
rect 79512 791944 79580 792000
rect 79636 791944 79704 792000
rect 79760 791944 79828 792000
rect 79884 791944 79952 792000
rect 80008 791944 80078 792000
rect 70130 791938 80078 791944
rect 70000 791876 80078 791938
rect 70000 791870 79208 791876
rect 70000 791814 70074 791870
rect 70130 791820 79208 791870
rect 79264 791820 79332 791876
rect 79388 791820 79456 791876
rect 79512 791820 79580 791876
rect 79636 791820 79704 791876
rect 79760 791820 79828 791876
rect 79884 791820 79952 791876
rect 80008 791820 80078 791876
rect 70130 791814 80078 791820
rect 70000 791752 80078 791814
rect 70000 791746 79208 791752
rect 70000 791690 70074 791746
rect 70130 791696 79208 791746
rect 79264 791696 79332 791752
rect 79388 791696 79456 791752
rect 79512 791696 79580 791752
rect 79636 791696 79704 791752
rect 79760 791696 79828 791752
rect 79884 791696 79952 791752
rect 80008 791696 80078 791752
rect 70130 791690 80078 791696
rect 70000 791628 80078 791690
rect 70000 791622 79208 791628
rect 70000 791566 70074 791622
rect 70130 791572 79208 791622
rect 79264 791572 79332 791628
rect 79388 791572 79456 791628
rect 79512 791572 79580 791628
rect 79636 791572 79704 791628
rect 79760 791572 79828 791628
rect 79884 791572 79952 791628
rect 80008 791572 80078 791628
rect 70130 791566 80078 791572
rect 70000 791504 80078 791566
rect 70000 791498 79208 791504
rect 70000 791442 70074 791498
rect 70130 791448 79208 791498
rect 79264 791448 79332 791504
rect 79388 791448 79456 791504
rect 79512 791448 79580 791504
rect 79636 791448 79704 791504
rect 79760 791448 79828 791504
rect 79884 791448 79952 791504
rect 80008 791448 80078 791504
rect 70130 791442 80078 791448
rect 70000 791380 80078 791442
rect 70000 791374 79208 791380
rect 70000 791318 70074 791374
rect 70130 791324 79208 791374
rect 79264 791324 79332 791380
rect 79388 791324 79456 791380
rect 79512 791324 79580 791380
rect 79636 791324 79704 791380
rect 79760 791324 79828 791380
rect 79884 791324 79952 791380
rect 80008 791324 80078 791380
rect 70130 791318 80078 791324
rect 70000 791256 80078 791318
rect 70000 791250 79208 791256
rect 70000 791194 70074 791250
rect 70130 791200 79208 791250
rect 79264 791200 79332 791256
rect 79388 791200 79456 791256
rect 79512 791200 79580 791256
rect 79636 791200 79704 791256
rect 79760 791200 79828 791256
rect 79884 791200 79952 791256
rect 80008 791200 80078 791256
rect 70130 791194 80078 791200
rect 70000 791132 80078 791194
rect 70000 791126 79208 791132
rect 70000 791070 70074 791126
rect 70130 791076 79208 791126
rect 79264 791076 79332 791132
rect 79388 791076 79456 791132
rect 79512 791076 79580 791132
rect 79636 791076 79704 791132
rect 79760 791076 79828 791132
rect 79884 791076 79952 791132
rect 80008 791076 80078 791132
rect 70130 791070 80078 791076
rect 70000 791008 80078 791070
rect 70000 791002 79208 791008
rect 70000 790946 70074 791002
rect 70130 790952 79208 791002
rect 79264 790952 79332 791008
rect 79388 790952 79456 791008
rect 79512 790952 79580 791008
rect 79636 790952 79704 791008
rect 79760 790952 79828 791008
rect 79884 790952 79952 791008
rect 80008 790952 80078 791008
rect 70130 790946 80078 790952
rect 70000 790884 80078 790946
rect 70000 790878 79208 790884
rect 70000 790822 70074 790878
rect 70130 790828 79208 790878
rect 79264 790828 79332 790884
rect 79388 790828 79456 790884
rect 79512 790828 79580 790884
rect 79636 790828 79704 790884
rect 79760 790828 79828 790884
rect 79884 790828 79952 790884
rect 80008 790828 80078 790884
rect 699322 792746 699392 792802
rect 699448 792746 699516 792802
rect 699572 792746 699640 792802
rect 699696 792746 699764 792802
rect 699820 792746 699888 792802
rect 699944 792746 700012 792802
rect 700068 792746 700136 792802
rect 700192 792752 707870 792802
rect 707926 792752 708000 792808
rect 700192 792746 708000 792752
rect 699322 792684 708000 792746
rect 699322 792678 707870 792684
rect 699322 792622 699392 792678
rect 699448 792622 699516 792678
rect 699572 792622 699640 792678
rect 699696 792622 699764 792678
rect 699820 792622 699888 792678
rect 699944 792622 700012 792678
rect 700068 792622 700136 792678
rect 700192 792628 707870 792678
rect 707926 792628 708000 792684
rect 700192 792622 708000 792628
rect 699322 792560 708000 792622
rect 699322 792554 707870 792560
rect 699322 792498 699392 792554
rect 699448 792498 699516 792554
rect 699572 792498 699640 792554
rect 699696 792498 699764 792554
rect 699820 792498 699888 792554
rect 699944 792498 700012 792554
rect 700068 792498 700136 792554
rect 700192 792504 707870 792554
rect 707926 792504 708000 792560
rect 700192 792498 708000 792504
rect 699322 792436 708000 792498
rect 699322 792430 707870 792436
rect 699322 792374 699392 792430
rect 699448 792374 699516 792430
rect 699572 792374 699640 792430
rect 699696 792374 699764 792430
rect 699820 792374 699888 792430
rect 699944 792374 700012 792430
rect 700068 792374 700136 792430
rect 700192 792380 707870 792430
rect 707926 792380 708000 792436
rect 700192 792374 708000 792380
rect 699322 792312 708000 792374
rect 699322 792306 707870 792312
rect 699322 792250 699392 792306
rect 699448 792250 699516 792306
rect 699572 792250 699640 792306
rect 699696 792250 699764 792306
rect 699820 792250 699888 792306
rect 699944 792250 700012 792306
rect 700068 792250 700136 792306
rect 700192 792256 707870 792306
rect 707926 792256 708000 792312
rect 700192 792250 708000 792256
rect 699322 792188 708000 792250
rect 699322 792182 707870 792188
rect 699322 792126 699392 792182
rect 699448 792126 699516 792182
rect 699572 792126 699640 792182
rect 699696 792126 699764 792182
rect 699820 792126 699888 792182
rect 699944 792126 700012 792182
rect 700068 792126 700136 792182
rect 700192 792132 707870 792182
rect 707926 792132 708000 792188
rect 700192 792126 708000 792132
rect 699322 792064 708000 792126
rect 699322 792058 707870 792064
rect 699322 792002 699392 792058
rect 699448 792002 699516 792058
rect 699572 792002 699640 792058
rect 699696 792002 699764 792058
rect 699820 792002 699888 792058
rect 699944 792002 700012 792058
rect 700068 792002 700136 792058
rect 700192 792008 707870 792058
rect 707926 792008 708000 792064
rect 700192 792002 708000 792008
rect 699322 791940 708000 792002
rect 699322 791934 707870 791940
rect 699322 791878 699392 791934
rect 699448 791878 699516 791934
rect 699572 791878 699640 791934
rect 699696 791878 699764 791934
rect 699820 791878 699888 791934
rect 699944 791878 700012 791934
rect 700068 791878 700136 791934
rect 700192 791884 707870 791934
rect 707926 791884 708000 791940
rect 700192 791878 708000 791884
rect 699322 791816 708000 791878
rect 699322 791810 707870 791816
rect 699322 791754 699392 791810
rect 699448 791754 699516 791810
rect 699572 791754 699640 791810
rect 699696 791754 699764 791810
rect 699820 791754 699888 791810
rect 699944 791754 700012 791810
rect 700068 791754 700136 791810
rect 700192 791760 707870 791810
rect 707926 791760 708000 791816
rect 700192 791754 708000 791760
rect 699322 791692 708000 791754
rect 699322 791686 707870 791692
rect 699322 791630 699392 791686
rect 699448 791630 699516 791686
rect 699572 791630 699640 791686
rect 699696 791630 699764 791686
rect 699820 791630 699888 791686
rect 699944 791630 700012 791686
rect 700068 791630 700136 791686
rect 700192 791636 707870 791686
rect 707926 791636 708000 791692
rect 700192 791630 708000 791636
rect 699322 791568 708000 791630
rect 699322 791562 707870 791568
rect 699322 791506 699392 791562
rect 699448 791506 699516 791562
rect 699572 791506 699640 791562
rect 699696 791506 699764 791562
rect 699820 791506 699888 791562
rect 699944 791506 700012 791562
rect 700068 791506 700136 791562
rect 700192 791512 707870 791562
rect 707926 791512 708000 791568
rect 700192 791506 708000 791512
rect 699322 791444 708000 791506
rect 699322 791438 707870 791444
rect 699322 791382 699392 791438
rect 699448 791382 699516 791438
rect 699572 791382 699640 791438
rect 699696 791382 699764 791438
rect 699820 791382 699888 791438
rect 699944 791382 700012 791438
rect 700068 791382 700136 791438
rect 700192 791388 707870 791438
rect 707926 791388 708000 791444
rect 700192 791382 708000 791388
rect 699322 791320 708000 791382
rect 699322 791314 707870 791320
rect 699322 791258 699392 791314
rect 699448 791258 699516 791314
rect 699572 791258 699640 791314
rect 699696 791258 699764 791314
rect 699820 791258 699888 791314
rect 699944 791258 700012 791314
rect 700068 791258 700136 791314
rect 700192 791264 707870 791314
rect 707926 791264 708000 791320
rect 700192 791258 708000 791264
rect 699322 791196 708000 791258
rect 699322 791190 707870 791196
rect 699322 791134 699392 791190
rect 699448 791134 699516 791190
rect 699572 791134 699640 791190
rect 699696 791134 699764 791190
rect 699820 791134 699888 791190
rect 699944 791134 700012 791190
rect 700068 791134 700136 791190
rect 700192 791140 707870 791190
rect 707926 791140 708000 791196
rect 700192 791134 708000 791140
rect 699322 791072 708000 791134
rect 699322 791066 707870 791072
rect 699322 791010 699392 791066
rect 699448 791010 699516 791066
rect 699572 791010 699640 791066
rect 699696 791010 699764 791066
rect 699820 791010 699888 791066
rect 699944 791010 700012 791066
rect 700068 791010 700136 791066
rect 700192 791016 707870 791066
rect 707926 791016 708000 791072
rect 700192 791010 708000 791016
rect 699322 790948 708000 791010
rect 699322 790942 707870 790948
rect 699322 790886 699392 790942
rect 699448 790886 699516 790942
rect 699572 790886 699640 790942
rect 699696 790886 699764 790942
rect 699820 790886 699888 790942
rect 699944 790886 700012 790942
rect 700068 790886 700136 790942
rect 700192 790892 707870 790942
rect 707926 790892 708000 790948
rect 700192 790886 708000 790892
rect 699322 790828 708000 790886
rect 70130 790822 80078 790828
rect 70000 790752 80078 790822
rect 70000 790140 80078 790172
rect 70000 790134 79208 790140
rect 70000 790078 70074 790134
rect 70130 790084 79208 790134
rect 79264 790084 79332 790140
rect 79388 790084 79456 790140
rect 79512 790084 79580 790140
rect 79636 790084 79704 790140
rect 79760 790084 79828 790140
rect 79884 790084 79952 790140
rect 80008 790084 80078 790140
rect 70130 790078 80078 790084
rect 70000 790016 80078 790078
rect 70000 790010 79208 790016
rect 70000 789954 70074 790010
rect 70130 789960 79208 790010
rect 79264 789960 79332 790016
rect 79388 789960 79456 790016
rect 79512 789960 79580 790016
rect 79636 789960 79704 790016
rect 79760 789960 79828 790016
rect 79884 789960 79952 790016
rect 80008 789960 80078 790016
rect 70130 789954 80078 789960
rect 70000 789892 80078 789954
rect 70000 789886 79208 789892
rect 70000 789830 70074 789886
rect 70130 789836 79208 789886
rect 79264 789836 79332 789892
rect 79388 789836 79456 789892
rect 79512 789836 79580 789892
rect 79636 789836 79704 789892
rect 79760 789836 79828 789892
rect 79884 789836 79952 789892
rect 80008 789836 80078 789892
rect 70130 789830 80078 789836
rect 70000 789768 80078 789830
rect 70000 789762 79208 789768
rect 70000 789706 70074 789762
rect 70130 789712 79208 789762
rect 79264 789712 79332 789768
rect 79388 789712 79456 789768
rect 79512 789712 79580 789768
rect 79636 789712 79704 789768
rect 79760 789712 79828 789768
rect 79884 789712 79952 789768
rect 80008 789712 80078 789768
rect 70130 789706 80078 789712
rect 70000 789644 80078 789706
rect 70000 789638 79208 789644
rect 70000 789582 70074 789638
rect 70130 789588 79208 789638
rect 79264 789588 79332 789644
rect 79388 789588 79456 789644
rect 79512 789588 79580 789644
rect 79636 789588 79704 789644
rect 79760 789588 79828 789644
rect 79884 789588 79952 789644
rect 80008 789588 80078 789644
rect 70130 789582 80078 789588
rect 70000 789520 80078 789582
rect 70000 789514 79208 789520
rect 70000 789458 70074 789514
rect 70130 789464 79208 789514
rect 79264 789464 79332 789520
rect 79388 789464 79456 789520
rect 79512 789464 79580 789520
rect 79636 789464 79704 789520
rect 79760 789464 79828 789520
rect 79884 789464 79952 789520
rect 80008 789464 80078 789520
rect 70130 789458 80078 789464
rect 70000 789396 80078 789458
rect 70000 789390 79208 789396
rect 70000 789334 70074 789390
rect 70130 789340 79208 789390
rect 79264 789340 79332 789396
rect 79388 789340 79456 789396
rect 79512 789340 79580 789396
rect 79636 789340 79704 789396
rect 79760 789340 79828 789396
rect 79884 789340 79952 789396
rect 80008 789340 80078 789396
rect 70130 789334 80078 789340
rect 70000 789272 80078 789334
rect 70000 789266 79208 789272
rect 70000 789210 70074 789266
rect 70130 789216 79208 789266
rect 79264 789216 79332 789272
rect 79388 789216 79456 789272
rect 79512 789216 79580 789272
rect 79636 789216 79704 789272
rect 79760 789216 79828 789272
rect 79884 789216 79952 789272
rect 80008 789216 80078 789272
rect 70130 789210 80078 789216
rect 70000 789148 80078 789210
rect 70000 789142 79208 789148
rect 70000 789086 70074 789142
rect 70130 789092 79208 789142
rect 79264 789092 79332 789148
rect 79388 789092 79456 789148
rect 79512 789092 79580 789148
rect 79636 789092 79704 789148
rect 79760 789092 79828 789148
rect 79884 789092 79952 789148
rect 80008 789092 80078 789148
rect 70130 789086 80078 789092
rect 70000 789024 80078 789086
rect 70000 789018 79208 789024
rect 70000 788962 70074 789018
rect 70130 788968 79208 789018
rect 79264 788968 79332 789024
rect 79388 788968 79456 789024
rect 79512 788968 79580 789024
rect 79636 788968 79704 789024
rect 79760 788968 79828 789024
rect 79884 788968 79952 789024
rect 80008 788968 80078 789024
rect 70130 788962 80078 788968
rect 70000 788900 80078 788962
rect 70000 788894 79208 788900
rect 70000 788838 70074 788894
rect 70130 788844 79208 788894
rect 79264 788844 79332 788900
rect 79388 788844 79456 788900
rect 79512 788844 79580 788900
rect 79636 788844 79704 788900
rect 79760 788844 79828 788900
rect 79884 788844 79952 788900
rect 80008 788844 80078 788900
rect 70130 788838 80078 788844
rect 70000 788776 80078 788838
rect 70000 788770 79208 788776
rect 70000 788714 70074 788770
rect 70130 788720 79208 788770
rect 79264 788720 79332 788776
rect 79388 788720 79456 788776
rect 79512 788720 79580 788776
rect 79636 788720 79704 788776
rect 79760 788720 79828 788776
rect 79884 788720 79952 788776
rect 80008 788720 80078 788776
rect 70130 788714 80078 788720
rect 70000 788652 80078 788714
rect 70000 788646 79208 788652
rect 70000 788590 70074 788646
rect 70130 788596 79208 788646
rect 79264 788596 79332 788652
rect 79388 788596 79456 788652
rect 79512 788596 79580 788652
rect 79636 788596 79704 788652
rect 79760 788596 79828 788652
rect 79884 788596 79952 788652
rect 80008 788630 80078 788652
rect 699322 790102 708000 790172
rect 699322 790096 707870 790102
rect 699322 790040 699392 790096
rect 699448 790040 699516 790096
rect 699572 790040 699640 790096
rect 699696 790040 699764 790096
rect 699820 790040 699888 790096
rect 699944 790040 700012 790096
rect 700068 790040 700136 790096
rect 700192 790046 707870 790096
rect 707926 790046 708000 790102
rect 700192 790040 708000 790046
rect 699322 789978 708000 790040
rect 699322 789972 707870 789978
rect 699322 789916 699392 789972
rect 699448 789916 699516 789972
rect 699572 789916 699640 789972
rect 699696 789916 699764 789972
rect 699820 789916 699888 789972
rect 699944 789916 700012 789972
rect 700068 789916 700136 789972
rect 700192 789922 707870 789972
rect 707926 789922 708000 789978
rect 700192 789916 708000 789922
rect 699322 789854 708000 789916
rect 699322 789848 707870 789854
rect 699322 789792 699392 789848
rect 699448 789792 699516 789848
rect 699572 789792 699640 789848
rect 699696 789792 699764 789848
rect 699820 789792 699888 789848
rect 699944 789792 700012 789848
rect 700068 789792 700136 789848
rect 700192 789798 707870 789848
rect 707926 789798 708000 789854
rect 700192 789792 708000 789798
rect 699322 789730 708000 789792
rect 699322 789724 707870 789730
rect 699322 789668 699392 789724
rect 699448 789668 699516 789724
rect 699572 789668 699640 789724
rect 699696 789668 699764 789724
rect 699820 789668 699888 789724
rect 699944 789668 700012 789724
rect 700068 789668 700136 789724
rect 700192 789674 707870 789724
rect 707926 789674 708000 789730
rect 700192 789668 708000 789674
rect 699322 789606 708000 789668
rect 699322 789600 707870 789606
rect 699322 789544 699392 789600
rect 699448 789544 699516 789600
rect 699572 789544 699640 789600
rect 699696 789544 699764 789600
rect 699820 789544 699888 789600
rect 699944 789544 700012 789600
rect 700068 789544 700136 789600
rect 700192 789550 707870 789600
rect 707926 789550 708000 789606
rect 700192 789544 708000 789550
rect 699322 789482 708000 789544
rect 699322 789476 707870 789482
rect 699322 789420 699392 789476
rect 699448 789420 699516 789476
rect 699572 789420 699640 789476
rect 699696 789420 699764 789476
rect 699820 789420 699888 789476
rect 699944 789420 700012 789476
rect 700068 789420 700136 789476
rect 700192 789426 707870 789476
rect 707926 789426 708000 789482
rect 700192 789420 708000 789426
rect 699322 789358 708000 789420
rect 699322 789352 707870 789358
rect 699322 789296 699392 789352
rect 699448 789296 699516 789352
rect 699572 789296 699640 789352
rect 699696 789296 699764 789352
rect 699820 789296 699888 789352
rect 699944 789296 700012 789352
rect 700068 789296 700136 789352
rect 700192 789302 707870 789352
rect 707926 789302 708000 789358
rect 700192 789296 708000 789302
rect 699322 789234 708000 789296
rect 699322 789228 707870 789234
rect 699322 789172 699392 789228
rect 699448 789172 699516 789228
rect 699572 789172 699640 789228
rect 699696 789172 699764 789228
rect 699820 789172 699888 789228
rect 699944 789172 700012 789228
rect 700068 789172 700136 789228
rect 700192 789178 707870 789228
rect 707926 789178 708000 789234
rect 700192 789172 708000 789178
rect 699322 789110 708000 789172
rect 699322 789104 707870 789110
rect 699322 789048 699392 789104
rect 699448 789048 699516 789104
rect 699572 789048 699640 789104
rect 699696 789048 699764 789104
rect 699820 789048 699888 789104
rect 699944 789048 700012 789104
rect 700068 789048 700136 789104
rect 700192 789054 707870 789104
rect 707926 789054 708000 789110
rect 700192 789048 708000 789054
rect 699322 788986 708000 789048
rect 699322 788980 707870 788986
rect 699322 788924 699392 788980
rect 699448 788924 699516 788980
rect 699572 788924 699640 788980
rect 699696 788924 699764 788980
rect 699820 788924 699888 788980
rect 699944 788924 700012 788980
rect 700068 788924 700136 788980
rect 700192 788930 707870 788980
rect 707926 788930 708000 788986
rect 700192 788924 708000 788930
rect 699322 788862 708000 788924
rect 699322 788856 707870 788862
rect 699322 788800 699392 788856
rect 699448 788800 699516 788856
rect 699572 788800 699640 788856
rect 699696 788800 699764 788856
rect 699820 788800 699888 788856
rect 699944 788800 700012 788856
rect 700068 788800 700136 788856
rect 700192 788806 707870 788856
rect 707926 788806 708000 788862
rect 700192 788800 708000 788806
rect 699322 788738 708000 788800
rect 699322 788732 707870 788738
rect 699322 788676 699392 788732
rect 699448 788676 699516 788732
rect 699572 788676 699640 788732
rect 699696 788676 699764 788732
rect 699820 788676 699888 788732
rect 699944 788676 700012 788732
rect 700068 788676 700136 788732
rect 700192 788682 707870 788732
rect 707926 788682 708000 788738
rect 700192 788676 708000 788682
rect 80008 788596 83556 788630
rect 70130 788590 83556 788596
rect 70000 788528 83556 788590
rect 70000 788522 79208 788528
rect 70000 788466 70074 788522
rect 70130 788472 79208 788522
rect 79264 788472 79332 788528
rect 79388 788472 79456 788528
rect 79512 788472 79580 788528
rect 79636 788472 79704 788528
rect 79760 788472 79828 788528
rect 79884 788472 79952 788528
rect 80008 788472 83556 788528
rect 70130 788466 83556 788472
rect 70000 788404 83556 788466
rect 70000 788398 79208 788404
rect 70000 788342 70074 788398
rect 70130 788348 79208 788398
rect 79264 788348 79332 788404
rect 79388 788348 79456 788404
rect 79512 788348 79580 788404
rect 79636 788348 79704 788404
rect 79760 788348 79828 788404
rect 79884 788348 79952 788404
rect 80008 788348 83556 788404
rect 70130 788342 83556 788348
rect 70000 788272 83556 788342
rect 79078 788010 83556 788272
rect 699322 788614 708000 788676
rect 699322 788608 707870 788614
rect 699322 788552 699392 788608
rect 699448 788552 699516 788608
rect 699572 788552 699640 788608
rect 699696 788552 699764 788608
rect 699820 788552 699888 788608
rect 699944 788552 700012 788608
rect 700068 788552 700136 788608
rect 700192 788558 707870 788608
rect 707926 788558 708000 788614
rect 700192 788552 708000 788558
rect 699322 788490 708000 788552
rect 699322 788484 707870 788490
rect 699322 788428 699392 788484
rect 699448 788428 699516 788484
rect 699572 788428 699640 788484
rect 699696 788428 699764 788484
rect 699820 788428 699888 788484
rect 699944 788428 700012 788484
rect 700068 788428 700136 788484
rect 700192 788434 707870 788484
rect 707926 788434 708000 788490
rect 700192 788428 708000 788434
rect 699322 788366 708000 788428
rect 699322 788360 707870 788366
rect 699322 788304 699392 788360
rect 699448 788304 699516 788360
rect 699572 788304 699640 788360
rect 699696 788304 699764 788360
rect 699820 788304 699888 788360
rect 699944 788304 700012 788360
rect 700068 788304 700136 788360
rect 700192 788310 707870 788360
rect 707926 788310 708000 788366
rect 700192 788304 708000 788310
rect 699322 788242 708000 788304
rect 699322 788236 707870 788242
rect 699322 788180 699392 788236
rect 699448 788180 699516 788236
rect 699572 788180 699640 788236
rect 699696 788180 699764 788236
rect 699820 788180 699888 788236
rect 699944 788180 700012 788236
rect 700068 788180 700136 788236
rect 700192 788186 707870 788236
rect 707926 788186 708000 788242
rect 700192 788180 708000 788186
rect 699322 788122 708000 788180
rect 699322 787732 708000 787802
rect 699322 787726 707870 787732
rect 699322 787670 699392 787726
rect 699448 787670 699516 787726
rect 699572 787670 699640 787726
rect 699696 787670 699764 787726
rect 699820 787670 699888 787726
rect 699944 787670 700012 787726
rect 700068 787670 700136 787726
rect 700192 787676 707870 787726
rect 707926 787676 708000 787732
rect 700192 787670 708000 787676
rect 699322 787608 708000 787670
rect 699322 787602 707870 787608
rect 699322 787546 699392 787602
rect 699448 787546 699516 787602
rect 699572 787546 699640 787602
rect 699696 787546 699764 787602
rect 699820 787546 699888 787602
rect 699944 787546 700012 787602
rect 700068 787546 700136 787602
rect 700192 787552 707870 787602
rect 707926 787552 708000 787608
rect 700192 787546 708000 787552
rect 699322 787484 708000 787546
rect 699322 787478 707870 787484
rect 699322 787422 699392 787478
rect 699448 787422 699516 787478
rect 699572 787422 699640 787478
rect 699696 787422 699764 787478
rect 699820 787422 699888 787478
rect 699944 787422 700012 787478
rect 700068 787422 700136 787478
rect 700192 787428 707870 787478
rect 707926 787428 708000 787484
rect 700192 787422 708000 787428
rect 699322 787360 708000 787422
rect 699322 787354 707870 787360
rect 699322 787298 699392 787354
rect 699448 787298 699516 787354
rect 699572 787298 699640 787354
rect 699696 787298 699764 787354
rect 699820 787298 699888 787354
rect 699944 787298 700012 787354
rect 700068 787298 700136 787354
rect 700192 787304 707870 787354
rect 707926 787304 708000 787360
rect 700192 787298 708000 787304
rect 699322 787236 708000 787298
rect 699322 787230 707870 787236
rect 699322 787174 699392 787230
rect 699448 787174 699516 787230
rect 699572 787174 699640 787230
rect 699696 787174 699764 787230
rect 699820 787174 699888 787230
rect 699944 787174 700012 787230
rect 700068 787174 700136 787230
rect 700192 787180 707870 787230
rect 707926 787180 708000 787236
rect 700192 787174 708000 787180
rect 699322 787112 708000 787174
rect 699322 787106 707870 787112
rect 699322 787050 699392 787106
rect 699448 787050 699516 787106
rect 699572 787050 699640 787106
rect 699696 787050 699764 787106
rect 699820 787050 699888 787106
rect 699944 787050 700012 787106
rect 700068 787050 700136 787106
rect 700192 787056 707870 787106
rect 707926 787056 708000 787112
rect 700192 787050 708000 787056
rect 699322 786988 708000 787050
rect 699322 786982 707870 786988
rect 699322 786926 699392 786982
rect 699448 786926 699516 786982
rect 699572 786926 699640 786982
rect 699696 786926 699764 786982
rect 699820 786926 699888 786982
rect 699944 786926 700012 786982
rect 700068 786926 700136 786982
rect 700192 786932 707870 786982
rect 707926 786932 708000 786988
rect 700192 786926 708000 786932
rect 699322 786864 708000 786926
rect 699322 786858 707870 786864
rect 699322 786802 699392 786858
rect 699448 786802 699516 786858
rect 699572 786802 699640 786858
rect 699696 786802 699764 786858
rect 699820 786802 699888 786858
rect 699944 786802 700012 786858
rect 700068 786802 700136 786858
rect 700192 786808 707870 786858
rect 707926 786808 708000 786864
rect 700192 786802 708000 786808
rect 699322 786740 708000 786802
rect 699322 786734 707870 786740
rect 699322 786678 699392 786734
rect 699448 786678 699516 786734
rect 699572 786678 699640 786734
rect 699696 786678 699764 786734
rect 699820 786678 699888 786734
rect 699944 786678 700012 786734
rect 700068 786678 700136 786734
rect 700192 786684 707870 786734
rect 707926 786684 708000 786740
rect 700192 786678 708000 786684
rect 699322 786616 708000 786678
rect 699322 786610 707870 786616
rect 699322 786554 699392 786610
rect 699448 786554 699516 786610
rect 699572 786554 699640 786610
rect 699696 786554 699764 786610
rect 699820 786554 699888 786610
rect 699944 786554 700012 786610
rect 700068 786554 700136 786610
rect 700192 786560 707870 786610
rect 707926 786560 708000 786616
rect 700192 786554 708000 786560
rect 699322 786492 708000 786554
rect 699322 786486 707870 786492
rect 699322 786430 699392 786486
rect 699448 786430 699516 786486
rect 699572 786430 699640 786486
rect 699696 786430 699764 786486
rect 699820 786430 699888 786486
rect 699944 786430 700012 786486
rect 700068 786430 700136 786486
rect 700192 786436 707870 786486
rect 707926 786436 708000 786492
rect 700192 786430 708000 786436
rect 699322 786368 708000 786430
rect 699322 786362 707870 786368
rect 699322 786306 699392 786362
rect 699448 786306 699516 786362
rect 699572 786306 699640 786362
rect 699696 786306 699764 786362
rect 699820 786306 699888 786362
rect 699944 786306 700012 786362
rect 700068 786306 700136 786362
rect 700192 786312 707870 786362
rect 707926 786312 708000 786368
rect 700192 786306 708000 786312
rect 699322 786244 708000 786306
rect 699322 786238 707870 786244
rect 699322 786182 699392 786238
rect 699448 786182 699516 786238
rect 699572 786182 699640 786238
rect 699696 786182 699764 786238
rect 699820 786182 699888 786238
rect 699944 786182 700012 786238
rect 700068 786182 700136 786238
rect 700192 786188 707870 786238
rect 707926 786188 708000 786244
rect 700192 786182 708000 786188
rect 699322 786120 708000 786182
rect 699322 786114 707870 786120
rect 699322 786058 699392 786114
rect 699448 786058 699516 786114
rect 699572 786058 699640 786114
rect 699696 786058 699764 786114
rect 699820 786058 699888 786114
rect 699944 786058 700012 786114
rect 700068 786058 700136 786114
rect 700192 786064 707870 786114
rect 707926 786064 708000 786120
rect 700192 786058 708000 786064
rect 699322 785996 708000 786058
rect 699322 785990 707870 785996
rect 699322 785934 699392 785990
rect 699448 785934 699516 785990
rect 699572 785934 699640 785990
rect 699696 785934 699764 785990
rect 699820 785934 699888 785990
rect 699944 785934 700012 785990
rect 700068 785934 700136 785990
rect 700192 785940 707870 785990
rect 707926 785940 708000 785996
rect 700192 785934 708000 785940
rect 699322 785872 708000 785934
rect 699322 785866 707870 785872
rect 699322 785810 699392 785866
rect 699448 785810 699516 785866
rect 699572 785810 699640 785866
rect 699696 785810 699764 785866
rect 699820 785810 699888 785866
rect 699944 785810 700012 785866
rect 700068 785810 700136 785866
rect 700192 785816 707870 785866
rect 707926 785816 708000 785872
rect 700192 785810 708000 785816
rect 699322 785752 708000 785810
rect 699322 785134 708000 785172
rect 699322 785122 707870 785134
rect 699322 785066 699392 785122
rect 699448 785066 699516 785122
rect 699572 785066 699640 785122
rect 699696 785066 699764 785122
rect 699820 785066 699888 785122
rect 699944 785066 700012 785122
rect 700068 785066 700136 785122
rect 700192 785078 707870 785122
rect 707926 785078 708000 785134
rect 700192 785066 708000 785078
rect 699322 785010 708000 785066
rect 699322 784998 707870 785010
rect 699322 784942 699392 784998
rect 699448 784942 699516 784998
rect 699572 784942 699640 784998
rect 699696 784942 699764 784998
rect 699820 784942 699888 784998
rect 699944 784942 700012 784998
rect 700068 784942 700136 784998
rect 700192 784954 707870 784998
rect 707926 784954 708000 785010
rect 700192 784942 708000 784954
rect 699322 784886 708000 784942
rect 699322 784874 707870 784886
rect 699322 784818 699392 784874
rect 699448 784818 699516 784874
rect 699572 784818 699640 784874
rect 699696 784818 699764 784874
rect 699820 784818 699888 784874
rect 699944 784818 700012 784874
rect 700068 784818 700136 784874
rect 700192 784830 707870 784874
rect 707926 784830 708000 784886
rect 700192 784818 708000 784830
rect 699322 784762 708000 784818
rect 699322 784750 707870 784762
rect 699322 784694 699392 784750
rect 699448 784694 699516 784750
rect 699572 784694 699640 784750
rect 699696 784694 699764 784750
rect 699820 784694 699888 784750
rect 699944 784694 700012 784750
rect 700068 784694 700136 784750
rect 700192 784706 707870 784750
rect 707926 784706 708000 784762
rect 700192 784694 708000 784706
rect 699322 784638 708000 784694
rect 699322 784626 707870 784638
rect 699322 784570 699392 784626
rect 699448 784570 699516 784626
rect 699572 784570 699640 784626
rect 699696 784570 699764 784626
rect 699820 784570 699888 784626
rect 699944 784570 700012 784626
rect 700068 784570 700136 784626
rect 700192 784582 707870 784626
rect 707926 784582 708000 784638
rect 700192 784570 708000 784582
rect 699322 784514 708000 784570
rect 699322 784502 707870 784514
rect 699322 784446 699392 784502
rect 699448 784446 699516 784502
rect 699572 784446 699640 784502
rect 699696 784446 699764 784502
rect 699820 784446 699888 784502
rect 699944 784446 700012 784502
rect 700068 784446 700136 784502
rect 700192 784458 707870 784502
rect 707926 784458 708000 784514
rect 700192 784446 708000 784458
rect 699322 784390 708000 784446
rect 699322 784378 707870 784390
rect 699322 784322 699392 784378
rect 699448 784322 699516 784378
rect 699572 784322 699640 784378
rect 699696 784322 699764 784378
rect 699820 784322 699888 784378
rect 699944 784322 700012 784378
rect 700068 784322 700136 784378
rect 700192 784334 707870 784378
rect 707926 784334 708000 784390
rect 700192 784322 708000 784334
rect 699322 784266 708000 784322
rect 699322 784254 707870 784266
rect 699322 784198 699392 784254
rect 699448 784198 699516 784254
rect 699572 784198 699640 784254
rect 699696 784198 699764 784254
rect 699820 784198 699888 784254
rect 699944 784198 700012 784254
rect 700068 784198 700136 784254
rect 700192 784210 707870 784254
rect 707926 784210 708000 784266
rect 700192 784198 708000 784210
rect 699322 784142 708000 784198
rect 699322 784130 707870 784142
rect 699322 784074 699392 784130
rect 699448 784074 699516 784130
rect 699572 784074 699640 784130
rect 699696 784074 699764 784130
rect 699820 784074 699888 784130
rect 699944 784074 700012 784130
rect 700068 784074 700136 784130
rect 700192 784086 707870 784130
rect 707926 784086 708000 784142
rect 700192 784074 708000 784086
rect 699322 784018 708000 784074
rect 699322 784006 707870 784018
rect 699322 783950 699392 784006
rect 699448 783950 699516 784006
rect 699572 783950 699640 784006
rect 699696 783950 699764 784006
rect 699820 783950 699888 784006
rect 699944 783950 700012 784006
rect 700068 783950 700136 784006
rect 700192 783962 707870 784006
rect 707926 783962 708000 784018
rect 700192 783950 708000 783962
rect 699322 783894 708000 783950
rect 699322 783882 707870 783894
rect 699322 783826 699392 783882
rect 699448 783826 699516 783882
rect 699572 783826 699640 783882
rect 699696 783826 699764 783882
rect 699820 783826 699888 783882
rect 699944 783826 700012 783882
rect 700068 783826 700136 783882
rect 700192 783838 707870 783882
rect 707926 783838 708000 783894
rect 700192 783826 708000 783838
rect 699322 783770 708000 783826
rect 699322 783758 707870 783770
rect 699322 783702 699392 783758
rect 699448 783702 699516 783758
rect 699572 783702 699640 783758
rect 699696 783702 699764 783758
rect 699820 783702 699888 783758
rect 699944 783702 700012 783758
rect 700068 783702 700136 783758
rect 700192 783714 707870 783758
rect 707926 783714 708000 783770
rect 700192 783702 708000 783714
rect 699322 783646 708000 783702
rect 699322 783634 707870 783646
rect 699322 783578 699392 783634
rect 699448 783578 699516 783634
rect 699572 783578 699640 783634
rect 699696 783578 699764 783634
rect 699820 783578 699888 783634
rect 699944 783578 700012 783634
rect 700068 783578 700136 783634
rect 700192 783590 707870 783634
rect 707926 783590 708000 783646
rect 700192 783578 708000 783590
rect 699322 783522 708000 783578
rect 699322 783510 707870 783522
rect 699322 783454 699392 783510
rect 699448 783454 699516 783510
rect 699572 783454 699640 783510
rect 699696 783454 699764 783510
rect 699820 783454 699888 783510
rect 699944 783454 700012 783510
rect 700068 783454 700136 783510
rect 700192 783466 707870 783510
rect 707926 783466 708000 783522
rect 700192 783454 708000 783466
rect 699322 783398 708000 783454
rect 699322 783386 707870 783398
rect 699322 783330 699392 783386
rect 699448 783330 699516 783386
rect 699572 783330 699640 783386
rect 699696 783330 699764 783386
rect 699820 783330 699888 783386
rect 699944 783330 700012 783386
rect 700068 783330 700136 783386
rect 700192 783342 707870 783386
rect 707926 783342 708000 783398
rect 700192 783330 708000 783342
rect 699322 783272 708000 783330
rect 76115 782048 80078 782110
rect 76115 781992 79284 782048
rect 79340 781992 79584 782048
rect 79640 781992 79884 782048
rect 79940 781992 80078 782048
rect 76115 781910 80078 781992
rect 76115 781510 76435 781910
rect 76915 781633 78678 781710
rect 76915 781577 77847 781633
rect 77903 781577 78147 781633
rect 78203 781577 78447 781633
rect 78503 781577 78678 781633
rect 76915 781510 78678 781577
rect 77678 770429 84516 770630
rect 77678 770373 77800 770429
rect 77856 770373 78100 770429
rect 78156 770373 78400 770429
rect 78456 770373 84516 770429
rect 77678 770229 84516 770373
rect 77678 770173 77800 770229
rect 77856 770173 78100 770229
rect 78156 770173 78400 770229
rect 78456 770173 84516 770229
rect 77678 770010 84516 770173
rect 687412 770429 700322 770630
rect 687412 770373 699544 770429
rect 699600 770373 699844 770429
rect 699900 770373 700144 770429
rect 700200 770373 700322 770429
rect 687412 770229 700322 770373
rect 687412 770173 699544 770229
rect 699600 770173 699844 770229
rect 699900 770173 700144 770229
rect 700200 770173 700322 770229
rect 687412 770010 700322 770173
rect 75376 765622 80078 765744
rect 75376 765566 79300 765622
rect 79356 765566 79600 765622
rect 79656 765566 79900 765622
rect 79956 765566 80078 765622
rect 75376 765424 80078 765566
rect 75312 762102 78678 762244
rect 75312 762046 77900 762102
rect 77956 762046 78200 762102
rect 78256 762046 78500 762102
rect 78556 762046 78678 762102
rect 75312 761924 78678 762046
rect 75376 758622 80078 758744
rect 75376 758566 79300 758622
rect 79356 758566 79600 758622
rect 79656 758566 79900 758622
rect 79956 758566 80078 758622
rect 75376 758424 80078 758566
rect 75312 755102 78678 755244
rect 75312 755046 77900 755102
rect 77956 755046 78200 755102
rect 78256 755046 78500 755102
rect 78556 755046 78678 755102
rect 75312 754924 78678 755046
rect 699322 753954 702688 754076
rect 699322 753898 699444 753954
rect 699500 753898 699744 753954
rect 699800 753898 700044 753954
rect 700100 753898 702688 753954
rect 699322 753756 702688 753898
rect 79078 752429 83556 752630
rect 79078 752373 79200 752429
rect 79256 752373 79500 752429
rect 79556 752373 79800 752429
rect 79856 752373 83556 752429
rect 79078 752229 83556 752373
rect 79078 752173 79200 752229
rect 79256 752173 79500 752229
rect 79556 752173 79800 752229
rect 79856 752173 83556 752229
rect 79078 752010 83556 752173
rect 688372 752429 698922 752630
rect 688372 752373 698144 752429
rect 698200 752373 698444 752429
rect 698500 752373 698744 752429
rect 698800 752373 698922 752429
rect 688372 752229 698922 752373
rect 688372 752173 698144 752229
rect 698200 752173 698444 752229
rect 698500 752173 698744 752229
rect 698800 752173 698922 752229
rect 688372 752010 698922 752173
rect 75376 751622 80078 751744
rect 75376 751566 79300 751622
rect 79356 751566 79600 751622
rect 79656 751566 79900 751622
rect 79956 751566 80078 751622
rect 75376 751424 80078 751566
rect 697922 750434 702624 750576
rect 697922 750378 698044 750434
rect 698100 750378 698344 750434
rect 698400 750378 698644 750434
rect 698700 750378 702624 750434
rect 697922 750256 702624 750378
rect 75312 748102 78678 748244
rect 75312 748046 77900 748102
rect 77956 748046 78200 748102
rect 78256 748046 78500 748102
rect 78556 748046 78678 748102
rect 75312 747924 78678 748046
rect 699322 746954 702688 747076
rect 699322 746898 699444 746954
rect 699500 746898 699744 746954
rect 699800 746898 700044 746954
rect 700100 746898 702688 746954
rect 699322 746756 702688 746898
rect 697922 743434 702624 743576
rect 697922 743378 698044 743434
rect 698100 743378 698344 743434
rect 698400 743378 698644 743434
rect 698700 743378 702624 743434
rect 697922 743256 702624 743378
rect 76115 741048 80078 741110
rect 76115 740992 79284 741048
rect 79340 740992 79584 741048
rect 79640 740992 79884 741048
rect 79940 740992 80078 741048
rect 76115 740910 80078 740992
rect 76115 740510 76435 740910
rect 76915 740633 78678 740710
rect 76915 740577 77847 740633
rect 77903 740577 78147 740633
rect 78203 740577 78447 740633
rect 78503 740577 78678 740633
rect 76915 740510 78678 740577
rect 699322 739954 702688 740076
rect 699322 739898 699444 739954
rect 699500 739898 699744 739954
rect 699800 739898 700044 739954
rect 700100 739898 702688 739954
rect 699322 739756 702688 739898
rect 697922 736434 702624 736576
rect 697922 736378 698044 736434
rect 698100 736378 698344 736434
rect 698400 736378 698644 736434
rect 698700 736378 702624 736434
rect 697922 736256 702624 736378
rect 77678 734429 84516 734630
rect 77678 734373 77800 734429
rect 77856 734373 78100 734429
rect 78156 734373 78400 734429
rect 78456 734373 84516 734429
rect 77678 734229 84516 734373
rect 77678 734173 77800 734229
rect 77856 734173 78100 734229
rect 78156 734173 78400 734229
rect 78456 734173 84516 734229
rect 77678 734010 84516 734173
rect 687412 734429 700322 734630
rect 687412 734373 699544 734429
rect 699600 734373 699844 734429
rect 699900 734373 700144 734429
rect 700200 734373 700322 734429
rect 687412 734229 700322 734373
rect 687412 734173 699544 734229
rect 699600 734173 699844 734229
rect 699900 734173 700144 734229
rect 700200 734173 700322 734229
rect 687412 734010 700322 734173
rect 75376 724622 80078 724744
rect 75376 724566 79300 724622
rect 79356 724566 79600 724622
rect 79656 724566 79900 724622
rect 79956 724566 80078 724622
rect 75376 724424 80078 724566
rect 75312 721102 78678 721244
rect 75312 721046 77900 721102
rect 77956 721046 78200 721102
rect 78256 721046 78500 721102
rect 78556 721046 78678 721102
rect 75312 720924 78678 721046
rect 699322 720423 701085 720490
rect 699322 720367 699497 720423
rect 699553 720367 699797 720423
rect 699853 720367 700097 720423
rect 700153 720367 701085 720423
rect 699322 720290 701085 720367
rect 701565 720090 701885 720490
rect 697922 720008 701885 720090
rect 697922 719952 698060 720008
rect 698116 719952 698360 720008
rect 698416 719952 698660 720008
rect 698716 719952 701885 720008
rect 697922 719890 701885 719952
rect 75376 717622 80078 717744
rect 75376 717566 79300 717622
rect 79356 717566 79600 717622
rect 79656 717566 79900 717622
rect 79956 717566 80078 717622
rect 75376 717424 80078 717566
rect 79078 716429 83556 716630
rect 79078 716373 79200 716429
rect 79256 716373 79500 716429
rect 79556 716373 79800 716429
rect 79856 716373 83556 716429
rect 79078 716229 83556 716373
rect 79078 716173 79200 716229
rect 79256 716173 79500 716229
rect 79556 716173 79800 716229
rect 79856 716173 83556 716229
rect 79078 716010 83556 716173
rect 688372 716429 698922 716630
rect 688372 716373 698144 716429
rect 698200 716373 698444 716429
rect 698500 716373 698744 716429
rect 698800 716373 698922 716429
rect 688372 716229 698922 716373
rect 688372 716173 698144 716229
rect 698200 716173 698444 716229
rect 698500 716173 698744 716229
rect 698800 716173 698922 716229
rect 688372 716010 698922 716173
rect 75312 714102 78678 714244
rect 75312 714046 77900 714102
rect 77956 714046 78200 714102
rect 78256 714046 78500 714102
rect 78556 714046 78678 714102
rect 75312 713924 78678 714046
rect 699322 710954 702688 711076
rect 699322 710898 699444 710954
rect 699500 710898 699744 710954
rect 699800 710898 700044 710954
rect 700100 710898 702688 710954
rect 699322 710756 702688 710898
rect 75376 710622 80078 710744
rect 75376 710566 79300 710622
rect 79356 710566 79600 710622
rect 79656 710566 79900 710622
rect 79956 710566 80078 710622
rect 75376 710424 80078 710566
rect 697922 707434 702624 707576
rect 697922 707378 698044 707434
rect 698100 707378 698344 707434
rect 698400 707378 698644 707434
rect 698700 707378 702624 707434
rect 697922 707256 702624 707378
rect 75312 707102 78678 707244
rect 75312 707046 77900 707102
rect 77956 707046 78200 707102
rect 78256 707046 78500 707102
rect 78556 707046 78678 707102
rect 75312 706924 78678 707046
rect 699322 703954 702688 704076
rect 699322 703898 699444 703954
rect 699500 703898 699744 703954
rect 699800 703898 700044 703954
rect 700100 703898 702688 703954
rect 699322 703756 702688 703898
rect 697922 700434 702624 700576
rect 697922 700378 698044 700434
rect 698100 700378 698344 700434
rect 698400 700378 698644 700434
rect 698700 700378 702624 700434
rect 697922 700256 702624 700378
rect 76115 700048 80078 700110
rect 76115 699992 79284 700048
rect 79340 699992 79584 700048
rect 79640 699992 79884 700048
rect 79940 699992 80078 700048
rect 76115 699910 80078 699992
rect 76115 699510 76435 699910
rect 76915 699633 78678 699710
rect 76915 699577 77847 699633
rect 77903 699577 78147 699633
rect 78203 699577 78447 699633
rect 78503 699577 78678 699633
rect 76915 699510 78678 699577
rect 77678 698429 84516 698630
rect 77678 698373 77800 698429
rect 77856 698373 78100 698429
rect 78156 698373 78400 698429
rect 78456 698373 84516 698429
rect 77678 698229 84516 698373
rect 77678 698173 77800 698229
rect 77856 698173 78100 698229
rect 78156 698173 78400 698229
rect 78456 698173 84516 698229
rect 77678 698010 84516 698173
rect 687412 698429 700322 698630
rect 687412 698373 699544 698429
rect 699600 698373 699844 698429
rect 699900 698373 700144 698429
rect 700200 698373 700322 698429
rect 687412 698229 700322 698373
rect 687412 698173 699544 698229
rect 699600 698173 699844 698229
rect 699900 698173 700144 698229
rect 700200 698173 700322 698229
rect 687412 698010 700322 698173
rect 699322 696954 702688 697076
rect 699322 696898 699444 696954
rect 699500 696898 699744 696954
rect 699800 696898 700044 696954
rect 700100 696898 702688 696954
rect 699322 696756 702688 696898
rect 697922 693434 702624 693576
rect 697922 693378 698044 693434
rect 698100 693378 698344 693434
rect 698400 693378 698644 693434
rect 698700 693378 702624 693434
rect 697922 693256 702624 693378
rect 75376 683622 80078 683744
rect 75376 683566 79300 683622
rect 79356 683566 79600 683622
rect 79656 683566 79900 683622
rect 79956 683566 80078 683622
rect 75376 683424 80078 683566
rect 79078 680429 83556 680630
rect 79078 680373 79200 680429
rect 79256 680373 79500 680429
rect 79556 680373 79800 680429
rect 79856 680373 83556 680429
rect 75312 680102 78678 680244
rect 75312 680046 77900 680102
rect 77956 680046 78200 680102
rect 78256 680046 78500 680102
rect 78556 680046 78678 680102
rect 75312 679924 78678 680046
rect 79078 680229 83556 680373
rect 79078 680173 79200 680229
rect 79256 680173 79500 680229
rect 79556 680173 79800 680229
rect 79856 680173 83556 680229
rect 79078 680010 83556 680173
rect 688372 680429 698922 680630
rect 688372 680373 698144 680429
rect 698200 680373 698444 680429
rect 698500 680373 698744 680429
rect 698800 680373 698922 680429
rect 688372 680229 698922 680373
rect 688372 680173 698144 680229
rect 698200 680173 698444 680229
rect 698500 680173 698744 680229
rect 698800 680173 698922 680229
rect 688372 680010 698922 680173
rect 699322 677423 701085 677490
rect 699322 677367 699497 677423
rect 699553 677367 699797 677423
rect 699853 677367 700097 677423
rect 700153 677367 701085 677423
rect 699322 677290 701085 677367
rect 701565 677090 701885 677490
rect 697922 677008 701885 677090
rect 697922 676952 698060 677008
rect 698116 676952 698360 677008
rect 698416 676952 698660 677008
rect 698716 676952 701885 677008
rect 697922 676890 701885 676952
rect 75376 676622 80078 676744
rect 75376 676566 79300 676622
rect 79356 676566 79600 676622
rect 79656 676566 79900 676622
rect 79956 676566 80078 676622
rect 75376 676424 80078 676566
rect 75312 673102 78678 673244
rect 75312 673046 77900 673102
rect 77956 673046 78200 673102
rect 78256 673046 78500 673102
rect 78556 673046 78678 673102
rect 75312 672924 78678 673046
rect 75376 669622 80078 669744
rect 75376 669566 79300 669622
rect 79356 669566 79600 669622
rect 79656 669566 79900 669622
rect 79956 669566 80078 669622
rect 75376 669424 80078 669566
rect 699322 667954 702688 668076
rect 699322 667898 699444 667954
rect 699500 667898 699744 667954
rect 699800 667898 700044 667954
rect 700100 667898 702688 667954
rect 699322 667756 702688 667898
rect 75312 666102 78678 666244
rect 75312 666046 77900 666102
rect 77956 666046 78200 666102
rect 78256 666046 78500 666102
rect 78556 666046 78678 666102
rect 75312 665924 78678 666046
rect 697922 664434 702624 664576
rect 697922 664378 698044 664434
rect 698100 664378 698344 664434
rect 698400 664378 698644 664434
rect 698700 664378 702624 664434
rect 697922 664256 702624 664378
rect 77678 662429 84516 662630
rect 77678 662373 77800 662429
rect 77856 662373 78100 662429
rect 78156 662373 78400 662429
rect 78456 662373 84516 662429
rect 77678 662229 84516 662373
rect 77678 662173 77800 662229
rect 77856 662173 78100 662229
rect 78156 662173 78400 662229
rect 78456 662173 84516 662229
rect 77678 662010 84516 662173
rect 687412 662429 700322 662630
rect 687412 662373 699544 662429
rect 699600 662373 699844 662429
rect 699900 662373 700144 662429
rect 700200 662373 700322 662429
rect 687412 662229 700322 662373
rect 687412 662173 699544 662229
rect 699600 662173 699844 662229
rect 699900 662173 700144 662229
rect 700200 662173 700322 662229
rect 687412 662010 700322 662173
rect 699322 660954 702688 661076
rect 699322 660898 699444 660954
rect 699500 660898 699744 660954
rect 699800 660898 700044 660954
rect 700100 660898 702688 660954
rect 699322 660756 702688 660898
rect 76115 659048 80078 659110
rect 76115 658992 79284 659048
rect 79340 658992 79584 659048
rect 79640 658992 79884 659048
rect 79940 658992 80078 659048
rect 76115 658910 80078 658992
rect 76115 658510 76435 658910
rect 76915 658633 78678 658710
rect 76915 658577 77847 658633
rect 77903 658577 78147 658633
rect 78203 658577 78447 658633
rect 78503 658577 78678 658633
rect 76915 658510 78678 658577
rect 697922 657434 702624 657576
rect 697922 657378 698044 657434
rect 698100 657378 698344 657434
rect 698400 657378 698644 657434
rect 698700 657378 702624 657434
rect 697922 657256 702624 657378
rect 699322 653954 702688 654076
rect 699322 653898 699444 653954
rect 699500 653898 699744 653954
rect 699800 653898 700044 653954
rect 700100 653898 702688 653954
rect 699322 653756 702688 653898
rect 697922 650434 702624 650576
rect 697922 650378 698044 650434
rect 698100 650378 698344 650434
rect 698400 650378 698644 650434
rect 698700 650378 702624 650434
rect 697922 650256 702624 650378
rect 79078 644429 83556 644630
rect 79078 644373 79200 644429
rect 79256 644373 79500 644429
rect 79556 644373 79800 644429
rect 79856 644373 83556 644429
rect 79078 644229 83556 644373
rect 79078 644173 79200 644229
rect 79256 644173 79500 644229
rect 79556 644173 79800 644229
rect 79856 644173 83556 644229
rect 79078 644010 83556 644173
rect 688372 644429 698922 644630
rect 688372 644373 698144 644429
rect 698200 644373 698444 644429
rect 698500 644373 698744 644429
rect 698800 644373 698922 644429
rect 688372 644229 698922 644373
rect 688372 644173 698144 644229
rect 698200 644173 698444 644229
rect 698500 644173 698744 644229
rect 698800 644173 698922 644229
rect 688372 644010 698922 644173
rect 75376 642622 80078 642744
rect 75376 642566 79300 642622
rect 79356 642566 79600 642622
rect 79656 642566 79900 642622
rect 79956 642566 80078 642622
rect 75376 642424 80078 642566
rect 75312 639102 78678 639244
rect 75312 639046 77900 639102
rect 77956 639046 78200 639102
rect 78256 639046 78500 639102
rect 78556 639046 78678 639102
rect 75312 638924 78678 639046
rect 75376 635622 80078 635744
rect 75376 635566 79300 635622
rect 79356 635566 79600 635622
rect 79656 635566 79900 635622
rect 79956 635566 80078 635622
rect 75376 635424 80078 635566
rect 699322 634423 701085 634490
rect 699322 634367 699497 634423
rect 699553 634367 699797 634423
rect 699853 634367 700097 634423
rect 700153 634367 701085 634423
rect 699322 634290 701085 634367
rect 701565 634090 701885 634490
rect 697922 634008 701885 634090
rect 697922 633952 698060 634008
rect 698116 633952 698360 634008
rect 698416 633952 698660 634008
rect 698716 633952 701885 634008
rect 697922 633890 701885 633952
rect 75312 632102 78678 632244
rect 75312 632046 77900 632102
rect 77956 632046 78200 632102
rect 78256 632046 78500 632102
rect 78556 632046 78678 632102
rect 75312 631924 78678 632046
rect 75376 628622 80078 628744
rect 75376 628566 79300 628622
rect 79356 628566 79600 628622
rect 79656 628566 79900 628622
rect 79956 628566 80078 628622
rect 75376 628424 80078 628566
rect 77678 626429 84516 626630
rect 77678 626373 77800 626429
rect 77856 626373 78100 626429
rect 78156 626373 78400 626429
rect 78456 626373 84516 626429
rect 77678 626229 84516 626373
rect 77678 626173 77800 626229
rect 77856 626173 78100 626229
rect 78156 626173 78400 626229
rect 78456 626173 84516 626229
rect 77678 626010 84516 626173
rect 687412 626429 700322 626630
rect 687412 626373 699544 626429
rect 699600 626373 699844 626429
rect 699900 626373 700144 626429
rect 700200 626373 700322 626429
rect 687412 626229 700322 626373
rect 687412 626173 699544 626229
rect 699600 626173 699844 626229
rect 699900 626173 700144 626229
rect 700200 626173 700322 626229
rect 687412 626010 700322 626173
rect 75312 625102 78678 625244
rect 75312 625046 77900 625102
rect 77956 625046 78200 625102
rect 78256 625046 78500 625102
rect 78556 625046 78678 625102
rect 75312 624924 78678 625046
rect 699322 624954 702688 625076
rect 699322 624898 699444 624954
rect 699500 624898 699744 624954
rect 699800 624898 700044 624954
rect 700100 624898 702688 624954
rect 699322 624756 702688 624898
rect 697922 621434 702624 621576
rect 697922 621378 698044 621434
rect 698100 621378 698344 621434
rect 698400 621378 698644 621434
rect 698700 621378 702624 621434
rect 697922 621256 702624 621378
rect 76115 618048 80078 618110
rect 76115 617992 79284 618048
rect 79340 617992 79584 618048
rect 79640 617992 79884 618048
rect 79940 617992 80078 618048
rect 76115 617910 80078 617992
rect 699322 617954 702688 618076
rect 76115 617510 76435 617910
rect 699322 617898 699444 617954
rect 699500 617898 699744 617954
rect 699800 617898 700044 617954
rect 700100 617898 702688 617954
rect 699322 617756 702688 617898
rect 76915 617633 78678 617710
rect 76915 617577 77847 617633
rect 77903 617577 78147 617633
rect 78203 617577 78447 617633
rect 78503 617577 78678 617633
rect 76915 617510 78678 617577
rect 697922 614434 702624 614576
rect 697922 614378 698044 614434
rect 698100 614378 698344 614434
rect 698400 614378 698644 614434
rect 698700 614378 702624 614434
rect 697922 614256 702624 614378
rect 699322 610954 702688 611076
rect 699322 610898 699444 610954
rect 699500 610898 699744 610954
rect 699800 610898 700044 610954
rect 700100 610898 702688 610954
rect 699322 610756 702688 610898
rect 79078 608429 83556 608630
rect 79078 608373 79200 608429
rect 79256 608373 79500 608429
rect 79556 608373 79800 608429
rect 79856 608373 83556 608429
rect 79078 608229 83556 608373
rect 79078 608173 79200 608229
rect 79256 608173 79500 608229
rect 79556 608173 79800 608229
rect 79856 608173 83556 608229
rect 79078 608010 83556 608173
rect 688372 608429 698922 608630
rect 688372 608373 698144 608429
rect 698200 608373 698444 608429
rect 698500 608373 698744 608429
rect 698800 608373 698922 608429
rect 688372 608229 698922 608373
rect 688372 608173 698144 608229
rect 698200 608173 698444 608229
rect 698500 608173 698744 608229
rect 698800 608173 698922 608229
rect 688372 608010 698922 608173
rect 697922 607434 702624 607576
rect 697922 607378 698044 607434
rect 698100 607378 698344 607434
rect 698400 607378 698644 607434
rect 698700 607378 702624 607434
rect 697922 607256 702624 607378
rect 75376 601622 80078 601744
rect 75376 601566 79300 601622
rect 79356 601566 79600 601622
rect 79656 601566 79900 601622
rect 79956 601566 80078 601622
rect 75376 601424 80078 601566
rect 75312 598102 78678 598244
rect 75312 598046 77900 598102
rect 77956 598046 78200 598102
rect 78256 598046 78500 598102
rect 78556 598046 78678 598102
rect 75312 597924 78678 598046
rect 75376 594622 80078 594744
rect 75376 594566 79300 594622
rect 79356 594566 79600 594622
rect 79656 594566 79900 594622
rect 79956 594566 80078 594622
rect 75376 594424 80078 594566
rect 699322 591423 701085 591490
rect 699322 591367 699497 591423
rect 699553 591367 699797 591423
rect 699853 591367 700097 591423
rect 700153 591367 701085 591423
rect 699322 591290 701085 591367
rect 75312 591102 78678 591244
rect 75312 591046 77900 591102
rect 77956 591046 78200 591102
rect 78256 591046 78500 591102
rect 78556 591046 78678 591102
rect 701565 591090 701885 591490
rect 75312 590924 78678 591046
rect 697922 591008 701885 591090
rect 697922 590952 698060 591008
rect 698116 590952 698360 591008
rect 698416 590952 698660 591008
rect 698716 590952 701885 591008
rect 697922 590890 701885 590952
rect 77678 590429 84516 590630
rect 77678 590373 77800 590429
rect 77856 590373 78100 590429
rect 78156 590373 78400 590429
rect 78456 590373 84516 590429
rect 77678 590229 84516 590373
rect 77678 590173 77800 590229
rect 77856 590173 78100 590229
rect 78156 590173 78400 590229
rect 78456 590173 84516 590229
rect 77678 590010 84516 590173
rect 687412 590429 700322 590630
rect 687412 590373 699544 590429
rect 699600 590373 699844 590429
rect 699900 590373 700144 590429
rect 700200 590373 700322 590429
rect 687412 590229 700322 590373
rect 687412 590173 699544 590229
rect 699600 590173 699844 590229
rect 699900 590173 700144 590229
rect 700200 590173 700322 590229
rect 687412 590010 700322 590173
rect 75376 587622 80078 587744
rect 75376 587566 79300 587622
rect 79356 587566 79600 587622
rect 79656 587566 79900 587622
rect 79956 587566 80078 587622
rect 75376 587424 80078 587566
rect 75312 584102 78678 584244
rect 75312 584046 77900 584102
rect 77956 584046 78200 584102
rect 78256 584046 78500 584102
rect 78556 584046 78678 584102
rect 75312 583924 78678 584046
rect 699322 581954 702688 582076
rect 699322 581898 699444 581954
rect 699500 581898 699744 581954
rect 699800 581898 700044 581954
rect 700100 581898 702688 581954
rect 699322 581756 702688 581898
rect 697922 578434 702624 578576
rect 697922 578378 698044 578434
rect 698100 578378 698344 578434
rect 698400 578378 698644 578434
rect 698700 578378 702624 578434
rect 697922 578256 702624 578378
rect 76115 577048 80078 577110
rect 76115 576992 79284 577048
rect 79340 576992 79584 577048
rect 79640 576992 79884 577048
rect 79940 576992 80078 577048
rect 76115 576910 80078 576992
rect 76115 576510 76435 576910
rect 76915 576633 78678 576710
rect 76915 576577 77847 576633
rect 77903 576577 78147 576633
rect 78203 576577 78447 576633
rect 78503 576577 78678 576633
rect 76915 576510 78678 576577
rect 699322 574954 702688 575076
rect 699322 574898 699444 574954
rect 699500 574898 699744 574954
rect 699800 574898 700044 574954
rect 700100 574898 702688 574954
rect 699322 574756 702688 574898
rect 79078 572429 83556 572630
rect 79078 572373 79200 572429
rect 79256 572373 79500 572429
rect 79556 572373 79800 572429
rect 79856 572373 83556 572429
rect 79078 572229 83556 572373
rect 79078 572173 79200 572229
rect 79256 572173 79500 572229
rect 79556 572173 79800 572229
rect 79856 572173 83556 572229
rect 79078 572010 83556 572173
rect 688372 572429 698922 572630
rect 688372 572373 698144 572429
rect 698200 572373 698444 572429
rect 698500 572373 698744 572429
rect 698800 572373 698922 572429
rect 688372 572229 698922 572373
rect 688372 572173 698144 572229
rect 698200 572173 698444 572229
rect 698500 572173 698744 572229
rect 698800 572173 698922 572229
rect 688372 572010 698922 572173
rect 697922 571434 702624 571576
rect 697922 571378 698044 571434
rect 698100 571378 698344 571434
rect 698400 571378 698644 571434
rect 698700 571378 702624 571434
rect 697922 571256 702624 571378
rect 699322 567954 702688 568076
rect 699322 567898 699444 567954
rect 699500 567898 699744 567954
rect 699800 567898 700044 567954
rect 700100 567898 702688 567954
rect 699322 567756 702688 567898
rect 697922 564434 702624 564576
rect 697922 564378 698044 564434
rect 698100 564378 698344 564434
rect 698400 564378 698644 564434
rect 698700 564378 702624 564434
rect 697922 564256 702624 564378
rect 75376 560622 80078 560744
rect 75376 560566 79300 560622
rect 79356 560566 79600 560622
rect 79656 560566 79900 560622
rect 79956 560566 80078 560622
rect 75376 560424 80078 560566
rect 75312 557102 78678 557244
rect 75312 557046 77900 557102
rect 77956 557046 78200 557102
rect 78256 557046 78500 557102
rect 78556 557046 78678 557102
rect 75312 556924 78678 557046
rect 77678 554429 84516 554630
rect 77678 554373 77800 554429
rect 77856 554373 78100 554429
rect 78156 554373 78400 554429
rect 78456 554373 84516 554429
rect 77678 554229 84516 554373
rect 77678 554173 77800 554229
rect 77856 554173 78100 554229
rect 78156 554173 78400 554229
rect 78456 554173 84516 554229
rect 77678 554010 84516 554173
rect 687412 554429 700322 554630
rect 687412 554373 699544 554429
rect 699600 554373 699844 554429
rect 699900 554373 700144 554429
rect 700200 554373 700322 554429
rect 687412 554229 700322 554373
rect 687412 554173 699544 554229
rect 699600 554173 699844 554229
rect 699900 554173 700144 554229
rect 700200 554173 700322 554229
rect 687412 554010 700322 554173
rect 75376 553622 80078 553744
rect 75376 553566 79300 553622
rect 79356 553566 79600 553622
rect 79656 553566 79900 553622
rect 79956 553566 80078 553622
rect 75376 553424 80078 553566
rect 75312 550102 78678 550244
rect 75312 550046 77900 550102
rect 77956 550046 78200 550102
rect 78256 550046 78500 550102
rect 78556 550046 78678 550102
rect 75312 549924 78678 550046
rect 699322 548423 701085 548490
rect 699322 548367 699497 548423
rect 699553 548367 699797 548423
rect 699853 548367 700097 548423
rect 700153 548367 701085 548423
rect 699322 548290 701085 548367
rect 701565 548090 701885 548490
rect 697922 548008 701885 548090
rect 697922 547952 698060 548008
rect 698116 547952 698360 548008
rect 698416 547952 698660 548008
rect 698716 547952 701885 548008
rect 697922 547890 701885 547952
rect 75376 546622 80078 546744
rect 75376 546566 79300 546622
rect 79356 546566 79600 546622
rect 79656 546566 79900 546622
rect 79956 546566 80078 546622
rect 75376 546424 80078 546566
rect 75312 543102 78678 543244
rect 75312 543046 77900 543102
rect 77956 543046 78200 543102
rect 78256 543046 78500 543102
rect 78556 543046 78678 543102
rect 75312 542924 78678 543046
rect 699322 538954 702688 539076
rect 699322 538898 699444 538954
rect 699500 538898 699744 538954
rect 699800 538898 700044 538954
rect 700100 538898 702688 538954
rect 699322 538756 702688 538898
rect 79078 536429 83556 536630
rect 79078 536373 79200 536429
rect 79256 536373 79500 536429
rect 79556 536373 79800 536429
rect 79856 536373 83556 536429
rect 79078 536229 83556 536373
rect 79078 536173 79200 536229
rect 79256 536173 79500 536229
rect 79556 536173 79800 536229
rect 79856 536173 83556 536229
rect 79078 536110 83556 536173
rect 76115 536048 83556 536110
rect 76115 535992 79284 536048
rect 79340 535992 79584 536048
rect 79640 535992 79884 536048
rect 79940 536010 83556 536048
rect 688372 536429 698922 536630
rect 688372 536373 698144 536429
rect 698200 536373 698444 536429
rect 698500 536373 698744 536429
rect 698800 536373 698922 536429
rect 688372 536229 698922 536373
rect 688372 536173 698144 536229
rect 698200 536173 698444 536229
rect 698500 536173 698744 536229
rect 698800 536173 698922 536229
rect 688372 536010 698922 536173
rect 79940 535992 80078 536010
rect 76115 535910 80078 535992
rect 76115 535510 76435 535910
rect 76915 535633 78678 535710
rect 76915 535577 77847 535633
rect 77903 535577 78147 535633
rect 78203 535577 78447 535633
rect 78503 535577 78678 535633
rect 76915 535510 78678 535577
rect 697922 535434 702624 535576
rect 697922 535378 698044 535434
rect 698100 535378 698344 535434
rect 698400 535378 698644 535434
rect 698700 535378 702624 535434
rect 697922 535256 702624 535378
rect 699322 531954 702688 532076
rect 699322 531898 699444 531954
rect 699500 531898 699744 531954
rect 699800 531898 700044 531954
rect 700100 531898 702688 531954
rect 699322 531756 702688 531898
rect 697922 528434 702624 528576
rect 697922 528378 698044 528434
rect 698100 528378 698344 528434
rect 698400 528378 698644 528434
rect 698700 528378 702624 528434
rect 697922 528256 702624 528378
rect 699322 524954 702688 525076
rect 699322 524898 699444 524954
rect 699500 524898 699744 524954
rect 699800 524898 700044 524954
rect 700100 524898 702688 524954
rect 699322 524756 702688 524898
rect 697922 521434 702624 521576
rect 697922 521378 698044 521434
rect 698100 521378 698344 521434
rect 698400 521378 698644 521434
rect 698700 521378 702624 521434
rect 697922 521256 702624 521378
rect 75376 519622 80078 519744
rect 75376 519566 79300 519622
rect 79356 519566 79600 519622
rect 79656 519566 79900 519622
rect 79956 519566 80078 519622
rect 75376 519424 80078 519566
rect 77678 518429 84516 518630
rect 77678 518373 77800 518429
rect 77856 518373 78100 518429
rect 78156 518373 78400 518429
rect 78456 518373 84516 518429
rect 77678 518229 84516 518373
rect 77678 518173 77800 518229
rect 77856 518173 78100 518229
rect 78156 518173 78400 518229
rect 78456 518173 84516 518229
rect 77678 518010 84516 518173
rect 687412 518429 700322 518630
rect 687412 518373 699544 518429
rect 699600 518373 699844 518429
rect 699900 518373 700144 518429
rect 700200 518373 700322 518429
rect 687412 518229 700322 518373
rect 687412 518173 699544 518229
rect 699600 518173 699844 518229
rect 699900 518173 700144 518229
rect 700200 518173 700322 518229
rect 687412 518010 700322 518173
rect 75312 516102 78678 516244
rect 75312 516046 77900 516102
rect 77956 516046 78200 516102
rect 78256 516046 78500 516102
rect 78556 516046 78678 516102
rect 75312 515924 78678 516046
rect 75376 512622 80078 512744
rect 75376 512566 79300 512622
rect 79356 512566 79600 512622
rect 79656 512566 79900 512622
rect 79956 512566 80078 512622
rect 75376 512424 80078 512566
rect 75312 509102 78678 509244
rect 75312 509046 77900 509102
rect 77956 509046 78200 509102
rect 78256 509046 78500 509102
rect 78556 509046 78678 509102
rect 75312 508924 78678 509046
rect 75376 505622 80078 505744
rect 75376 505566 79300 505622
rect 79356 505566 79600 505622
rect 79656 505566 79900 505622
rect 79956 505566 80078 505622
rect 75376 505424 80078 505566
rect 699322 505423 701085 505490
rect 699322 505367 699497 505423
rect 699553 505367 699797 505423
rect 699853 505367 700097 505423
rect 700153 505367 701085 505423
rect 699322 505290 701085 505367
rect 701565 505090 701885 505490
rect 697922 505008 701885 505090
rect 697922 504952 698060 505008
rect 698116 504952 698360 505008
rect 698416 504952 698660 505008
rect 698716 504952 701885 505008
rect 697922 504890 701885 504952
rect 75312 502102 78678 502244
rect 75312 502046 77900 502102
rect 77956 502046 78200 502102
rect 78256 502046 78500 502102
rect 78556 502046 78678 502102
rect 75312 501924 78678 502046
rect 79078 500429 83556 500630
rect 79078 500373 79200 500429
rect 79256 500373 79500 500429
rect 79556 500373 79800 500429
rect 79856 500373 83556 500429
rect 79078 500229 83556 500373
rect 79078 500173 79200 500229
rect 79256 500173 79500 500229
rect 79556 500173 79800 500229
rect 79856 500173 83556 500229
rect 79078 500010 83556 500173
rect 688372 500429 698922 500630
rect 688372 500373 698144 500429
rect 698200 500373 698444 500429
rect 698500 500373 698744 500429
rect 698800 500373 698922 500429
rect 688372 500229 698922 500373
rect 688372 500173 698144 500229
rect 698200 500173 698444 500229
rect 698500 500173 698744 500229
rect 698800 500173 698922 500229
rect 688372 500010 698922 500173
rect 699322 496658 708000 496728
rect 699322 496652 707870 496658
rect 699322 496596 699392 496652
rect 699448 496596 699516 496652
rect 699572 496596 699640 496652
rect 699696 496596 699764 496652
rect 699820 496596 699888 496652
rect 699944 496596 700012 496652
rect 700068 496596 700136 496652
rect 700192 496602 707870 496652
rect 707926 496602 708000 496658
rect 700192 496596 708000 496602
rect 699322 496534 708000 496596
rect 699322 496528 707870 496534
rect 699322 496472 699392 496528
rect 699448 496472 699516 496528
rect 699572 496472 699640 496528
rect 699696 496472 699764 496528
rect 699820 496472 699888 496528
rect 699944 496472 700012 496528
rect 700068 496472 700136 496528
rect 700192 496478 707870 496528
rect 707926 496478 708000 496534
rect 700192 496472 708000 496478
rect 699322 496410 708000 496472
rect 699322 496404 707870 496410
rect 699322 496348 699392 496404
rect 699448 496348 699516 496404
rect 699572 496348 699640 496404
rect 699696 496348 699764 496404
rect 699820 496348 699888 496404
rect 699944 496348 700012 496404
rect 700068 496348 700136 496404
rect 700192 496354 707870 496404
rect 707926 496354 708000 496410
rect 700192 496348 708000 496354
rect 699322 496286 708000 496348
rect 699322 496280 707870 496286
rect 699322 496224 699392 496280
rect 699448 496224 699516 496280
rect 699572 496224 699640 496280
rect 699696 496224 699764 496280
rect 699820 496224 699888 496280
rect 699944 496224 700012 496280
rect 700068 496224 700136 496280
rect 700192 496230 707870 496280
rect 707926 496230 708000 496286
rect 700192 496224 708000 496230
rect 699322 496162 708000 496224
rect 699322 496156 707870 496162
rect 699322 496100 699392 496156
rect 699448 496100 699516 496156
rect 699572 496100 699640 496156
rect 699696 496100 699764 496156
rect 699820 496100 699888 496156
rect 699944 496100 700012 496156
rect 700068 496100 700136 496156
rect 700192 496106 707870 496156
rect 707926 496106 708000 496162
rect 700192 496100 708000 496106
rect 699322 496038 708000 496100
rect 699322 496032 707870 496038
rect 699322 495976 699392 496032
rect 699448 495976 699516 496032
rect 699572 495976 699640 496032
rect 699696 495976 699764 496032
rect 699820 495976 699888 496032
rect 699944 495976 700012 496032
rect 700068 495976 700136 496032
rect 700192 495982 707870 496032
rect 707926 495982 708000 496038
rect 700192 495976 708000 495982
rect 699322 495914 708000 495976
rect 699322 495908 707870 495914
rect 699322 495852 699392 495908
rect 699448 495852 699516 495908
rect 699572 495852 699640 495908
rect 699696 495852 699764 495908
rect 699820 495852 699888 495908
rect 699944 495852 700012 495908
rect 700068 495852 700136 495908
rect 700192 495858 707870 495908
rect 707926 495858 708000 495914
rect 700192 495852 708000 495858
rect 699322 495790 708000 495852
rect 699322 495784 707870 495790
rect 699322 495728 699392 495784
rect 699448 495728 699516 495784
rect 699572 495728 699640 495784
rect 699696 495728 699764 495784
rect 699820 495728 699888 495784
rect 699944 495728 700012 495784
rect 700068 495728 700136 495784
rect 700192 495734 707870 495784
rect 707926 495734 708000 495790
rect 700192 495728 708000 495734
rect 699322 495666 708000 495728
rect 699322 495660 707870 495666
rect 699322 495604 699392 495660
rect 699448 495604 699516 495660
rect 699572 495604 699640 495660
rect 699696 495604 699764 495660
rect 699820 495604 699888 495660
rect 699944 495604 700012 495660
rect 700068 495604 700136 495660
rect 700192 495610 707870 495660
rect 707926 495610 708000 495666
rect 700192 495604 708000 495610
rect 699322 495542 708000 495604
rect 699322 495536 707870 495542
rect 699322 495480 699392 495536
rect 699448 495480 699516 495536
rect 699572 495480 699640 495536
rect 699696 495480 699764 495536
rect 699820 495480 699888 495536
rect 699944 495480 700012 495536
rect 700068 495480 700136 495536
rect 700192 495486 707870 495536
rect 707926 495486 708000 495542
rect 700192 495480 708000 495486
rect 699322 495418 708000 495480
rect 699322 495412 707870 495418
rect 699322 495356 699392 495412
rect 699448 495356 699516 495412
rect 699572 495356 699640 495412
rect 699696 495356 699764 495412
rect 699820 495356 699888 495412
rect 699944 495356 700012 495412
rect 700068 495356 700136 495412
rect 700192 495362 707870 495412
rect 707926 495362 708000 495418
rect 700192 495356 708000 495362
rect 699322 495294 708000 495356
rect 699322 495288 707870 495294
rect 699322 495232 699392 495288
rect 699448 495232 699516 495288
rect 699572 495232 699640 495288
rect 699696 495232 699764 495288
rect 699820 495232 699888 495288
rect 699944 495232 700012 495288
rect 700068 495232 700136 495288
rect 700192 495238 707870 495288
rect 707926 495238 708000 495294
rect 700192 495232 708000 495238
rect 699322 495170 708000 495232
rect 699322 495164 707870 495170
rect 699322 495108 699392 495164
rect 699448 495108 699516 495164
rect 699572 495108 699640 495164
rect 699696 495108 699764 495164
rect 699820 495108 699888 495164
rect 699944 495108 700012 495164
rect 700068 495108 700136 495164
rect 700192 495114 707870 495164
rect 707926 495114 708000 495170
rect 700192 495108 708000 495114
rect 699322 495046 708000 495108
rect 699322 495040 707870 495046
rect 699322 494984 699392 495040
rect 699448 494984 699516 495040
rect 699572 494984 699640 495040
rect 699696 494984 699764 495040
rect 699820 494984 699888 495040
rect 699944 494984 700012 495040
rect 700068 494984 700136 495040
rect 700192 494990 707870 495040
rect 707926 494990 708000 495046
rect 700192 494984 708000 494990
rect 699322 494922 708000 494984
rect 699322 494916 707870 494922
rect 699322 494860 699392 494916
rect 699448 494860 699516 494916
rect 699572 494860 699640 494916
rect 699696 494860 699764 494916
rect 699820 494860 699888 494916
rect 699944 494860 700012 494916
rect 700068 494860 700136 494916
rect 700192 494866 707870 494916
rect 707926 494866 708000 494922
rect 700192 494860 708000 494866
rect 699322 494828 708000 494860
rect 699322 494178 708000 494248
rect 699322 494172 707870 494178
rect 699322 494116 699392 494172
rect 699448 494116 699516 494172
rect 699572 494116 699640 494172
rect 699696 494116 699764 494172
rect 699820 494116 699888 494172
rect 699944 494116 700012 494172
rect 700068 494116 700136 494172
rect 700192 494122 707870 494172
rect 707926 494122 708000 494178
rect 700192 494116 708000 494122
rect 699322 494054 708000 494116
rect 699322 494048 707870 494054
rect 699322 493992 699392 494048
rect 699448 493992 699516 494048
rect 699572 493992 699640 494048
rect 699696 493992 699764 494048
rect 699820 493992 699888 494048
rect 699944 493992 700012 494048
rect 700068 493992 700136 494048
rect 700192 493998 707870 494048
rect 707926 493998 708000 494054
rect 700192 493992 708000 493998
rect 699322 493930 708000 493992
rect 699322 493924 707870 493930
rect 699322 493868 699392 493924
rect 699448 493868 699516 493924
rect 699572 493868 699640 493924
rect 699696 493868 699764 493924
rect 699820 493868 699888 493924
rect 699944 493868 700012 493924
rect 700068 493868 700136 493924
rect 700192 493874 707870 493924
rect 707926 493874 708000 493930
rect 700192 493868 708000 493874
rect 699322 493806 708000 493868
rect 699322 493800 707870 493806
rect 699322 493744 699392 493800
rect 699448 493744 699516 493800
rect 699572 493744 699640 493800
rect 699696 493744 699764 493800
rect 699820 493744 699888 493800
rect 699944 493744 700012 493800
rect 700068 493744 700136 493800
rect 700192 493750 707870 493800
rect 707926 493750 708000 493806
rect 700192 493744 708000 493750
rect 699322 493682 708000 493744
rect 699322 493676 707870 493682
rect 699322 493620 699392 493676
rect 699448 493620 699516 493676
rect 699572 493620 699640 493676
rect 699696 493620 699764 493676
rect 699820 493620 699888 493676
rect 699944 493620 700012 493676
rect 700068 493620 700136 493676
rect 700192 493626 707870 493676
rect 707926 493626 708000 493682
rect 700192 493620 708000 493626
rect 699322 493558 708000 493620
rect 699322 493552 707870 493558
rect 699322 493496 699392 493552
rect 699448 493496 699516 493552
rect 699572 493496 699640 493552
rect 699696 493496 699764 493552
rect 699820 493496 699888 493552
rect 699944 493496 700012 493552
rect 700068 493496 700136 493552
rect 700192 493502 707870 493552
rect 707926 493502 708000 493558
rect 700192 493496 708000 493502
rect 699322 493434 708000 493496
rect 699322 493428 707870 493434
rect 699322 493372 699392 493428
rect 699448 493372 699516 493428
rect 699572 493372 699640 493428
rect 699696 493372 699764 493428
rect 699820 493372 699888 493428
rect 699944 493372 700012 493428
rect 700068 493372 700136 493428
rect 700192 493378 707870 493428
rect 707926 493378 708000 493434
rect 700192 493372 708000 493378
rect 699322 493310 708000 493372
rect 699322 493304 707870 493310
rect 699322 493248 699392 493304
rect 699448 493248 699516 493304
rect 699572 493248 699640 493304
rect 699696 493248 699764 493304
rect 699820 493248 699888 493304
rect 699944 493248 700012 493304
rect 700068 493248 700136 493304
rect 700192 493254 707870 493304
rect 707926 493254 708000 493310
rect 700192 493248 708000 493254
rect 699322 493186 708000 493248
rect 699322 493180 707870 493186
rect 699322 493124 699392 493180
rect 699448 493124 699516 493180
rect 699572 493124 699640 493180
rect 699696 493124 699764 493180
rect 699820 493124 699888 493180
rect 699944 493124 700012 493180
rect 700068 493124 700136 493180
rect 700192 493130 707870 493180
rect 707926 493130 708000 493186
rect 700192 493124 708000 493130
rect 699322 493062 708000 493124
rect 699322 493056 707870 493062
rect 699322 493000 699392 493056
rect 699448 493000 699516 493056
rect 699572 493000 699640 493056
rect 699696 493000 699764 493056
rect 699820 493000 699888 493056
rect 699944 493000 700012 493056
rect 700068 493000 700136 493056
rect 700192 493006 707870 493056
rect 707926 493006 708000 493062
rect 700192 493000 708000 493006
rect 699322 492938 708000 493000
rect 699322 492932 707870 492938
rect 699322 492876 699392 492932
rect 699448 492876 699516 492932
rect 699572 492876 699640 492932
rect 699696 492876 699764 492932
rect 699820 492876 699888 492932
rect 699944 492876 700012 492932
rect 700068 492876 700136 492932
rect 700192 492882 707870 492932
rect 707926 492882 708000 492938
rect 700192 492876 708000 492882
rect 699322 492814 708000 492876
rect 699322 492808 707870 492814
rect 699322 492752 699392 492808
rect 699448 492752 699516 492808
rect 699572 492752 699640 492808
rect 699696 492752 699764 492808
rect 699820 492752 699888 492808
rect 699944 492752 700012 492808
rect 700068 492752 700136 492808
rect 700192 492758 707870 492808
rect 707926 492758 708000 492814
rect 700192 492752 708000 492758
rect 699322 492690 708000 492752
rect 699322 492684 707870 492690
rect 699322 492628 699392 492684
rect 699448 492628 699516 492684
rect 699572 492628 699640 492684
rect 699696 492628 699764 492684
rect 699820 492628 699888 492684
rect 699944 492628 700012 492684
rect 700068 492628 700136 492684
rect 700192 492634 707870 492684
rect 707926 492634 708000 492690
rect 700192 492628 708000 492634
rect 699322 492566 708000 492628
rect 699322 492560 707870 492566
rect 699322 492504 699392 492560
rect 699448 492504 699516 492560
rect 699572 492504 699640 492560
rect 699696 492504 699764 492560
rect 699820 492504 699888 492560
rect 699944 492504 700012 492560
rect 700068 492504 700136 492560
rect 700192 492510 707870 492560
rect 707926 492510 708000 492566
rect 700192 492504 708000 492510
rect 699322 492442 708000 492504
rect 699322 492436 707870 492442
rect 699322 492380 699392 492436
rect 699448 492380 699516 492436
rect 699572 492380 699640 492436
rect 699696 492380 699764 492436
rect 699820 492380 699888 492436
rect 699944 492380 700012 492436
rect 700068 492380 700136 492436
rect 700192 492386 707870 492436
rect 707926 492386 708000 492442
rect 700192 492380 708000 492386
rect 699322 492318 708000 492380
rect 699322 492312 707870 492318
rect 699322 492256 699392 492312
rect 699448 492256 699516 492312
rect 699572 492256 699640 492312
rect 699696 492256 699764 492312
rect 699820 492256 699888 492312
rect 699944 492256 700012 492312
rect 700068 492256 700136 492312
rect 700192 492262 707870 492312
rect 707926 492262 708000 492318
rect 700192 492256 708000 492262
rect 699322 492198 708000 492256
rect 699322 491808 708000 491878
rect 699322 491802 707870 491808
rect 699322 491746 699392 491802
rect 699448 491746 699516 491802
rect 699572 491746 699640 491802
rect 699696 491746 699764 491802
rect 699820 491746 699888 491802
rect 699944 491746 700012 491802
rect 700068 491746 700136 491802
rect 700192 491752 707870 491802
rect 707926 491752 708000 491808
rect 700192 491746 708000 491752
rect 699322 491684 708000 491746
rect 699322 491678 707870 491684
rect 699322 491622 699392 491678
rect 699448 491622 699516 491678
rect 699572 491622 699640 491678
rect 699696 491622 699764 491678
rect 699820 491622 699888 491678
rect 699944 491622 700012 491678
rect 700068 491622 700136 491678
rect 700192 491628 707870 491678
rect 707926 491628 708000 491684
rect 700192 491622 708000 491628
rect 699322 491560 708000 491622
rect 699322 491554 707870 491560
rect 699322 491498 699392 491554
rect 699448 491498 699516 491554
rect 699572 491498 699640 491554
rect 699696 491498 699764 491554
rect 699820 491498 699888 491554
rect 699944 491498 700012 491554
rect 700068 491498 700136 491554
rect 700192 491504 707870 491554
rect 707926 491504 708000 491560
rect 700192 491498 708000 491504
rect 699322 491436 708000 491498
rect 699322 491430 707870 491436
rect 699322 491374 699392 491430
rect 699448 491374 699516 491430
rect 699572 491374 699640 491430
rect 699696 491374 699764 491430
rect 699820 491374 699888 491430
rect 699944 491374 700012 491430
rect 700068 491374 700136 491430
rect 700192 491380 707870 491430
rect 707926 491380 708000 491436
rect 700192 491374 708000 491380
rect 699322 491312 708000 491374
rect 699322 491306 707870 491312
rect 699322 491250 699392 491306
rect 699448 491250 699516 491306
rect 699572 491250 699640 491306
rect 699696 491250 699764 491306
rect 699820 491250 699888 491306
rect 699944 491250 700012 491306
rect 700068 491250 700136 491306
rect 700192 491256 707870 491306
rect 707926 491256 708000 491312
rect 700192 491250 708000 491256
rect 699322 491188 708000 491250
rect 699322 491182 707870 491188
rect 699322 491126 699392 491182
rect 699448 491126 699516 491182
rect 699572 491126 699640 491182
rect 699696 491126 699764 491182
rect 699820 491126 699888 491182
rect 699944 491126 700012 491182
rect 700068 491126 700136 491182
rect 700192 491132 707870 491182
rect 707926 491132 708000 491188
rect 700192 491126 708000 491132
rect 699322 491064 708000 491126
rect 699322 491058 707870 491064
rect 699322 491002 699392 491058
rect 699448 491002 699516 491058
rect 699572 491002 699640 491058
rect 699696 491002 699764 491058
rect 699820 491002 699888 491058
rect 699944 491002 700012 491058
rect 700068 491002 700136 491058
rect 700192 491008 707870 491058
rect 707926 491008 708000 491064
rect 700192 491002 708000 491008
rect 699322 490940 708000 491002
rect 699322 490934 707870 490940
rect 699322 490878 699392 490934
rect 699448 490878 699516 490934
rect 699572 490878 699640 490934
rect 699696 490878 699764 490934
rect 699820 490878 699888 490934
rect 699944 490878 700012 490934
rect 700068 490878 700136 490934
rect 700192 490884 707870 490934
rect 707926 490884 708000 490940
rect 700192 490878 708000 490884
rect 699322 490816 708000 490878
rect 699322 490810 707870 490816
rect 699322 490754 699392 490810
rect 699448 490754 699516 490810
rect 699572 490754 699640 490810
rect 699696 490754 699764 490810
rect 699820 490754 699888 490810
rect 699944 490754 700012 490810
rect 700068 490754 700136 490810
rect 700192 490760 707870 490810
rect 707926 490760 708000 490816
rect 700192 490754 708000 490760
rect 699322 490692 708000 490754
rect 699322 490686 707870 490692
rect 699322 490630 699392 490686
rect 699448 490630 699516 490686
rect 699572 490630 699640 490686
rect 699696 490630 699764 490686
rect 699820 490630 699888 490686
rect 699944 490630 700012 490686
rect 700068 490630 700136 490686
rect 700192 490636 707870 490686
rect 707926 490636 708000 490692
rect 700192 490630 708000 490636
rect 699322 490568 708000 490630
rect 699322 490562 707870 490568
rect 699322 490506 699392 490562
rect 699448 490506 699516 490562
rect 699572 490506 699640 490562
rect 699696 490506 699764 490562
rect 699820 490506 699888 490562
rect 699944 490506 700012 490562
rect 700068 490506 700136 490562
rect 700192 490512 707870 490562
rect 707926 490512 708000 490568
rect 700192 490506 708000 490512
rect 699322 490444 708000 490506
rect 699322 490438 707870 490444
rect 699322 490382 699392 490438
rect 699448 490382 699516 490438
rect 699572 490382 699640 490438
rect 699696 490382 699764 490438
rect 699820 490382 699888 490438
rect 699944 490382 700012 490438
rect 700068 490382 700136 490438
rect 700192 490388 707870 490438
rect 707926 490388 708000 490444
rect 700192 490382 708000 490388
rect 699322 490320 708000 490382
rect 699322 490314 707870 490320
rect 699322 490258 699392 490314
rect 699448 490258 699516 490314
rect 699572 490258 699640 490314
rect 699696 490258 699764 490314
rect 699820 490258 699888 490314
rect 699944 490258 700012 490314
rect 700068 490258 700136 490314
rect 700192 490264 707870 490314
rect 707926 490264 708000 490320
rect 700192 490258 708000 490264
rect 699322 490196 708000 490258
rect 699322 490190 707870 490196
rect 699322 490134 699392 490190
rect 699448 490134 699516 490190
rect 699572 490134 699640 490190
rect 699696 490134 699764 490190
rect 699820 490134 699888 490190
rect 699944 490134 700012 490190
rect 700068 490134 700136 490190
rect 700192 490140 707870 490190
rect 707926 490140 708000 490196
rect 700192 490134 708000 490140
rect 699322 490072 708000 490134
rect 699322 490066 707870 490072
rect 699322 490010 699392 490066
rect 699448 490010 699516 490066
rect 699572 490010 699640 490066
rect 699696 490010 699764 490066
rect 699820 490010 699888 490066
rect 699944 490010 700012 490066
rect 700068 490010 700136 490066
rect 700192 490016 707870 490066
rect 707926 490016 708000 490072
rect 700192 490010 708000 490016
rect 699322 489948 708000 490010
rect 699322 489942 707870 489948
rect 699322 489886 699392 489942
rect 699448 489886 699516 489942
rect 699572 489886 699640 489942
rect 699696 489886 699764 489942
rect 699820 489886 699888 489942
rect 699944 489886 700012 489942
rect 700068 489886 700136 489942
rect 700192 489892 707870 489942
rect 707926 489892 708000 489948
rect 700192 489886 708000 489892
rect 699322 489828 708000 489886
rect 699322 489102 708000 489172
rect 699322 489096 707870 489102
rect 699322 489040 699392 489096
rect 699448 489040 699516 489096
rect 699572 489040 699640 489096
rect 699696 489040 699764 489096
rect 699820 489040 699888 489096
rect 699944 489040 700012 489096
rect 700068 489040 700136 489096
rect 700192 489046 707870 489096
rect 707926 489046 708000 489102
rect 700192 489040 708000 489046
rect 699322 488978 708000 489040
rect 699322 488972 707870 488978
rect 699322 488916 699392 488972
rect 699448 488916 699516 488972
rect 699572 488916 699640 488972
rect 699696 488916 699764 488972
rect 699820 488916 699888 488972
rect 699944 488916 700012 488972
rect 700068 488916 700136 488972
rect 700192 488922 707870 488972
rect 707926 488922 708000 488978
rect 700192 488916 708000 488922
rect 699322 488854 708000 488916
rect 699322 488848 707870 488854
rect 699322 488792 699392 488848
rect 699448 488792 699516 488848
rect 699572 488792 699640 488848
rect 699696 488792 699764 488848
rect 699820 488792 699888 488848
rect 699944 488792 700012 488848
rect 700068 488792 700136 488848
rect 700192 488798 707870 488848
rect 707926 488798 708000 488854
rect 700192 488792 708000 488798
rect 699322 488730 708000 488792
rect 699322 488724 707870 488730
rect 699322 488668 699392 488724
rect 699448 488668 699516 488724
rect 699572 488668 699640 488724
rect 699696 488668 699764 488724
rect 699820 488668 699888 488724
rect 699944 488668 700012 488724
rect 700068 488668 700136 488724
rect 700192 488674 707870 488724
rect 707926 488674 708000 488730
rect 700192 488668 708000 488674
rect 699322 488606 708000 488668
rect 699322 488600 707870 488606
rect 699322 488544 699392 488600
rect 699448 488544 699516 488600
rect 699572 488544 699640 488600
rect 699696 488544 699764 488600
rect 699820 488544 699888 488600
rect 699944 488544 700012 488600
rect 700068 488544 700136 488600
rect 700192 488550 707870 488600
rect 707926 488550 708000 488606
rect 700192 488544 708000 488550
rect 699322 488482 708000 488544
rect 699322 488476 707870 488482
rect 699322 488420 699392 488476
rect 699448 488420 699516 488476
rect 699572 488420 699640 488476
rect 699696 488420 699764 488476
rect 699820 488420 699888 488476
rect 699944 488420 700012 488476
rect 700068 488420 700136 488476
rect 700192 488426 707870 488476
rect 707926 488426 708000 488482
rect 700192 488420 708000 488426
rect 699322 488358 708000 488420
rect 699322 488352 707870 488358
rect 699322 488296 699392 488352
rect 699448 488296 699516 488352
rect 699572 488296 699640 488352
rect 699696 488296 699764 488352
rect 699820 488296 699888 488352
rect 699944 488296 700012 488352
rect 700068 488296 700136 488352
rect 700192 488302 707870 488352
rect 707926 488302 708000 488358
rect 700192 488296 708000 488302
rect 699322 488234 708000 488296
rect 699322 488228 707870 488234
rect 699322 488172 699392 488228
rect 699448 488172 699516 488228
rect 699572 488172 699640 488228
rect 699696 488172 699764 488228
rect 699820 488172 699888 488228
rect 699944 488172 700012 488228
rect 700068 488172 700136 488228
rect 700192 488178 707870 488228
rect 707926 488178 708000 488234
rect 700192 488172 708000 488178
rect 699322 488110 708000 488172
rect 699322 488104 707870 488110
rect 699322 488048 699392 488104
rect 699448 488048 699516 488104
rect 699572 488048 699640 488104
rect 699696 488048 699764 488104
rect 699820 488048 699888 488104
rect 699944 488048 700012 488104
rect 700068 488048 700136 488104
rect 700192 488054 707870 488104
rect 707926 488054 708000 488110
rect 700192 488048 708000 488054
rect 699322 487986 708000 488048
rect 699322 487980 707870 487986
rect 699322 487924 699392 487980
rect 699448 487924 699516 487980
rect 699572 487924 699640 487980
rect 699696 487924 699764 487980
rect 699820 487924 699888 487980
rect 699944 487924 700012 487980
rect 700068 487924 700136 487980
rect 700192 487930 707870 487980
rect 707926 487930 708000 487986
rect 700192 487924 708000 487930
rect 699322 487862 708000 487924
rect 699322 487856 707870 487862
rect 699322 487800 699392 487856
rect 699448 487800 699516 487856
rect 699572 487800 699640 487856
rect 699696 487800 699764 487856
rect 699820 487800 699888 487856
rect 699944 487800 700012 487856
rect 700068 487800 700136 487856
rect 700192 487806 707870 487856
rect 707926 487806 708000 487862
rect 700192 487800 708000 487806
rect 699322 487738 708000 487800
rect 699322 487732 707870 487738
rect 699322 487676 699392 487732
rect 699448 487676 699516 487732
rect 699572 487676 699640 487732
rect 699696 487676 699764 487732
rect 699820 487676 699888 487732
rect 699944 487676 700012 487732
rect 700068 487676 700136 487732
rect 700192 487682 707870 487732
rect 707926 487682 708000 487738
rect 700192 487676 708000 487682
rect 699322 487614 708000 487676
rect 699322 487608 707870 487614
rect 699322 487552 699392 487608
rect 699448 487552 699516 487608
rect 699572 487552 699640 487608
rect 699696 487552 699764 487608
rect 699820 487552 699888 487608
rect 699944 487552 700012 487608
rect 700068 487552 700136 487608
rect 700192 487558 707870 487608
rect 707926 487558 708000 487614
rect 700192 487552 708000 487558
rect 699322 487490 708000 487552
rect 699322 487484 707870 487490
rect 699322 487428 699392 487484
rect 699448 487428 699516 487484
rect 699572 487428 699640 487484
rect 699696 487428 699764 487484
rect 699820 487428 699888 487484
rect 699944 487428 700012 487484
rect 700068 487428 700136 487484
rect 700192 487434 707870 487484
rect 707926 487434 708000 487490
rect 700192 487428 708000 487434
rect 699322 487366 708000 487428
rect 699322 487360 707870 487366
rect 699322 487304 699392 487360
rect 699448 487304 699516 487360
rect 699572 487304 699640 487360
rect 699696 487304 699764 487360
rect 699820 487304 699888 487360
rect 699944 487304 700012 487360
rect 700068 487304 700136 487360
rect 700192 487310 707870 487360
rect 707926 487310 708000 487366
rect 700192 487304 708000 487310
rect 699322 487242 708000 487304
rect 699322 487236 707870 487242
rect 699322 487180 699392 487236
rect 699448 487180 699516 487236
rect 699572 487180 699640 487236
rect 699696 487180 699764 487236
rect 699820 487180 699888 487236
rect 699944 487180 700012 487236
rect 700068 487180 700136 487236
rect 700192 487186 707870 487236
rect 707926 487186 708000 487242
rect 700192 487180 708000 487186
rect 699322 487122 708000 487180
rect 699322 486732 708000 486802
rect 699322 486726 707870 486732
rect 699322 486670 699392 486726
rect 699448 486670 699516 486726
rect 699572 486670 699640 486726
rect 699696 486670 699764 486726
rect 699820 486670 699888 486726
rect 699944 486670 700012 486726
rect 700068 486670 700136 486726
rect 700192 486676 707870 486726
rect 707926 486676 708000 486732
rect 700192 486670 708000 486676
rect 699322 486608 708000 486670
rect 699322 486602 707870 486608
rect 699322 486546 699392 486602
rect 699448 486546 699516 486602
rect 699572 486546 699640 486602
rect 699696 486546 699764 486602
rect 699820 486546 699888 486602
rect 699944 486546 700012 486602
rect 700068 486546 700136 486602
rect 700192 486552 707870 486602
rect 707926 486552 708000 486608
rect 700192 486546 708000 486552
rect 699322 486484 708000 486546
rect 699322 486478 707870 486484
rect 699322 486422 699392 486478
rect 699448 486422 699516 486478
rect 699572 486422 699640 486478
rect 699696 486422 699764 486478
rect 699820 486422 699888 486478
rect 699944 486422 700012 486478
rect 700068 486422 700136 486478
rect 700192 486428 707870 486478
rect 707926 486428 708000 486484
rect 700192 486422 708000 486428
rect 699322 486360 708000 486422
rect 699322 486354 707870 486360
rect 699322 486298 699392 486354
rect 699448 486298 699516 486354
rect 699572 486298 699640 486354
rect 699696 486298 699764 486354
rect 699820 486298 699888 486354
rect 699944 486298 700012 486354
rect 700068 486298 700136 486354
rect 700192 486304 707870 486354
rect 707926 486304 708000 486360
rect 700192 486298 708000 486304
rect 699322 486236 708000 486298
rect 699322 486230 707870 486236
rect 699322 486174 699392 486230
rect 699448 486174 699516 486230
rect 699572 486174 699640 486230
rect 699696 486174 699764 486230
rect 699820 486174 699888 486230
rect 699944 486174 700012 486230
rect 700068 486174 700136 486230
rect 700192 486180 707870 486230
rect 707926 486180 708000 486236
rect 700192 486174 708000 486180
rect 699322 486112 708000 486174
rect 699322 486106 707870 486112
rect 699322 486050 699392 486106
rect 699448 486050 699516 486106
rect 699572 486050 699640 486106
rect 699696 486050 699764 486106
rect 699820 486050 699888 486106
rect 699944 486050 700012 486106
rect 700068 486050 700136 486106
rect 700192 486056 707870 486106
rect 707926 486056 708000 486112
rect 700192 486050 708000 486056
rect 699322 485988 708000 486050
rect 699322 485982 707870 485988
rect 699322 485926 699392 485982
rect 699448 485926 699516 485982
rect 699572 485926 699640 485982
rect 699696 485926 699764 485982
rect 699820 485926 699888 485982
rect 699944 485926 700012 485982
rect 700068 485926 700136 485982
rect 700192 485932 707870 485982
rect 707926 485932 708000 485988
rect 700192 485926 708000 485932
rect 699322 485864 708000 485926
rect 699322 485858 707870 485864
rect 699322 485802 699392 485858
rect 699448 485802 699516 485858
rect 699572 485802 699640 485858
rect 699696 485802 699764 485858
rect 699820 485802 699888 485858
rect 699944 485802 700012 485858
rect 700068 485802 700136 485858
rect 700192 485808 707870 485858
rect 707926 485808 708000 485864
rect 700192 485802 708000 485808
rect 699322 485740 708000 485802
rect 699322 485734 707870 485740
rect 699322 485678 699392 485734
rect 699448 485678 699516 485734
rect 699572 485678 699640 485734
rect 699696 485678 699764 485734
rect 699820 485678 699888 485734
rect 699944 485678 700012 485734
rect 700068 485678 700136 485734
rect 700192 485684 707870 485734
rect 707926 485684 708000 485740
rect 700192 485678 708000 485684
rect 699322 485616 708000 485678
rect 699322 485610 707870 485616
rect 699322 485554 699392 485610
rect 699448 485554 699516 485610
rect 699572 485554 699640 485610
rect 699696 485554 699764 485610
rect 699820 485554 699888 485610
rect 699944 485554 700012 485610
rect 700068 485554 700136 485610
rect 700192 485560 707870 485610
rect 707926 485560 708000 485616
rect 700192 485554 708000 485560
rect 699322 485492 708000 485554
rect 699322 485486 707870 485492
rect 699322 485430 699392 485486
rect 699448 485430 699516 485486
rect 699572 485430 699640 485486
rect 699696 485430 699764 485486
rect 699820 485430 699888 485486
rect 699944 485430 700012 485486
rect 700068 485430 700136 485486
rect 700192 485436 707870 485486
rect 707926 485436 708000 485492
rect 700192 485430 708000 485436
rect 699322 485368 708000 485430
rect 699322 485362 707870 485368
rect 699322 485306 699392 485362
rect 699448 485306 699516 485362
rect 699572 485306 699640 485362
rect 699696 485306 699764 485362
rect 699820 485306 699888 485362
rect 699944 485306 700012 485362
rect 700068 485306 700136 485362
rect 700192 485312 707870 485362
rect 707926 485312 708000 485368
rect 700192 485306 708000 485312
rect 699322 485244 708000 485306
rect 699322 485238 707870 485244
rect 699322 485182 699392 485238
rect 699448 485182 699516 485238
rect 699572 485182 699640 485238
rect 699696 485182 699764 485238
rect 699820 485182 699888 485238
rect 699944 485182 700012 485238
rect 700068 485182 700136 485238
rect 700192 485188 707870 485238
rect 707926 485188 708000 485244
rect 700192 485182 708000 485188
rect 699322 485120 708000 485182
rect 699322 485114 707870 485120
rect 699322 485058 699392 485114
rect 699448 485058 699516 485114
rect 699572 485058 699640 485114
rect 699696 485058 699764 485114
rect 699820 485058 699888 485114
rect 699944 485058 700012 485114
rect 700068 485058 700136 485114
rect 700192 485064 707870 485114
rect 707926 485064 708000 485120
rect 700192 485058 708000 485064
rect 699322 484996 708000 485058
rect 699322 484990 707870 484996
rect 699322 484934 699392 484990
rect 699448 484934 699516 484990
rect 699572 484934 699640 484990
rect 699696 484934 699764 484990
rect 699820 484934 699888 484990
rect 699944 484934 700012 484990
rect 700068 484934 700136 484990
rect 700192 484940 707870 484990
rect 707926 484940 708000 484996
rect 700192 484934 708000 484940
rect 699322 484872 708000 484934
rect 699322 484866 707870 484872
rect 699322 484810 699392 484866
rect 699448 484810 699516 484866
rect 699572 484810 699640 484866
rect 699696 484810 699764 484866
rect 699820 484810 699888 484866
rect 699944 484810 700012 484866
rect 700068 484810 700136 484866
rect 700192 484816 707870 484866
rect 707926 484816 708000 484872
rect 700192 484810 708000 484816
rect 699322 484752 708000 484810
rect 699322 484134 708000 484172
rect 699322 484122 707870 484134
rect 699322 484066 699392 484122
rect 699448 484066 699516 484122
rect 699572 484066 699640 484122
rect 699696 484066 699764 484122
rect 699820 484066 699888 484122
rect 699944 484066 700012 484122
rect 700068 484066 700136 484122
rect 700192 484078 707870 484122
rect 707926 484078 708000 484134
rect 700192 484066 708000 484078
rect 699322 484010 708000 484066
rect 699322 483998 707870 484010
rect 699322 483942 699392 483998
rect 699448 483942 699516 483998
rect 699572 483942 699640 483998
rect 699696 483942 699764 483998
rect 699820 483942 699888 483998
rect 699944 483942 700012 483998
rect 700068 483942 700136 483998
rect 700192 483954 707870 483998
rect 707926 483954 708000 484010
rect 700192 483942 708000 483954
rect 699322 483886 708000 483942
rect 699322 483874 707870 483886
rect 699322 483818 699392 483874
rect 699448 483818 699516 483874
rect 699572 483818 699640 483874
rect 699696 483818 699764 483874
rect 699820 483818 699888 483874
rect 699944 483818 700012 483874
rect 700068 483818 700136 483874
rect 700192 483830 707870 483874
rect 707926 483830 708000 483886
rect 700192 483818 708000 483830
rect 699322 483762 708000 483818
rect 699322 483750 707870 483762
rect 699322 483694 699392 483750
rect 699448 483694 699516 483750
rect 699572 483694 699640 483750
rect 699696 483694 699764 483750
rect 699820 483694 699888 483750
rect 699944 483694 700012 483750
rect 700068 483694 700136 483750
rect 700192 483706 707870 483750
rect 707926 483706 708000 483762
rect 700192 483694 708000 483706
rect 699322 483638 708000 483694
rect 699322 483626 707870 483638
rect 699322 483570 699392 483626
rect 699448 483570 699516 483626
rect 699572 483570 699640 483626
rect 699696 483570 699764 483626
rect 699820 483570 699888 483626
rect 699944 483570 700012 483626
rect 700068 483570 700136 483626
rect 700192 483582 707870 483626
rect 707926 483582 708000 483638
rect 700192 483570 708000 483582
rect 699322 483514 708000 483570
rect 699322 483502 707870 483514
rect 699322 483446 699392 483502
rect 699448 483446 699516 483502
rect 699572 483446 699640 483502
rect 699696 483446 699764 483502
rect 699820 483446 699888 483502
rect 699944 483446 700012 483502
rect 700068 483446 700136 483502
rect 700192 483458 707870 483502
rect 707926 483458 708000 483514
rect 700192 483446 708000 483458
rect 699322 483390 708000 483446
rect 699322 483378 707870 483390
rect 699322 483322 699392 483378
rect 699448 483322 699516 483378
rect 699572 483322 699640 483378
rect 699696 483322 699764 483378
rect 699820 483322 699888 483378
rect 699944 483322 700012 483378
rect 700068 483322 700136 483378
rect 700192 483334 707870 483378
rect 707926 483334 708000 483390
rect 700192 483322 708000 483334
rect 699322 483266 708000 483322
rect 699322 483254 707870 483266
rect 699322 483198 699392 483254
rect 699448 483198 699516 483254
rect 699572 483198 699640 483254
rect 699696 483198 699764 483254
rect 699820 483198 699888 483254
rect 699944 483198 700012 483254
rect 700068 483198 700136 483254
rect 700192 483210 707870 483254
rect 707926 483210 708000 483266
rect 700192 483198 708000 483210
rect 699322 483142 708000 483198
rect 699322 483130 707870 483142
rect 699322 483074 699392 483130
rect 699448 483074 699516 483130
rect 699572 483074 699640 483130
rect 699696 483074 699764 483130
rect 699820 483074 699888 483130
rect 699944 483074 700012 483130
rect 700068 483074 700136 483130
rect 700192 483086 707870 483130
rect 707926 483086 708000 483142
rect 700192 483074 708000 483086
rect 699322 483018 708000 483074
rect 699322 483006 707870 483018
rect 699322 482950 699392 483006
rect 699448 482950 699516 483006
rect 699572 482950 699640 483006
rect 699696 482950 699764 483006
rect 699820 482950 699888 483006
rect 699944 482950 700012 483006
rect 700068 482950 700136 483006
rect 700192 482962 707870 483006
rect 707926 482962 708000 483018
rect 700192 482950 708000 482962
rect 699322 482894 708000 482950
rect 699322 482882 707870 482894
rect 699322 482826 699392 482882
rect 699448 482826 699516 482882
rect 699572 482826 699640 482882
rect 699696 482826 699764 482882
rect 699820 482826 699888 482882
rect 699944 482826 700012 482882
rect 700068 482826 700136 482882
rect 700192 482838 707870 482882
rect 707926 482838 708000 482894
rect 700192 482826 708000 482838
rect 699322 482770 708000 482826
rect 699322 482758 707870 482770
rect 699322 482702 699392 482758
rect 699448 482702 699516 482758
rect 699572 482702 699640 482758
rect 699696 482702 699764 482758
rect 699820 482702 699888 482758
rect 699944 482702 700012 482758
rect 700068 482702 700136 482758
rect 700192 482714 707870 482758
rect 707926 482714 708000 482770
rect 700192 482702 708000 482714
rect 699322 482646 708000 482702
rect 699322 482634 707870 482646
rect 699322 482630 699392 482634
rect 77678 482429 84516 482630
rect 77678 482373 77800 482429
rect 77856 482373 78100 482429
rect 78156 482373 78400 482429
rect 78456 482373 84516 482429
rect 77678 482229 84516 482373
rect 77678 482173 77800 482229
rect 77856 482173 78100 482229
rect 78156 482173 78400 482229
rect 78456 482173 84516 482229
rect 77678 482010 84516 482173
rect 687412 482578 699392 482630
rect 699448 482578 699516 482634
rect 699572 482578 699640 482634
rect 699696 482578 699764 482634
rect 699820 482578 699888 482634
rect 699944 482578 700012 482634
rect 700068 482578 700136 482634
rect 700192 482590 707870 482634
rect 707926 482590 708000 482646
rect 700192 482578 708000 482590
rect 687412 482522 708000 482578
rect 687412 482510 707870 482522
rect 687412 482454 699392 482510
rect 699448 482454 699516 482510
rect 699572 482454 699640 482510
rect 699696 482454 699764 482510
rect 699820 482454 699888 482510
rect 699944 482454 700012 482510
rect 700068 482454 700136 482510
rect 700192 482466 707870 482510
rect 707926 482466 708000 482522
rect 700192 482454 708000 482466
rect 687412 482398 708000 482454
rect 687412 482386 707870 482398
rect 687412 482330 699392 482386
rect 699448 482330 699516 482386
rect 699572 482330 699640 482386
rect 699696 482330 699764 482386
rect 699820 482330 699888 482386
rect 699944 482330 700012 482386
rect 700068 482330 700136 482386
rect 700192 482342 707870 482386
rect 707926 482342 708000 482398
rect 700192 482330 708000 482342
rect 687412 482272 708000 482330
rect 687412 482010 700322 482272
rect 70000 474670 78678 474728
rect 70000 474658 77808 474670
rect 70000 474602 70074 474658
rect 70130 474614 77808 474658
rect 77864 474614 77932 474670
rect 77988 474614 78056 474670
rect 78112 474614 78180 474670
rect 78236 474614 78304 474670
rect 78360 474614 78428 474670
rect 78484 474614 78552 474670
rect 78608 474614 78678 474670
rect 70130 474602 78678 474614
rect 70000 474546 78678 474602
rect 70000 474534 77808 474546
rect 70000 474478 70074 474534
rect 70130 474490 77808 474534
rect 77864 474490 77932 474546
rect 77988 474490 78056 474546
rect 78112 474490 78180 474546
rect 78236 474490 78304 474546
rect 78360 474490 78428 474546
rect 78484 474490 78552 474546
rect 78608 474490 78678 474546
rect 70130 474478 78678 474490
rect 70000 474422 78678 474478
rect 70000 474410 77808 474422
rect 70000 474354 70074 474410
rect 70130 474366 77808 474410
rect 77864 474366 77932 474422
rect 77988 474366 78056 474422
rect 78112 474366 78180 474422
rect 78236 474366 78304 474422
rect 78360 474366 78428 474422
rect 78484 474366 78552 474422
rect 78608 474366 78678 474422
rect 70130 474354 78678 474366
rect 70000 474298 78678 474354
rect 70000 474286 77808 474298
rect 70000 474230 70074 474286
rect 70130 474242 77808 474286
rect 77864 474242 77932 474298
rect 77988 474242 78056 474298
rect 78112 474242 78180 474298
rect 78236 474242 78304 474298
rect 78360 474242 78428 474298
rect 78484 474242 78552 474298
rect 78608 474242 78678 474298
rect 70130 474230 78678 474242
rect 70000 474174 78678 474230
rect 70000 474162 77808 474174
rect 70000 474106 70074 474162
rect 70130 474118 77808 474162
rect 77864 474118 77932 474174
rect 77988 474118 78056 474174
rect 78112 474118 78180 474174
rect 78236 474118 78304 474174
rect 78360 474118 78428 474174
rect 78484 474118 78552 474174
rect 78608 474118 78678 474174
rect 70130 474106 78678 474118
rect 70000 474050 78678 474106
rect 70000 474038 77808 474050
rect 70000 473982 70074 474038
rect 70130 473994 77808 474038
rect 77864 473994 77932 474050
rect 77988 473994 78056 474050
rect 78112 473994 78180 474050
rect 78236 473994 78304 474050
rect 78360 473994 78428 474050
rect 78484 473994 78552 474050
rect 78608 473994 78678 474050
rect 70130 473982 78678 473994
rect 70000 473926 78678 473982
rect 70000 473914 77808 473926
rect 70000 473858 70074 473914
rect 70130 473870 77808 473914
rect 77864 473870 77932 473926
rect 77988 473870 78056 473926
rect 78112 473870 78180 473926
rect 78236 473870 78304 473926
rect 78360 473870 78428 473926
rect 78484 473870 78552 473926
rect 78608 473870 78678 473926
rect 70130 473858 78678 473870
rect 70000 473802 78678 473858
rect 70000 473790 77808 473802
rect 70000 473734 70074 473790
rect 70130 473746 77808 473790
rect 77864 473746 77932 473802
rect 77988 473746 78056 473802
rect 78112 473746 78180 473802
rect 78236 473746 78304 473802
rect 78360 473746 78428 473802
rect 78484 473746 78552 473802
rect 78608 473746 78678 473802
rect 70130 473734 78678 473746
rect 70000 473678 78678 473734
rect 70000 473666 77808 473678
rect 70000 473610 70074 473666
rect 70130 473622 77808 473666
rect 77864 473622 77932 473678
rect 77988 473622 78056 473678
rect 78112 473622 78180 473678
rect 78236 473622 78304 473678
rect 78360 473622 78428 473678
rect 78484 473622 78552 473678
rect 78608 473622 78678 473678
rect 70130 473610 78678 473622
rect 70000 473554 78678 473610
rect 70000 473542 77808 473554
rect 70000 473486 70074 473542
rect 70130 473498 77808 473542
rect 77864 473498 77932 473554
rect 77988 473498 78056 473554
rect 78112 473498 78180 473554
rect 78236 473498 78304 473554
rect 78360 473498 78428 473554
rect 78484 473498 78552 473554
rect 78608 473498 78678 473554
rect 70130 473486 78678 473498
rect 70000 473430 78678 473486
rect 70000 473418 77808 473430
rect 70000 473362 70074 473418
rect 70130 473374 77808 473418
rect 77864 473374 77932 473430
rect 77988 473374 78056 473430
rect 78112 473374 78180 473430
rect 78236 473374 78304 473430
rect 78360 473374 78428 473430
rect 78484 473374 78552 473430
rect 78608 473374 78678 473430
rect 70130 473362 78678 473374
rect 70000 473306 78678 473362
rect 70000 473294 77808 473306
rect 70000 473238 70074 473294
rect 70130 473250 77808 473294
rect 77864 473250 77932 473306
rect 77988 473250 78056 473306
rect 78112 473250 78180 473306
rect 78236 473250 78304 473306
rect 78360 473250 78428 473306
rect 78484 473250 78552 473306
rect 78608 473250 78678 473306
rect 70130 473238 78678 473250
rect 70000 473182 78678 473238
rect 70000 473170 77808 473182
rect 70000 473114 70074 473170
rect 70130 473126 77808 473170
rect 77864 473126 77932 473182
rect 77988 473126 78056 473182
rect 78112 473126 78180 473182
rect 78236 473126 78304 473182
rect 78360 473126 78428 473182
rect 78484 473126 78552 473182
rect 78608 473126 78678 473182
rect 70130 473114 78678 473126
rect 70000 473058 78678 473114
rect 70000 473046 77808 473058
rect 70000 472990 70074 473046
rect 70130 473002 77808 473046
rect 77864 473002 77932 473058
rect 77988 473002 78056 473058
rect 78112 473002 78180 473058
rect 78236 473002 78304 473058
rect 78360 473002 78428 473058
rect 78484 473002 78552 473058
rect 78608 473002 78678 473058
rect 70130 472990 78678 473002
rect 70000 472934 78678 472990
rect 70000 472922 77808 472934
rect 70000 472866 70074 472922
rect 70130 472878 77808 472922
rect 77864 472878 77932 472934
rect 77988 472878 78056 472934
rect 78112 472878 78180 472934
rect 78236 472878 78304 472934
rect 78360 472878 78428 472934
rect 78484 472878 78552 472934
rect 78608 472878 78678 472934
rect 70130 472866 78678 472878
rect 70000 472828 78678 472866
rect 70000 472190 78678 472248
rect 70000 472184 77808 472190
rect 70000 472128 70074 472184
rect 70130 472134 77808 472184
rect 77864 472134 77932 472190
rect 77988 472134 78056 472190
rect 78112 472134 78180 472190
rect 78236 472134 78304 472190
rect 78360 472134 78428 472190
rect 78484 472134 78552 472190
rect 78608 472134 78678 472190
rect 70130 472128 78678 472134
rect 70000 472066 78678 472128
rect 70000 472060 77808 472066
rect 70000 472004 70074 472060
rect 70130 472010 77808 472060
rect 77864 472010 77932 472066
rect 77988 472010 78056 472066
rect 78112 472010 78180 472066
rect 78236 472010 78304 472066
rect 78360 472010 78428 472066
rect 78484 472010 78552 472066
rect 78608 472010 78678 472066
rect 70130 472004 78678 472010
rect 70000 471942 78678 472004
rect 70000 471936 77808 471942
rect 70000 471880 70074 471936
rect 70130 471886 77808 471936
rect 77864 471886 77932 471942
rect 77988 471886 78056 471942
rect 78112 471886 78180 471942
rect 78236 471886 78304 471942
rect 78360 471886 78428 471942
rect 78484 471886 78552 471942
rect 78608 471886 78678 471942
rect 70130 471880 78678 471886
rect 70000 471818 78678 471880
rect 70000 471812 77808 471818
rect 70000 471756 70074 471812
rect 70130 471762 77808 471812
rect 77864 471762 77932 471818
rect 77988 471762 78056 471818
rect 78112 471762 78180 471818
rect 78236 471762 78304 471818
rect 78360 471762 78428 471818
rect 78484 471762 78552 471818
rect 78608 471762 78678 471818
rect 70130 471756 78678 471762
rect 70000 471694 78678 471756
rect 70000 471688 77808 471694
rect 70000 471632 70074 471688
rect 70130 471638 77808 471688
rect 77864 471638 77932 471694
rect 77988 471638 78056 471694
rect 78112 471638 78180 471694
rect 78236 471638 78304 471694
rect 78360 471638 78428 471694
rect 78484 471638 78552 471694
rect 78608 471638 78678 471694
rect 70130 471632 78678 471638
rect 70000 471570 78678 471632
rect 70000 471564 77808 471570
rect 70000 471508 70074 471564
rect 70130 471514 77808 471564
rect 77864 471514 77932 471570
rect 77988 471514 78056 471570
rect 78112 471514 78180 471570
rect 78236 471514 78304 471570
rect 78360 471514 78428 471570
rect 78484 471514 78552 471570
rect 78608 471514 78678 471570
rect 70130 471508 78678 471514
rect 70000 471446 78678 471508
rect 70000 471440 77808 471446
rect 70000 471384 70074 471440
rect 70130 471390 77808 471440
rect 77864 471390 77932 471446
rect 77988 471390 78056 471446
rect 78112 471390 78180 471446
rect 78236 471390 78304 471446
rect 78360 471390 78428 471446
rect 78484 471390 78552 471446
rect 78608 471390 78678 471446
rect 70130 471384 78678 471390
rect 70000 471322 78678 471384
rect 70000 471316 77808 471322
rect 70000 471260 70074 471316
rect 70130 471266 77808 471316
rect 77864 471266 77932 471322
rect 77988 471266 78056 471322
rect 78112 471266 78180 471322
rect 78236 471266 78304 471322
rect 78360 471266 78428 471322
rect 78484 471266 78552 471322
rect 78608 471266 78678 471322
rect 70130 471260 78678 471266
rect 70000 471198 78678 471260
rect 70000 471192 77808 471198
rect 70000 471136 70074 471192
rect 70130 471142 77808 471192
rect 77864 471142 77932 471198
rect 77988 471142 78056 471198
rect 78112 471142 78180 471198
rect 78236 471142 78304 471198
rect 78360 471142 78428 471198
rect 78484 471142 78552 471198
rect 78608 471142 78678 471198
rect 70130 471136 78678 471142
rect 70000 471074 78678 471136
rect 70000 471068 77808 471074
rect 70000 471012 70074 471068
rect 70130 471018 77808 471068
rect 77864 471018 77932 471074
rect 77988 471018 78056 471074
rect 78112 471018 78180 471074
rect 78236 471018 78304 471074
rect 78360 471018 78428 471074
rect 78484 471018 78552 471074
rect 78608 471018 78678 471074
rect 70130 471012 78678 471018
rect 70000 470950 78678 471012
rect 70000 470944 77808 470950
rect 70000 470888 70074 470944
rect 70130 470894 77808 470944
rect 77864 470894 77932 470950
rect 77988 470894 78056 470950
rect 78112 470894 78180 470950
rect 78236 470894 78304 470950
rect 78360 470894 78428 470950
rect 78484 470894 78552 470950
rect 78608 470894 78678 470950
rect 70130 470888 78678 470894
rect 70000 470826 78678 470888
rect 70000 470820 77808 470826
rect 70000 470764 70074 470820
rect 70130 470770 77808 470820
rect 77864 470770 77932 470826
rect 77988 470770 78056 470826
rect 78112 470770 78180 470826
rect 78236 470770 78304 470826
rect 78360 470770 78428 470826
rect 78484 470770 78552 470826
rect 78608 470770 78678 470826
rect 70130 470764 78678 470770
rect 70000 470702 78678 470764
rect 70000 470696 77808 470702
rect 70000 470640 70074 470696
rect 70130 470646 77808 470696
rect 77864 470646 77932 470702
rect 77988 470646 78056 470702
rect 78112 470646 78180 470702
rect 78236 470646 78304 470702
rect 78360 470646 78428 470702
rect 78484 470646 78552 470702
rect 78608 470646 78678 470702
rect 70130 470640 78678 470646
rect 70000 470578 78678 470640
rect 70000 470572 77808 470578
rect 70000 470516 70074 470572
rect 70130 470522 77808 470572
rect 77864 470522 77932 470578
rect 77988 470522 78056 470578
rect 78112 470522 78180 470578
rect 78236 470522 78304 470578
rect 78360 470522 78428 470578
rect 78484 470522 78552 470578
rect 78608 470522 78678 470578
rect 70130 470516 78678 470522
rect 70000 470454 78678 470516
rect 70000 470448 77808 470454
rect 70000 470392 70074 470448
rect 70130 470398 77808 470448
rect 77864 470398 77932 470454
rect 77988 470398 78056 470454
rect 78112 470398 78180 470454
rect 78236 470398 78304 470454
rect 78360 470398 78428 470454
rect 78484 470398 78552 470454
rect 78608 470398 78678 470454
rect 70130 470392 78678 470398
rect 70000 470330 78678 470392
rect 70000 470324 77808 470330
rect 70000 470268 70074 470324
rect 70130 470274 77808 470324
rect 77864 470274 77932 470330
rect 77988 470274 78056 470330
rect 78112 470274 78180 470330
rect 78236 470274 78304 470330
rect 78360 470274 78428 470330
rect 78484 470274 78552 470330
rect 78608 470274 78678 470330
rect 70130 470268 78678 470274
rect 70000 470198 78678 470268
rect 70000 469820 78678 469878
rect 70000 469814 77808 469820
rect 70000 469758 70074 469814
rect 70130 469764 77808 469814
rect 77864 469764 77932 469820
rect 77988 469764 78056 469820
rect 78112 469764 78180 469820
rect 78236 469764 78304 469820
rect 78360 469764 78428 469820
rect 78484 469764 78552 469820
rect 78608 469764 78678 469820
rect 70130 469758 78678 469764
rect 70000 469696 78678 469758
rect 70000 469690 77808 469696
rect 70000 469634 70074 469690
rect 70130 469640 77808 469690
rect 77864 469640 77932 469696
rect 77988 469640 78056 469696
rect 78112 469640 78180 469696
rect 78236 469640 78304 469696
rect 78360 469640 78428 469696
rect 78484 469640 78552 469696
rect 78608 469640 78678 469696
rect 70130 469634 78678 469640
rect 70000 469572 78678 469634
rect 70000 469566 77808 469572
rect 70000 469510 70074 469566
rect 70130 469516 77808 469566
rect 77864 469516 77932 469572
rect 77988 469516 78056 469572
rect 78112 469516 78180 469572
rect 78236 469516 78304 469572
rect 78360 469516 78428 469572
rect 78484 469516 78552 469572
rect 78608 469516 78678 469572
rect 70130 469510 78678 469516
rect 70000 469448 78678 469510
rect 70000 469442 77808 469448
rect 70000 469386 70074 469442
rect 70130 469392 77808 469442
rect 77864 469392 77932 469448
rect 77988 469392 78056 469448
rect 78112 469392 78180 469448
rect 78236 469392 78304 469448
rect 78360 469392 78428 469448
rect 78484 469392 78552 469448
rect 78608 469392 78678 469448
rect 70130 469386 78678 469392
rect 70000 469324 78678 469386
rect 70000 469318 77808 469324
rect 70000 469262 70074 469318
rect 70130 469268 77808 469318
rect 77864 469268 77932 469324
rect 77988 469268 78056 469324
rect 78112 469268 78180 469324
rect 78236 469268 78304 469324
rect 78360 469268 78428 469324
rect 78484 469268 78552 469324
rect 78608 469268 78678 469324
rect 70130 469262 78678 469268
rect 70000 469200 78678 469262
rect 70000 469194 77808 469200
rect 70000 469138 70074 469194
rect 70130 469144 77808 469194
rect 77864 469144 77932 469200
rect 77988 469144 78056 469200
rect 78112 469144 78180 469200
rect 78236 469144 78304 469200
rect 78360 469144 78428 469200
rect 78484 469144 78552 469200
rect 78608 469144 78678 469200
rect 70130 469138 78678 469144
rect 70000 469076 78678 469138
rect 70000 469070 77808 469076
rect 70000 469014 70074 469070
rect 70130 469020 77808 469070
rect 77864 469020 77932 469076
rect 77988 469020 78056 469076
rect 78112 469020 78180 469076
rect 78236 469020 78304 469076
rect 78360 469020 78428 469076
rect 78484 469020 78552 469076
rect 78608 469020 78678 469076
rect 70130 469014 78678 469020
rect 70000 468952 78678 469014
rect 70000 468946 77808 468952
rect 70000 468890 70074 468946
rect 70130 468896 77808 468946
rect 77864 468896 77932 468952
rect 77988 468896 78056 468952
rect 78112 468896 78180 468952
rect 78236 468896 78304 468952
rect 78360 468896 78428 468952
rect 78484 468896 78552 468952
rect 78608 468896 78678 468952
rect 70130 468890 78678 468896
rect 70000 468828 78678 468890
rect 70000 468822 77808 468828
rect 70000 468766 70074 468822
rect 70130 468772 77808 468822
rect 77864 468772 77932 468828
rect 77988 468772 78056 468828
rect 78112 468772 78180 468828
rect 78236 468772 78304 468828
rect 78360 468772 78428 468828
rect 78484 468772 78552 468828
rect 78608 468772 78678 468828
rect 70130 468766 78678 468772
rect 70000 468704 78678 468766
rect 70000 468698 77808 468704
rect 70000 468642 70074 468698
rect 70130 468648 77808 468698
rect 77864 468648 77932 468704
rect 77988 468648 78056 468704
rect 78112 468648 78180 468704
rect 78236 468648 78304 468704
rect 78360 468648 78428 468704
rect 78484 468648 78552 468704
rect 78608 468648 78678 468704
rect 70130 468642 78678 468648
rect 70000 468580 78678 468642
rect 70000 468574 77808 468580
rect 70000 468518 70074 468574
rect 70130 468524 77808 468574
rect 77864 468524 77932 468580
rect 77988 468524 78056 468580
rect 78112 468524 78180 468580
rect 78236 468524 78304 468580
rect 78360 468524 78428 468580
rect 78484 468524 78552 468580
rect 78608 468524 78678 468580
rect 70130 468518 78678 468524
rect 70000 468456 78678 468518
rect 70000 468450 77808 468456
rect 70000 468394 70074 468450
rect 70130 468400 77808 468450
rect 77864 468400 77932 468456
rect 77988 468400 78056 468456
rect 78112 468400 78180 468456
rect 78236 468400 78304 468456
rect 78360 468400 78428 468456
rect 78484 468400 78552 468456
rect 78608 468400 78678 468456
rect 70130 468394 78678 468400
rect 70000 468332 78678 468394
rect 70000 468326 77808 468332
rect 70000 468270 70074 468326
rect 70130 468276 77808 468326
rect 77864 468276 77932 468332
rect 77988 468276 78056 468332
rect 78112 468276 78180 468332
rect 78236 468276 78304 468332
rect 78360 468276 78428 468332
rect 78484 468276 78552 468332
rect 78608 468276 78678 468332
rect 70130 468270 78678 468276
rect 70000 468208 78678 468270
rect 70000 468202 77808 468208
rect 70000 468146 70074 468202
rect 70130 468152 77808 468202
rect 77864 468152 77932 468208
rect 77988 468152 78056 468208
rect 78112 468152 78180 468208
rect 78236 468152 78304 468208
rect 78360 468152 78428 468208
rect 78484 468152 78552 468208
rect 78608 468152 78678 468208
rect 70130 468146 78678 468152
rect 70000 468084 78678 468146
rect 70000 468078 77808 468084
rect 70000 468022 70074 468078
rect 70130 468028 77808 468078
rect 77864 468028 77932 468084
rect 77988 468028 78056 468084
rect 78112 468028 78180 468084
rect 78236 468028 78304 468084
rect 78360 468028 78428 468084
rect 78484 468028 78552 468084
rect 78608 468028 78678 468084
rect 70130 468022 78678 468028
rect 70000 467960 78678 468022
rect 70000 467954 77808 467960
rect 70000 467898 70074 467954
rect 70130 467904 77808 467954
rect 77864 467904 77932 467960
rect 77988 467904 78056 467960
rect 78112 467904 78180 467960
rect 78236 467904 78304 467960
rect 78360 467904 78428 467960
rect 78484 467904 78552 467960
rect 78608 467904 78678 467960
rect 70130 467898 78678 467904
rect 70000 467828 78678 467898
rect 70000 467114 78678 467172
rect 70000 467108 77808 467114
rect 70000 467052 70074 467108
rect 70130 467058 77808 467108
rect 77864 467058 77932 467114
rect 77988 467058 78056 467114
rect 78112 467058 78180 467114
rect 78236 467058 78304 467114
rect 78360 467058 78428 467114
rect 78484 467058 78552 467114
rect 78608 467058 78678 467114
rect 70130 467052 78678 467058
rect 70000 466990 78678 467052
rect 70000 466984 77808 466990
rect 70000 466928 70074 466984
rect 70130 466934 77808 466984
rect 77864 466934 77932 466990
rect 77988 466934 78056 466990
rect 78112 466934 78180 466990
rect 78236 466934 78304 466990
rect 78360 466934 78428 466990
rect 78484 466934 78552 466990
rect 78608 466934 78678 466990
rect 70130 466928 78678 466934
rect 70000 466866 78678 466928
rect 70000 466860 77808 466866
rect 70000 466804 70074 466860
rect 70130 466810 77808 466860
rect 77864 466810 77932 466866
rect 77988 466810 78056 466866
rect 78112 466810 78180 466866
rect 78236 466810 78304 466866
rect 78360 466810 78428 466866
rect 78484 466810 78552 466866
rect 78608 466810 78678 466866
rect 70130 466804 78678 466810
rect 70000 466742 78678 466804
rect 70000 466736 77808 466742
rect 70000 466680 70074 466736
rect 70130 466686 77808 466736
rect 77864 466686 77932 466742
rect 77988 466686 78056 466742
rect 78112 466686 78180 466742
rect 78236 466686 78304 466742
rect 78360 466686 78428 466742
rect 78484 466686 78552 466742
rect 78608 466686 78678 466742
rect 70130 466680 78678 466686
rect 70000 466618 78678 466680
rect 70000 466612 77808 466618
rect 70000 466556 70074 466612
rect 70130 466562 77808 466612
rect 77864 466562 77932 466618
rect 77988 466562 78056 466618
rect 78112 466562 78180 466618
rect 78236 466562 78304 466618
rect 78360 466562 78428 466618
rect 78484 466562 78552 466618
rect 78608 466562 78678 466618
rect 70130 466556 78678 466562
rect 70000 466494 78678 466556
rect 70000 466488 77808 466494
rect 70000 466432 70074 466488
rect 70130 466438 77808 466488
rect 77864 466438 77932 466494
rect 77988 466438 78056 466494
rect 78112 466438 78180 466494
rect 78236 466438 78304 466494
rect 78360 466438 78428 466494
rect 78484 466438 78552 466494
rect 78608 466438 78678 466494
rect 70130 466432 78678 466438
rect 70000 466370 78678 466432
rect 70000 466364 77808 466370
rect 70000 466308 70074 466364
rect 70130 466314 77808 466364
rect 77864 466314 77932 466370
rect 77988 466314 78056 466370
rect 78112 466314 78180 466370
rect 78236 466314 78304 466370
rect 78360 466314 78428 466370
rect 78484 466314 78552 466370
rect 78608 466314 78678 466370
rect 70130 466308 78678 466314
rect 70000 466246 78678 466308
rect 70000 466240 77808 466246
rect 70000 466184 70074 466240
rect 70130 466190 77808 466240
rect 77864 466190 77932 466246
rect 77988 466190 78056 466246
rect 78112 466190 78180 466246
rect 78236 466190 78304 466246
rect 78360 466190 78428 466246
rect 78484 466190 78552 466246
rect 78608 466190 78678 466246
rect 70130 466184 78678 466190
rect 70000 466122 78678 466184
rect 70000 466116 77808 466122
rect 70000 466060 70074 466116
rect 70130 466066 77808 466116
rect 77864 466066 77932 466122
rect 77988 466066 78056 466122
rect 78112 466066 78180 466122
rect 78236 466066 78304 466122
rect 78360 466066 78428 466122
rect 78484 466066 78552 466122
rect 78608 466066 78678 466122
rect 70130 466060 78678 466066
rect 70000 465998 78678 466060
rect 70000 465992 77808 465998
rect 70000 465936 70074 465992
rect 70130 465942 77808 465992
rect 77864 465942 77932 465998
rect 77988 465942 78056 465998
rect 78112 465942 78180 465998
rect 78236 465942 78304 465998
rect 78360 465942 78428 465998
rect 78484 465942 78552 465998
rect 78608 465942 78678 465998
rect 70130 465936 78678 465942
rect 70000 465874 78678 465936
rect 70000 465868 77808 465874
rect 70000 465812 70074 465868
rect 70130 465818 77808 465868
rect 77864 465818 77932 465874
rect 77988 465818 78056 465874
rect 78112 465818 78180 465874
rect 78236 465818 78304 465874
rect 78360 465818 78428 465874
rect 78484 465818 78552 465874
rect 78608 465818 78678 465874
rect 70130 465812 78678 465818
rect 70000 465750 78678 465812
rect 70000 465744 77808 465750
rect 70000 465688 70074 465744
rect 70130 465694 77808 465744
rect 77864 465694 77932 465750
rect 77988 465694 78056 465750
rect 78112 465694 78180 465750
rect 78236 465694 78304 465750
rect 78360 465694 78428 465750
rect 78484 465694 78552 465750
rect 78608 465694 78678 465750
rect 70130 465688 78678 465694
rect 70000 465626 78678 465688
rect 70000 465620 77808 465626
rect 70000 465564 70074 465620
rect 70130 465570 77808 465620
rect 77864 465570 77932 465626
rect 77988 465570 78056 465626
rect 78112 465570 78180 465626
rect 78236 465570 78304 465626
rect 78360 465570 78428 465626
rect 78484 465570 78552 465626
rect 78608 465570 78678 465626
rect 70130 465564 78678 465570
rect 70000 465502 78678 465564
rect 70000 465496 77808 465502
rect 70000 465440 70074 465496
rect 70130 465446 77808 465496
rect 77864 465446 77932 465502
rect 77988 465446 78056 465502
rect 78112 465446 78180 465502
rect 78236 465446 78304 465502
rect 78360 465446 78428 465502
rect 78484 465446 78552 465502
rect 78608 465446 78678 465502
rect 70130 465440 78678 465446
rect 70000 465378 78678 465440
rect 70000 465372 77808 465378
rect 70000 465316 70074 465372
rect 70130 465322 77808 465372
rect 77864 465322 77932 465378
rect 77988 465322 78056 465378
rect 78112 465322 78180 465378
rect 78236 465322 78304 465378
rect 78360 465322 78428 465378
rect 78484 465322 78552 465378
rect 78608 465322 78678 465378
rect 70130 465316 78678 465322
rect 70000 465254 78678 465316
rect 70000 465248 77808 465254
rect 70000 465192 70074 465248
rect 70130 465198 77808 465248
rect 77864 465198 77932 465254
rect 77988 465198 78056 465254
rect 78112 465198 78180 465254
rect 78236 465198 78304 465254
rect 78360 465198 78428 465254
rect 78484 465198 78552 465254
rect 78608 465198 78678 465254
rect 70130 465192 78678 465198
rect 70000 465122 78678 465192
rect 70000 464744 78678 464802
rect 70000 464738 77808 464744
rect 70000 464682 70074 464738
rect 70130 464688 77808 464738
rect 77864 464688 77932 464744
rect 77988 464688 78056 464744
rect 78112 464688 78180 464744
rect 78236 464688 78304 464744
rect 78360 464688 78428 464744
rect 78484 464688 78552 464744
rect 78608 464688 78678 464744
rect 70130 464682 78678 464688
rect 70000 464620 78678 464682
rect 70000 464614 77808 464620
rect 70000 464558 70074 464614
rect 70130 464564 77808 464614
rect 77864 464564 77932 464620
rect 77988 464564 78056 464620
rect 78112 464564 78180 464620
rect 78236 464564 78304 464620
rect 78360 464564 78428 464620
rect 78484 464564 78552 464620
rect 78608 464564 78678 464620
rect 70130 464558 78678 464564
rect 70000 464496 78678 464558
rect 70000 464490 77808 464496
rect 70000 464434 70074 464490
rect 70130 464440 77808 464490
rect 77864 464440 77932 464496
rect 77988 464440 78056 464496
rect 78112 464440 78180 464496
rect 78236 464440 78304 464496
rect 78360 464440 78428 464496
rect 78484 464440 78552 464496
rect 78608 464440 78678 464496
rect 70130 464434 78678 464440
rect 70000 464372 78678 464434
rect 70000 464366 77808 464372
rect 70000 464310 70074 464366
rect 70130 464316 77808 464366
rect 77864 464316 77932 464372
rect 77988 464316 78056 464372
rect 78112 464316 78180 464372
rect 78236 464316 78304 464372
rect 78360 464316 78428 464372
rect 78484 464316 78552 464372
rect 78608 464316 78678 464372
rect 70130 464310 78678 464316
rect 70000 464248 78678 464310
rect 70000 464242 77808 464248
rect 70000 464186 70074 464242
rect 70130 464192 77808 464242
rect 77864 464192 77932 464248
rect 77988 464192 78056 464248
rect 78112 464192 78180 464248
rect 78236 464192 78304 464248
rect 78360 464192 78428 464248
rect 78484 464192 78552 464248
rect 78608 464192 78678 464248
rect 70130 464186 78678 464192
rect 70000 464124 78678 464186
rect 70000 464118 77808 464124
rect 70000 464062 70074 464118
rect 70130 464068 77808 464118
rect 77864 464068 77932 464124
rect 77988 464068 78056 464124
rect 78112 464068 78180 464124
rect 78236 464068 78304 464124
rect 78360 464068 78428 464124
rect 78484 464068 78552 464124
rect 78608 464068 78678 464124
rect 70130 464062 78678 464068
rect 70000 464000 78678 464062
rect 688372 464429 698922 464630
rect 688372 464373 698144 464429
rect 698200 464373 698444 464429
rect 698500 464373 698744 464429
rect 698800 464373 698922 464429
rect 688372 464229 698922 464373
rect 688372 464173 698144 464229
rect 698200 464173 698444 464229
rect 698500 464173 698744 464229
rect 698800 464173 698922 464229
rect 688372 464010 698922 464173
rect 70000 463994 77808 464000
rect 70000 463938 70074 463994
rect 70130 463944 77808 463994
rect 77864 463944 77932 464000
rect 77988 463944 78056 464000
rect 78112 463944 78180 464000
rect 78236 463944 78304 464000
rect 78360 463944 78428 464000
rect 78484 463944 78552 464000
rect 78608 463944 78678 464000
rect 70130 463938 78678 463944
rect 70000 463876 78678 463938
rect 70000 463870 77808 463876
rect 70000 463814 70074 463870
rect 70130 463820 77808 463870
rect 77864 463820 77932 463876
rect 77988 463820 78056 463876
rect 78112 463820 78180 463876
rect 78236 463820 78304 463876
rect 78360 463820 78428 463876
rect 78484 463820 78552 463876
rect 78608 463820 78678 463876
rect 70130 463814 78678 463820
rect 70000 463752 78678 463814
rect 70000 463746 77808 463752
rect 70000 463690 70074 463746
rect 70130 463696 77808 463746
rect 77864 463696 77932 463752
rect 77988 463696 78056 463752
rect 78112 463696 78180 463752
rect 78236 463696 78304 463752
rect 78360 463696 78428 463752
rect 78484 463696 78552 463752
rect 78608 463696 78678 463752
rect 70130 463690 78678 463696
rect 70000 463628 78678 463690
rect 70000 463622 77808 463628
rect 70000 463566 70074 463622
rect 70130 463572 77808 463622
rect 77864 463572 77932 463628
rect 77988 463572 78056 463628
rect 78112 463572 78180 463628
rect 78236 463572 78304 463628
rect 78360 463572 78428 463628
rect 78484 463572 78552 463628
rect 78608 463572 78678 463628
rect 70130 463566 78678 463572
rect 70000 463504 78678 463566
rect 70000 463498 77808 463504
rect 70000 463442 70074 463498
rect 70130 463448 77808 463498
rect 77864 463448 77932 463504
rect 77988 463448 78056 463504
rect 78112 463448 78180 463504
rect 78236 463448 78304 463504
rect 78360 463448 78428 463504
rect 78484 463448 78552 463504
rect 78608 463448 78678 463504
rect 70130 463442 78678 463448
rect 70000 463380 78678 463442
rect 70000 463374 77808 463380
rect 70000 463318 70074 463374
rect 70130 463324 77808 463374
rect 77864 463324 77932 463380
rect 77988 463324 78056 463380
rect 78112 463324 78180 463380
rect 78236 463324 78304 463380
rect 78360 463324 78428 463380
rect 78484 463324 78552 463380
rect 78608 463324 78678 463380
rect 70130 463318 78678 463324
rect 70000 463256 78678 463318
rect 70000 463250 77808 463256
rect 70000 463194 70074 463250
rect 70130 463200 77808 463250
rect 77864 463200 77932 463256
rect 77988 463200 78056 463256
rect 78112 463200 78180 463256
rect 78236 463200 78304 463256
rect 78360 463200 78428 463256
rect 78484 463200 78552 463256
rect 78608 463200 78678 463256
rect 70130 463194 78678 463200
rect 70000 463132 78678 463194
rect 70000 463126 77808 463132
rect 70000 463070 70074 463126
rect 70130 463076 77808 463126
rect 77864 463076 77932 463132
rect 77988 463076 78056 463132
rect 78112 463076 78180 463132
rect 78236 463076 78304 463132
rect 78360 463076 78428 463132
rect 78484 463076 78552 463132
rect 78608 463076 78678 463132
rect 70130 463070 78678 463076
rect 70000 463008 78678 463070
rect 70000 463002 77808 463008
rect 70000 462946 70074 463002
rect 70130 462952 77808 463002
rect 77864 462952 77932 463008
rect 77988 462952 78056 463008
rect 78112 462952 78180 463008
rect 78236 462952 78304 463008
rect 78360 462952 78428 463008
rect 78484 462952 78552 463008
rect 78608 462952 78678 463008
rect 70130 462946 78678 462952
rect 70000 462884 78678 462946
rect 70000 462878 77808 462884
rect 70000 462822 70074 462878
rect 70130 462828 77808 462878
rect 77864 462828 77932 462884
rect 77988 462828 78056 462884
rect 78112 462828 78180 462884
rect 78236 462828 78304 462884
rect 78360 462828 78428 462884
rect 78484 462828 78552 462884
rect 78608 462828 78678 462884
rect 70130 462822 78678 462828
rect 70000 462752 78678 462822
rect 70000 462140 78678 462172
rect 70000 462134 77808 462140
rect 70000 462078 70074 462134
rect 70130 462084 77808 462134
rect 77864 462084 77932 462140
rect 77988 462084 78056 462140
rect 78112 462084 78180 462140
rect 78236 462084 78304 462140
rect 78360 462084 78428 462140
rect 78484 462084 78552 462140
rect 78608 462084 78678 462140
rect 70130 462078 78678 462084
rect 70000 462016 78678 462078
rect 70000 462010 77808 462016
rect 70000 461954 70074 462010
rect 70130 461960 77808 462010
rect 77864 461960 77932 462016
rect 77988 461960 78056 462016
rect 78112 461960 78180 462016
rect 78236 461960 78304 462016
rect 78360 461960 78428 462016
rect 78484 461960 78552 462016
rect 78608 461960 78678 462016
rect 70130 461954 78678 461960
rect 70000 461892 78678 461954
rect 70000 461886 77808 461892
rect 70000 461830 70074 461886
rect 70130 461836 77808 461886
rect 77864 461836 77932 461892
rect 77988 461836 78056 461892
rect 78112 461836 78180 461892
rect 78236 461836 78304 461892
rect 78360 461836 78428 461892
rect 78484 461836 78552 461892
rect 78608 461836 78678 461892
rect 70130 461830 78678 461836
rect 70000 461768 78678 461830
rect 70000 461762 77808 461768
rect 70000 461706 70074 461762
rect 70130 461712 77808 461762
rect 77864 461712 77932 461768
rect 77988 461712 78056 461768
rect 78112 461712 78180 461768
rect 78236 461712 78304 461768
rect 78360 461712 78428 461768
rect 78484 461712 78552 461768
rect 78608 461712 78678 461768
rect 70130 461706 78678 461712
rect 70000 461644 78678 461706
rect 70000 461638 77808 461644
rect 70000 461582 70074 461638
rect 70130 461588 77808 461638
rect 77864 461588 77932 461644
rect 77988 461588 78056 461644
rect 78112 461588 78180 461644
rect 78236 461588 78304 461644
rect 78360 461588 78428 461644
rect 78484 461588 78552 461644
rect 78608 461588 78678 461644
rect 70130 461582 78678 461588
rect 70000 461520 78678 461582
rect 70000 461514 77808 461520
rect 70000 461458 70074 461514
rect 70130 461464 77808 461514
rect 77864 461464 77932 461520
rect 77988 461464 78056 461520
rect 78112 461464 78180 461520
rect 78236 461464 78304 461520
rect 78360 461464 78428 461520
rect 78484 461464 78552 461520
rect 78608 461464 78678 461520
rect 70130 461458 78678 461464
rect 70000 461396 78678 461458
rect 70000 461390 77808 461396
rect 70000 461334 70074 461390
rect 70130 461340 77808 461390
rect 77864 461340 77932 461396
rect 77988 461340 78056 461396
rect 78112 461340 78180 461396
rect 78236 461340 78304 461396
rect 78360 461340 78428 461396
rect 78484 461340 78552 461396
rect 78608 461340 78678 461396
rect 70130 461334 78678 461340
rect 70000 461272 78678 461334
rect 70000 461266 77808 461272
rect 70000 461210 70074 461266
rect 70130 461216 77808 461266
rect 77864 461216 77932 461272
rect 77988 461216 78056 461272
rect 78112 461216 78180 461272
rect 78236 461216 78304 461272
rect 78360 461216 78428 461272
rect 78484 461216 78552 461272
rect 78608 461216 78678 461272
rect 70130 461210 78678 461216
rect 70000 461148 78678 461210
rect 70000 461142 77808 461148
rect 70000 461086 70074 461142
rect 70130 461092 77808 461142
rect 77864 461092 77932 461148
rect 77988 461092 78056 461148
rect 78112 461092 78180 461148
rect 78236 461092 78304 461148
rect 78360 461092 78428 461148
rect 78484 461092 78552 461148
rect 78608 461092 78678 461148
rect 70130 461086 78678 461092
rect 70000 461024 78678 461086
rect 70000 461018 77808 461024
rect 70000 460962 70074 461018
rect 70130 460968 77808 461018
rect 77864 460968 77932 461024
rect 77988 460968 78056 461024
rect 78112 460968 78180 461024
rect 78236 460968 78304 461024
rect 78360 460968 78428 461024
rect 78484 460968 78552 461024
rect 78608 460968 78678 461024
rect 70130 460962 78678 460968
rect 70000 460900 78678 460962
rect 70000 460894 77808 460900
rect 70000 460838 70074 460894
rect 70130 460844 77808 460894
rect 77864 460844 77932 460900
rect 77988 460844 78056 460900
rect 78112 460844 78180 460900
rect 78236 460844 78304 460900
rect 78360 460844 78428 460900
rect 78484 460844 78552 460900
rect 78608 460844 78678 460900
rect 70130 460838 78678 460844
rect 70000 460776 78678 460838
rect 70000 460770 77808 460776
rect 70000 460714 70074 460770
rect 70130 460720 77808 460770
rect 77864 460720 77932 460776
rect 77988 460720 78056 460776
rect 78112 460720 78180 460776
rect 78236 460720 78304 460776
rect 78360 460720 78428 460776
rect 78484 460720 78552 460776
rect 78608 460720 78678 460776
rect 70130 460714 78678 460720
rect 70000 460652 78678 460714
rect 70000 460646 77808 460652
rect 70000 460590 70074 460646
rect 70130 460596 77808 460646
rect 77864 460596 77932 460652
rect 77988 460596 78056 460652
rect 78112 460596 78180 460652
rect 78236 460596 78304 460652
rect 78360 460596 78428 460652
rect 78484 460596 78552 460652
rect 78608 460596 78678 460652
rect 70130 460590 78678 460596
rect 70000 460528 78678 460590
rect 70000 460522 77808 460528
rect 70000 460466 70074 460522
rect 70130 460472 77808 460522
rect 77864 460472 77932 460528
rect 77988 460472 78056 460528
rect 78112 460472 78180 460528
rect 78236 460472 78304 460528
rect 78360 460472 78428 460528
rect 78484 460472 78552 460528
rect 78608 460472 78678 460528
rect 70130 460466 78678 460472
rect 70000 460404 78678 460466
rect 70000 460398 77808 460404
rect 70000 460342 70074 460398
rect 70130 460348 77808 460398
rect 77864 460348 77932 460404
rect 77988 460348 78056 460404
rect 78112 460348 78180 460404
rect 78236 460348 78304 460404
rect 78360 460348 78428 460404
rect 78484 460348 78552 460404
rect 78608 460348 78678 460404
rect 70130 460342 78678 460348
rect 70000 460272 78678 460342
rect 697922 453658 708000 453728
rect 697922 453652 707870 453658
rect 697922 453596 697992 453652
rect 698048 453596 698116 453652
rect 698172 453596 698240 453652
rect 698296 453596 698364 453652
rect 698420 453596 698488 453652
rect 698544 453596 698612 453652
rect 698668 453596 698736 453652
rect 698792 453602 707870 453652
rect 707926 453602 708000 453658
rect 698792 453596 708000 453602
rect 697922 453534 708000 453596
rect 697922 453528 707870 453534
rect 697922 453472 697992 453528
rect 698048 453472 698116 453528
rect 698172 453472 698240 453528
rect 698296 453472 698364 453528
rect 698420 453472 698488 453528
rect 698544 453472 698612 453528
rect 698668 453472 698736 453528
rect 698792 453478 707870 453528
rect 707926 453478 708000 453534
rect 698792 453472 708000 453478
rect 697922 453410 708000 453472
rect 697922 453404 707870 453410
rect 697922 453348 697992 453404
rect 698048 453348 698116 453404
rect 698172 453348 698240 453404
rect 698296 453348 698364 453404
rect 698420 453348 698488 453404
rect 698544 453348 698612 453404
rect 698668 453348 698736 453404
rect 698792 453354 707870 453404
rect 707926 453354 708000 453410
rect 698792 453348 708000 453354
rect 697922 453286 708000 453348
rect 697922 453280 707870 453286
rect 697922 453224 697992 453280
rect 698048 453224 698116 453280
rect 698172 453224 698240 453280
rect 698296 453224 698364 453280
rect 698420 453224 698488 453280
rect 698544 453224 698612 453280
rect 698668 453224 698736 453280
rect 698792 453230 707870 453280
rect 707926 453230 708000 453286
rect 698792 453224 708000 453230
rect 697922 453162 708000 453224
rect 697922 453156 707870 453162
rect 697922 453100 697992 453156
rect 698048 453100 698116 453156
rect 698172 453100 698240 453156
rect 698296 453100 698364 453156
rect 698420 453100 698488 453156
rect 698544 453100 698612 453156
rect 698668 453100 698736 453156
rect 698792 453106 707870 453156
rect 707926 453106 708000 453162
rect 698792 453100 708000 453106
rect 697922 453038 708000 453100
rect 697922 453032 707870 453038
rect 697922 452976 697992 453032
rect 698048 452976 698116 453032
rect 698172 452976 698240 453032
rect 698296 452976 698364 453032
rect 698420 452976 698488 453032
rect 698544 452976 698612 453032
rect 698668 452976 698736 453032
rect 698792 452982 707870 453032
rect 707926 452982 708000 453038
rect 698792 452976 708000 452982
rect 697922 452914 708000 452976
rect 697922 452908 707870 452914
rect 697922 452852 697992 452908
rect 698048 452852 698116 452908
rect 698172 452852 698240 452908
rect 698296 452852 698364 452908
rect 698420 452852 698488 452908
rect 698544 452852 698612 452908
rect 698668 452852 698736 452908
rect 698792 452858 707870 452908
rect 707926 452858 708000 452914
rect 698792 452852 708000 452858
rect 697922 452790 708000 452852
rect 697922 452784 707870 452790
rect 697922 452728 697992 452784
rect 698048 452728 698116 452784
rect 698172 452728 698240 452784
rect 698296 452728 698364 452784
rect 698420 452728 698488 452784
rect 698544 452728 698612 452784
rect 698668 452728 698736 452784
rect 698792 452734 707870 452784
rect 707926 452734 708000 452790
rect 698792 452728 708000 452734
rect 697922 452666 708000 452728
rect 697922 452660 707870 452666
rect 697922 452604 697992 452660
rect 698048 452604 698116 452660
rect 698172 452604 698240 452660
rect 698296 452604 698364 452660
rect 698420 452604 698488 452660
rect 698544 452604 698612 452660
rect 698668 452604 698736 452660
rect 698792 452610 707870 452660
rect 707926 452610 708000 452666
rect 698792 452604 708000 452610
rect 697922 452542 708000 452604
rect 697922 452536 707870 452542
rect 697922 452480 697992 452536
rect 698048 452480 698116 452536
rect 698172 452480 698240 452536
rect 698296 452480 698364 452536
rect 698420 452480 698488 452536
rect 698544 452480 698612 452536
rect 698668 452480 698736 452536
rect 698792 452486 707870 452536
rect 707926 452486 708000 452542
rect 698792 452480 708000 452486
rect 697922 452418 708000 452480
rect 697922 452412 707870 452418
rect 697922 452356 697992 452412
rect 698048 452356 698116 452412
rect 698172 452356 698240 452412
rect 698296 452356 698364 452412
rect 698420 452356 698488 452412
rect 698544 452356 698612 452412
rect 698668 452356 698736 452412
rect 698792 452362 707870 452412
rect 707926 452362 708000 452418
rect 698792 452356 708000 452362
rect 697922 452294 708000 452356
rect 697922 452288 707870 452294
rect 697922 452232 697992 452288
rect 698048 452232 698116 452288
rect 698172 452232 698240 452288
rect 698296 452232 698364 452288
rect 698420 452232 698488 452288
rect 698544 452232 698612 452288
rect 698668 452232 698736 452288
rect 698792 452238 707870 452288
rect 707926 452238 708000 452294
rect 698792 452232 708000 452238
rect 697922 452170 708000 452232
rect 697922 452164 707870 452170
rect 697922 452108 697992 452164
rect 698048 452108 698116 452164
rect 698172 452108 698240 452164
rect 698296 452108 698364 452164
rect 698420 452108 698488 452164
rect 698544 452108 698612 452164
rect 698668 452108 698736 452164
rect 698792 452114 707870 452164
rect 707926 452114 708000 452170
rect 698792 452108 708000 452114
rect 697922 452046 708000 452108
rect 697922 452040 707870 452046
rect 697922 451984 697992 452040
rect 698048 451984 698116 452040
rect 698172 451984 698240 452040
rect 698296 451984 698364 452040
rect 698420 451984 698488 452040
rect 698544 451984 698612 452040
rect 698668 451984 698736 452040
rect 698792 451990 707870 452040
rect 707926 451990 708000 452046
rect 698792 451984 708000 451990
rect 697922 451922 708000 451984
rect 697922 451916 707870 451922
rect 697922 451860 697992 451916
rect 698048 451860 698116 451916
rect 698172 451860 698240 451916
rect 698296 451860 698364 451916
rect 698420 451860 698488 451916
rect 698544 451860 698612 451916
rect 698668 451860 698736 451916
rect 698792 451866 707870 451916
rect 707926 451866 708000 451922
rect 698792 451860 708000 451866
rect 697922 451828 708000 451860
rect 697922 451178 708000 451248
rect 697922 451172 707870 451178
rect 697922 451116 697992 451172
rect 698048 451116 698116 451172
rect 698172 451116 698240 451172
rect 698296 451116 698364 451172
rect 698420 451116 698488 451172
rect 698544 451116 698612 451172
rect 698668 451116 698736 451172
rect 698792 451122 707870 451172
rect 707926 451122 708000 451178
rect 698792 451116 708000 451122
rect 697922 451054 708000 451116
rect 697922 451048 707870 451054
rect 697922 450992 697992 451048
rect 698048 450992 698116 451048
rect 698172 450992 698240 451048
rect 698296 450992 698364 451048
rect 698420 450992 698488 451048
rect 698544 450992 698612 451048
rect 698668 450992 698736 451048
rect 698792 450998 707870 451048
rect 707926 450998 708000 451054
rect 698792 450992 708000 450998
rect 697922 450930 708000 450992
rect 697922 450924 707870 450930
rect 697922 450868 697992 450924
rect 698048 450868 698116 450924
rect 698172 450868 698240 450924
rect 698296 450868 698364 450924
rect 698420 450868 698488 450924
rect 698544 450868 698612 450924
rect 698668 450868 698736 450924
rect 698792 450874 707870 450924
rect 707926 450874 708000 450930
rect 698792 450868 708000 450874
rect 697922 450806 708000 450868
rect 697922 450800 707870 450806
rect 697922 450744 697992 450800
rect 698048 450744 698116 450800
rect 698172 450744 698240 450800
rect 698296 450744 698364 450800
rect 698420 450744 698488 450800
rect 698544 450744 698612 450800
rect 698668 450744 698736 450800
rect 698792 450750 707870 450800
rect 707926 450750 708000 450806
rect 698792 450744 708000 450750
rect 697922 450682 708000 450744
rect 697922 450676 707870 450682
rect 697922 450620 697992 450676
rect 698048 450620 698116 450676
rect 698172 450620 698240 450676
rect 698296 450620 698364 450676
rect 698420 450620 698488 450676
rect 698544 450620 698612 450676
rect 698668 450620 698736 450676
rect 698792 450626 707870 450676
rect 707926 450626 708000 450682
rect 698792 450620 708000 450626
rect 697922 450558 708000 450620
rect 697922 450552 707870 450558
rect 697922 450496 697992 450552
rect 698048 450496 698116 450552
rect 698172 450496 698240 450552
rect 698296 450496 698364 450552
rect 698420 450496 698488 450552
rect 698544 450496 698612 450552
rect 698668 450496 698736 450552
rect 698792 450502 707870 450552
rect 707926 450502 708000 450558
rect 698792 450496 708000 450502
rect 697922 450434 708000 450496
rect 697922 450428 707870 450434
rect 697922 450372 697992 450428
rect 698048 450372 698116 450428
rect 698172 450372 698240 450428
rect 698296 450372 698364 450428
rect 698420 450372 698488 450428
rect 698544 450372 698612 450428
rect 698668 450372 698736 450428
rect 698792 450378 707870 450428
rect 707926 450378 708000 450434
rect 698792 450372 708000 450378
rect 697922 450310 708000 450372
rect 697922 450304 707870 450310
rect 697922 450248 697992 450304
rect 698048 450248 698116 450304
rect 698172 450248 698240 450304
rect 698296 450248 698364 450304
rect 698420 450248 698488 450304
rect 698544 450248 698612 450304
rect 698668 450248 698736 450304
rect 698792 450254 707870 450304
rect 707926 450254 708000 450310
rect 698792 450248 708000 450254
rect 697922 450186 708000 450248
rect 697922 450180 707870 450186
rect 697922 450124 697992 450180
rect 698048 450124 698116 450180
rect 698172 450124 698240 450180
rect 698296 450124 698364 450180
rect 698420 450124 698488 450180
rect 698544 450124 698612 450180
rect 698668 450124 698736 450180
rect 698792 450130 707870 450180
rect 707926 450130 708000 450186
rect 698792 450124 708000 450130
rect 697922 450062 708000 450124
rect 697922 450056 707870 450062
rect 697922 450000 697992 450056
rect 698048 450000 698116 450056
rect 698172 450000 698240 450056
rect 698296 450000 698364 450056
rect 698420 450000 698488 450056
rect 698544 450000 698612 450056
rect 698668 450000 698736 450056
rect 698792 450006 707870 450056
rect 707926 450006 708000 450062
rect 698792 450000 708000 450006
rect 697922 449938 708000 450000
rect 697922 449932 707870 449938
rect 697922 449876 697992 449932
rect 698048 449876 698116 449932
rect 698172 449876 698240 449932
rect 698296 449876 698364 449932
rect 698420 449876 698488 449932
rect 698544 449876 698612 449932
rect 698668 449876 698736 449932
rect 698792 449882 707870 449932
rect 707926 449882 708000 449938
rect 698792 449876 708000 449882
rect 697922 449814 708000 449876
rect 697922 449808 707870 449814
rect 697922 449752 697992 449808
rect 698048 449752 698116 449808
rect 698172 449752 698240 449808
rect 698296 449752 698364 449808
rect 698420 449752 698488 449808
rect 698544 449752 698612 449808
rect 698668 449752 698736 449808
rect 698792 449758 707870 449808
rect 707926 449758 708000 449814
rect 698792 449752 708000 449758
rect 697922 449690 708000 449752
rect 697922 449684 707870 449690
rect 697922 449628 697992 449684
rect 698048 449628 698116 449684
rect 698172 449628 698240 449684
rect 698296 449628 698364 449684
rect 698420 449628 698488 449684
rect 698544 449628 698612 449684
rect 698668 449628 698736 449684
rect 698792 449634 707870 449684
rect 707926 449634 708000 449690
rect 698792 449628 708000 449634
rect 697922 449566 708000 449628
rect 697922 449560 707870 449566
rect 697922 449504 697992 449560
rect 698048 449504 698116 449560
rect 698172 449504 698240 449560
rect 698296 449504 698364 449560
rect 698420 449504 698488 449560
rect 698544 449504 698612 449560
rect 698668 449504 698736 449560
rect 698792 449510 707870 449560
rect 707926 449510 708000 449566
rect 698792 449504 708000 449510
rect 697922 449442 708000 449504
rect 697922 449436 707870 449442
rect 697922 449380 697992 449436
rect 698048 449380 698116 449436
rect 698172 449380 698240 449436
rect 698296 449380 698364 449436
rect 698420 449380 698488 449436
rect 698544 449380 698612 449436
rect 698668 449380 698736 449436
rect 698792 449386 707870 449436
rect 707926 449386 708000 449442
rect 698792 449380 708000 449386
rect 697922 449318 708000 449380
rect 697922 449312 707870 449318
rect 697922 449256 697992 449312
rect 698048 449256 698116 449312
rect 698172 449256 698240 449312
rect 698296 449256 698364 449312
rect 698420 449256 698488 449312
rect 698544 449256 698612 449312
rect 698668 449256 698736 449312
rect 698792 449262 707870 449312
rect 707926 449262 708000 449318
rect 698792 449256 708000 449262
rect 697922 449198 708000 449256
rect 697922 448808 708000 448878
rect 697922 448802 707870 448808
rect 697922 448746 697992 448802
rect 698048 448746 698116 448802
rect 698172 448746 698240 448802
rect 698296 448746 698364 448802
rect 698420 448746 698488 448802
rect 698544 448746 698612 448802
rect 698668 448746 698736 448802
rect 698792 448752 707870 448802
rect 707926 448752 708000 448808
rect 698792 448746 708000 448752
rect 697922 448684 708000 448746
rect 697922 448678 707870 448684
rect 697922 448622 697992 448678
rect 698048 448622 698116 448678
rect 698172 448622 698240 448678
rect 698296 448622 698364 448678
rect 698420 448622 698488 448678
rect 698544 448622 698612 448678
rect 698668 448622 698736 448678
rect 698792 448628 707870 448678
rect 707926 448628 708000 448684
rect 698792 448622 708000 448628
rect 697922 448560 708000 448622
rect 697922 448554 707870 448560
rect 697922 448498 697992 448554
rect 698048 448498 698116 448554
rect 698172 448498 698240 448554
rect 698296 448498 698364 448554
rect 698420 448498 698488 448554
rect 698544 448498 698612 448554
rect 698668 448498 698736 448554
rect 698792 448504 707870 448554
rect 707926 448504 708000 448560
rect 698792 448498 708000 448504
rect 697922 448436 708000 448498
rect 697922 448430 707870 448436
rect 697922 448374 697992 448430
rect 698048 448374 698116 448430
rect 698172 448374 698240 448430
rect 698296 448374 698364 448430
rect 698420 448374 698488 448430
rect 698544 448374 698612 448430
rect 698668 448374 698736 448430
rect 698792 448380 707870 448430
rect 707926 448380 708000 448436
rect 698792 448374 708000 448380
rect 697922 448312 708000 448374
rect 697922 448306 707870 448312
rect 697922 448250 697992 448306
rect 698048 448250 698116 448306
rect 698172 448250 698240 448306
rect 698296 448250 698364 448306
rect 698420 448250 698488 448306
rect 698544 448250 698612 448306
rect 698668 448250 698736 448306
rect 698792 448256 707870 448306
rect 707926 448256 708000 448312
rect 698792 448250 708000 448256
rect 697922 448188 708000 448250
rect 697922 448182 707870 448188
rect 697922 448126 697992 448182
rect 698048 448126 698116 448182
rect 698172 448126 698240 448182
rect 698296 448126 698364 448182
rect 698420 448126 698488 448182
rect 698544 448126 698612 448182
rect 698668 448126 698736 448182
rect 698792 448132 707870 448182
rect 707926 448132 708000 448188
rect 698792 448126 708000 448132
rect 697922 448064 708000 448126
rect 697922 448058 707870 448064
rect 697922 448002 697992 448058
rect 698048 448002 698116 448058
rect 698172 448002 698240 448058
rect 698296 448002 698364 448058
rect 698420 448002 698488 448058
rect 698544 448002 698612 448058
rect 698668 448002 698736 448058
rect 698792 448008 707870 448058
rect 707926 448008 708000 448064
rect 698792 448002 708000 448008
rect 697922 447940 708000 448002
rect 697922 447934 707870 447940
rect 697922 447878 697992 447934
rect 698048 447878 698116 447934
rect 698172 447878 698240 447934
rect 698296 447878 698364 447934
rect 698420 447878 698488 447934
rect 698544 447878 698612 447934
rect 698668 447878 698736 447934
rect 698792 447884 707870 447934
rect 707926 447884 708000 447940
rect 698792 447878 708000 447884
rect 697922 447816 708000 447878
rect 697922 447810 707870 447816
rect 697922 447754 697992 447810
rect 698048 447754 698116 447810
rect 698172 447754 698240 447810
rect 698296 447754 698364 447810
rect 698420 447754 698488 447810
rect 698544 447754 698612 447810
rect 698668 447754 698736 447810
rect 698792 447760 707870 447810
rect 707926 447760 708000 447816
rect 698792 447754 708000 447760
rect 697922 447692 708000 447754
rect 697922 447686 707870 447692
rect 697922 447630 697992 447686
rect 698048 447630 698116 447686
rect 698172 447630 698240 447686
rect 698296 447630 698364 447686
rect 698420 447630 698488 447686
rect 698544 447630 698612 447686
rect 698668 447630 698736 447686
rect 698792 447636 707870 447686
rect 707926 447636 708000 447692
rect 698792 447630 708000 447636
rect 697922 447568 708000 447630
rect 697922 447562 707870 447568
rect 697922 447506 697992 447562
rect 698048 447506 698116 447562
rect 698172 447506 698240 447562
rect 698296 447506 698364 447562
rect 698420 447506 698488 447562
rect 698544 447506 698612 447562
rect 698668 447506 698736 447562
rect 698792 447512 707870 447562
rect 707926 447512 708000 447568
rect 698792 447506 708000 447512
rect 697922 447444 708000 447506
rect 697922 447438 707870 447444
rect 697922 447382 697992 447438
rect 698048 447382 698116 447438
rect 698172 447382 698240 447438
rect 698296 447382 698364 447438
rect 698420 447382 698488 447438
rect 698544 447382 698612 447438
rect 698668 447382 698736 447438
rect 698792 447388 707870 447438
rect 707926 447388 708000 447444
rect 698792 447382 708000 447388
rect 697922 447320 708000 447382
rect 697922 447314 707870 447320
rect 697922 447258 697992 447314
rect 698048 447258 698116 447314
rect 698172 447258 698240 447314
rect 698296 447258 698364 447314
rect 698420 447258 698488 447314
rect 698544 447258 698612 447314
rect 698668 447258 698736 447314
rect 698792 447264 707870 447314
rect 707926 447264 708000 447320
rect 698792 447258 708000 447264
rect 697922 447196 708000 447258
rect 697922 447190 707870 447196
rect 697922 447134 697992 447190
rect 698048 447134 698116 447190
rect 698172 447134 698240 447190
rect 698296 447134 698364 447190
rect 698420 447134 698488 447190
rect 698544 447134 698612 447190
rect 698668 447134 698736 447190
rect 698792 447140 707870 447190
rect 707926 447140 708000 447196
rect 698792 447134 708000 447140
rect 697922 447072 708000 447134
rect 697922 447066 707870 447072
rect 697922 447010 697992 447066
rect 698048 447010 698116 447066
rect 698172 447010 698240 447066
rect 698296 447010 698364 447066
rect 698420 447010 698488 447066
rect 698544 447010 698612 447066
rect 698668 447010 698736 447066
rect 698792 447016 707870 447066
rect 707926 447016 708000 447072
rect 698792 447010 708000 447016
rect 697922 446948 708000 447010
rect 697922 446942 707870 446948
rect 697922 446886 697992 446942
rect 698048 446886 698116 446942
rect 698172 446886 698240 446942
rect 698296 446886 698364 446942
rect 698420 446886 698488 446942
rect 698544 446886 698612 446942
rect 698668 446886 698736 446942
rect 698792 446892 707870 446942
rect 707926 446892 708000 446948
rect 698792 446886 708000 446892
rect 697922 446828 708000 446886
rect 77678 446429 84516 446630
rect 77678 446373 77800 446429
rect 77856 446373 78100 446429
rect 78156 446373 78400 446429
rect 78456 446373 84516 446429
rect 77678 446229 84516 446373
rect 77678 446173 77800 446229
rect 77856 446173 78100 446229
rect 78156 446173 78400 446229
rect 78456 446173 84516 446229
rect 77678 446010 84516 446173
rect 697922 446102 708000 446172
rect 697922 446096 707870 446102
rect 697922 446040 697992 446096
rect 698048 446040 698116 446096
rect 698172 446040 698240 446096
rect 698296 446040 698364 446096
rect 698420 446040 698488 446096
rect 698544 446040 698612 446096
rect 698668 446040 698736 446096
rect 698792 446046 707870 446096
rect 707926 446046 708000 446102
rect 698792 446040 708000 446046
rect 697922 445978 708000 446040
rect 697922 445972 707870 445978
rect 697922 445916 697992 445972
rect 698048 445916 698116 445972
rect 698172 445916 698240 445972
rect 698296 445916 698364 445972
rect 698420 445916 698488 445972
rect 698544 445916 698612 445972
rect 698668 445916 698736 445972
rect 698792 445922 707870 445972
rect 707926 445922 708000 445978
rect 698792 445916 708000 445922
rect 697922 445854 708000 445916
rect 697922 445848 707870 445854
rect 697922 445792 697992 445848
rect 698048 445792 698116 445848
rect 698172 445792 698240 445848
rect 698296 445792 698364 445848
rect 698420 445792 698488 445848
rect 698544 445792 698612 445848
rect 698668 445792 698736 445848
rect 698792 445798 707870 445848
rect 707926 445798 708000 445854
rect 698792 445792 708000 445798
rect 697922 445730 708000 445792
rect 697922 445724 707870 445730
rect 697922 445668 697992 445724
rect 698048 445668 698116 445724
rect 698172 445668 698240 445724
rect 698296 445668 698364 445724
rect 698420 445668 698488 445724
rect 698544 445668 698612 445724
rect 698668 445668 698736 445724
rect 698792 445674 707870 445724
rect 707926 445674 708000 445730
rect 698792 445668 708000 445674
rect 697922 445606 708000 445668
rect 697922 445600 707870 445606
rect 697922 445544 697992 445600
rect 698048 445544 698116 445600
rect 698172 445544 698240 445600
rect 698296 445544 698364 445600
rect 698420 445544 698488 445600
rect 698544 445544 698612 445600
rect 698668 445544 698736 445600
rect 698792 445550 707870 445600
rect 707926 445550 708000 445606
rect 698792 445544 708000 445550
rect 697922 445482 708000 445544
rect 697922 445476 707870 445482
rect 697922 445420 697992 445476
rect 698048 445420 698116 445476
rect 698172 445420 698240 445476
rect 698296 445420 698364 445476
rect 698420 445420 698488 445476
rect 698544 445420 698612 445476
rect 698668 445420 698736 445476
rect 698792 445426 707870 445476
rect 707926 445426 708000 445482
rect 698792 445420 708000 445426
rect 697922 445358 708000 445420
rect 697922 445352 707870 445358
rect 697922 445296 697992 445352
rect 698048 445296 698116 445352
rect 698172 445296 698240 445352
rect 698296 445296 698364 445352
rect 698420 445296 698488 445352
rect 698544 445296 698612 445352
rect 698668 445296 698736 445352
rect 698792 445302 707870 445352
rect 707926 445302 708000 445358
rect 698792 445296 708000 445302
rect 697922 445234 708000 445296
rect 697922 445228 707870 445234
rect 697922 445172 697992 445228
rect 698048 445172 698116 445228
rect 698172 445172 698240 445228
rect 698296 445172 698364 445228
rect 698420 445172 698488 445228
rect 698544 445172 698612 445228
rect 698668 445172 698736 445228
rect 698792 445178 707870 445228
rect 707926 445178 708000 445234
rect 698792 445172 708000 445178
rect 697922 445110 708000 445172
rect 697922 445104 707870 445110
rect 697922 445048 697992 445104
rect 698048 445048 698116 445104
rect 698172 445048 698240 445104
rect 698296 445048 698364 445104
rect 698420 445048 698488 445104
rect 698544 445048 698612 445104
rect 698668 445048 698736 445104
rect 698792 445054 707870 445104
rect 707926 445054 708000 445110
rect 698792 445048 708000 445054
rect 697922 444986 708000 445048
rect 697922 444980 707870 444986
rect 697922 444924 697992 444980
rect 698048 444924 698116 444980
rect 698172 444924 698240 444980
rect 698296 444924 698364 444980
rect 698420 444924 698488 444980
rect 698544 444924 698612 444980
rect 698668 444924 698736 444980
rect 698792 444930 707870 444980
rect 707926 444930 708000 444986
rect 698792 444924 708000 444930
rect 697922 444862 708000 444924
rect 697922 444856 707870 444862
rect 697922 444800 697992 444856
rect 698048 444800 698116 444856
rect 698172 444800 698240 444856
rect 698296 444800 698364 444856
rect 698420 444800 698488 444856
rect 698544 444800 698612 444856
rect 698668 444800 698736 444856
rect 698792 444806 707870 444856
rect 707926 444806 708000 444862
rect 698792 444800 708000 444806
rect 697922 444738 708000 444800
rect 697922 444732 707870 444738
rect 697922 444676 697992 444732
rect 698048 444676 698116 444732
rect 698172 444676 698240 444732
rect 698296 444676 698364 444732
rect 698420 444676 698488 444732
rect 698544 444676 698612 444732
rect 698668 444676 698736 444732
rect 698792 444682 707870 444732
rect 707926 444682 708000 444738
rect 698792 444676 708000 444682
rect 697922 444614 708000 444676
rect 697922 444608 707870 444614
rect 697922 444552 697992 444608
rect 698048 444552 698116 444608
rect 698172 444552 698240 444608
rect 698296 444552 698364 444608
rect 698420 444552 698488 444608
rect 698544 444552 698612 444608
rect 698668 444552 698736 444608
rect 698792 444558 707870 444608
rect 707926 444558 708000 444614
rect 698792 444552 708000 444558
rect 697922 444490 708000 444552
rect 697922 444484 707870 444490
rect 697922 444428 697992 444484
rect 698048 444428 698116 444484
rect 698172 444428 698240 444484
rect 698296 444428 698364 444484
rect 698420 444428 698488 444484
rect 698544 444428 698612 444484
rect 698668 444428 698736 444484
rect 698792 444434 707870 444484
rect 707926 444434 708000 444490
rect 698792 444428 708000 444434
rect 697922 444366 708000 444428
rect 697922 444360 707870 444366
rect 697922 444304 697992 444360
rect 698048 444304 698116 444360
rect 698172 444304 698240 444360
rect 698296 444304 698364 444360
rect 698420 444304 698488 444360
rect 698544 444304 698612 444360
rect 698668 444304 698736 444360
rect 698792 444310 707870 444360
rect 707926 444310 708000 444366
rect 698792 444304 708000 444310
rect 697922 444242 708000 444304
rect 697922 444236 707870 444242
rect 697922 444180 697992 444236
rect 698048 444180 698116 444236
rect 698172 444180 698240 444236
rect 698296 444180 698364 444236
rect 698420 444180 698488 444236
rect 698544 444180 698612 444236
rect 698668 444180 698736 444236
rect 698792 444186 707870 444236
rect 707926 444186 708000 444242
rect 698792 444180 708000 444186
rect 697922 444122 708000 444180
rect 697922 443732 708000 443802
rect 697922 443726 707870 443732
rect 697922 443670 697992 443726
rect 698048 443670 698116 443726
rect 698172 443670 698240 443726
rect 698296 443670 698364 443726
rect 698420 443670 698488 443726
rect 698544 443670 698612 443726
rect 698668 443670 698736 443726
rect 698792 443676 707870 443726
rect 707926 443676 708000 443732
rect 698792 443670 708000 443676
rect 697922 443608 708000 443670
rect 697922 443602 707870 443608
rect 697922 443546 697992 443602
rect 698048 443546 698116 443602
rect 698172 443546 698240 443602
rect 698296 443546 698364 443602
rect 698420 443546 698488 443602
rect 698544 443546 698612 443602
rect 698668 443546 698736 443602
rect 698792 443552 707870 443602
rect 707926 443552 708000 443608
rect 698792 443546 708000 443552
rect 697922 443484 708000 443546
rect 697922 443478 707870 443484
rect 697922 443422 697992 443478
rect 698048 443422 698116 443478
rect 698172 443422 698240 443478
rect 698296 443422 698364 443478
rect 698420 443422 698488 443478
rect 698544 443422 698612 443478
rect 698668 443422 698736 443478
rect 698792 443428 707870 443478
rect 707926 443428 708000 443484
rect 698792 443422 708000 443428
rect 697922 443360 708000 443422
rect 697922 443354 707870 443360
rect 697922 443298 697992 443354
rect 698048 443298 698116 443354
rect 698172 443298 698240 443354
rect 698296 443298 698364 443354
rect 698420 443298 698488 443354
rect 698544 443298 698612 443354
rect 698668 443298 698736 443354
rect 698792 443304 707870 443354
rect 707926 443304 708000 443360
rect 698792 443298 708000 443304
rect 697922 443236 708000 443298
rect 697922 443230 707870 443236
rect 697922 443174 697992 443230
rect 698048 443174 698116 443230
rect 698172 443174 698240 443230
rect 698296 443174 698364 443230
rect 698420 443174 698488 443230
rect 698544 443174 698612 443230
rect 698668 443174 698736 443230
rect 698792 443180 707870 443230
rect 707926 443180 708000 443236
rect 698792 443174 708000 443180
rect 697922 443112 708000 443174
rect 697922 443106 707870 443112
rect 697922 443050 697992 443106
rect 698048 443050 698116 443106
rect 698172 443050 698240 443106
rect 698296 443050 698364 443106
rect 698420 443050 698488 443106
rect 698544 443050 698612 443106
rect 698668 443050 698736 443106
rect 698792 443056 707870 443106
rect 707926 443056 708000 443112
rect 698792 443050 708000 443056
rect 697922 442988 708000 443050
rect 697922 442982 707870 442988
rect 697922 442926 697992 442982
rect 698048 442926 698116 442982
rect 698172 442926 698240 442982
rect 698296 442926 698364 442982
rect 698420 442926 698488 442982
rect 698544 442926 698612 442982
rect 698668 442926 698736 442982
rect 698792 442932 707870 442982
rect 707926 442932 708000 442988
rect 698792 442926 708000 442932
rect 697922 442864 708000 442926
rect 697922 442858 707870 442864
rect 697922 442802 697992 442858
rect 698048 442802 698116 442858
rect 698172 442802 698240 442858
rect 698296 442802 698364 442858
rect 698420 442802 698488 442858
rect 698544 442802 698612 442858
rect 698668 442802 698736 442858
rect 698792 442808 707870 442858
rect 707926 442808 708000 442864
rect 698792 442802 708000 442808
rect 697922 442740 708000 442802
rect 697922 442734 707870 442740
rect 697922 442678 697992 442734
rect 698048 442678 698116 442734
rect 698172 442678 698240 442734
rect 698296 442678 698364 442734
rect 698420 442678 698488 442734
rect 698544 442678 698612 442734
rect 698668 442678 698736 442734
rect 698792 442684 707870 442734
rect 707926 442684 708000 442740
rect 698792 442678 708000 442684
rect 697922 442616 708000 442678
rect 697922 442610 707870 442616
rect 697922 442554 697992 442610
rect 698048 442554 698116 442610
rect 698172 442554 698240 442610
rect 698296 442554 698364 442610
rect 698420 442554 698488 442610
rect 698544 442554 698612 442610
rect 698668 442554 698736 442610
rect 698792 442560 707870 442610
rect 707926 442560 708000 442616
rect 698792 442554 708000 442560
rect 697922 442492 708000 442554
rect 697922 442486 707870 442492
rect 697922 442430 697992 442486
rect 698048 442430 698116 442486
rect 698172 442430 698240 442486
rect 698296 442430 698364 442486
rect 698420 442430 698488 442486
rect 698544 442430 698612 442486
rect 698668 442430 698736 442486
rect 698792 442436 707870 442486
rect 707926 442436 708000 442492
rect 698792 442430 708000 442436
rect 697922 442368 708000 442430
rect 697922 442362 707870 442368
rect 697922 442306 697992 442362
rect 698048 442306 698116 442362
rect 698172 442306 698240 442362
rect 698296 442306 698364 442362
rect 698420 442306 698488 442362
rect 698544 442306 698612 442362
rect 698668 442306 698736 442362
rect 698792 442312 707870 442362
rect 707926 442312 708000 442368
rect 698792 442306 708000 442312
rect 697922 442244 708000 442306
rect 697922 442238 707870 442244
rect 697922 442182 697992 442238
rect 698048 442182 698116 442238
rect 698172 442182 698240 442238
rect 698296 442182 698364 442238
rect 698420 442182 698488 442238
rect 698544 442182 698612 442238
rect 698668 442182 698736 442238
rect 698792 442188 707870 442238
rect 707926 442188 708000 442244
rect 698792 442182 708000 442188
rect 697922 442120 708000 442182
rect 697922 442114 707870 442120
rect 697922 442058 697992 442114
rect 698048 442058 698116 442114
rect 698172 442058 698240 442114
rect 698296 442058 698364 442114
rect 698420 442058 698488 442114
rect 698544 442058 698612 442114
rect 698668 442058 698736 442114
rect 698792 442064 707870 442114
rect 707926 442064 708000 442120
rect 698792 442058 708000 442064
rect 697922 441996 708000 442058
rect 697922 441990 707870 441996
rect 697922 441934 697992 441990
rect 698048 441934 698116 441990
rect 698172 441934 698240 441990
rect 698296 441934 698364 441990
rect 698420 441934 698488 441990
rect 698544 441934 698612 441990
rect 698668 441934 698736 441990
rect 698792 441940 707870 441990
rect 707926 441940 708000 441996
rect 698792 441934 708000 441940
rect 697922 441872 708000 441934
rect 697922 441866 707870 441872
rect 697922 441810 697992 441866
rect 698048 441810 698116 441866
rect 698172 441810 698240 441866
rect 698296 441810 698364 441866
rect 698420 441810 698488 441866
rect 698544 441810 698612 441866
rect 698668 441810 698736 441866
rect 698792 441816 707870 441866
rect 707926 441816 708000 441872
rect 698792 441810 708000 441816
rect 697922 441752 708000 441810
rect 697922 441134 708000 441172
rect 697922 441122 707870 441134
rect 697922 441066 697992 441122
rect 698048 441066 698116 441122
rect 698172 441066 698240 441122
rect 698296 441066 698364 441122
rect 698420 441066 698488 441122
rect 698544 441066 698612 441122
rect 698668 441066 698736 441122
rect 698792 441078 707870 441122
rect 707926 441078 708000 441134
rect 698792 441066 708000 441078
rect 697922 441010 708000 441066
rect 697922 440998 707870 441010
rect 697922 440942 697992 440998
rect 698048 440942 698116 440998
rect 698172 440942 698240 440998
rect 698296 440942 698364 440998
rect 698420 440942 698488 440998
rect 698544 440942 698612 440998
rect 698668 440942 698736 440998
rect 698792 440954 707870 440998
rect 707926 440954 708000 441010
rect 698792 440942 708000 440954
rect 697922 440886 708000 440942
rect 697922 440874 707870 440886
rect 697922 440818 697992 440874
rect 698048 440818 698116 440874
rect 698172 440818 698240 440874
rect 698296 440818 698364 440874
rect 698420 440818 698488 440874
rect 698544 440818 698612 440874
rect 698668 440818 698736 440874
rect 698792 440830 707870 440874
rect 707926 440830 708000 440886
rect 698792 440818 708000 440830
rect 697922 440762 708000 440818
rect 697922 440750 707870 440762
rect 697922 440694 697992 440750
rect 698048 440694 698116 440750
rect 698172 440694 698240 440750
rect 698296 440694 698364 440750
rect 698420 440694 698488 440750
rect 698544 440694 698612 440750
rect 698668 440694 698736 440750
rect 698792 440706 707870 440750
rect 707926 440706 708000 440762
rect 698792 440694 708000 440706
rect 697922 440638 708000 440694
rect 697922 440626 707870 440638
rect 697922 440570 697992 440626
rect 698048 440570 698116 440626
rect 698172 440570 698240 440626
rect 698296 440570 698364 440626
rect 698420 440570 698488 440626
rect 698544 440570 698612 440626
rect 698668 440570 698736 440626
rect 698792 440582 707870 440626
rect 707926 440582 708000 440638
rect 698792 440570 708000 440582
rect 697922 440514 708000 440570
rect 697922 440502 707870 440514
rect 697922 440446 697992 440502
rect 698048 440446 698116 440502
rect 698172 440446 698240 440502
rect 698296 440446 698364 440502
rect 698420 440446 698488 440502
rect 698544 440446 698612 440502
rect 698668 440446 698736 440502
rect 698792 440458 707870 440502
rect 707926 440458 708000 440514
rect 698792 440446 708000 440458
rect 697922 440390 708000 440446
rect 697922 440378 707870 440390
rect 697922 440322 697992 440378
rect 698048 440322 698116 440378
rect 698172 440322 698240 440378
rect 698296 440322 698364 440378
rect 698420 440322 698488 440378
rect 698544 440322 698612 440378
rect 698668 440322 698736 440378
rect 698792 440334 707870 440378
rect 707926 440334 708000 440390
rect 698792 440322 708000 440334
rect 697922 440266 708000 440322
rect 697922 440254 707870 440266
rect 697922 440198 697992 440254
rect 698048 440198 698116 440254
rect 698172 440198 698240 440254
rect 698296 440198 698364 440254
rect 698420 440198 698488 440254
rect 698544 440198 698612 440254
rect 698668 440198 698736 440254
rect 698792 440210 707870 440254
rect 707926 440210 708000 440266
rect 698792 440198 708000 440210
rect 697922 440142 708000 440198
rect 697922 440130 707870 440142
rect 697922 440074 697992 440130
rect 698048 440074 698116 440130
rect 698172 440074 698240 440130
rect 698296 440074 698364 440130
rect 698420 440074 698488 440130
rect 698544 440074 698612 440130
rect 698668 440074 698736 440130
rect 698792 440086 707870 440130
rect 707926 440086 708000 440142
rect 698792 440074 708000 440086
rect 697922 440018 708000 440074
rect 697922 440006 707870 440018
rect 697922 439950 697992 440006
rect 698048 439950 698116 440006
rect 698172 439950 698240 440006
rect 698296 439950 698364 440006
rect 698420 439950 698488 440006
rect 698544 439950 698612 440006
rect 698668 439950 698736 440006
rect 698792 439962 707870 440006
rect 707926 439962 708000 440018
rect 698792 439950 708000 439962
rect 697922 439894 708000 439950
rect 697922 439882 707870 439894
rect 697922 439826 697992 439882
rect 698048 439826 698116 439882
rect 698172 439826 698240 439882
rect 698296 439826 698364 439882
rect 698420 439826 698488 439882
rect 698544 439826 698612 439882
rect 698668 439826 698736 439882
rect 698792 439838 707870 439882
rect 707926 439838 708000 439894
rect 698792 439826 708000 439838
rect 697922 439770 708000 439826
rect 697922 439758 707870 439770
rect 697922 439702 697992 439758
rect 698048 439702 698116 439758
rect 698172 439702 698240 439758
rect 698296 439702 698364 439758
rect 698420 439702 698488 439758
rect 698544 439702 698612 439758
rect 698668 439702 698736 439758
rect 698792 439714 707870 439758
rect 707926 439714 708000 439770
rect 698792 439702 708000 439714
rect 697922 439646 708000 439702
rect 697922 439634 707870 439646
rect 697922 439578 697992 439634
rect 698048 439578 698116 439634
rect 698172 439578 698240 439634
rect 698296 439578 698364 439634
rect 698420 439578 698488 439634
rect 698544 439578 698612 439634
rect 698668 439578 698736 439634
rect 698792 439590 707870 439634
rect 707926 439590 708000 439646
rect 698792 439578 708000 439590
rect 697922 439522 708000 439578
rect 697922 439510 707870 439522
rect 697922 439454 697992 439510
rect 698048 439454 698116 439510
rect 698172 439454 698240 439510
rect 698296 439454 698364 439510
rect 698420 439454 698488 439510
rect 698544 439454 698612 439510
rect 698668 439454 698736 439510
rect 698792 439466 707870 439510
rect 707926 439466 708000 439522
rect 698792 439454 708000 439466
rect 697922 439398 708000 439454
rect 697922 439386 707870 439398
rect 697922 439330 697992 439386
rect 698048 439330 698116 439386
rect 698172 439330 698240 439386
rect 698296 439330 698364 439386
rect 698420 439330 698488 439386
rect 698544 439330 698612 439386
rect 698668 439330 698736 439386
rect 698792 439342 707870 439386
rect 707926 439342 708000 439398
rect 698792 439330 708000 439342
rect 697922 439272 708000 439330
rect 70000 433670 80078 433728
rect 70000 433658 79208 433670
rect 70000 433602 70074 433658
rect 70130 433614 79208 433658
rect 79264 433614 79332 433670
rect 79388 433614 79456 433670
rect 79512 433614 79580 433670
rect 79636 433614 79704 433670
rect 79760 433614 79828 433670
rect 79884 433614 79952 433670
rect 80008 433614 80078 433670
rect 70130 433602 80078 433614
rect 70000 433546 80078 433602
rect 70000 433534 79208 433546
rect 70000 433478 70074 433534
rect 70130 433490 79208 433534
rect 79264 433490 79332 433546
rect 79388 433490 79456 433546
rect 79512 433490 79580 433546
rect 79636 433490 79704 433546
rect 79760 433490 79828 433546
rect 79884 433490 79952 433546
rect 80008 433490 80078 433546
rect 70130 433478 80078 433490
rect 70000 433422 80078 433478
rect 70000 433410 79208 433422
rect 70000 433354 70074 433410
rect 70130 433366 79208 433410
rect 79264 433366 79332 433422
rect 79388 433366 79456 433422
rect 79512 433366 79580 433422
rect 79636 433366 79704 433422
rect 79760 433366 79828 433422
rect 79884 433366 79952 433422
rect 80008 433366 80078 433422
rect 70130 433354 80078 433366
rect 70000 433298 80078 433354
rect 70000 433286 79208 433298
rect 70000 433230 70074 433286
rect 70130 433242 79208 433286
rect 79264 433242 79332 433298
rect 79388 433242 79456 433298
rect 79512 433242 79580 433298
rect 79636 433242 79704 433298
rect 79760 433242 79828 433298
rect 79884 433242 79952 433298
rect 80008 433242 80078 433298
rect 70130 433230 80078 433242
rect 70000 433174 80078 433230
rect 70000 433162 79208 433174
rect 70000 433106 70074 433162
rect 70130 433118 79208 433162
rect 79264 433118 79332 433174
rect 79388 433118 79456 433174
rect 79512 433118 79580 433174
rect 79636 433118 79704 433174
rect 79760 433118 79828 433174
rect 79884 433118 79952 433174
rect 80008 433118 80078 433174
rect 70130 433106 80078 433118
rect 70000 433050 80078 433106
rect 70000 433038 79208 433050
rect 70000 432982 70074 433038
rect 70130 432994 79208 433038
rect 79264 432994 79332 433050
rect 79388 432994 79456 433050
rect 79512 432994 79580 433050
rect 79636 432994 79704 433050
rect 79760 432994 79828 433050
rect 79884 432994 79952 433050
rect 80008 432994 80078 433050
rect 70130 432982 80078 432994
rect 70000 432926 80078 432982
rect 70000 432914 79208 432926
rect 70000 432858 70074 432914
rect 70130 432870 79208 432914
rect 79264 432870 79332 432926
rect 79388 432870 79456 432926
rect 79512 432870 79580 432926
rect 79636 432870 79704 432926
rect 79760 432870 79828 432926
rect 79884 432870 79952 432926
rect 80008 432870 80078 432926
rect 70130 432858 80078 432870
rect 70000 432802 80078 432858
rect 70000 432790 79208 432802
rect 70000 432734 70074 432790
rect 70130 432746 79208 432790
rect 79264 432746 79332 432802
rect 79388 432746 79456 432802
rect 79512 432746 79580 432802
rect 79636 432746 79704 432802
rect 79760 432746 79828 432802
rect 79884 432746 79952 432802
rect 80008 432746 80078 432802
rect 70130 432734 80078 432746
rect 70000 432678 80078 432734
rect 70000 432666 79208 432678
rect 70000 432610 70074 432666
rect 70130 432622 79208 432666
rect 79264 432622 79332 432678
rect 79388 432622 79456 432678
rect 79512 432622 79580 432678
rect 79636 432622 79704 432678
rect 79760 432622 79828 432678
rect 79884 432622 79952 432678
rect 80008 432622 80078 432678
rect 70130 432610 80078 432622
rect 70000 432554 80078 432610
rect 70000 432542 79208 432554
rect 70000 432486 70074 432542
rect 70130 432498 79208 432542
rect 79264 432498 79332 432554
rect 79388 432498 79456 432554
rect 79512 432498 79580 432554
rect 79636 432498 79704 432554
rect 79760 432498 79828 432554
rect 79884 432498 79952 432554
rect 80008 432498 80078 432554
rect 70130 432486 80078 432498
rect 70000 432430 80078 432486
rect 70000 432418 79208 432430
rect 70000 432362 70074 432418
rect 70130 432374 79208 432418
rect 79264 432374 79332 432430
rect 79388 432374 79456 432430
rect 79512 432374 79580 432430
rect 79636 432374 79704 432430
rect 79760 432374 79828 432430
rect 79884 432374 79952 432430
rect 80008 432374 80078 432430
rect 70130 432362 80078 432374
rect 70000 432306 80078 432362
rect 70000 432294 79208 432306
rect 70000 432238 70074 432294
rect 70130 432250 79208 432294
rect 79264 432250 79332 432306
rect 79388 432250 79456 432306
rect 79512 432250 79580 432306
rect 79636 432250 79704 432306
rect 79760 432250 79828 432306
rect 79884 432250 79952 432306
rect 80008 432250 80078 432306
rect 70130 432238 80078 432250
rect 70000 432182 80078 432238
rect 70000 432170 79208 432182
rect 70000 432114 70074 432170
rect 70130 432126 79208 432170
rect 79264 432126 79332 432182
rect 79388 432126 79456 432182
rect 79512 432126 79580 432182
rect 79636 432126 79704 432182
rect 79760 432126 79828 432182
rect 79884 432126 79952 432182
rect 80008 432126 80078 432182
rect 70130 432114 80078 432126
rect 70000 432058 80078 432114
rect 70000 432046 79208 432058
rect 70000 431990 70074 432046
rect 70130 432002 79208 432046
rect 79264 432002 79332 432058
rect 79388 432002 79456 432058
rect 79512 432002 79580 432058
rect 79636 432002 79704 432058
rect 79760 432002 79828 432058
rect 79884 432002 79952 432058
rect 80008 432002 80078 432058
rect 70130 431990 80078 432002
rect 70000 431934 80078 431990
rect 70000 431922 79208 431934
rect 70000 431866 70074 431922
rect 70130 431878 79208 431922
rect 79264 431878 79332 431934
rect 79388 431878 79456 431934
rect 79512 431878 79580 431934
rect 79636 431878 79704 431934
rect 79760 431878 79828 431934
rect 79884 431878 79952 431934
rect 80008 431878 80078 431934
rect 70130 431866 80078 431878
rect 70000 431828 80078 431866
rect 70000 431190 80078 431248
rect 70000 431184 79208 431190
rect 70000 431128 70074 431184
rect 70130 431134 79208 431184
rect 79264 431134 79332 431190
rect 79388 431134 79456 431190
rect 79512 431134 79580 431190
rect 79636 431134 79704 431190
rect 79760 431134 79828 431190
rect 79884 431134 79952 431190
rect 80008 431134 80078 431190
rect 70130 431128 80078 431134
rect 70000 431066 80078 431128
rect 70000 431060 79208 431066
rect 70000 431004 70074 431060
rect 70130 431010 79208 431060
rect 79264 431010 79332 431066
rect 79388 431010 79456 431066
rect 79512 431010 79580 431066
rect 79636 431010 79704 431066
rect 79760 431010 79828 431066
rect 79884 431010 79952 431066
rect 80008 431010 80078 431066
rect 70130 431004 80078 431010
rect 70000 430942 80078 431004
rect 70000 430936 79208 430942
rect 70000 430880 70074 430936
rect 70130 430886 79208 430936
rect 79264 430886 79332 430942
rect 79388 430886 79456 430942
rect 79512 430886 79580 430942
rect 79636 430886 79704 430942
rect 79760 430886 79828 430942
rect 79884 430886 79952 430942
rect 80008 430886 80078 430942
rect 70130 430880 80078 430886
rect 70000 430818 80078 430880
rect 70000 430812 79208 430818
rect 70000 430756 70074 430812
rect 70130 430762 79208 430812
rect 79264 430762 79332 430818
rect 79388 430762 79456 430818
rect 79512 430762 79580 430818
rect 79636 430762 79704 430818
rect 79760 430762 79828 430818
rect 79884 430762 79952 430818
rect 80008 430762 80078 430818
rect 70130 430756 80078 430762
rect 70000 430694 80078 430756
rect 70000 430688 79208 430694
rect 70000 430632 70074 430688
rect 70130 430638 79208 430688
rect 79264 430638 79332 430694
rect 79388 430638 79456 430694
rect 79512 430638 79580 430694
rect 79636 430638 79704 430694
rect 79760 430638 79828 430694
rect 79884 430638 79952 430694
rect 80008 430638 80078 430694
rect 70130 430632 80078 430638
rect 70000 430570 80078 430632
rect 70000 430564 79208 430570
rect 70000 430508 70074 430564
rect 70130 430514 79208 430564
rect 79264 430514 79332 430570
rect 79388 430514 79456 430570
rect 79512 430514 79580 430570
rect 79636 430514 79704 430570
rect 79760 430514 79828 430570
rect 79884 430514 79952 430570
rect 80008 430514 80078 430570
rect 70130 430508 80078 430514
rect 70000 430446 80078 430508
rect 70000 430440 79208 430446
rect 70000 430384 70074 430440
rect 70130 430390 79208 430440
rect 79264 430390 79332 430446
rect 79388 430390 79456 430446
rect 79512 430390 79580 430446
rect 79636 430390 79704 430446
rect 79760 430390 79828 430446
rect 79884 430390 79952 430446
rect 80008 430390 80078 430446
rect 70130 430384 80078 430390
rect 70000 430322 80078 430384
rect 70000 430316 79208 430322
rect 70000 430260 70074 430316
rect 70130 430266 79208 430316
rect 79264 430266 79332 430322
rect 79388 430266 79456 430322
rect 79512 430266 79580 430322
rect 79636 430266 79704 430322
rect 79760 430266 79828 430322
rect 79884 430266 79952 430322
rect 80008 430266 80078 430322
rect 70130 430260 80078 430266
rect 70000 430198 80078 430260
rect 70000 430192 79208 430198
rect 70000 430136 70074 430192
rect 70130 430142 79208 430192
rect 79264 430142 79332 430198
rect 79388 430142 79456 430198
rect 79512 430142 79580 430198
rect 79636 430142 79704 430198
rect 79760 430142 79828 430198
rect 79884 430142 79952 430198
rect 80008 430142 80078 430198
rect 70130 430136 80078 430142
rect 70000 430074 80078 430136
rect 70000 430068 79208 430074
rect 70000 430012 70074 430068
rect 70130 430018 79208 430068
rect 79264 430018 79332 430074
rect 79388 430018 79456 430074
rect 79512 430018 79580 430074
rect 79636 430018 79704 430074
rect 79760 430018 79828 430074
rect 79884 430018 79952 430074
rect 80008 430018 80078 430074
rect 70130 430012 80078 430018
rect 70000 429950 80078 430012
rect 70000 429944 79208 429950
rect 70000 429888 70074 429944
rect 70130 429894 79208 429944
rect 79264 429894 79332 429950
rect 79388 429894 79456 429950
rect 79512 429894 79580 429950
rect 79636 429894 79704 429950
rect 79760 429894 79828 429950
rect 79884 429894 79952 429950
rect 80008 429894 80078 429950
rect 70130 429888 80078 429894
rect 70000 429826 80078 429888
rect 70000 429820 79208 429826
rect 70000 429764 70074 429820
rect 70130 429770 79208 429820
rect 79264 429770 79332 429826
rect 79388 429770 79456 429826
rect 79512 429770 79580 429826
rect 79636 429770 79704 429826
rect 79760 429770 79828 429826
rect 79884 429770 79952 429826
rect 80008 429770 80078 429826
rect 70130 429764 80078 429770
rect 70000 429702 80078 429764
rect 70000 429696 79208 429702
rect 70000 429640 70074 429696
rect 70130 429646 79208 429696
rect 79264 429646 79332 429702
rect 79388 429646 79456 429702
rect 79512 429646 79580 429702
rect 79636 429646 79704 429702
rect 79760 429646 79828 429702
rect 79884 429646 79952 429702
rect 80008 429646 80078 429702
rect 70130 429640 80078 429646
rect 70000 429578 80078 429640
rect 70000 429572 79208 429578
rect 70000 429516 70074 429572
rect 70130 429522 79208 429572
rect 79264 429522 79332 429578
rect 79388 429522 79456 429578
rect 79512 429522 79580 429578
rect 79636 429522 79704 429578
rect 79760 429522 79828 429578
rect 79884 429522 79952 429578
rect 80008 429522 80078 429578
rect 70130 429516 80078 429522
rect 70000 429454 80078 429516
rect 70000 429448 79208 429454
rect 70000 429392 70074 429448
rect 70130 429398 79208 429448
rect 79264 429398 79332 429454
rect 79388 429398 79456 429454
rect 79512 429398 79580 429454
rect 79636 429398 79704 429454
rect 79760 429398 79828 429454
rect 79884 429398 79952 429454
rect 80008 429398 80078 429454
rect 70130 429392 80078 429398
rect 70000 429330 80078 429392
rect 70000 429324 79208 429330
rect 70000 429268 70074 429324
rect 70130 429274 79208 429324
rect 79264 429274 79332 429330
rect 79388 429274 79456 429330
rect 79512 429274 79580 429330
rect 79636 429274 79704 429330
rect 79760 429274 79828 429330
rect 79884 429274 79952 429330
rect 80008 429274 80078 429330
rect 70130 429268 80078 429274
rect 70000 429198 80078 429268
rect 70000 428820 80078 428878
rect 70000 428814 79208 428820
rect 70000 428758 70074 428814
rect 70130 428764 79208 428814
rect 79264 428764 79332 428820
rect 79388 428764 79456 428820
rect 79512 428764 79580 428820
rect 79636 428764 79704 428820
rect 79760 428764 79828 428820
rect 79884 428764 79952 428820
rect 80008 428764 80078 428820
rect 70130 428758 80078 428764
rect 70000 428696 80078 428758
rect 70000 428690 79208 428696
rect 70000 428634 70074 428690
rect 70130 428640 79208 428690
rect 79264 428640 79332 428696
rect 79388 428640 79456 428696
rect 79512 428640 79580 428696
rect 79636 428640 79704 428696
rect 79760 428640 79828 428696
rect 79884 428640 79952 428696
rect 80008 428640 80078 428696
rect 70130 428634 80078 428640
rect 70000 428572 80078 428634
rect 70000 428566 79208 428572
rect 70000 428510 70074 428566
rect 70130 428516 79208 428566
rect 79264 428516 79332 428572
rect 79388 428516 79456 428572
rect 79512 428516 79580 428572
rect 79636 428516 79704 428572
rect 79760 428516 79828 428572
rect 79884 428516 79952 428572
rect 80008 428516 80078 428572
rect 70130 428510 80078 428516
rect 70000 428448 80078 428510
rect 70000 428442 79208 428448
rect 70000 428386 70074 428442
rect 70130 428392 79208 428442
rect 79264 428392 79332 428448
rect 79388 428392 79456 428448
rect 79512 428392 79580 428448
rect 79636 428392 79704 428448
rect 79760 428392 79828 428448
rect 79884 428392 79952 428448
rect 80008 428392 80078 428448
rect 70130 428386 80078 428392
rect 70000 428324 80078 428386
rect 70000 428318 79208 428324
rect 70000 428262 70074 428318
rect 70130 428268 79208 428318
rect 79264 428268 79332 428324
rect 79388 428268 79456 428324
rect 79512 428268 79580 428324
rect 79636 428268 79704 428324
rect 79760 428268 79828 428324
rect 79884 428268 79952 428324
rect 80008 428268 80078 428324
rect 70130 428262 80078 428268
rect 70000 428200 80078 428262
rect 70000 428194 79208 428200
rect 70000 428138 70074 428194
rect 70130 428144 79208 428194
rect 79264 428144 79332 428200
rect 79388 428144 79456 428200
rect 79512 428144 79580 428200
rect 79636 428144 79704 428200
rect 79760 428144 79828 428200
rect 79884 428144 79952 428200
rect 80008 428144 80078 428200
rect 70130 428138 80078 428144
rect 70000 428076 80078 428138
rect 70000 428070 79208 428076
rect 70000 428014 70074 428070
rect 70130 428020 79208 428070
rect 79264 428020 79332 428076
rect 79388 428020 79456 428076
rect 79512 428020 79580 428076
rect 79636 428020 79704 428076
rect 79760 428020 79828 428076
rect 79884 428020 79952 428076
rect 80008 428020 80078 428076
rect 70130 428014 80078 428020
rect 70000 427952 80078 428014
rect 688372 428429 698922 428630
rect 688372 428373 698144 428429
rect 698200 428373 698444 428429
rect 698500 428373 698744 428429
rect 698800 428373 698922 428429
rect 688372 428229 698922 428373
rect 688372 428173 698144 428229
rect 698200 428173 698444 428229
rect 698500 428173 698744 428229
rect 698800 428173 698922 428229
rect 688372 428010 698922 428173
rect 70000 427946 79208 427952
rect 70000 427890 70074 427946
rect 70130 427896 79208 427946
rect 79264 427896 79332 427952
rect 79388 427896 79456 427952
rect 79512 427896 79580 427952
rect 79636 427896 79704 427952
rect 79760 427896 79828 427952
rect 79884 427896 79952 427952
rect 80008 427896 80078 427952
rect 70130 427890 80078 427896
rect 70000 427828 80078 427890
rect 70000 427822 79208 427828
rect 70000 427766 70074 427822
rect 70130 427772 79208 427822
rect 79264 427772 79332 427828
rect 79388 427772 79456 427828
rect 79512 427772 79580 427828
rect 79636 427772 79704 427828
rect 79760 427772 79828 427828
rect 79884 427772 79952 427828
rect 80008 427772 80078 427828
rect 70130 427766 80078 427772
rect 70000 427704 80078 427766
rect 70000 427698 79208 427704
rect 70000 427642 70074 427698
rect 70130 427648 79208 427698
rect 79264 427648 79332 427704
rect 79388 427648 79456 427704
rect 79512 427648 79580 427704
rect 79636 427648 79704 427704
rect 79760 427648 79828 427704
rect 79884 427648 79952 427704
rect 80008 427648 80078 427704
rect 70130 427642 80078 427648
rect 70000 427580 80078 427642
rect 70000 427574 79208 427580
rect 70000 427518 70074 427574
rect 70130 427524 79208 427574
rect 79264 427524 79332 427580
rect 79388 427524 79456 427580
rect 79512 427524 79580 427580
rect 79636 427524 79704 427580
rect 79760 427524 79828 427580
rect 79884 427524 79952 427580
rect 80008 427524 80078 427580
rect 70130 427518 80078 427524
rect 70000 427456 80078 427518
rect 70000 427450 79208 427456
rect 70000 427394 70074 427450
rect 70130 427400 79208 427450
rect 79264 427400 79332 427456
rect 79388 427400 79456 427456
rect 79512 427400 79580 427456
rect 79636 427400 79704 427456
rect 79760 427400 79828 427456
rect 79884 427400 79952 427456
rect 80008 427400 80078 427456
rect 70130 427394 80078 427400
rect 70000 427332 80078 427394
rect 70000 427326 79208 427332
rect 70000 427270 70074 427326
rect 70130 427276 79208 427326
rect 79264 427276 79332 427332
rect 79388 427276 79456 427332
rect 79512 427276 79580 427332
rect 79636 427276 79704 427332
rect 79760 427276 79828 427332
rect 79884 427276 79952 427332
rect 80008 427276 80078 427332
rect 70130 427270 80078 427276
rect 70000 427208 80078 427270
rect 70000 427202 79208 427208
rect 70000 427146 70074 427202
rect 70130 427152 79208 427202
rect 79264 427152 79332 427208
rect 79388 427152 79456 427208
rect 79512 427152 79580 427208
rect 79636 427152 79704 427208
rect 79760 427152 79828 427208
rect 79884 427152 79952 427208
rect 80008 427152 80078 427208
rect 70130 427146 80078 427152
rect 70000 427084 80078 427146
rect 70000 427078 79208 427084
rect 70000 427022 70074 427078
rect 70130 427028 79208 427078
rect 79264 427028 79332 427084
rect 79388 427028 79456 427084
rect 79512 427028 79580 427084
rect 79636 427028 79704 427084
rect 79760 427028 79828 427084
rect 79884 427028 79952 427084
rect 80008 427028 80078 427084
rect 70130 427022 80078 427028
rect 70000 426960 80078 427022
rect 70000 426954 79208 426960
rect 70000 426898 70074 426954
rect 70130 426904 79208 426954
rect 79264 426904 79332 426960
rect 79388 426904 79456 426960
rect 79512 426904 79580 426960
rect 79636 426904 79704 426960
rect 79760 426904 79828 426960
rect 79884 426904 79952 426960
rect 80008 426904 80078 426960
rect 70130 426898 80078 426904
rect 70000 426828 80078 426898
rect 70000 426114 80078 426172
rect 70000 426108 79208 426114
rect 70000 426052 70074 426108
rect 70130 426058 79208 426108
rect 79264 426058 79332 426114
rect 79388 426058 79456 426114
rect 79512 426058 79580 426114
rect 79636 426058 79704 426114
rect 79760 426058 79828 426114
rect 79884 426058 79952 426114
rect 80008 426058 80078 426114
rect 70130 426052 80078 426058
rect 70000 425990 80078 426052
rect 70000 425984 79208 425990
rect 70000 425928 70074 425984
rect 70130 425934 79208 425984
rect 79264 425934 79332 425990
rect 79388 425934 79456 425990
rect 79512 425934 79580 425990
rect 79636 425934 79704 425990
rect 79760 425934 79828 425990
rect 79884 425934 79952 425990
rect 80008 425934 80078 425990
rect 70130 425928 80078 425934
rect 70000 425866 80078 425928
rect 70000 425860 79208 425866
rect 70000 425804 70074 425860
rect 70130 425810 79208 425860
rect 79264 425810 79332 425866
rect 79388 425810 79456 425866
rect 79512 425810 79580 425866
rect 79636 425810 79704 425866
rect 79760 425810 79828 425866
rect 79884 425810 79952 425866
rect 80008 425810 80078 425866
rect 70130 425804 80078 425810
rect 70000 425742 80078 425804
rect 70000 425736 79208 425742
rect 70000 425680 70074 425736
rect 70130 425686 79208 425736
rect 79264 425686 79332 425742
rect 79388 425686 79456 425742
rect 79512 425686 79580 425742
rect 79636 425686 79704 425742
rect 79760 425686 79828 425742
rect 79884 425686 79952 425742
rect 80008 425686 80078 425742
rect 70130 425680 80078 425686
rect 70000 425618 80078 425680
rect 70000 425612 79208 425618
rect 70000 425556 70074 425612
rect 70130 425562 79208 425612
rect 79264 425562 79332 425618
rect 79388 425562 79456 425618
rect 79512 425562 79580 425618
rect 79636 425562 79704 425618
rect 79760 425562 79828 425618
rect 79884 425562 79952 425618
rect 80008 425562 80078 425618
rect 70130 425556 80078 425562
rect 70000 425494 80078 425556
rect 70000 425488 79208 425494
rect 70000 425432 70074 425488
rect 70130 425438 79208 425488
rect 79264 425438 79332 425494
rect 79388 425438 79456 425494
rect 79512 425438 79580 425494
rect 79636 425438 79704 425494
rect 79760 425438 79828 425494
rect 79884 425438 79952 425494
rect 80008 425438 80078 425494
rect 70130 425432 80078 425438
rect 70000 425370 80078 425432
rect 70000 425364 79208 425370
rect 70000 425308 70074 425364
rect 70130 425314 79208 425364
rect 79264 425314 79332 425370
rect 79388 425314 79456 425370
rect 79512 425314 79580 425370
rect 79636 425314 79704 425370
rect 79760 425314 79828 425370
rect 79884 425314 79952 425370
rect 80008 425314 80078 425370
rect 70130 425308 80078 425314
rect 70000 425246 80078 425308
rect 70000 425240 79208 425246
rect 70000 425184 70074 425240
rect 70130 425190 79208 425240
rect 79264 425190 79332 425246
rect 79388 425190 79456 425246
rect 79512 425190 79580 425246
rect 79636 425190 79704 425246
rect 79760 425190 79828 425246
rect 79884 425190 79952 425246
rect 80008 425190 80078 425246
rect 70130 425184 80078 425190
rect 70000 425122 80078 425184
rect 70000 425116 79208 425122
rect 70000 425060 70074 425116
rect 70130 425066 79208 425116
rect 79264 425066 79332 425122
rect 79388 425066 79456 425122
rect 79512 425066 79580 425122
rect 79636 425066 79704 425122
rect 79760 425066 79828 425122
rect 79884 425066 79952 425122
rect 80008 425066 80078 425122
rect 70130 425060 80078 425066
rect 70000 424998 80078 425060
rect 70000 424992 79208 424998
rect 70000 424936 70074 424992
rect 70130 424942 79208 424992
rect 79264 424942 79332 424998
rect 79388 424942 79456 424998
rect 79512 424942 79580 424998
rect 79636 424942 79704 424998
rect 79760 424942 79828 424998
rect 79884 424942 79952 424998
rect 80008 424942 80078 424998
rect 70130 424936 80078 424942
rect 70000 424874 80078 424936
rect 70000 424868 79208 424874
rect 70000 424812 70074 424868
rect 70130 424818 79208 424868
rect 79264 424818 79332 424874
rect 79388 424818 79456 424874
rect 79512 424818 79580 424874
rect 79636 424818 79704 424874
rect 79760 424818 79828 424874
rect 79884 424818 79952 424874
rect 80008 424818 80078 424874
rect 70130 424812 80078 424818
rect 70000 424750 80078 424812
rect 70000 424744 79208 424750
rect 70000 424688 70074 424744
rect 70130 424694 79208 424744
rect 79264 424694 79332 424750
rect 79388 424694 79456 424750
rect 79512 424694 79580 424750
rect 79636 424694 79704 424750
rect 79760 424694 79828 424750
rect 79884 424694 79952 424750
rect 80008 424694 80078 424750
rect 70130 424688 80078 424694
rect 70000 424626 80078 424688
rect 70000 424620 79208 424626
rect 70000 424564 70074 424620
rect 70130 424570 79208 424620
rect 79264 424570 79332 424626
rect 79388 424570 79456 424626
rect 79512 424570 79580 424626
rect 79636 424570 79704 424626
rect 79760 424570 79828 424626
rect 79884 424570 79952 424626
rect 80008 424570 80078 424626
rect 70130 424564 80078 424570
rect 70000 424502 80078 424564
rect 70000 424496 79208 424502
rect 70000 424440 70074 424496
rect 70130 424446 79208 424496
rect 79264 424446 79332 424502
rect 79388 424446 79456 424502
rect 79512 424446 79580 424502
rect 79636 424446 79704 424502
rect 79760 424446 79828 424502
rect 79884 424446 79952 424502
rect 80008 424446 80078 424502
rect 70130 424440 80078 424446
rect 70000 424378 80078 424440
rect 70000 424372 79208 424378
rect 70000 424316 70074 424372
rect 70130 424322 79208 424372
rect 79264 424322 79332 424378
rect 79388 424322 79456 424378
rect 79512 424322 79580 424378
rect 79636 424322 79704 424378
rect 79760 424322 79828 424378
rect 79884 424322 79952 424378
rect 80008 424322 80078 424378
rect 70130 424316 80078 424322
rect 70000 424254 80078 424316
rect 70000 424248 79208 424254
rect 70000 424192 70074 424248
rect 70130 424198 79208 424248
rect 79264 424198 79332 424254
rect 79388 424198 79456 424254
rect 79512 424198 79580 424254
rect 79636 424198 79704 424254
rect 79760 424198 79828 424254
rect 79884 424198 79952 424254
rect 80008 424198 80078 424254
rect 70130 424192 80078 424198
rect 70000 424122 80078 424192
rect 70000 423744 80078 423802
rect 70000 423738 79208 423744
rect 70000 423682 70074 423738
rect 70130 423688 79208 423738
rect 79264 423688 79332 423744
rect 79388 423688 79456 423744
rect 79512 423688 79580 423744
rect 79636 423688 79704 423744
rect 79760 423688 79828 423744
rect 79884 423688 79952 423744
rect 80008 423688 80078 423744
rect 70130 423682 80078 423688
rect 70000 423620 80078 423682
rect 70000 423614 79208 423620
rect 70000 423558 70074 423614
rect 70130 423564 79208 423614
rect 79264 423564 79332 423620
rect 79388 423564 79456 423620
rect 79512 423564 79580 423620
rect 79636 423564 79704 423620
rect 79760 423564 79828 423620
rect 79884 423564 79952 423620
rect 80008 423564 80078 423620
rect 70130 423558 80078 423564
rect 70000 423496 80078 423558
rect 70000 423490 79208 423496
rect 70000 423434 70074 423490
rect 70130 423440 79208 423490
rect 79264 423440 79332 423496
rect 79388 423440 79456 423496
rect 79512 423440 79580 423496
rect 79636 423440 79704 423496
rect 79760 423440 79828 423496
rect 79884 423440 79952 423496
rect 80008 423440 80078 423496
rect 70130 423434 80078 423440
rect 70000 423372 80078 423434
rect 70000 423366 79208 423372
rect 70000 423310 70074 423366
rect 70130 423316 79208 423366
rect 79264 423316 79332 423372
rect 79388 423316 79456 423372
rect 79512 423316 79580 423372
rect 79636 423316 79704 423372
rect 79760 423316 79828 423372
rect 79884 423316 79952 423372
rect 80008 423316 80078 423372
rect 70130 423310 80078 423316
rect 70000 423248 80078 423310
rect 70000 423242 79208 423248
rect 70000 423186 70074 423242
rect 70130 423192 79208 423242
rect 79264 423192 79332 423248
rect 79388 423192 79456 423248
rect 79512 423192 79580 423248
rect 79636 423192 79704 423248
rect 79760 423192 79828 423248
rect 79884 423192 79952 423248
rect 80008 423192 80078 423248
rect 70130 423186 80078 423192
rect 70000 423124 80078 423186
rect 70000 423118 79208 423124
rect 70000 423062 70074 423118
rect 70130 423068 79208 423118
rect 79264 423068 79332 423124
rect 79388 423068 79456 423124
rect 79512 423068 79580 423124
rect 79636 423068 79704 423124
rect 79760 423068 79828 423124
rect 79884 423068 79952 423124
rect 80008 423068 80078 423124
rect 70130 423062 80078 423068
rect 70000 423000 80078 423062
rect 70000 422994 79208 423000
rect 70000 422938 70074 422994
rect 70130 422944 79208 422994
rect 79264 422944 79332 423000
rect 79388 422944 79456 423000
rect 79512 422944 79580 423000
rect 79636 422944 79704 423000
rect 79760 422944 79828 423000
rect 79884 422944 79952 423000
rect 80008 422944 80078 423000
rect 70130 422938 80078 422944
rect 70000 422876 80078 422938
rect 70000 422870 79208 422876
rect 70000 422814 70074 422870
rect 70130 422820 79208 422870
rect 79264 422820 79332 422876
rect 79388 422820 79456 422876
rect 79512 422820 79580 422876
rect 79636 422820 79704 422876
rect 79760 422820 79828 422876
rect 79884 422820 79952 422876
rect 80008 422820 80078 422876
rect 70130 422814 80078 422820
rect 70000 422752 80078 422814
rect 70000 422746 79208 422752
rect 70000 422690 70074 422746
rect 70130 422696 79208 422746
rect 79264 422696 79332 422752
rect 79388 422696 79456 422752
rect 79512 422696 79580 422752
rect 79636 422696 79704 422752
rect 79760 422696 79828 422752
rect 79884 422696 79952 422752
rect 80008 422696 80078 422752
rect 70130 422690 80078 422696
rect 70000 422628 80078 422690
rect 70000 422622 79208 422628
rect 70000 422566 70074 422622
rect 70130 422572 79208 422622
rect 79264 422572 79332 422628
rect 79388 422572 79456 422628
rect 79512 422572 79580 422628
rect 79636 422572 79704 422628
rect 79760 422572 79828 422628
rect 79884 422572 79952 422628
rect 80008 422572 80078 422628
rect 70130 422566 80078 422572
rect 70000 422504 80078 422566
rect 70000 422498 79208 422504
rect 70000 422442 70074 422498
rect 70130 422448 79208 422498
rect 79264 422448 79332 422504
rect 79388 422448 79456 422504
rect 79512 422448 79580 422504
rect 79636 422448 79704 422504
rect 79760 422448 79828 422504
rect 79884 422448 79952 422504
rect 80008 422448 80078 422504
rect 70130 422442 80078 422448
rect 70000 422380 80078 422442
rect 70000 422374 79208 422380
rect 70000 422318 70074 422374
rect 70130 422324 79208 422374
rect 79264 422324 79332 422380
rect 79388 422324 79456 422380
rect 79512 422324 79580 422380
rect 79636 422324 79704 422380
rect 79760 422324 79828 422380
rect 79884 422324 79952 422380
rect 80008 422324 80078 422380
rect 70130 422318 80078 422324
rect 70000 422256 80078 422318
rect 70000 422250 79208 422256
rect 70000 422194 70074 422250
rect 70130 422200 79208 422250
rect 79264 422200 79332 422256
rect 79388 422200 79456 422256
rect 79512 422200 79580 422256
rect 79636 422200 79704 422256
rect 79760 422200 79828 422256
rect 79884 422200 79952 422256
rect 80008 422200 80078 422256
rect 70130 422194 80078 422200
rect 70000 422132 80078 422194
rect 70000 422126 79208 422132
rect 70000 422070 70074 422126
rect 70130 422076 79208 422126
rect 79264 422076 79332 422132
rect 79388 422076 79456 422132
rect 79512 422076 79580 422132
rect 79636 422076 79704 422132
rect 79760 422076 79828 422132
rect 79884 422076 79952 422132
rect 80008 422076 80078 422132
rect 70130 422070 80078 422076
rect 70000 422008 80078 422070
rect 70000 422002 79208 422008
rect 70000 421946 70074 422002
rect 70130 421952 79208 422002
rect 79264 421952 79332 422008
rect 79388 421952 79456 422008
rect 79512 421952 79580 422008
rect 79636 421952 79704 422008
rect 79760 421952 79828 422008
rect 79884 421952 79952 422008
rect 80008 421952 80078 422008
rect 70130 421946 80078 421952
rect 70000 421884 80078 421946
rect 70000 421878 79208 421884
rect 70000 421822 70074 421878
rect 70130 421828 79208 421878
rect 79264 421828 79332 421884
rect 79388 421828 79456 421884
rect 79512 421828 79580 421884
rect 79636 421828 79704 421884
rect 79760 421828 79828 421884
rect 79884 421828 79952 421884
rect 80008 421828 80078 421884
rect 70130 421822 80078 421828
rect 70000 421752 80078 421822
rect 70000 421140 80078 421172
rect 70000 421134 79208 421140
rect 70000 421078 70074 421134
rect 70130 421084 79208 421134
rect 79264 421084 79332 421140
rect 79388 421084 79456 421140
rect 79512 421084 79580 421140
rect 79636 421084 79704 421140
rect 79760 421084 79828 421140
rect 79884 421084 79952 421140
rect 80008 421084 80078 421140
rect 70130 421078 80078 421084
rect 70000 421016 80078 421078
rect 70000 421010 79208 421016
rect 70000 420954 70074 421010
rect 70130 420960 79208 421010
rect 79264 420960 79332 421016
rect 79388 420960 79456 421016
rect 79512 420960 79580 421016
rect 79636 420960 79704 421016
rect 79760 420960 79828 421016
rect 79884 420960 79952 421016
rect 80008 420960 80078 421016
rect 70130 420954 80078 420960
rect 70000 420892 80078 420954
rect 70000 420886 79208 420892
rect 70000 420830 70074 420886
rect 70130 420836 79208 420886
rect 79264 420836 79332 420892
rect 79388 420836 79456 420892
rect 79512 420836 79580 420892
rect 79636 420836 79704 420892
rect 79760 420836 79828 420892
rect 79884 420836 79952 420892
rect 80008 420836 80078 420892
rect 70130 420830 80078 420836
rect 70000 420768 80078 420830
rect 70000 420762 79208 420768
rect 70000 420706 70074 420762
rect 70130 420712 79208 420762
rect 79264 420712 79332 420768
rect 79388 420712 79456 420768
rect 79512 420712 79580 420768
rect 79636 420712 79704 420768
rect 79760 420712 79828 420768
rect 79884 420712 79952 420768
rect 80008 420712 80078 420768
rect 70130 420706 80078 420712
rect 70000 420644 80078 420706
rect 70000 420638 79208 420644
rect 70000 420582 70074 420638
rect 70130 420588 79208 420638
rect 79264 420588 79332 420644
rect 79388 420588 79456 420644
rect 79512 420588 79580 420644
rect 79636 420588 79704 420644
rect 79760 420588 79828 420644
rect 79884 420588 79952 420644
rect 80008 420588 80078 420644
rect 70130 420582 80078 420588
rect 70000 420520 80078 420582
rect 70000 420514 79208 420520
rect 70000 420458 70074 420514
rect 70130 420464 79208 420514
rect 79264 420464 79332 420520
rect 79388 420464 79456 420520
rect 79512 420464 79580 420520
rect 79636 420464 79704 420520
rect 79760 420464 79828 420520
rect 79884 420464 79952 420520
rect 80008 420464 80078 420520
rect 70130 420458 80078 420464
rect 70000 420396 80078 420458
rect 70000 420390 79208 420396
rect 70000 420334 70074 420390
rect 70130 420340 79208 420390
rect 79264 420340 79332 420396
rect 79388 420340 79456 420396
rect 79512 420340 79580 420396
rect 79636 420340 79704 420396
rect 79760 420340 79828 420396
rect 79884 420340 79952 420396
rect 80008 420340 80078 420396
rect 70130 420334 80078 420340
rect 70000 420272 80078 420334
rect 70000 420266 79208 420272
rect 70000 420210 70074 420266
rect 70130 420216 79208 420266
rect 79264 420216 79332 420272
rect 79388 420216 79456 420272
rect 79512 420216 79580 420272
rect 79636 420216 79704 420272
rect 79760 420216 79828 420272
rect 79884 420216 79952 420272
rect 80008 420216 80078 420272
rect 70130 420210 80078 420216
rect 70000 420148 80078 420210
rect 70000 420142 79208 420148
rect 70000 420086 70074 420142
rect 70130 420092 79208 420142
rect 79264 420092 79332 420148
rect 79388 420092 79456 420148
rect 79512 420092 79580 420148
rect 79636 420092 79704 420148
rect 79760 420092 79828 420148
rect 79884 420092 79952 420148
rect 80008 420092 80078 420148
rect 70130 420086 80078 420092
rect 70000 420024 80078 420086
rect 70000 420018 79208 420024
rect 70000 419962 70074 420018
rect 70130 419968 79208 420018
rect 79264 419968 79332 420024
rect 79388 419968 79456 420024
rect 79512 419968 79580 420024
rect 79636 419968 79704 420024
rect 79760 419968 79828 420024
rect 79884 419968 79952 420024
rect 80008 419968 80078 420024
rect 70130 419962 80078 419968
rect 70000 419900 80078 419962
rect 70000 419894 79208 419900
rect 70000 419838 70074 419894
rect 70130 419844 79208 419894
rect 79264 419844 79332 419900
rect 79388 419844 79456 419900
rect 79512 419844 79580 419900
rect 79636 419844 79704 419900
rect 79760 419844 79828 419900
rect 79884 419844 79952 419900
rect 80008 419844 80078 419900
rect 70130 419838 80078 419844
rect 70000 419776 80078 419838
rect 70000 419770 79208 419776
rect 70000 419714 70074 419770
rect 70130 419720 79208 419770
rect 79264 419720 79332 419776
rect 79388 419720 79456 419776
rect 79512 419720 79580 419776
rect 79636 419720 79704 419776
rect 79760 419720 79828 419776
rect 79884 419720 79952 419776
rect 80008 419720 80078 419776
rect 70130 419714 80078 419720
rect 70000 419652 80078 419714
rect 70000 419646 79208 419652
rect 70000 419590 70074 419646
rect 70130 419596 79208 419646
rect 79264 419596 79332 419652
rect 79388 419596 79456 419652
rect 79512 419596 79580 419652
rect 79636 419596 79704 419652
rect 79760 419596 79828 419652
rect 79884 419596 79952 419652
rect 80008 419596 80078 419652
rect 70130 419590 80078 419596
rect 70000 419528 80078 419590
rect 70000 419522 79208 419528
rect 70000 419466 70074 419522
rect 70130 419472 79208 419522
rect 79264 419472 79332 419528
rect 79388 419472 79456 419528
rect 79512 419472 79580 419528
rect 79636 419472 79704 419528
rect 79760 419472 79828 419528
rect 79884 419472 79952 419528
rect 80008 419472 80078 419528
rect 70130 419466 80078 419472
rect 70000 419404 80078 419466
rect 70000 419398 79208 419404
rect 70000 419342 70074 419398
rect 70130 419348 79208 419398
rect 79264 419348 79332 419404
rect 79388 419348 79456 419404
rect 79512 419348 79580 419404
rect 79636 419348 79704 419404
rect 79760 419348 79828 419404
rect 79884 419348 79952 419404
rect 80008 419348 80078 419404
rect 70130 419342 80078 419348
rect 70000 419272 80078 419342
rect 76115 413048 80078 413110
rect 76115 412992 79284 413048
rect 79340 412992 79584 413048
rect 79640 412992 79884 413048
rect 79940 412992 80078 413048
rect 76115 412910 80078 412992
rect 76115 412510 76435 412910
rect 76915 412633 78678 412710
rect 76915 412577 77847 412633
rect 77903 412577 78147 412633
rect 78203 412577 78447 412633
rect 78503 412577 78678 412633
rect 76915 412510 78678 412577
rect 697922 410658 708000 410728
rect 697922 410652 707870 410658
rect 77678 410429 84516 410630
rect 77678 410373 77800 410429
rect 77856 410373 78100 410429
rect 78156 410373 78400 410429
rect 78456 410373 84516 410429
rect 77678 410229 84516 410373
rect 77678 410173 77800 410229
rect 77856 410173 78100 410229
rect 78156 410173 78400 410229
rect 78456 410173 84516 410229
rect 77678 410010 84516 410173
rect 697922 410596 697992 410652
rect 698048 410596 698116 410652
rect 698172 410596 698240 410652
rect 698296 410596 698364 410652
rect 698420 410596 698488 410652
rect 698544 410596 698612 410652
rect 698668 410596 698736 410652
rect 698792 410602 707870 410652
rect 707926 410602 708000 410658
rect 698792 410596 708000 410602
rect 697922 410534 708000 410596
rect 697922 410528 707870 410534
rect 697922 410472 697992 410528
rect 698048 410472 698116 410528
rect 698172 410472 698240 410528
rect 698296 410472 698364 410528
rect 698420 410472 698488 410528
rect 698544 410472 698612 410528
rect 698668 410472 698736 410528
rect 698792 410478 707870 410528
rect 707926 410478 708000 410534
rect 698792 410472 708000 410478
rect 697922 410410 708000 410472
rect 697922 410404 707870 410410
rect 697922 410348 697992 410404
rect 698048 410348 698116 410404
rect 698172 410348 698240 410404
rect 698296 410348 698364 410404
rect 698420 410348 698488 410404
rect 698544 410348 698612 410404
rect 698668 410348 698736 410404
rect 698792 410354 707870 410404
rect 707926 410354 708000 410410
rect 698792 410348 708000 410354
rect 697922 410286 708000 410348
rect 697922 410280 707870 410286
rect 697922 410224 697992 410280
rect 698048 410224 698116 410280
rect 698172 410224 698240 410280
rect 698296 410224 698364 410280
rect 698420 410224 698488 410280
rect 698544 410224 698612 410280
rect 698668 410224 698736 410280
rect 698792 410230 707870 410280
rect 707926 410230 708000 410286
rect 698792 410224 708000 410230
rect 697922 410162 708000 410224
rect 697922 410156 707870 410162
rect 697922 410100 697992 410156
rect 698048 410100 698116 410156
rect 698172 410100 698240 410156
rect 698296 410100 698364 410156
rect 698420 410100 698488 410156
rect 698544 410100 698612 410156
rect 698668 410100 698736 410156
rect 698792 410106 707870 410156
rect 707926 410106 708000 410162
rect 698792 410100 708000 410106
rect 697922 410038 708000 410100
rect 697922 410032 707870 410038
rect 697922 409976 697992 410032
rect 698048 409976 698116 410032
rect 698172 409976 698240 410032
rect 698296 409976 698364 410032
rect 698420 409976 698488 410032
rect 698544 409976 698612 410032
rect 698668 409976 698736 410032
rect 698792 409982 707870 410032
rect 707926 409982 708000 410038
rect 698792 409976 708000 409982
rect 697922 409914 708000 409976
rect 697922 409908 707870 409914
rect 697922 409852 697992 409908
rect 698048 409852 698116 409908
rect 698172 409852 698240 409908
rect 698296 409852 698364 409908
rect 698420 409852 698488 409908
rect 698544 409852 698612 409908
rect 698668 409852 698736 409908
rect 698792 409858 707870 409908
rect 707926 409858 708000 409914
rect 698792 409852 708000 409858
rect 697922 409790 708000 409852
rect 697922 409784 707870 409790
rect 697922 409728 697992 409784
rect 698048 409728 698116 409784
rect 698172 409728 698240 409784
rect 698296 409728 698364 409784
rect 698420 409728 698488 409784
rect 698544 409728 698612 409784
rect 698668 409728 698736 409784
rect 698792 409734 707870 409784
rect 707926 409734 708000 409790
rect 698792 409728 708000 409734
rect 697922 409666 708000 409728
rect 697922 409660 707870 409666
rect 697922 409604 697992 409660
rect 698048 409604 698116 409660
rect 698172 409604 698240 409660
rect 698296 409604 698364 409660
rect 698420 409604 698488 409660
rect 698544 409604 698612 409660
rect 698668 409604 698736 409660
rect 698792 409610 707870 409660
rect 707926 409610 708000 409666
rect 698792 409604 708000 409610
rect 697922 409542 708000 409604
rect 697922 409536 707870 409542
rect 697922 409480 697992 409536
rect 698048 409480 698116 409536
rect 698172 409480 698240 409536
rect 698296 409480 698364 409536
rect 698420 409480 698488 409536
rect 698544 409480 698612 409536
rect 698668 409480 698736 409536
rect 698792 409486 707870 409536
rect 707926 409486 708000 409542
rect 698792 409480 708000 409486
rect 697922 409418 708000 409480
rect 697922 409412 707870 409418
rect 697922 409356 697992 409412
rect 698048 409356 698116 409412
rect 698172 409356 698240 409412
rect 698296 409356 698364 409412
rect 698420 409356 698488 409412
rect 698544 409356 698612 409412
rect 698668 409356 698736 409412
rect 698792 409362 707870 409412
rect 707926 409362 708000 409418
rect 698792 409356 708000 409362
rect 697922 409294 708000 409356
rect 697922 409288 707870 409294
rect 697922 409232 697992 409288
rect 698048 409232 698116 409288
rect 698172 409232 698240 409288
rect 698296 409232 698364 409288
rect 698420 409232 698488 409288
rect 698544 409232 698612 409288
rect 698668 409232 698736 409288
rect 698792 409238 707870 409288
rect 707926 409238 708000 409294
rect 698792 409232 708000 409238
rect 697922 409170 708000 409232
rect 697922 409164 707870 409170
rect 697922 409108 697992 409164
rect 698048 409108 698116 409164
rect 698172 409108 698240 409164
rect 698296 409108 698364 409164
rect 698420 409108 698488 409164
rect 698544 409108 698612 409164
rect 698668 409108 698736 409164
rect 698792 409114 707870 409164
rect 707926 409114 708000 409170
rect 698792 409108 708000 409114
rect 697922 409046 708000 409108
rect 697922 409040 707870 409046
rect 697922 408984 697992 409040
rect 698048 408984 698116 409040
rect 698172 408984 698240 409040
rect 698296 408984 698364 409040
rect 698420 408984 698488 409040
rect 698544 408984 698612 409040
rect 698668 408984 698736 409040
rect 698792 408990 707870 409040
rect 707926 408990 708000 409046
rect 698792 408984 708000 408990
rect 697922 408922 708000 408984
rect 697922 408916 707870 408922
rect 697922 408860 697992 408916
rect 698048 408860 698116 408916
rect 698172 408860 698240 408916
rect 698296 408860 698364 408916
rect 698420 408860 698488 408916
rect 698544 408860 698612 408916
rect 698668 408860 698736 408916
rect 698792 408866 707870 408916
rect 707926 408866 708000 408922
rect 698792 408860 708000 408866
rect 697922 408828 708000 408860
rect 697922 408178 708000 408248
rect 697922 408172 707870 408178
rect 697922 408116 697992 408172
rect 698048 408116 698116 408172
rect 698172 408116 698240 408172
rect 698296 408116 698364 408172
rect 698420 408116 698488 408172
rect 698544 408116 698612 408172
rect 698668 408116 698736 408172
rect 698792 408122 707870 408172
rect 707926 408122 708000 408178
rect 698792 408116 708000 408122
rect 697922 408054 708000 408116
rect 697922 408048 707870 408054
rect 697922 407992 697992 408048
rect 698048 407992 698116 408048
rect 698172 407992 698240 408048
rect 698296 407992 698364 408048
rect 698420 407992 698488 408048
rect 698544 407992 698612 408048
rect 698668 407992 698736 408048
rect 698792 407998 707870 408048
rect 707926 407998 708000 408054
rect 698792 407992 708000 407998
rect 697922 407930 708000 407992
rect 697922 407924 707870 407930
rect 697922 407868 697992 407924
rect 698048 407868 698116 407924
rect 698172 407868 698240 407924
rect 698296 407868 698364 407924
rect 698420 407868 698488 407924
rect 698544 407868 698612 407924
rect 698668 407868 698736 407924
rect 698792 407874 707870 407924
rect 707926 407874 708000 407930
rect 698792 407868 708000 407874
rect 697922 407806 708000 407868
rect 697922 407800 707870 407806
rect 697922 407744 697992 407800
rect 698048 407744 698116 407800
rect 698172 407744 698240 407800
rect 698296 407744 698364 407800
rect 698420 407744 698488 407800
rect 698544 407744 698612 407800
rect 698668 407744 698736 407800
rect 698792 407750 707870 407800
rect 707926 407750 708000 407806
rect 698792 407744 708000 407750
rect 697922 407682 708000 407744
rect 697922 407676 707870 407682
rect 697922 407620 697992 407676
rect 698048 407620 698116 407676
rect 698172 407620 698240 407676
rect 698296 407620 698364 407676
rect 698420 407620 698488 407676
rect 698544 407620 698612 407676
rect 698668 407620 698736 407676
rect 698792 407626 707870 407676
rect 707926 407626 708000 407682
rect 698792 407620 708000 407626
rect 697922 407558 708000 407620
rect 697922 407552 707870 407558
rect 697922 407496 697992 407552
rect 698048 407496 698116 407552
rect 698172 407496 698240 407552
rect 698296 407496 698364 407552
rect 698420 407496 698488 407552
rect 698544 407496 698612 407552
rect 698668 407496 698736 407552
rect 698792 407502 707870 407552
rect 707926 407502 708000 407558
rect 698792 407496 708000 407502
rect 697922 407434 708000 407496
rect 697922 407428 707870 407434
rect 697922 407372 697992 407428
rect 698048 407372 698116 407428
rect 698172 407372 698240 407428
rect 698296 407372 698364 407428
rect 698420 407372 698488 407428
rect 698544 407372 698612 407428
rect 698668 407372 698736 407428
rect 698792 407378 707870 407428
rect 707926 407378 708000 407434
rect 698792 407372 708000 407378
rect 697922 407310 708000 407372
rect 697922 407304 707870 407310
rect 697922 407248 697992 407304
rect 698048 407248 698116 407304
rect 698172 407248 698240 407304
rect 698296 407248 698364 407304
rect 698420 407248 698488 407304
rect 698544 407248 698612 407304
rect 698668 407248 698736 407304
rect 698792 407254 707870 407304
rect 707926 407254 708000 407310
rect 698792 407248 708000 407254
rect 697922 407186 708000 407248
rect 697922 407180 707870 407186
rect 697922 407124 697992 407180
rect 698048 407124 698116 407180
rect 698172 407124 698240 407180
rect 698296 407124 698364 407180
rect 698420 407124 698488 407180
rect 698544 407124 698612 407180
rect 698668 407124 698736 407180
rect 698792 407130 707870 407180
rect 707926 407130 708000 407186
rect 698792 407124 708000 407130
rect 697922 407062 708000 407124
rect 697922 407056 707870 407062
rect 697922 407000 697992 407056
rect 698048 407000 698116 407056
rect 698172 407000 698240 407056
rect 698296 407000 698364 407056
rect 698420 407000 698488 407056
rect 698544 407000 698612 407056
rect 698668 407000 698736 407056
rect 698792 407006 707870 407056
rect 707926 407006 708000 407062
rect 698792 407000 708000 407006
rect 697922 406938 708000 407000
rect 697922 406932 707870 406938
rect 697922 406876 697992 406932
rect 698048 406876 698116 406932
rect 698172 406876 698240 406932
rect 698296 406876 698364 406932
rect 698420 406876 698488 406932
rect 698544 406876 698612 406932
rect 698668 406876 698736 406932
rect 698792 406882 707870 406932
rect 707926 406882 708000 406938
rect 698792 406876 708000 406882
rect 697922 406814 708000 406876
rect 697922 406808 707870 406814
rect 697922 406752 697992 406808
rect 698048 406752 698116 406808
rect 698172 406752 698240 406808
rect 698296 406752 698364 406808
rect 698420 406752 698488 406808
rect 698544 406752 698612 406808
rect 698668 406752 698736 406808
rect 698792 406758 707870 406808
rect 707926 406758 708000 406814
rect 698792 406752 708000 406758
rect 697922 406690 708000 406752
rect 697922 406684 707870 406690
rect 697922 406628 697992 406684
rect 698048 406628 698116 406684
rect 698172 406628 698240 406684
rect 698296 406628 698364 406684
rect 698420 406628 698488 406684
rect 698544 406628 698612 406684
rect 698668 406628 698736 406684
rect 698792 406634 707870 406684
rect 707926 406634 708000 406690
rect 698792 406628 708000 406634
rect 697922 406566 708000 406628
rect 697922 406560 707870 406566
rect 697922 406504 697992 406560
rect 698048 406504 698116 406560
rect 698172 406504 698240 406560
rect 698296 406504 698364 406560
rect 698420 406504 698488 406560
rect 698544 406504 698612 406560
rect 698668 406504 698736 406560
rect 698792 406510 707870 406560
rect 707926 406510 708000 406566
rect 698792 406504 708000 406510
rect 697922 406442 708000 406504
rect 697922 406436 707870 406442
rect 697922 406380 697992 406436
rect 698048 406380 698116 406436
rect 698172 406380 698240 406436
rect 698296 406380 698364 406436
rect 698420 406380 698488 406436
rect 698544 406380 698612 406436
rect 698668 406380 698736 406436
rect 698792 406386 707870 406436
rect 707926 406386 708000 406442
rect 698792 406380 708000 406386
rect 697922 406318 708000 406380
rect 697922 406312 707870 406318
rect 697922 406256 697992 406312
rect 698048 406256 698116 406312
rect 698172 406256 698240 406312
rect 698296 406256 698364 406312
rect 698420 406256 698488 406312
rect 698544 406256 698612 406312
rect 698668 406256 698736 406312
rect 698792 406262 707870 406312
rect 707926 406262 708000 406318
rect 698792 406256 708000 406262
rect 697922 406198 708000 406256
rect 697922 405808 708000 405878
rect 697922 405802 707870 405808
rect 697922 405746 697992 405802
rect 698048 405746 698116 405802
rect 698172 405746 698240 405802
rect 698296 405746 698364 405802
rect 698420 405746 698488 405802
rect 698544 405746 698612 405802
rect 698668 405746 698736 405802
rect 698792 405752 707870 405802
rect 707926 405752 708000 405808
rect 698792 405746 708000 405752
rect 697922 405684 708000 405746
rect 697922 405678 707870 405684
rect 697922 405622 697992 405678
rect 698048 405622 698116 405678
rect 698172 405622 698240 405678
rect 698296 405622 698364 405678
rect 698420 405622 698488 405678
rect 698544 405622 698612 405678
rect 698668 405622 698736 405678
rect 698792 405628 707870 405678
rect 707926 405628 708000 405684
rect 698792 405622 708000 405628
rect 697922 405560 708000 405622
rect 697922 405554 707870 405560
rect 697922 405498 697992 405554
rect 698048 405498 698116 405554
rect 698172 405498 698240 405554
rect 698296 405498 698364 405554
rect 698420 405498 698488 405554
rect 698544 405498 698612 405554
rect 698668 405498 698736 405554
rect 698792 405504 707870 405554
rect 707926 405504 708000 405560
rect 698792 405498 708000 405504
rect 697922 405436 708000 405498
rect 697922 405430 707870 405436
rect 697922 405374 697992 405430
rect 698048 405374 698116 405430
rect 698172 405374 698240 405430
rect 698296 405374 698364 405430
rect 698420 405374 698488 405430
rect 698544 405374 698612 405430
rect 698668 405374 698736 405430
rect 698792 405380 707870 405430
rect 707926 405380 708000 405436
rect 698792 405374 708000 405380
rect 697922 405312 708000 405374
rect 697922 405306 707870 405312
rect 697922 405250 697992 405306
rect 698048 405250 698116 405306
rect 698172 405250 698240 405306
rect 698296 405250 698364 405306
rect 698420 405250 698488 405306
rect 698544 405250 698612 405306
rect 698668 405250 698736 405306
rect 698792 405256 707870 405306
rect 707926 405256 708000 405312
rect 698792 405250 708000 405256
rect 697922 405188 708000 405250
rect 697922 405182 707870 405188
rect 697922 405126 697992 405182
rect 698048 405126 698116 405182
rect 698172 405126 698240 405182
rect 698296 405126 698364 405182
rect 698420 405126 698488 405182
rect 698544 405126 698612 405182
rect 698668 405126 698736 405182
rect 698792 405132 707870 405182
rect 707926 405132 708000 405188
rect 698792 405126 708000 405132
rect 697922 405064 708000 405126
rect 697922 405058 707870 405064
rect 697922 405002 697992 405058
rect 698048 405002 698116 405058
rect 698172 405002 698240 405058
rect 698296 405002 698364 405058
rect 698420 405002 698488 405058
rect 698544 405002 698612 405058
rect 698668 405002 698736 405058
rect 698792 405008 707870 405058
rect 707926 405008 708000 405064
rect 698792 405002 708000 405008
rect 697922 404940 708000 405002
rect 697922 404934 707870 404940
rect 697922 404878 697992 404934
rect 698048 404878 698116 404934
rect 698172 404878 698240 404934
rect 698296 404878 698364 404934
rect 698420 404878 698488 404934
rect 698544 404878 698612 404934
rect 698668 404878 698736 404934
rect 698792 404884 707870 404934
rect 707926 404884 708000 404940
rect 698792 404878 708000 404884
rect 697922 404816 708000 404878
rect 697922 404810 707870 404816
rect 697922 404754 697992 404810
rect 698048 404754 698116 404810
rect 698172 404754 698240 404810
rect 698296 404754 698364 404810
rect 698420 404754 698488 404810
rect 698544 404754 698612 404810
rect 698668 404754 698736 404810
rect 698792 404760 707870 404810
rect 707926 404760 708000 404816
rect 698792 404754 708000 404760
rect 697922 404692 708000 404754
rect 697922 404686 707870 404692
rect 697922 404630 697992 404686
rect 698048 404630 698116 404686
rect 698172 404630 698240 404686
rect 698296 404630 698364 404686
rect 698420 404630 698488 404686
rect 698544 404630 698612 404686
rect 698668 404630 698736 404686
rect 698792 404636 707870 404686
rect 707926 404636 708000 404692
rect 698792 404630 708000 404636
rect 697922 404568 708000 404630
rect 697922 404562 707870 404568
rect 697922 404506 697992 404562
rect 698048 404506 698116 404562
rect 698172 404506 698240 404562
rect 698296 404506 698364 404562
rect 698420 404506 698488 404562
rect 698544 404506 698612 404562
rect 698668 404506 698736 404562
rect 698792 404512 707870 404562
rect 707926 404512 708000 404568
rect 698792 404506 708000 404512
rect 697922 404444 708000 404506
rect 697922 404438 707870 404444
rect 697922 404382 697992 404438
rect 698048 404382 698116 404438
rect 698172 404382 698240 404438
rect 698296 404382 698364 404438
rect 698420 404382 698488 404438
rect 698544 404382 698612 404438
rect 698668 404382 698736 404438
rect 698792 404388 707870 404438
rect 707926 404388 708000 404444
rect 698792 404382 708000 404388
rect 697922 404320 708000 404382
rect 697922 404314 707870 404320
rect 697922 404258 697992 404314
rect 698048 404258 698116 404314
rect 698172 404258 698240 404314
rect 698296 404258 698364 404314
rect 698420 404258 698488 404314
rect 698544 404258 698612 404314
rect 698668 404258 698736 404314
rect 698792 404264 707870 404314
rect 707926 404264 708000 404320
rect 698792 404258 708000 404264
rect 697922 404196 708000 404258
rect 697922 404190 707870 404196
rect 697922 404134 697992 404190
rect 698048 404134 698116 404190
rect 698172 404134 698240 404190
rect 698296 404134 698364 404190
rect 698420 404134 698488 404190
rect 698544 404134 698612 404190
rect 698668 404134 698736 404190
rect 698792 404140 707870 404190
rect 707926 404140 708000 404196
rect 698792 404134 708000 404140
rect 697922 404072 708000 404134
rect 697922 404066 707870 404072
rect 697922 404010 697992 404066
rect 698048 404010 698116 404066
rect 698172 404010 698240 404066
rect 698296 404010 698364 404066
rect 698420 404010 698488 404066
rect 698544 404010 698612 404066
rect 698668 404010 698736 404066
rect 698792 404016 707870 404066
rect 707926 404016 708000 404072
rect 698792 404010 708000 404016
rect 697922 403948 708000 404010
rect 697922 403942 707870 403948
rect 697922 403886 697992 403942
rect 698048 403886 698116 403942
rect 698172 403886 698240 403942
rect 698296 403886 698364 403942
rect 698420 403886 698488 403942
rect 698544 403886 698612 403942
rect 698668 403886 698736 403942
rect 698792 403892 707870 403942
rect 707926 403892 708000 403948
rect 698792 403886 708000 403892
rect 697922 403828 708000 403886
rect 697922 403102 708000 403172
rect 697922 403096 707870 403102
rect 697922 403040 697992 403096
rect 698048 403040 698116 403096
rect 698172 403040 698240 403096
rect 698296 403040 698364 403096
rect 698420 403040 698488 403096
rect 698544 403040 698612 403096
rect 698668 403040 698736 403096
rect 698792 403046 707870 403096
rect 707926 403046 708000 403102
rect 698792 403040 708000 403046
rect 697922 402978 708000 403040
rect 697922 402972 707870 402978
rect 697922 402916 697992 402972
rect 698048 402916 698116 402972
rect 698172 402916 698240 402972
rect 698296 402916 698364 402972
rect 698420 402916 698488 402972
rect 698544 402916 698612 402972
rect 698668 402916 698736 402972
rect 698792 402922 707870 402972
rect 707926 402922 708000 402978
rect 698792 402916 708000 402922
rect 697922 402854 708000 402916
rect 697922 402848 707870 402854
rect 697922 402792 697992 402848
rect 698048 402792 698116 402848
rect 698172 402792 698240 402848
rect 698296 402792 698364 402848
rect 698420 402792 698488 402848
rect 698544 402792 698612 402848
rect 698668 402792 698736 402848
rect 698792 402798 707870 402848
rect 707926 402798 708000 402854
rect 698792 402792 708000 402798
rect 697922 402730 708000 402792
rect 697922 402724 707870 402730
rect 697922 402668 697992 402724
rect 698048 402668 698116 402724
rect 698172 402668 698240 402724
rect 698296 402668 698364 402724
rect 698420 402668 698488 402724
rect 698544 402668 698612 402724
rect 698668 402668 698736 402724
rect 698792 402674 707870 402724
rect 707926 402674 708000 402730
rect 698792 402668 708000 402674
rect 697922 402606 708000 402668
rect 697922 402600 707870 402606
rect 697922 402544 697992 402600
rect 698048 402544 698116 402600
rect 698172 402544 698240 402600
rect 698296 402544 698364 402600
rect 698420 402544 698488 402600
rect 698544 402544 698612 402600
rect 698668 402544 698736 402600
rect 698792 402550 707870 402600
rect 707926 402550 708000 402606
rect 698792 402544 708000 402550
rect 697922 402482 708000 402544
rect 697922 402476 707870 402482
rect 697922 402420 697992 402476
rect 698048 402420 698116 402476
rect 698172 402420 698240 402476
rect 698296 402420 698364 402476
rect 698420 402420 698488 402476
rect 698544 402420 698612 402476
rect 698668 402420 698736 402476
rect 698792 402426 707870 402476
rect 707926 402426 708000 402482
rect 698792 402420 708000 402426
rect 697922 402358 708000 402420
rect 697922 402352 707870 402358
rect 697922 402296 697992 402352
rect 698048 402296 698116 402352
rect 698172 402296 698240 402352
rect 698296 402296 698364 402352
rect 698420 402296 698488 402352
rect 698544 402296 698612 402352
rect 698668 402296 698736 402352
rect 698792 402302 707870 402352
rect 707926 402302 708000 402358
rect 698792 402296 708000 402302
rect 697922 402234 708000 402296
rect 697922 402228 707870 402234
rect 697922 402172 697992 402228
rect 698048 402172 698116 402228
rect 698172 402172 698240 402228
rect 698296 402172 698364 402228
rect 698420 402172 698488 402228
rect 698544 402172 698612 402228
rect 698668 402172 698736 402228
rect 698792 402178 707870 402228
rect 707926 402178 708000 402234
rect 698792 402172 708000 402178
rect 697922 402110 708000 402172
rect 697922 402104 707870 402110
rect 697922 402048 697992 402104
rect 698048 402048 698116 402104
rect 698172 402048 698240 402104
rect 698296 402048 698364 402104
rect 698420 402048 698488 402104
rect 698544 402048 698612 402104
rect 698668 402048 698736 402104
rect 698792 402054 707870 402104
rect 707926 402054 708000 402110
rect 698792 402048 708000 402054
rect 697922 401986 708000 402048
rect 697922 401980 707870 401986
rect 697922 401924 697992 401980
rect 698048 401924 698116 401980
rect 698172 401924 698240 401980
rect 698296 401924 698364 401980
rect 698420 401924 698488 401980
rect 698544 401924 698612 401980
rect 698668 401924 698736 401980
rect 698792 401930 707870 401980
rect 707926 401930 708000 401986
rect 698792 401924 708000 401930
rect 697922 401862 708000 401924
rect 697922 401856 707870 401862
rect 697922 401800 697992 401856
rect 698048 401800 698116 401856
rect 698172 401800 698240 401856
rect 698296 401800 698364 401856
rect 698420 401800 698488 401856
rect 698544 401800 698612 401856
rect 698668 401800 698736 401856
rect 698792 401806 707870 401856
rect 707926 401806 708000 401862
rect 698792 401800 708000 401806
rect 697922 401738 708000 401800
rect 697922 401732 707870 401738
rect 697922 401676 697992 401732
rect 698048 401676 698116 401732
rect 698172 401676 698240 401732
rect 698296 401676 698364 401732
rect 698420 401676 698488 401732
rect 698544 401676 698612 401732
rect 698668 401676 698736 401732
rect 698792 401682 707870 401732
rect 707926 401682 708000 401738
rect 698792 401676 708000 401682
rect 697922 401614 708000 401676
rect 697922 401608 707870 401614
rect 697922 401552 697992 401608
rect 698048 401552 698116 401608
rect 698172 401552 698240 401608
rect 698296 401552 698364 401608
rect 698420 401552 698488 401608
rect 698544 401552 698612 401608
rect 698668 401552 698736 401608
rect 698792 401558 707870 401608
rect 707926 401558 708000 401614
rect 698792 401552 708000 401558
rect 697922 401490 708000 401552
rect 697922 401484 707870 401490
rect 697922 401428 697992 401484
rect 698048 401428 698116 401484
rect 698172 401428 698240 401484
rect 698296 401428 698364 401484
rect 698420 401428 698488 401484
rect 698544 401428 698612 401484
rect 698668 401428 698736 401484
rect 698792 401434 707870 401484
rect 707926 401434 708000 401490
rect 698792 401428 708000 401434
rect 697922 401366 708000 401428
rect 697922 401360 707870 401366
rect 697922 401304 697992 401360
rect 698048 401304 698116 401360
rect 698172 401304 698240 401360
rect 698296 401304 698364 401360
rect 698420 401304 698488 401360
rect 698544 401304 698612 401360
rect 698668 401304 698736 401360
rect 698792 401310 707870 401360
rect 707926 401310 708000 401366
rect 698792 401304 708000 401310
rect 697922 401242 708000 401304
rect 697922 401236 707870 401242
rect 697922 401180 697992 401236
rect 698048 401180 698116 401236
rect 698172 401180 698240 401236
rect 698296 401180 698364 401236
rect 698420 401180 698488 401236
rect 698544 401180 698612 401236
rect 698668 401180 698736 401236
rect 698792 401186 707870 401236
rect 707926 401186 708000 401242
rect 698792 401180 708000 401186
rect 697922 401122 708000 401180
rect 697922 400732 708000 400802
rect 697922 400726 707870 400732
rect 697922 400670 697992 400726
rect 698048 400670 698116 400726
rect 698172 400670 698240 400726
rect 698296 400670 698364 400726
rect 698420 400670 698488 400726
rect 698544 400670 698612 400726
rect 698668 400670 698736 400726
rect 698792 400676 707870 400726
rect 707926 400676 708000 400732
rect 698792 400670 708000 400676
rect 697922 400608 708000 400670
rect 697922 400602 707870 400608
rect 697922 400546 697992 400602
rect 698048 400546 698116 400602
rect 698172 400546 698240 400602
rect 698296 400546 698364 400602
rect 698420 400546 698488 400602
rect 698544 400546 698612 400602
rect 698668 400546 698736 400602
rect 698792 400552 707870 400602
rect 707926 400552 708000 400608
rect 698792 400546 708000 400552
rect 697922 400484 708000 400546
rect 697922 400478 707870 400484
rect 697922 400422 697992 400478
rect 698048 400422 698116 400478
rect 698172 400422 698240 400478
rect 698296 400422 698364 400478
rect 698420 400422 698488 400478
rect 698544 400422 698612 400478
rect 698668 400422 698736 400478
rect 698792 400428 707870 400478
rect 707926 400428 708000 400484
rect 698792 400422 708000 400428
rect 697922 400360 708000 400422
rect 697922 400354 707870 400360
rect 697922 400298 697992 400354
rect 698048 400298 698116 400354
rect 698172 400298 698240 400354
rect 698296 400298 698364 400354
rect 698420 400298 698488 400354
rect 698544 400298 698612 400354
rect 698668 400298 698736 400354
rect 698792 400304 707870 400354
rect 707926 400304 708000 400360
rect 698792 400298 708000 400304
rect 697922 400236 708000 400298
rect 697922 400230 707870 400236
rect 697922 400174 697992 400230
rect 698048 400174 698116 400230
rect 698172 400174 698240 400230
rect 698296 400174 698364 400230
rect 698420 400174 698488 400230
rect 698544 400174 698612 400230
rect 698668 400174 698736 400230
rect 698792 400180 707870 400230
rect 707926 400180 708000 400236
rect 698792 400174 708000 400180
rect 697922 400112 708000 400174
rect 697922 400106 707870 400112
rect 697922 400050 697992 400106
rect 698048 400050 698116 400106
rect 698172 400050 698240 400106
rect 698296 400050 698364 400106
rect 698420 400050 698488 400106
rect 698544 400050 698612 400106
rect 698668 400050 698736 400106
rect 698792 400056 707870 400106
rect 707926 400056 708000 400112
rect 698792 400050 708000 400056
rect 697922 399988 708000 400050
rect 697922 399982 707870 399988
rect 697922 399926 697992 399982
rect 698048 399926 698116 399982
rect 698172 399926 698240 399982
rect 698296 399926 698364 399982
rect 698420 399926 698488 399982
rect 698544 399926 698612 399982
rect 698668 399926 698736 399982
rect 698792 399932 707870 399982
rect 707926 399932 708000 399988
rect 698792 399926 708000 399932
rect 697922 399864 708000 399926
rect 697922 399858 707870 399864
rect 697922 399802 697992 399858
rect 698048 399802 698116 399858
rect 698172 399802 698240 399858
rect 698296 399802 698364 399858
rect 698420 399802 698488 399858
rect 698544 399802 698612 399858
rect 698668 399802 698736 399858
rect 698792 399808 707870 399858
rect 707926 399808 708000 399864
rect 698792 399802 708000 399808
rect 697922 399740 708000 399802
rect 697922 399734 707870 399740
rect 697922 399678 697992 399734
rect 698048 399678 698116 399734
rect 698172 399678 698240 399734
rect 698296 399678 698364 399734
rect 698420 399678 698488 399734
rect 698544 399678 698612 399734
rect 698668 399678 698736 399734
rect 698792 399684 707870 399734
rect 707926 399684 708000 399740
rect 698792 399678 708000 399684
rect 697922 399616 708000 399678
rect 697922 399610 707870 399616
rect 697922 399554 697992 399610
rect 698048 399554 698116 399610
rect 698172 399554 698240 399610
rect 698296 399554 698364 399610
rect 698420 399554 698488 399610
rect 698544 399554 698612 399610
rect 698668 399554 698736 399610
rect 698792 399560 707870 399610
rect 707926 399560 708000 399616
rect 698792 399554 708000 399560
rect 697922 399492 708000 399554
rect 697922 399486 707870 399492
rect 697922 399430 697992 399486
rect 698048 399430 698116 399486
rect 698172 399430 698240 399486
rect 698296 399430 698364 399486
rect 698420 399430 698488 399486
rect 698544 399430 698612 399486
rect 698668 399430 698736 399486
rect 698792 399436 707870 399486
rect 707926 399436 708000 399492
rect 698792 399430 708000 399436
rect 697922 399368 708000 399430
rect 697922 399362 707870 399368
rect 697922 399306 697992 399362
rect 698048 399306 698116 399362
rect 698172 399306 698240 399362
rect 698296 399306 698364 399362
rect 698420 399306 698488 399362
rect 698544 399306 698612 399362
rect 698668 399306 698736 399362
rect 698792 399312 707870 399362
rect 707926 399312 708000 399368
rect 698792 399306 708000 399312
rect 697922 399244 708000 399306
rect 697922 399238 707870 399244
rect 697922 399182 697992 399238
rect 698048 399182 698116 399238
rect 698172 399182 698240 399238
rect 698296 399182 698364 399238
rect 698420 399182 698488 399238
rect 698544 399182 698612 399238
rect 698668 399182 698736 399238
rect 698792 399188 707870 399238
rect 707926 399188 708000 399244
rect 698792 399182 708000 399188
rect 697922 399120 708000 399182
rect 697922 399114 707870 399120
rect 697922 399058 697992 399114
rect 698048 399058 698116 399114
rect 698172 399058 698240 399114
rect 698296 399058 698364 399114
rect 698420 399058 698488 399114
rect 698544 399058 698612 399114
rect 698668 399058 698736 399114
rect 698792 399064 707870 399114
rect 707926 399064 708000 399120
rect 698792 399058 708000 399064
rect 697922 398996 708000 399058
rect 697922 398990 707870 398996
rect 697922 398934 697992 398990
rect 698048 398934 698116 398990
rect 698172 398934 698240 398990
rect 698296 398934 698364 398990
rect 698420 398934 698488 398990
rect 698544 398934 698612 398990
rect 698668 398934 698736 398990
rect 698792 398940 707870 398990
rect 707926 398940 708000 398996
rect 698792 398934 708000 398940
rect 697922 398872 708000 398934
rect 697922 398866 707870 398872
rect 697922 398810 697992 398866
rect 698048 398810 698116 398866
rect 698172 398810 698240 398866
rect 698296 398810 698364 398866
rect 698420 398810 698488 398866
rect 698544 398810 698612 398866
rect 698668 398810 698736 398866
rect 698792 398816 707870 398866
rect 707926 398816 708000 398872
rect 698792 398810 708000 398816
rect 697922 398752 708000 398810
rect 697922 398134 708000 398172
rect 697922 398122 707870 398134
rect 697922 398066 697992 398122
rect 698048 398066 698116 398122
rect 698172 398066 698240 398122
rect 698296 398066 698364 398122
rect 698420 398066 698488 398122
rect 698544 398066 698612 398122
rect 698668 398066 698736 398122
rect 698792 398078 707870 398122
rect 707926 398078 708000 398134
rect 698792 398066 708000 398078
rect 697922 398010 708000 398066
rect 697922 397998 707870 398010
rect 697922 397942 697992 397998
rect 698048 397942 698116 397998
rect 698172 397942 698240 397998
rect 698296 397942 698364 397998
rect 698420 397942 698488 397998
rect 698544 397942 698612 397998
rect 698668 397942 698736 397998
rect 698792 397954 707870 397998
rect 707926 397954 708000 398010
rect 698792 397942 708000 397954
rect 697922 397886 708000 397942
rect 697922 397874 707870 397886
rect 697922 397818 697992 397874
rect 698048 397818 698116 397874
rect 698172 397818 698240 397874
rect 698296 397818 698364 397874
rect 698420 397818 698488 397874
rect 698544 397818 698612 397874
rect 698668 397818 698736 397874
rect 698792 397830 707870 397874
rect 707926 397830 708000 397886
rect 698792 397818 708000 397830
rect 697922 397762 708000 397818
rect 697922 397750 707870 397762
rect 697922 397694 697992 397750
rect 698048 397694 698116 397750
rect 698172 397694 698240 397750
rect 698296 397694 698364 397750
rect 698420 397694 698488 397750
rect 698544 397694 698612 397750
rect 698668 397694 698736 397750
rect 698792 397706 707870 397750
rect 707926 397706 708000 397762
rect 698792 397694 708000 397706
rect 697922 397638 708000 397694
rect 697922 397626 707870 397638
rect 697922 397570 697992 397626
rect 698048 397570 698116 397626
rect 698172 397570 698240 397626
rect 698296 397570 698364 397626
rect 698420 397570 698488 397626
rect 698544 397570 698612 397626
rect 698668 397570 698736 397626
rect 698792 397582 707870 397626
rect 707926 397582 708000 397638
rect 698792 397570 708000 397582
rect 697922 397514 708000 397570
rect 697922 397502 707870 397514
rect 697922 397446 697992 397502
rect 698048 397446 698116 397502
rect 698172 397446 698240 397502
rect 698296 397446 698364 397502
rect 698420 397446 698488 397502
rect 698544 397446 698612 397502
rect 698668 397446 698736 397502
rect 698792 397458 707870 397502
rect 707926 397458 708000 397514
rect 698792 397446 708000 397458
rect 697922 397390 708000 397446
rect 697922 397378 707870 397390
rect 697922 397322 697992 397378
rect 698048 397322 698116 397378
rect 698172 397322 698240 397378
rect 698296 397322 698364 397378
rect 698420 397322 698488 397378
rect 698544 397322 698612 397378
rect 698668 397322 698736 397378
rect 698792 397334 707870 397378
rect 707926 397334 708000 397390
rect 698792 397322 708000 397334
rect 697922 397266 708000 397322
rect 697922 397254 707870 397266
rect 697922 397198 697992 397254
rect 698048 397198 698116 397254
rect 698172 397198 698240 397254
rect 698296 397198 698364 397254
rect 698420 397198 698488 397254
rect 698544 397198 698612 397254
rect 698668 397198 698736 397254
rect 698792 397210 707870 397254
rect 707926 397210 708000 397266
rect 698792 397198 708000 397210
rect 697922 397142 708000 397198
rect 697922 397130 707870 397142
rect 697922 397074 697992 397130
rect 698048 397074 698116 397130
rect 698172 397074 698240 397130
rect 698296 397074 698364 397130
rect 698420 397074 698488 397130
rect 698544 397074 698612 397130
rect 698668 397074 698736 397130
rect 698792 397086 707870 397130
rect 707926 397086 708000 397142
rect 698792 397074 708000 397086
rect 697922 397018 708000 397074
rect 697922 397006 707870 397018
rect 697922 396950 697992 397006
rect 698048 396950 698116 397006
rect 698172 396950 698240 397006
rect 698296 396950 698364 397006
rect 698420 396950 698488 397006
rect 698544 396950 698612 397006
rect 698668 396950 698736 397006
rect 698792 396962 707870 397006
rect 707926 396962 708000 397018
rect 698792 396950 708000 396962
rect 697922 396894 708000 396950
rect 697922 396882 707870 396894
rect 697922 396826 697992 396882
rect 698048 396826 698116 396882
rect 698172 396826 698240 396882
rect 698296 396826 698364 396882
rect 698420 396826 698488 396882
rect 698544 396826 698612 396882
rect 698668 396826 698736 396882
rect 698792 396838 707870 396882
rect 707926 396838 708000 396894
rect 698792 396826 708000 396838
rect 697922 396770 708000 396826
rect 697922 396758 707870 396770
rect 75376 396622 80078 396744
rect 75376 396566 79300 396622
rect 79356 396566 79600 396622
rect 79656 396566 79900 396622
rect 79956 396566 80078 396622
rect 75376 396424 80078 396566
rect 697922 396702 697992 396758
rect 698048 396702 698116 396758
rect 698172 396702 698240 396758
rect 698296 396702 698364 396758
rect 698420 396702 698488 396758
rect 698544 396702 698612 396758
rect 698668 396702 698736 396758
rect 698792 396714 707870 396758
rect 707926 396714 708000 396770
rect 698792 396702 708000 396714
rect 697922 396646 708000 396702
rect 697922 396634 707870 396646
rect 697922 396578 697992 396634
rect 698048 396578 698116 396634
rect 698172 396578 698240 396634
rect 698296 396578 698364 396634
rect 698420 396578 698488 396634
rect 698544 396578 698612 396634
rect 698668 396578 698736 396634
rect 698792 396590 707870 396634
rect 707926 396590 708000 396646
rect 698792 396578 708000 396590
rect 697922 396522 708000 396578
rect 697922 396510 707870 396522
rect 697922 396454 697992 396510
rect 698048 396454 698116 396510
rect 698172 396454 698240 396510
rect 698296 396454 698364 396510
rect 698420 396454 698488 396510
rect 698544 396454 698612 396510
rect 698668 396454 698736 396510
rect 698792 396466 707870 396510
rect 707926 396466 708000 396522
rect 698792 396454 708000 396466
rect 697922 396398 708000 396454
rect 697922 396386 707870 396398
rect 697922 396330 697992 396386
rect 698048 396330 698116 396386
rect 698172 396330 698240 396386
rect 698296 396330 698364 396386
rect 698420 396330 698488 396386
rect 698544 396330 698612 396386
rect 698668 396330 698736 396386
rect 698792 396342 707870 396386
rect 707926 396342 708000 396398
rect 698792 396330 708000 396342
rect 697922 396272 708000 396330
rect 75312 393102 78678 393244
rect 75312 393046 77900 393102
rect 77956 393046 78200 393102
rect 78256 393046 78500 393102
rect 78556 393046 78678 393102
rect 75312 392924 78678 393046
rect 79078 392429 83556 392630
rect 79078 392373 79200 392429
rect 79256 392373 79500 392429
rect 79556 392373 79800 392429
rect 79856 392373 83556 392429
rect 79078 392229 83556 392373
rect 79078 392173 79200 392229
rect 79256 392173 79500 392229
rect 79556 392173 79800 392229
rect 79856 392173 83556 392229
rect 79078 392010 83556 392173
rect 688372 392429 698922 392630
rect 688372 392373 698144 392429
rect 698200 392373 698444 392429
rect 698500 392373 698744 392429
rect 698800 392373 698922 392429
rect 688372 392229 698922 392373
rect 688372 392173 698144 392229
rect 698200 392173 698444 392229
rect 698500 392173 698744 392229
rect 698800 392173 698922 392229
rect 688372 392010 698922 392173
rect 75376 389622 80078 389744
rect 75376 389566 79300 389622
rect 79356 389566 79600 389622
rect 79656 389566 79900 389622
rect 79956 389566 80078 389622
rect 75376 389424 80078 389566
rect 75312 386102 78678 386244
rect 75312 386046 77900 386102
rect 77956 386046 78200 386102
rect 78256 386046 78500 386102
rect 78556 386046 78678 386102
rect 75312 385924 78678 386046
rect 75376 382622 80078 382744
rect 75376 382566 79300 382622
rect 79356 382566 79600 382622
rect 79656 382566 79900 382622
rect 79956 382566 80078 382622
rect 75376 382424 80078 382566
rect 75312 379102 78678 379244
rect 75312 379046 77900 379102
rect 77956 379046 78200 379102
rect 78256 379046 78500 379102
rect 78556 379046 78678 379102
rect 75312 378924 78678 379046
rect 77678 374429 84516 374630
rect 77678 374373 77800 374429
rect 77856 374373 78100 374429
rect 78156 374373 78400 374429
rect 78456 374373 84516 374429
rect 77678 374229 84516 374373
rect 77678 374173 77800 374229
rect 77856 374173 78100 374229
rect 78156 374173 78400 374229
rect 78456 374173 84516 374229
rect 77678 374010 84516 374173
rect 687412 374429 700322 374630
rect 687412 374373 699544 374429
rect 699600 374373 699844 374429
rect 699900 374373 700144 374429
rect 700200 374373 700322 374429
rect 687412 374229 700322 374373
rect 687412 374173 699544 374229
rect 699600 374173 699844 374229
rect 699900 374173 700144 374229
rect 700200 374173 700322 374229
rect 687412 374010 700322 374173
rect 76115 372048 80078 372110
rect 76115 371992 79284 372048
rect 79340 371992 79584 372048
rect 79640 371992 79884 372048
rect 79940 371992 80078 372048
rect 76115 371910 80078 371992
rect 76115 371510 76435 371910
rect 76915 371633 78678 371710
rect 76915 371577 77847 371633
rect 77903 371577 78147 371633
rect 78203 371577 78447 371633
rect 78503 371577 78678 371633
rect 76915 371510 78678 371577
rect 699322 366954 702688 367076
rect 699322 366898 699444 366954
rect 699500 366898 699744 366954
rect 699800 366898 700044 366954
rect 700100 366898 702688 366954
rect 699322 366756 702688 366898
rect 697922 363434 702624 363576
rect 697922 363378 698044 363434
rect 698100 363378 698344 363434
rect 698400 363378 698644 363434
rect 698700 363378 702624 363434
rect 697922 363256 702624 363378
rect 699322 359954 702688 360076
rect 699322 359898 699444 359954
rect 699500 359898 699744 359954
rect 699800 359898 700044 359954
rect 700100 359898 702688 359954
rect 699322 359756 702688 359898
rect 79078 356429 83556 356630
rect 79078 356373 79200 356429
rect 79256 356373 79500 356429
rect 79556 356373 79800 356429
rect 79856 356373 83556 356429
rect 79078 356229 83556 356373
rect 79078 356173 79200 356229
rect 79256 356173 79500 356229
rect 79556 356173 79800 356229
rect 79856 356173 83556 356229
rect 79078 356010 83556 356173
rect 688372 356576 698922 356630
rect 688372 356429 702624 356576
rect 688372 356373 698144 356429
rect 698200 356373 698444 356429
rect 698500 356373 698744 356429
rect 698800 356373 702624 356429
rect 688372 356256 702624 356373
rect 688372 356229 698922 356256
rect 688372 356173 698144 356229
rect 698200 356173 698444 356229
rect 698500 356173 698744 356229
rect 698800 356173 698922 356229
rect 688372 356010 698922 356173
rect 75376 355622 80078 355744
rect 75376 355566 79300 355622
rect 79356 355566 79600 355622
rect 79656 355566 79900 355622
rect 79956 355566 80078 355622
rect 75376 355424 80078 355566
rect 699322 352954 702688 353076
rect 699322 352898 699444 352954
rect 699500 352898 699744 352954
rect 699800 352898 700044 352954
rect 700100 352898 702688 352954
rect 699322 352756 702688 352898
rect 75312 352102 78678 352244
rect 75312 352046 77900 352102
rect 77956 352046 78200 352102
rect 78256 352046 78500 352102
rect 78556 352046 78678 352102
rect 75312 351924 78678 352046
rect 697922 349434 702624 349576
rect 697922 349378 698044 349434
rect 698100 349378 698344 349434
rect 698400 349378 698644 349434
rect 698700 349378 702624 349434
rect 697922 349256 702624 349378
rect 75376 348622 80078 348744
rect 75376 348566 79300 348622
rect 79356 348566 79600 348622
rect 79656 348566 79900 348622
rect 79956 348566 80078 348622
rect 75376 348424 80078 348566
rect 75312 345102 78678 345244
rect 75312 345046 77900 345102
rect 77956 345046 78200 345102
rect 78256 345046 78500 345102
rect 78556 345046 78678 345102
rect 75312 344924 78678 345046
rect 75376 341622 80078 341744
rect 75376 341566 79300 341622
rect 79356 341566 79600 341622
rect 79656 341566 79900 341622
rect 79956 341566 80078 341622
rect 75376 341424 80078 341566
rect 77678 338429 84516 338630
rect 77678 338373 77800 338429
rect 77856 338373 78100 338429
rect 78156 338373 78400 338429
rect 78456 338373 84516 338429
rect 77678 338244 84516 338373
rect 75312 338229 84516 338244
rect 75312 338173 77800 338229
rect 77856 338173 78100 338229
rect 78156 338173 78400 338229
rect 78456 338173 84516 338229
rect 75312 338102 84516 338173
rect 75312 338046 77900 338102
rect 77956 338046 78200 338102
rect 78256 338046 78500 338102
rect 78556 338046 84516 338102
rect 75312 338010 84516 338046
rect 687412 338429 700322 338630
rect 687412 338373 699544 338429
rect 699600 338373 699844 338429
rect 699900 338373 700144 338429
rect 700200 338373 700322 338429
rect 687412 338229 700322 338373
rect 687412 338173 699544 338229
rect 699600 338173 699844 338229
rect 699900 338173 700144 338229
rect 700200 338173 700322 338229
rect 687412 338010 700322 338173
rect 75312 337924 78678 338010
rect 699322 333423 701085 333490
rect 699322 333367 699497 333423
rect 699553 333367 699797 333423
rect 699853 333367 700097 333423
rect 700153 333367 701085 333423
rect 699322 333290 701085 333367
rect 701565 333090 701885 333490
rect 697922 333008 701885 333090
rect 697922 332952 698060 333008
rect 698116 332952 698360 333008
rect 698416 332952 698660 333008
rect 698716 332952 701885 333008
rect 697922 332890 701885 332952
rect 76115 331040 698922 331110
rect 76115 330984 79208 331040
rect 79264 330984 79332 331040
rect 79388 330984 79456 331040
rect 79512 330984 79580 331040
rect 79636 330984 79704 331040
rect 79760 330984 79828 331040
rect 79884 330984 79952 331040
rect 80008 330984 158178 331040
rect 158234 330984 158302 331040
rect 158358 330984 158426 331040
rect 158482 330984 158550 331040
rect 158606 330984 381310 331040
rect 381366 330984 381434 331040
rect 381490 330984 381558 331040
rect 381614 330984 381682 331040
rect 381738 330984 698052 331040
rect 698108 330984 698176 331040
rect 698232 330984 698300 331040
rect 698356 330984 698424 331040
rect 698480 330984 698548 331040
rect 698604 330984 698672 331040
rect 698728 330984 698796 331040
rect 698852 330984 698922 331040
rect 76115 330916 698922 330984
rect 76115 330910 79208 330916
rect 76115 330510 76435 330910
rect 79078 330860 79208 330910
rect 79264 330860 79332 330916
rect 79388 330860 79456 330916
rect 79512 330860 79580 330916
rect 79636 330860 79704 330916
rect 79760 330860 79828 330916
rect 79884 330860 79952 330916
rect 80008 330888 158178 330916
rect 80008 330860 106207 330888
rect 79078 330832 106207 330860
rect 106263 330832 106407 330888
rect 106463 330832 142207 330888
rect 142263 330832 142407 330888
rect 142463 330860 158178 330888
rect 158234 330860 158302 330916
rect 158358 330860 158426 330916
rect 158482 330860 158550 330916
rect 158606 330888 381310 330916
rect 158606 330860 178207 330888
rect 142463 330832 178207 330860
rect 178263 330832 178407 330888
rect 178463 330832 214207 330888
rect 214263 330832 214407 330888
rect 214463 330832 250207 330888
rect 250263 330832 250407 330888
rect 250463 330832 286207 330888
rect 286263 330832 286407 330888
rect 286463 330832 322207 330888
rect 322263 330832 322407 330888
rect 322463 330832 358207 330888
rect 358263 330832 358407 330888
rect 358463 330860 381310 330888
rect 381366 330860 381434 330916
rect 381490 330860 381558 330916
rect 381614 330860 381682 330916
rect 381738 330888 698052 330916
rect 381738 330860 394207 330888
rect 358463 330832 394207 330860
rect 394263 330832 394407 330888
rect 394463 330832 430207 330888
rect 430263 330832 430407 330888
rect 430463 330832 466207 330888
rect 466263 330832 466407 330888
rect 466463 330832 502207 330888
rect 502263 330832 502407 330888
rect 502463 330832 538207 330888
rect 538263 330832 538407 330888
rect 538463 330832 574207 330888
rect 574263 330832 574407 330888
rect 574463 330832 610207 330888
rect 610263 330832 610407 330888
rect 610463 330832 646207 330888
rect 646263 330832 646407 330888
rect 646463 330832 682207 330888
rect 682263 330832 682407 330888
rect 682463 330860 698052 330888
rect 698108 330860 698176 330916
rect 698232 330860 698300 330916
rect 698356 330860 698424 330916
rect 698480 330860 698548 330916
rect 698604 330860 698672 330916
rect 698728 330860 698796 330916
rect 698852 330860 698922 330916
rect 682463 330832 698922 330860
rect 79078 330792 698922 330832
rect 79078 330736 79208 330792
rect 79264 330736 79332 330792
rect 79388 330736 79456 330792
rect 79512 330736 79580 330792
rect 79636 330736 79704 330792
rect 79760 330736 79828 330792
rect 79884 330736 79952 330792
rect 80008 330736 158178 330792
rect 158234 330736 158302 330792
rect 158358 330736 158426 330792
rect 158482 330736 158550 330792
rect 158606 330736 381310 330792
rect 381366 330736 381434 330792
rect 381490 330736 381558 330792
rect 381614 330736 381682 330792
rect 381738 330736 698052 330792
rect 698108 330736 698176 330792
rect 698232 330736 698300 330792
rect 698356 330736 698424 330792
rect 698480 330736 698548 330792
rect 698604 330736 698672 330792
rect 698728 330736 698796 330792
rect 698852 330736 698922 330792
rect 76915 330633 78678 330710
rect 76915 330577 77847 330633
rect 77903 330577 78147 330633
rect 78203 330577 78447 330633
rect 78503 330577 78678 330633
rect 76915 330510 78678 330577
rect 79078 330668 698922 330736
rect 79078 330612 79208 330668
rect 79264 330612 79332 330668
rect 79388 330612 79456 330668
rect 79512 330612 79580 330668
rect 79636 330612 79704 330668
rect 79760 330612 79828 330668
rect 79884 330612 79952 330668
rect 80008 330612 158178 330668
rect 158234 330612 158302 330668
rect 158358 330612 158426 330668
rect 158482 330612 158550 330668
rect 158606 330612 381310 330668
rect 381366 330612 381434 330668
rect 381490 330612 381558 330668
rect 381614 330612 381682 330668
rect 381738 330612 698052 330668
rect 698108 330612 698176 330668
rect 698232 330612 698300 330668
rect 698356 330612 698424 330668
rect 698480 330612 698548 330668
rect 698604 330612 698672 330668
rect 698728 330612 698796 330668
rect 698852 330612 698922 330668
rect 79078 330588 698922 330612
rect 79078 330544 106207 330588
rect 79078 330488 79208 330544
rect 79264 330488 79332 330544
rect 79388 330488 79456 330544
rect 79512 330488 79580 330544
rect 79636 330488 79704 330544
rect 79760 330488 79828 330544
rect 79884 330488 79952 330544
rect 80008 330532 106207 330544
rect 106263 330532 106407 330588
rect 106463 330532 142207 330588
rect 142263 330532 142407 330588
rect 142463 330544 178207 330588
rect 142463 330532 158178 330544
rect 80008 330488 158178 330532
rect 158234 330488 158302 330544
rect 158358 330488 158426 330544
rect 158482 330488 158550 330544
rect 158606 330532 178207 330544
rect 178263 330532 178407 330588
rect 178463 330532 214207 330588
rect 214263 330532 214407 330588
rect 214463 330532 250207 330588
rect 250263 330532 250407 330588
rect 250463 330532 286207 330588
rect 286263 330532 286407 330588
rect 286463 330532 322207 330588
rect 322263 330532 322407 330588
rect 322463 330532 358207 330588
rect 358263 330532 358407 330588
rect 358463 330544 394207 330588
rect 358463 330532 381310 330544
rect 158606 330488 381310 330532
rect 381366 330488 381434 330544
rect 381490 330488 381558 330544
rect 381614 330488 381682 330544
rect 381738 330532 394207 330544
rect 394263 330532 394407 330588
rect 394463 330532 430207 330588
rect 430263 330532 430407 330588
rect 430463 330532 466207 330588
rect 466263 330532 466407 330588
rect 466463 330532 502207 330588
rect 502263 330532 502407 330588
rect 502463 330532 538207 330588
rect 538263 330532 538407 330588
rect 538463 330532 574207 330588
rect 574263 330532 574407 330588
rect 574463 330532 610207 330588
rect 610263 330532 610407 330588
rect 610463 330532 646207 330588
rect 646263 330532 646407 330588
rect 646463 330532 682207 330588
rect 682263 330532 682407 330588
rect 682463 330544 698922 330588
rect 682463 330532 698052 330544
rect 381738 330488 698052 330532
rect 698108 330488 698176 330544
rect 698232 330488 698300 330544
rect 698356 330488 698424 330544
rect 698480 330488 698548 330544
rect 698604 330488 698672 330544
rect 698728 330488 698796 330544
rect 698852 330488 698922 330544
rect 79078 330420 698922 330488
rect 79078 330364 79208 330420
rect 79264 330364 79332 330420
rect 79388 330364 79456 330420
rect 79512 330364 79580 330420
rect 79636 330364 79704 330420
rect 79760 330364 79828 330420
rect 79884 330364 79952 330420
rect 80008 330364 158178 330420
rect 158234 330364 158302 330420
rect 158358 330364 158426 330420
rect 158482 330364 158550 330420
rect 158606 330364 381310 330420
rect 381366 330364 381434 330420
rect 381490 330364 381558 330420
rect 381614 330364 381682 330420
rect 381738 330364 698052 330420
rect 698108 330364 698176 330420
rect 698232 330364 698300 330420
rect 698356 330364 698424 330420
rect 698480 330364 698548 330420
rect 698604 330364 698672 330420
rect 698728 330364 698796 330420
rect 698852 330364 698922 330420
rect 79078 330296 698922 330364
rect 79078 330240 79208 330296
rect 79264 330240 79332 330296
rect 79388 330240 79456 330296
rect 79512 330240 79580 330296
rect 79636 330240 79704 330296
rect 79760 330240 79828 330296
rect 79884 330240 79952 330296
rect 80008 330288 158178 330296
rect 80008 330240 106207 330288
rect 79078 330232 106207 330240
rect 106263 330232 106407 330288
rect 106463 330232 142207 330288
rect 142263 330232 142407 330288
rect 142463 330240 158178 330288
rect 158234 330240 158302 330296
rect 158358 330240 158426 330296
rect 158482 330240 158550 330296
rect 158606 330288 381310 330296
rect 158606 330240 178207 330288
rect 142463 330232 178207 330240
rect 178263 330232 178407 330288
rect 178463 330232 214207 330288
rect 214263 330232 214407 330288
rect 214463 330232 250207 330288
rect 250263 330232 250407 330288
rect 250463 330232 286207 330288
rect 286263 330232 286407 330288
rect 286463 330232 322207 330288
rect 322263 330232 322407 330288
rect 322463 330232 358207 330288
rect 358263 330232 358407 330288
rect 358463 330240 381310 330288
rect 381366 330240 381434 330296
rect 381490 330240 381558 330296
rect 381614 330240 381682 330296
rect 381738 330288 698052 330296
rect 381738 330240 394207 330288
rect 358463 330232 394207 330240
rect 394263 330232 394407 330288
rect 394463 330232 430207 330288
rect 430263 330232 430407 330288
rect 430463 330232 466207 330288
rect 466263 330232 466407 330288
rect 466463 330232 502207 330288
rect 502263 330232 502407 330288
rect 502463 330232 538207 330288
rect 538263 330232 538407 330288
rect 538463 330232 574207 330288
rect 574263 330232 574407 330288
rect 574463 330232 610207 330288
rect 610263 330232 610407 330288
rect 610463 330232 646207 330288
rect 646263 330232 646407 330288
rect 646463 330232 682207 330288
rect 682263 330232 682407 330288
rect 682463 330240 698052 330288
rect 698108 330240 698176 330296
rect 698232 330240 698300 330296
rect 698356 330240 698424 330296
rect 698480 330240 698548 330296
rect 698604 330240 698672 330296
rect 698728 330240 698796 330296
rect 698852 330240 698922 330296
rect 682463 330232 698922 330240
rect 79078 330110 698922 330232
rect 77678 329640 700322 329710
rect 77678 329584 77808 329640
rect 77864 329584 77932 329640
rect 77988 329584 78056 329640
rect 78112 329584 78180 329640
rect 78236 329584 78304 329640
rect 78360 329584 78428 329640
rect 78484 329584 78552 329640
rect 78608 329584 157158 329640
rect 157214 329584 157282 329640
rect 157338 329584 157406 329640
rect 157462 329584 157530 329640
rect 157586 329584 382330 329640
rect 382386 329584 382454 329640
rect 382510 329584 382578 329640
rect 382634 329584 382702 329640
rect 382758 329584 699452 329640
rect 699508 329584 699576 329640
rect 699632 329584 699700 329640
rect 699756 329584 699824 329640
rect 699880 329584 699948 329640
rect 700004 329584 700072 329640
rect 700128 329584 700196 329640
rect 700252 329584 700322 329640
rect 77678 329516 700322 329584
rect 77678 329460 77808 329516
rect 77864 329460 77932 329516
rect 77988 329460 78056 329516
rect 78112 329460 78180 329516
rect 78236 329460 78304 329516
rect 78360 329460 78428 329516
rect 78484 329460 78552 329516
rect 78608 329488 157158 329516
rect 78608 329460 88207 329488
rect 77678 329432 88207 329460
rect 88263 329432 88407 329488
rect 88463 329432 124207 329488
rect 124263 329432 124407 329488
rect 124463 329460 157158 329488
rect 157214 329460 157282 329516
rect 157338 329460 157406 329516
rect 157462 329460 157530 329516
rect 157586 329488 382330 329516
rect 157586 329460 160207 329488
rect 124463 329432 160207 329460
rect 160263 329432 160407 329488
rect 160463 329432 196207 329488
rect 196263 329432 196407 329488
rect 196463 329432 232207 329488
rect 232263 329432 232407 329488
rect 232463 329432 268207 329488
rect 268263 329432 268407 329488
rect 268463 329432 304207 329488
rect 304263 329432 304407 329488
rect 304463 329432 340207 329488
rect 340263 329432 340407 329488
rect 340463 329432 376207 329488
rect 376263 329432 376407 329488
rect 376463 329460 382330 329488
rect 382386 329460 382454 329516
rect 382510 329460 382578 329516
rect 382634 329460 382702 329516
rect 382758 329488 699452 329516
rect 382758 329460 412207 329488
rect 376463 329432 412207 329460
rect 412263 329432 412407 329488
rect 412463 329432 448207 329488
rect 448263 329432 448407 329488
rect 448463 329432 484207 329488
rect 484263 329432 484407 329488
rect 484463 329432 520207 329488
rect 520263 329432 520407 329488
rect 520463 329432 556207 329488
rect 556263 329432 556407 329488
rect 556463 329432 592207 329488
rect 592263 329432 592407 329488
rect 592463 329432 628207 329488
rect 628263 329432 628407 329488
rect 628463 329432 664207 329488
rect 664263 329432 664407 329488
rect 664463 329460 699452 329488
rect 699508 329460 699576 329516
rect 699632 329460 699700 329516
rect 699756 329460 699824 329516
rect 699880 329460 699948 329516
rect 700004 329460 700072 329516
rect 700128 329460 700196 329516
rect 700252 329460 700322 329516
rect 664463 329432 700322 329460
rect 77678 329392 700322 329432
rect 77678 329336 77808 329392
rect 77864 329336 77932 329392
rect 77988 329336 78056 329392
rect 78112 329336 78180 329392
rect 78236 329336 78304 329392
rect 78360 329336 78428 329392
rect 78484 329336 78552 329392
rect 78608 329336 157158 329392
rect 157214 329336 157282 329392
rect 157338 329336 157406 329392
rect 157462 329336 157530 329392
rect 157586 329336 382330 329392
rect 382386 329336 382454 329392
rect 382510 329336 382578 329392
rect 382634 329336 382702 329392
rect 382758 329336 699452 329392
rect 699508 329336 699576 329392
rect 699632 329336 699700 329392
rect 699756 329336 699824 329392
rect 699880 329336 699948 329392
rect 700004 329336 700072 329392
rect 700128 329336 700196 329392
rect 700252 329336 700322 329392
rect 77678 329268 700322 329336
rect 77678 329212 77808 329268
rect 77864 329212 77932 329268
rect 77988 329212 78056 329268
rect 78112 329212 78180 329268
rect 78236 329212 78304 329268
rect 78360 329212 78428 329268
rect 78484 329212 78552 329268
rect 78608 329212 157158 329268
rect 157214 329212 157282 329268
rect 157338 329212 157406 329268
rect 157462 329212 157530 329268
rect 157586 329212 382330 329268
rect 382386 329212 382454 329268
rect 382510 329212 382578 329268
rect 382634 329212 382702 329268
rect 382758 329212 699452 329268
rect 699508 329212 699576 329268
rect 699632 329212 699700 329268
rect 699756 329212 699824 329268
rect 699880 329212 699948 329268
rect 700004 329212 700072 329268
rect 700128 329212 700196 329268
rect 700252 329212 700322 329268
rect 77678 329188 700322 329212
rect 77678 329144 88207 329188
rect 77678 329088 77808 329144
rect 77864 329088 77932 329144
rect 77988 329088 78056 329144
rect 78112 329088 78180 329144
rect 78236 329088 78304 329144
rect 78360 329088 78428 329144
rect 78484 329088 78552 329144
rect 78608 329132 88207 329144
rect 88263 329132 88407 329188
rect 88463 329132 124207 329188
rect 124263 329132 124407 329188
rect 124463 329144 160207 329188
rect 124463 329132 157158 329144
rect 78608 329088 157158 329132
rect 157214 329088 157282 329144
rect 157338 329088 157406 329144
rect 157462 329088 157530 329144
rect 157586 329132 160207 329144
rect 160263 329132 160407 329188
rect 160463 329132 196207 329188
rect 196263 329132 196407 329188
rect 196463 329132 232207 329188
rect 232263 329132 232407 329188
rect 232463 329132 268207 329188
rect 268263 329132 268407 329188
rect 268463 329132 304207 329188
rect 304263 329132 304407 329188
rect 304463 329132 340207 329188
rect 340263 329132 340407 329188
rect 340463 329132 376207 329188
rect 376263 329132 376407 329188
rect 376463 329144 412207 329188
rect 376463 329132 382330 329144
rect 157586 329088 382330 329132
rect 382386 329088 382454 329144
rect 382510 329088 382578 329144
rect 382634 329088 382702 329144
rect 382758 329132 412207 329144
rect 412263 329132 412407 329188
rect 412463 329132 448207 329188
rect 448263 329132 448407 329188
rect 448463 329132 484207 329188
rect 484263 329132 484407 329188
rect 484463 329132 520207 329188
rect 520263 329132 520407 329188
rect 520463 329132 556207 329188
rect 556263 329132 556407 329188
rect 556463 329132 592207 329188
rect 592263 329132 592407 329188
rect 592463 329132 628207 329188
rect 628263 329132 628407 329188
rect 628463 329132 664207 329188
rect 664263 329132 664407 329188
rect 664463 329144 700322 329188
rect 664463 329132 699452 329144
rect 382758 329088 699452 329132
rect 699508 329088 699576 329144
rect 699632 329088 699700 329144
rect 699756 329088 699824 329144
rect 699880 329088 699948 329144
rect 700004 329088 700072 329144
rect 700128 329088 700196 329144
rect 700252 329088 700322 329144
rect 77678 329020 700322 329088
rect 77678 328964 77808 329020
rect 77864 328964 77932 329020
rect 77988 328964 78056 329020
rect 78112 328964 78180 329020
rect 78236 328964 78304 329020
rect 78360 328964 78428 329020
rect 78484 328964 78552 329020
rect 78608 328964 157158 329020
rect 157214 328964 157282 329020
rect 157338 328964 157406 329020
rect 157462 328964 157530 329020
rect 157586 328964 382330 329020
rect 382386 328964 382454 329020
rect 382510 328964 382578 329020
rect 382634 328964 382702 329020
rect 382758 328964 699452 329020
rect 699508 328964 699576 329020
rect 699632 328964 699700 329020
rect 699756 328964 699824 329020
rect 699880 328964 699948 329020
rect 700004 328964 700072 329020
rect 700128 328964 700196 329020
rect 700252 328964 700322 329020
rect 77678 328896 700322 328964
rect 77678 328840 77808 328896
rect 77864 328840 77932 328896
rect 77988 328840 78056 328896
rect 78112 328840 78180 328896
rect 78236 328840 78304 328896
rect 78360 328840 78428 328896
rect 78484 328840 78552 328896
rect 78608 328888 157158 328896
rect 78608 328840 88207 328888
rect 77678 328832 88207 328840
rect 88263 328832 88407 328888
rect 88463 328832 124207 328888
rect 124263 328832 124407 328888
rect 124463 328840 157158 328888
rect 157214 328840 157282 328896
rect 157338 328840 157406 328896
rect 157462 328840 157530 328896
rect 157586 328888 382330 328896
rect 157586 328840 160207 328888
rect 124463 328832 160207 328840
rect 160263 328832 160407 328888
rect 160463 328832 196207 328888
rect 196263 328832 196407 328888
rect 196463 328832 232207 328888
rect 232263 328832 232407 328888
rect 232463 328832 268207 328888
rect 268263 328832 268407 328888
rect 268463 328832 304207 328888
rect 304263 328832 304407 328888
rect 304463 328832 340207 328888
rect 340263 328832 340407 328888
rect 340463 328832 376207 328888
rect 376263 328832 376407 328888
rect 376463 328840 382330 328888
rect 382386 328840 382454 328896
rect 382510 328840 382578 328896
rect 382634 328840 382702 328896
rect 382758 328888 699452 328896
rect 382758 328840 412207 328888
rect 376463 328832 412207 328840
rect 412263 328832 412407 328888
rect 412463 328832 448207 328888
rect 448263 328832 448407 328888
rect 448463 328832 484207 328888
rect 484263 328832 484407 328888
rect 484463 328832 520207 328888
rect 520263 328832 520407 328888
rect 520463 328832 556207 328888
rect 556263 328832 556407 328888
rect 556463 328832 592207 328888
rect 592263 328832 592407 328888
rect 592463 328832 628207 328888
rect 628263 328832 628407 328888
rect 628463 328832 664207 328888
rect 664263 328832 664407 328888
rect 664463 328840 699452 328888
rect 699508 328840 699576 328896
rect 699632 328840 699700 328896
rect 699756 328840 699824 328896
rect 699880 328840 699948 328896
rect 700004 328840 700072 328896
rect 700128 328840 700196 328896
rect 700252 328840 700322 328896
rect 664463 328832 700322 328840
rect 77678 328710 700322 328832
rect 699322 323954 702688 324076
rect 699322 323898 699444 323954
rect 699500 323898 699744 323954
rect 699800 323898 700044 323954
rect 700100 323898 702688 323954
rect 699322 323756 702688 323898
rect 697922 320434 702624 320576
rect 697922 320378 698044 320434
rect 698100 320378 698344 320434
rect 698400 320378 698644 320434
rect 698700 320378 702624 320434
rect 697922 320256 702624 320378
rect 157088 318424 161684 318557
rect 157088 318368 157210 318424
rect 157266 318368 157510 318424
rect 157566 318368 161684 318424
rect 157088 318237 161684 318368
rect 378284 318426 382880 318557
rect 378284 318370 382402 318426
rect 382458 318370 382702 318426
rect 382758 318370 382880 318426
rect 378284 318237 382880 318370
rect 158108 317725 161684 317858
rect 158108 317669 158230 317725
rect 158286 317669 158530 317725
rect 158586 317669 161684 317725
rect 158108 317538 161684 317669
rect 378284 317727 381860 317858
rect 378284 317671 381382 317727
rect 381438 317671 381682 317727
rect 381738 317671 381860 317727
rect 378284 317538 381860 317671
rect 157088 317026 161684 317159
rect 157088 316970 157210 317026
rect 157266 316970 157510 317026
rect 157566 316970 161684 317026
rect 157088 316839 161684 316970
rect 378284 317028 382880 317159
rect 378284 316972 382402 317028
rect 382458 316972 382702 317028
rect 382758 316972 382880 317028
rect 378284 316839 382880 316972
rect 699322 316954 702688 317076
rect 699322 316898 699444 316954
rect 699500 316898 699744 316954
rect 699800 316898 700044 316954
rect 700100 316898 702688 316954
rect 699322 316756 702688 316898
rect 158108 316327 161684 316460
rect 158108 316271 158230 316327
rect 158286 316271 158530 316327
rect 158586 316271 161684 316327
rect 158108 316140 161684 316271
rect 378284 316329 381860 316460
rect 378284 316273 381382 316329
rect 381438 316273 381682 316329
rect 381738 316273 381860 316329
rect 378284 316140 381860 316273
rect 157088 315628 161684 315761
rect 157088 315572 157210 315628
rect 157266 315572 157510 315628
rect 157566 315572 161684 315628
rect 157088 315441 161684 315572
rect 378284 315630 382880 315761
rect 378284 315574 382402 315630
rect 382458 315574 382702 315630
rect 382758 315574 382880 315630
rect 378284 315441 382880 315574
rect 158108 314929 161684 315062
rect 158108 314873 158230 314929
rect 158286 314873 158530 314929
rect 158586 314873 161684 314929
rect 75376 314622 80078 314744
rect 158108 314742 161684 314873
rect 378284 314931 381860 315062
rect 378284 314875 381382 314931
rect 381438 314875 381682 314931
rect 381738 314875 381860 314931
rect 378284 314742 381860 314875
rect 75376 314566 79300 314622
rect 79356 314566 79600 314622
rect 79656 314566 79900 314622
rect 79956 314566 80078 314622
rect 75376 314424 80078 314566
rect 157088 314230 161684 314363
rect 157088 314174 157210 314230
rect 157266 314174 157510 314230
rect 157566 314174 161684 314230
rect 157088 314043 161684 314174
rect 378284 314232 382880 314363
rect 378284 314176 382402 314232
rect 382458 314176 382702 314232
rect 382758 314176 382880 314232
rect 378284 314043 382880 314176
rect 697922 313434 702624 313576
rect 697922 313378 698044 313434
rect 698100 313378 698344 313434
rect 698400 313378 698644 313434
rect 698700 313378 702624 313434
rect 697922 313256 702624 313378
rect 75312 311102 78678 311244
rect 75312 311046 77900 311102
rect 77956 311046 78200 311102
rect 78256 311046 78500 311102
rect 78556 311046 78678 311102
rect 75312 310924 78678 311046
rect 699322 309954 702688 310076
rect 699322 309898 699444 309954
rect 699500 309898 699744 309954
rect 699800 309898 700044 309954
rect 700100 309898 702688 309954
rect 699322 309756 702688 309898
rect 75376 307622 80078 307744
rect 75376 307566 79300 307622
rect 79356 307566 79600 307622
rect 79656 307566 79900 307622
rect 79956 307566 80078 307622
rect 75376 307424 80078 307566
rect 79078 307186 698922 307256
rect 79078 307130 79208 307186
rect 79264 307130 79332 307186
rect 79388 307130 79456 307186
rect 79512 307130 79580 307186
rect 79636 307130 79704 307186
rect 79760 307130 79828 307186
rect 79884 307130 79952 307186
rect 80008 307130 116220 307186
rect 116276 307130 116344 307186
rect 116400 307130 119410 307186
rect 119466 307130 119534 307186
rect 119590 307130 122600 307186
rect 122656 307130 122724 307186
rect 122780 307130 390220 307186
rect 390276 307130 390344 307186
rect 390400 307130 393410 307186
rect 393466 307130 393534 307186
rect 393590 307130 396600 307186
rect 396656 307130 396724 307186
rect 396780 307130 490220 307186
rect 490276 307130 490344 307186
rect 490400 307130 493410 307186
rect 493466 307130 493534 307186
rect 493590 307130 496600 307186
rect 496656 307130 496724 307186
rect 496780 307130 634860 307186
rect 634916 307130 634984 307186
rect 635040 307130 638050 307186
rect 638106 307130 638174 307186
rect 638230 307130 641240 307186
rect 641296 307130 641364 307186
rect 641420 307130 698052 307186
rect 698108 307130 698176 307186
rect 698232 307130 698300 307186
rect 698356 307130 698424 307186
rect 698480 307130 698548 307186
rect 698604 307130 698672 307186
rect 698728 307130 698796 307186
rect 698852 307130 698922 307186
rect 79078 307126 698922 307130
rect 79078 307070 158178 307126
rect 158234 307070 158302 307126
rect 158358 307070 158426 307126
rect 158482 307070 158550 307126
rect 158606 307070 381310 307126
rect 381366 307070 381434 307126
rect 381490 307070 381558 307126
rect 381614 307070 381682 307126
rect 381738 307070 590910 307126
rect 590966 307070 591034 307126
rect 591090 307070 591158 307126
rect 591214 307070 591282 307126
rect 591338 307070 591406 307126
rect 591462 307070 591530 307126
rect 591586 307070 591654 307126
rect 591710 307070 698922 307126
rect 79078 307062 698922 307070
rect 79078 307006 79208 307062
rect 79264 307006 79332 307062
rect 79388 307006 79456 307062
rect 79512 307006 79580 307062
rect 79636 307006 79704 307062
rect 79760 307006 79828 307062
rect 79884 307006 79952 307062
rect 80008 307006 116220 307062
rect 116276 307006 116344 307062
rect 116400 307006 119410 307062
rect 119466 307006 119534 307062
rect 119590 307006 122600 307062
rect 122656 307006 122724 307062
rect 122780 307006 390220 307062
rect 390276 307006 390344 307062
rect 390400 307006 393410 307062
rect 393466 307006 393534 307062
rect 393590 307006 396600 307062
rect 396656 307006 396724 307062
rect 396780 307006 490220 307062
rect 490276 307006 490344 307062
rect 490400 307006 493410 307062
rect 493466 307006 493534 307062
rect 493590 307006 496600 307062
rect 496656 307006 496724 307062
rect 496780 307006 634860 307062
rect 634916 307006 634984 307062
rect 635040 307006 638050 307062
rect 638106 307006 638174 307062
rect 638230 307006 641240 307062
rect 641296 307006 641364 307062
rect 641420 307006 698052 307062
rect 698108 307006 698176 307062
rect 698232 307006 698300 307062
rect 698356 307006 698424 307062
rect 698480 307006 698548 307062
rect 698604 307006 698672 307062
rect 698728 307006 698796 307062
rect 698852 307006 698922 307062
rect 79078 307002 698922 307006
rect 79078 306946 158178 307002
rect 158234 306946 158302 307002
rect 158358 306946 158426 307002
rect 158482 306946 158550 307002
rect 158606 306946 381310 307002
rect 381366 306946 381434 307002
rect 381490 306946 381558 307002
rect 381614 306946 381682 307002
rect 381738 306946 590910 307002
rect 590966 306946 591034 307002
rect 591090 306946 591158 307002
rect 591214 306946 591282 307002
rect 591338 306946 591406 307002
rect 591462 306946 591530 307002
rect 591586 306946 591654 307002
rect 591710 306946 698922 307002
rect 79078 306938 698922 306946
rect 79078 306882 79208 306938
rect 79264 306882 79332 306938
rect 79388 306882 79456 306938
rect 79512 306882 79580 306938
rect 79636 306882 79704 306938
rect 79760 306882 79828 306938
rect 79884 306882 79952 306938
rect 80008 306882 116220 306938
rect 116276 306882 116344 306938
rect 116400 306882 119410 306938
rect 119466 306882 119534 306938
rect 119590 306882 122600 306938
rect 122656 306882 122724 306938
rect 122780 306882 390220 306938
rect 390276 306882 390344 306938
rect 390400 306882 393410 306938
rect 393466 306882 393534 306938
rect 393590 306882 396600 306938
rect 396656 306882 396724 306938
rect 396780 306882 490220 306938
rect 490276 306882 490344 306938
rect 490400 306882 493410 306938
rect 493466 306882 493534 306938
rect 493590 306882 496600 306938
rect 496656 306882 496724 306938
rect 496780 306882 634860 306938
rect 634916 306882 634984 306938
rect 635040 306882 638050 306938
rect 638106 306882 638174 306938
rect 638230 306882 641240 306938
rect 641296 306882 641364 306938
rect 641420 306882 698052 306938
rect 698108 306882 698176 306938
rect 698232 306882 698300 306938
rect 698356 306882 698424 306938
rect 698480 306882 698548 306938
rect 698604 306882 698672 306938
rect 698728 306882 698796 306938
rect 698852 306882 698922 306938
rect 79078 306878 698922 306882
rect 79078 306822 158178 306878
rect 158234 306822 158302 306878
rect 158358 306822 158426 306878
rect 158482 306822 158550 306878
rect 158606 306822 381310 306878
rect 381366 306822 381434 306878
rect 381490 306822 381558 306878
rect 381614 306822 381682 306878
rect 381738 306822 590910 306878
rect 590966 306822 591034 306878
rect 591090 306822 591158 306878
rect 591214 306822 591282 306878
rect 591338 306822 591406 306878
rect 591462 306822 591530 306878
rect 591586 306822 591654 306878
rect 591710 306822 698922 306878
rect 79078 306814 698922 306822
rect 79078 306758 79208 306814
rect 79264 306758 79332 306814
rect 79388 306758 79456 306814
rect 79512 306758 79580 306814
rect 79636 306758 79704 306814
rect 79760 306758 79828 306814
rect 79884 306758 79952 306814
rect 80008 306758 116220 306814
rect 116276 306758 116344 306814
rect 116400 306758 119410 306814
rect 119466 306758 119534 306814
rect 119590 306758 122600 306814
rect 122656 306758 122724 306814
rect 122780 306758 390220 306814
rect 390276 306758 390344 306814
rect 390400 306758 393410 306814
rect 393466 306758 393534 306814
rect 393590 306758 396600 306814
rect 396656 306758 396724 306814
rect 396780 306758 490220 306814
rect 490276 306758 490344 306814
rect 490400 306758 493410 306814
rect 493466 306758 493534 306814
rect 493590 306758 496600 306814
rect 496656 306758 496724 306814
rect 496780 306758 634860 306814
rect 634916 306758 634984 306814
rect 635040 306758 638050 306814
rect 638106 306758 638174 306814
rect 638230 306758 641240 306814
rect 641296 306758 641364 306814
rect 641420 306758 698052 306814
rect 698108 306758 698176 306814
rect 698232 306758 698300 306814
rect 698356 306758 698424 306814
rect 698480 306758 698548 306814
rect 698604 306758 698672 306814
rect 698728 306758 698796 306814
rect 698852 306758 698922 306814
rect 79078 306754 698922 306758
rect 79078 306698 158178 306754
rect 158234 306698 158302 306754
rect 158358 306698 158426 306754
rect 158482 306698 158550 306754
rect 158606 306698 381310 306754
rect 381366 306698 381434 306754
rect 381490 306698 381558 306754
rect 381614 306698 381682 306754
rect 381738 306698 590910 306754
rect 590966 306698 591034 306754
rect 591090 306698 591158 306754
rect 591214 306698 591282 306754
rect 591338 306698 591406 306754
rect 591462 306698 591530 306754
rect 591586 306698 591654 306754
rect 591710 306698 698922 306754
rect 79078 306690 698922 306698
rect 79078 306634 79208 306690
rect 79264 306634 79332 306690
rect 79388 306634 79456 306690
rect 79512 306634 79580 306690
rect 79636 306634 79704 306690
rect 79760 306634 79828 306690
rect 79884 306634 79952 306690
rect 80008 306634 116220 306690
rect 116276 306634 116344 306690
rect 116400 306634 119410 306690
rect 119466 306634 119534 306690
rect 119590 306634 122600 306690
rect 122656 306634 122724 306690
rect 122780 306634 390220 306690
rect 390276 306634 390344 306690
rect 390400 306634 393410 306690
rect 393466 306634 393534 306690
rect 393590 306634 396600 306690
rect 396656 306634 396724 306690
rect 396780 306634 490220 306690
rect 490276 306634 490344 306690
rect 490400 306634 493410 306690
rect 493466 306634 493534 306690
rect 493590 306634 496600 306690
rect 496656 306634 496724 306690
rect 496780 306634 634860 306690
rect 634916 306634 634984 306690
rect 635040 306634 638050 306690
rect 638106 306634 638174 306690
rect 638230 306634 641240 306690
rect 641296 306634 641364 306690
rect 641420 306634 698052 306690
rect 698108 306634 698176 306690
rect 698232 306634 698300 306690
rect 698356 306634 698424 306690
rect 698480 306634 698548 306690
rect 698604 306634 698672 306690
rect 698728 306634 698796 306690
rect 698852 306634 698922 306690
rect 79078 306630 698922 306634
rect 79078 306574 158178 306630
rect 158234 306574 158302 306630
rect 158358 306574 158426 306630
rect 158482 306574 158550 306630
rect 158606 306574 381310 306630
rect 381366 306574 381434 306630
rect 381490 306574 381558 306630
rect 381614 306574 381682 306630
rect 381738 306574 590910 306630
rect 590966 306574 591034 306630
rect 591090 306574 591158 306630
rect 591214 306574 591282 306630
rect 591338 306574 591406 306630
rect 591462 306574 591530 306630
rect 591586 306574 591654 306630
rect 591710 306576 698922 306630
rect 591710 306574 702624 306576
rect 79078 306566 702624 306574
rect 79078 306510 79208 306566
rect 79264 306510 79332 306566
rect 79388 306510 79456 306566
rect 79512 306510 79580 306566
rect 79636 306510 79704 306566
rect 79760 306510 79828 306566
rect 79884 306510 79952 306566
rect 80008 306510 116220 306566
rect 116276 306510 116344 306566
rect 116400 306510 119410 306566
rect 119466 306510 119534 306566
rect 119590 306510 122600 306566
rect 122656 306510 122724 306566
rect 122780 306510 390220 306566
rect 390276 306510 390344 306566
rect 390400 306510 393410 306566
rect 393466 306510 393534 306566
rect 393590 306510 396600 306566
rect 396656 306510 396724 306566
rect 396780 306510 490220 306566
rect 490276 306510 490344 306566
rect 490400 306510 493410 306566
rect 493466 306510 493534 306566
rect 493590 306510 496600 306566
rect 496656 306510 496724 306566
rect 496780 306510 634860 306566
rect 634916 306510 634984 306566
rect 635040 306510 638050 306566
rect 638106 306510 638174 306566
rect 638230 306510 641240 306566
rect 641296 306510 641364 306566
rect 641420 306510 698052 306566
rect 698108 306510 698176 306566
rect 698232 306510 698300 306566
rect 698356 306510 698424 306566
rect 698480 306510 698548 306566
rect 698604 306510 698672 306566
rect 698728 306510 698796 306566
rect 698852 306510 702624 306566
rect 79078 306506 702624 306510
rect 79078 306450 158178 306506
rect 158234 306450 158302 306506
rect 158358 306450 158426 306506
rect 158482 306450 158550 306506
rect 158606 306450 381310 306506
rect 381366 306450 381434 306506
rect 381490 306450 381558 306506
rect 381614 306450 381682 306506
rect 381738 306450 590910 306506
rect 590966 306450 591034 306506
rect 591090 306450 591158 306506
rect 591214 306450 591282 306506
rect 591338 306450 591406 306506
rect 591462 306450 591530 306506
rect 591586 306450 591654 306506
rect 591710 306450 702624 306506
rect 79078 306442 702624 306450
rect 79078 306386 79208 306442
rect 79264 306386 79332 306442
rect 79388 306386 79456 306442
rect 79512 306386 79580 306442
rect 79636 306386 79704 306442
rect 79760 306386 79828 306442
rect 79884 306386 79952 306442
rect 80008 306386 116220 306442
rect 116276 306386 116344 306442
rect 116400 306386 119410 306442
rect 119466 306386 119534 306442
rect 119590 306386 122600 306442
rect 122656 306386 122724 306442
rect 122780 306386 390220 306442
rect 390276 306386 390344 306442
rect 390400 306386 393410 306442
rect 393466 306386 393534 306442
rect 393590 306386 396600 306442
rect 396656 306386 396724 306442
rect 396780 306386 490220 306442
rect 490276 306386 490344 306442
rect 490400 306386 493410 306442
rect 493466 306386 493534 306442
rect 493590 306386 496600 306442
rect 496656 306386 496724 306442
rect 496780 306386 634860 306442
rect 634916 306386 634984 306442
rect 635040 306386 638050 306442
rect 638106 306386 638174 306442
rect 638230 306386 641240 306442
rect 641296 306386 641364 306442
rect 641420 306386 698052 306442
rect 698108 306386 698176 306442
rect 698232 306386 698300 306442
rect 698356 306386 698424 306442
rect 698480 306386 698548 306442
rect 698604 306386 698672 306442
rect 698728 306386 698796 306442
rect 698852 306386 702624 306442
rect 79078 306382 702624 306386
rect 79078 306326 158178 306382
rect 158234 306326 158302 306382
rect 158358 306326 158426 306382
rect 158482 306326 158550 306382
rect 158606 306326 381310 306382
rect 381366 306326 381434 306382
rect 381490 306326 381558 306382
rect 381614 306326 381682 306382
rect 381738 306326 590910 306382
rect 590966 306326 591034 306382
rect 591090 306326 591158 306382
rect 591214 306326 591282 306382
rect 591338 306326 591406 306382
rect 591462 306326 591530 306382
rect 591586 306326 591654 306382
rect 591710 306326 702624 306382
rect 79078 306256 702624 306326
rect 77678 305786 700322 305856
rect 77678 305730 77808 305786
rect 77864 305730 77932 305786
rect 77988 305730 78056 305786
rect 78112 305730 78180 305786
rect 78236 305730 78304 305786
rect 78360 305730 78428 305786
rect 78484 305730 78552 305786
rect 78608 305730 114625 305786
rect 114681 305730 114749 305786
rect 114805 305730 117815 305786
rect 117871 305730 117939 305786
rect 117995 305730 121005 305786
rect 121061 305730 121129 305786
rect 121185 305730 124195 305786
rect 124251 305730 124319 305786
rect 124375 305730 388625 305786
rect 388681 305730 388749 305786
rect 388805 305730 391815 305786
rect 391871 305730 391939 305786
rect 391995 305730 395005 305786
rect 395061 305730 395129 305786
rect 395185 305730 398195 305786
rect 398251 305730 398319 305786
rect 398375 305730 488625 305786
rect 488681 305730 488749 305786
rect 488805 305730 491815 305786
rect 491871 305730 491939 305786
rect 491995 305730 495005 305786
rect 495061 305730 495129 305786
rect 495185 305730 498195 305786
rect 498251 305730 498319 305786
rect 498375 305730 633265 305786
rect 633321 305730 633389 305786
rect 633445 305730 636455 305786
rect 636511 305730 636579 305786
rect 636635 305730 639645 305786
rect 639701 305730 639769 305786
rect 639825 305730 642835 305786
rect 642891 305730 642959 305786
rect 643015 305730 699452 305786
rect 699508 305730 699576 305786
rect 699632 305730 699700 305786
rect 699756 305730 699824 305786
rect 699880 305730 699948 305786
rect 700004 305730 700072 305786
rect 700128 305730 700196 305786
rect 700252 305730 700322 305786
rect 77678 305726 700322 305730
rect 77678 305670 157158 305726
rect 157214 305670 157282 305726
rect 157338 305670 157406 305726
rect 157462 305670 157530 305726
rect 157586 305670 382330 305726
rect 382386 305670 382454 305726
rect 382510 305670 382578 305726
rect 382634 305670 382702 305726
rect 382758 305670 592310 305726
rect 592366 305670 592434 305726
rect 592490 305670 592558 305726
rect 592614 305670 592682 305726
rect 592738 305670 592806 305726
rect 592862 305670 592930 305726
rect 592986 305670 593054 305726
rect 593110 305670 700322 305726
rect 77678 305662 700322 305670
rect 77678 305606 77808 305662
rect 77864 305606 77932 305662
rect 77988 305606 78056 305662
rect 78112 305606 78180 305662
rect 78236 305606 78304 305662
rect 78360 305606 78428 305662
rect 78484 305606 78552 305662
rect 78608 305606 114625 305662
rect 114681 305606 114749 305662
rect 114805 305606 117815 305662
rect 117871 305606 117939 305662
rect 117995 305606 121005 305662
rect 121061 305606 121129 305662
rect 121185 305606 124195 305662
rect 124251 305606 124319 305662
rect 124375 305606 388625 305662
rect 388681 305606 388749 305662
rect 388805 305606 391815 305662
rect 391871 305606 391939 305662
rect 391995 305606 395005 305662
rect 395061 305606 395129 305662
rect 395185 305606 398195 305662
rect 398251 305606 398319 305662
rect 398375 305606 488625 305662
rect 488681 305606 488749 305662
rect 488805 305606 491815 305662
rect 491871 305606 491939 305662
rect 491995 305606 495005 305662
rect 495061 305606 495129 305662
rect 495185 305606 498195 305662
rect 498251 305606 498319 305662
rect 498375 305606 633265 305662
rect 633321 305606 633389 305662
rect 633445 305606 636455 305662
rect 636511 305606 636579 305662
rect 636635 305606 639645 305662
rect 639701 305606 639769 305662
rect 639825 305606 642835 305662
rect 642891 305606 642959 305662
rect 643015 305606 699452 305662
rect 699508 305606 699576 305662
rect 699632 305606 699700 305662
rect 699756 305606 699824 305662
rect 699880 305606 699948 305662
rect 700004 305606 700072 305662
rect 700128 305606 700196 305662
rect 700252 305606 700322 305662
rect 77678 305602 700322 305606
rect 77678 305546 157158 305602
rect 157214 305546 157282 305602
rect 157338 305546 157406 305602
rect 157462 305546 157530 305602
rect 157586 305546 382330 305602
rect 382386 305546 382454 305602
rect 382510 305546 382578 305602
rect 382634 305546 382702 305602
rect 382758 305546 592310 305602
rect 592366 305546 592434 305602
rect 592490 305546 592558 305602
rect 592614 305546 592682 305602
rect 592738 305546 592806 305602
rect 592862 305546 592930 305602
rect 592986 305546 593054 305602
rect 593110 305546 700322 305602
rect 77678 305538 700322 305546
rect 77678 305482 77808 305538
rect 77864 305482 77932 305538
rect 77988 305482 78056 305538
rect 78112 305482 78180 305538
rect 78236 305482 78304 305538
rect 78360 305482 78428 305538
rect 78484 305482 78552 305538
rect 78608 305482 114625 305538
rect 114681 305482 114749 305538
rect 114805 305482 117815 305538
rect 117871 305482 117939 305538
rect 117995 305482 121005 305538
rect 121061 305482 121129 305538
rect 121185 305482 124195 305538
rect 124251 305482 124319 305538
rect 124375 305482 388625 305538
rect 388681 305482 388749 305538
rect 388805 305482 391815 305538
rect 391871 305482 391939 305538
rect 391995 305482 395005 305538
rect 395061 305482 395129 305538
rect 395185 305482 398195 305538
rect 398251 305482 398319 305538
rect 398375 305482 488625 305538
rect 488681 305482 488749 305538
rect 488805 305482 491815 305538
rect 491871 305482 491939 305538
rect 491995 305482 495005 305538
rect 495061 305482 495129 305538
rect 495185 305482 498195 305538
rect 498251 305482 498319 305538
rect 498375 305482 633265 305538
rect 633321 305482 633389 305538
rect 633445 305482 636455 305538
rect 636511 305482 636579 305538
rect 636635 305482 639645 305538
rect 639701 305482 639769 305538
rect 639825 305482 642835 305538
rect 642891 305482 642959 305538
rect 643015 305482 699452 305538
rect 699508 305482 699576 305538
rect 699632 305482 699700 305538
rect 699756 305482 699824 305538
rect 699880 305482 699948 305538
rect 700004 305482 700072 305538
rect 700128 305482 700196 305538
rect 700252 305482 700322 305538
rect 77678 305478 700322 305482
rect 77678 305422 157158 305478
rect 157214 305422 157282 305478
rect 157338 305422 157406 305478
rect 157462 305422 157530 305478
rect 157586 305422 382330 305478
rect 382386 305422 382454 305478
rect 382510 305422 382578 305478
rect 382634 305422 382702 305478
rect 382758 305422 592310 305478
rect 592366 305422 592434 305478
rect 592490 305422 592558 305478
rect 592614 305422 592682 305478
rect 592738 305422 592806 305478
rect 592862 305422 592930 305478
rect 592986 305422 593054 305478
rect 593110 305422 700322 305478
rect 77678 305414 700322 305422
rect 77678 305358 77808 305414
rect 77864 305358 77932 305414
rect 77988 305358 78056 305414
rect 78112 305358 78180 305414
rect 78236 305358 78304 305414
rect 78360 305358 78428 305414
rect 78484 305358 78552 305414
rect 78608 305358 114625 305414
rect 114681 305358 114749 305414
rect 114805 305358 117815 305414
rect 117871 305358 117939 305414
rect 117995 305358 121005 305414
rect 121061 305358 121129 305414
rect 121185 305358 124195 305414
rect 124251 305358 124319 305414
rect 124375 305358 388625 305414
rect 388681 305358 388749 305414
rect 388805 305358 391815 305414
rect 391871 305358 391939 305414
rect 391995 305358 395005 305414
rect 395061 305358 395129 305414
rect 395185 305358 398195 305414
rect 398251 305358 398319 305414
rect 398375 305358 488625 305414
rect 488681 305358 488749 305414
rect 488805 305358 491815 305414
rect 491871 305358 491939 305414
rect 491995 305358 495005 305414
rect 495061 305358 495129 305414
rect 495185 305358 498195 305414
rect 498251 305358 498319 305414
rect 498375 305358 633265 305414
rect 633321 305358 633389 305414
rect 633445 305358 636455 305414
rect 636511 305358 636579 305414
rect 636635 305358 639645 305414
rect 639701 305358 639769 305414
rect 639825 305358 642835 305414
rect 642891 305358 642959 305414
rect 643015 305358 699452 305414
rect 699508 305358 699576 305414
rect 699632 305358 699700 305414
rect 699756 305358 699824 305414
rect 699880 305358 699948 305414
rect 700004 305358 700072 305414
rect 700128 305358 700196 305414
rect 700252 305358 700322 305414
rect 77678 305354 700322 305358
rect 77678 305298 157158 305354
rect 157214 305298 157282 305354
rect 157338 305298 157406 305354
rect 157462 305298 157530 305354
rect 157586 305298 382330 305354
rect 382386 305298 382454 305354
rect 382510 305298 382578 305354
rect 382634 305298 382702 305354
rect 382758 305298 592310 305354
rect 592366 305298 592434 305354
rect 592490 305298 592558 305354
rect 592614 305298 592682 305354
rect 592738 305298 592806 305354
rect 592862 305298 592930 305354
rect 592986 305298 593054 305354
rect 593110 305298 700322 305354
rect 77678 305290 700322 305298
rect 77678 305234 77808 305290
rect 77864 305234 77932 305290
rect 77988 305234 78056 305290
rect 78112 305234 78180 305290
rect 78236 305234 78304 305290
rect 78360 305234 78428 305290
rect 78484 305234 78552 305290
rect 78608 305234 114625 305290
rect 114681 305234 114749 305290
rect 114805 305234 117815 305290
rect 117871 305234 117939 305290
rect 117995 305234 121005 305290
rect 121061 305234 121129 305290
rect 121185 305234 124195 305290
rect 124251 305234 124319 305290
rect 124375 305234 388625 305290
rect 388681 305234 388749 305290
rect 388805 305234 391815 305290
rect 391871 305234 391939 305290
rect 391995 305234 395005 305290
rect 395061 305234 395129 305290
rect 395185 305234 398195 305290
rect 398251 305234 398319 305290
rect 398375 305234 488625 305290
rect 488681 305234 488749 305290
rect 488805 305234 491815 305290
rect 491871 305234 491939 305290
rect 491995 305234 495005 305290
rect 495061 305234 495129 305290
rect 495185 305234 498195 305290
rect 498251 305234 498319 305290
rect 498375 305234 633265 305290
rect 633321 305234 633389 305290
rect 633445 305234 636455 305290
rect 636511 305234 636579 305290
rect 636635 305234 639645 305290
rect 639701 305234 639769 305290
rect 639825 305234 642835 305290
rect 642891 305234 642959 305290
rect 643015 305234 699452 305290
rect 699508 305234 699576 305290
rect 699632 305234 699700 305290
rect 699756 305234 699824 305290
rect 699880 305234 699948 305290
rect 700004 305234 700072 305290
rect 700128 305234 700196 305290
rect 700252 305234 700322 305290
rect 77678 305230 700322 305234
rect 77678 305174 157158 305230
rect 157214 305174 157282 305230
rect 157338 305174 157406 305230
rect 157462 305174 157530 305230
rect 157586 305174 382330 305230
rect 382386 305174 382454 305230
rect 382510 305174 382578 305230
rect 382634 305174 382702 305230
rect 382758 305174 592310 305230
rect 592366 305174 592434 305230
rect 592490 305174 592558 305230
rect 592614 305174 592682 305230
rect 592738 305174 592806 305230
rect 592862 305174 592930 305230
rect 592986 305174 593054 305230
rect 593110 305174 700322 305230
rect 77678 305166 700322 305174
rect 77678 305110 77808 305166
rect 77864 305110 77932 305166
rect 77988 305110 78056 305166
rect 78112 305110 78180 305166
rect 78236 305110 78304 305166
rect 78360 305110 78428 305166
rect 78484 305110 78552 305166
rect 78608 305110 114625 305166
rect 114681 305110 114749 305166
rect 114805 305110 117815 305166
rect 117871 305110 117939 305166
rect 117995 305110 121005 305166
rect 121061 305110 121129 305166
rect 121185 305110 124195 305166
rect 124251 305110 124319 305166
rect 124375 305110 388625 305166
rect 388681 305110 388749 305166
rect 388805 305110 391815 305166
rect 391871 305110 391939 305166
rect 391995 305110 395005 305166
rect 395061 305110 395129 305166
rect 395185 305110 398195 305166
rect 398251 305110 398319 305166
rect 398375 305110 488625 305166
rect 488681 305110 488749 305166
rect 488805 305110 491815 305166
rect 491871 305110 491939 305166
rect 491995 305110 495005 305166
rect 495061 305110 495129 305166
rect 495185 305110 498195 305166
rect 498251 305110 498319 305166
rect 498375 305110 633265 305166
rect 633321 305110 633389 305166
rect 633445 305110 636455 305166
rect 636511 305110 636579 305166
rect 636635 305110 639645 305166
rect 639701 305110 639769 305166
rect 639825 305110 642835 305166
rect 642891 305110 642959 305166
rect 643015 305110 699452 305166
rect 699508 305110 699576 305166
rect 699632 305110 699700 305166
rect 699756 305110 699824 305166
rect 699880 305110 699948 305166
rect 700004 305110 700072 305166
rect 700128 305110 700196 305166
rect 700252 305110 700322 305166
rect 77678 305106 700322 305110
rect 77678 305050 157158 305106
rect 157214 305050 157282 305106
rect 157338 305050 157406 305106
rect 157462 305050 157530 305106
rect 157586 305050 382330 305106
rect 382386 305050 382454 305106
rect 382510 305050 382578 305106
rect 382634 305050 382702 305106
rect 382758 305050 592310 305106
rect 592366 305050 592434 305106
rect 592490 305050 592558 305106
rect 592614 305050 592682 305106
rect 592738 305050 592806 305106
rect 592862 305050 592930 305106
rect 592986 305050 593054 305106
rect 593110 305050 700322 305106
rect 77678 305042 700322 305050
rect 77678 304986 77808 305042
rect 77864 304986 77932 305042
rect 77988 304986 78056 305042
rect 78112 304986 78180 305042
rect 78236 304986 78304 305042
rect 78360 304986 78428 305042
rect 78484 304986 78552 305042
rect 78608 304986 114625 305042
rect 114681 304986 114749 305042
rect 114805 304986 117815 305042
rect 117871 304986 117939 305042
rect 117995 304986 121005 305042
rect 121061 304986 121129 305042
rect 121185 304986 124195 305042
rect 124251 304986 124319 305042
rect 124375 304986 388625 305042
rect 388681 304986 388749 305042
rect 388805 304986 391815 305042
rect 391871 304986 391939 305042
rect 391995 304986 395005 305042
rect 395061 304986 395129 305042
rect 395185 304986 398195 305042
rect 398251 304986 398319 305042
rect 398375 304986 488625 305042
rect 488681 304986 488749 305042
rect 488805 304986 491815 305042
rect 491871 304986 491939 305042
rect 491995 304986 495005 305042
rect 495061 304986 495129 305042
rect 495185 304986 498195 305042
rect 498251 304986 498319 305042
rect 498375 304986 633265 305042
rect 633321 304986 633389 305042
rect 633445 304986 636455 305042
rect 636511 304986 636579 305042
rect 636635 304986 639645 305042
rect 639701 304986 639769 305042
rect 639825 304986 642835 305042
rect 642891 304986 642959 305042
rect 643015 304986 699452 305042
rect 699508 304986 699576 305042
rect 699632 304986 699700 305042
rect 699756 304986 699824 305042
rect 699880 304986 699948 305042
rect 700004 304986 700072 305042
rect 700128 304986 700196 305042
rect 700252 304986 700322 305042
rect 77678 304982 700322 304986
rect 77678 304926 157158 304982
rect 157214 304926 157282 304982
rect 157338 304926 157406 304982
rect 157462 304926 157530 304982
rect 157586 304926 382330 304982
rect 382386 304926 382454 304982
rect 382510 304926 382578 304982
rect 382634 304926 382702 304982
rect 382758 304926 592310 304982
rect 592366 304926 592434 304982
rect 592490 304926 592558 304982
rect 592614 304926 592682 304982
rect 592738 304926 592806 304982
rect 592862 304926 592930 304982
rect 592986 304926 593054 304982
rect 593110 304926 700322 304982
rect 77678 304856 700322 304926
rect 75312 304122 78678 304244
rect 75312 304066 77800 304122
rect 77856 304066 78100 304122
rect 78156 304066 78400 304122
rect 78456 304066 78678 304122
rect 75312 303924 78678 304066
rect 75376 300622 80078 300744
rect 75376 300566 79300 300622
rect 79356 300566 79600 300622
rect 79656 300566 79900 300622
rect 79956 300566 80078 300622
rect 75376 300424 80078 300566
rect 75312 297102 78678 297244
rect 75312 297046 77900 297102
rect 77956 297046 78200 297102
rect 78256 297046 78500 297102
rect 78556 297046 78678 297102
rect 75312 296924 78678 297046
rect 699322 290423 701085 290490
rect 699322 290367 699497 290423
rect 699553 290367 699797 290423
rect 699853 290367 700097 290423
rect 700153 290367 701085 290423
rect 699322 290290 701085 290367
rect 76115 290048 80078 290110
rect 701565 290090 701885 290490
rect 76115 289992 79284 290048
rect 79340 289992 79584 290048
rect 79640 289992 79884 290048
rect 79940 289992 80078 290048
rect 76115 289910 80078 289992
rect 697922 290008 701885 290090
rect 697922 289952 698060 290008
rect 698116 289952 698360 290008
rect 698416 289952 698660 290008
rect 698716 289952 701885 290008
rect 76115 289510 76435 289910
rect 697922 289890 701885 289952
rect 76915 289633 78678 289710
rect 76915 289577 77847 289633
rect 77903 289577 78147 289633
rect 78203 289577 78447 289633
rect 78503 289577 78678 289633
rect 76915 289510 78678 289577
rect 666132 283925 698922 284067
rect 666132 283869 698044 283925
rect 698100 283869 698344 283925
rect 698400 283869 698644 283925
rect 698700 283869 698922 283925
rect 666132 283747 698922 283869
rect 79078 283372 591840 283442
rect 79078 283316 79208 283372
rect 79264 283316 79332 283372
rect 79388 283316 79456 283372
rect 79512 283316 79580 283372
rect 79636 283316 79704 283372
rect 79760 283316 79828 283372
rect 79884 283316 79952 283372
rect 80008 283316 590970 283372
rect 591026 283316 591094 283372
rect 591150 283316 591218 283372
rect 591274 283316 591342 283372
rect 591398 283316 591466 283372
rect 591522 283316 591590 283372
rect 591646 283316 591714 283372
rect 591770 283316 591840 283372
rect 79078 283312 591840 283316
rect 79078 283256 99294 283312
rect 99350 283256 99418 283312
rect 99474 283256 109294 283312
rect 109350 283256 109418 283312
rect 109474 283256 119294 283312
rect 119350 283256 119418 283312
rect 119474 283256 129294 283312
rect 129350 283256 129418 283312
rect 129474 283256 139294 283312
rect 139350 283256 139418 283312
rect 139474 283256 149294 283312
rect 149350 283256 149418 283312
rect 149474 283256 159294 283312
rect 159350 283256 159418 283312
rect 159474 283256 169294 283312
rect 169350 283256 169418 283312
rect 169474 283256 179294 283312
rect 179350 283256 179418 283312
rect 179474 283256 189294 283312
rect 189350 283256 189418 283312
rect 189474 283256 199294 283312
rect 199350 283256 199418 283312
rect 199474 283256 209294 283312
rect 209350 283256 209418 283312
rect 209474 283256 219294 283312
rect 219350 283256 219418 283312
rect 219474 283256 229294 283312
rect 229350 283256 229418 283312
rect 229474 283256 239294 283312
rect 239350 283256 239418 283312
rect 239474 283256 249294 283312
rect 249350 283256 249418 283312
rect 249474 283256 259294 283312
rect 259350 283256 259418 283312
rect 259474 283256 269294 283312
rect 269350 283256 269418 283312
rect 269474 283256 279294 283312
rect 279350 283256 279418 283312
rect 279474 283256 289294 283312
rect 289350 283256 289418 283312
rect 289474 283256 299294 283312
rect 299350 283256 299418 283312
rect 299474 283256 309294 283312
rect 309350 283256 309418 283312
rect 309474 283256 319294 283312
rect 319350 283256 319418 283312
rect 319474 283256 329294 283312
rect 329350 283256 329418 283312
rect 329474 283256 339294 283312
rect 339350 283256 339418 283312
rect 339474 283256 349294 283312
rect 349350 283256 349418 283312
rect 349474 283256 359294 283312
rect 359350 283256 359418 283312
rect 359474 283256 369294 283312
rect 369350 283256 369418 283312
rect 369474 283256 379294 283312
rect 379350 283256 379418 283312
rect 379474 283256 389294 283312
rect 389350 283256 389418 283312
rect 389474 283256 399294 283312
rect 399350 283256 399418 283312
rect 399474 283256 409294 283312
rect 409350 283256 409418 283312
rect 409474 283256 419294 283312
rect 419350 283256 419418 283312
rect 419474 283256 429294 283312
rect 429350 283256 429418 283312
rect 429474 283256 439294 283312
rect 439350 283256 439418 283312
rect 439474 283256 449294 283312
rect 449350 283256 449418 283312
rect 449474 283256 459294 283312
rect 459350 283256 459418 283312
rect 459474 283256 469294 283312
rect 469350 283256 469418 283312
rect 469474 283256 479294 283312
rect 479350 283256 479418 283312
rect 479474 283256 489294 283312
rect 489350 283256 489418 283312
rect 489474 283256 499294 283312
rect 499350 283256 499418 283312
rect 499474 283256 509294 283312
rect 509350 283256 509418 283312
rect 509474 283256 519294 283312
rect 519350 283256 519418 283312
rect 519474 283256 529294 283312
rect 529350 283256 529418 283312
rect 529474 283256 539294 283312
rect 539350 283256 539418 283312
rect 539474 283256 549294 283312
rect 549350 283256 549418 283312
rect 549474 283256 591840 283312
rect 79078 283248 591840 283256
rect 79078 283192 79208 283248
rect 79264 283192 79332 283248
rect 79388 283192 79456 283248
rect 79512 283192 79580 283248
rect 79636 283192 79704 283248
rect 79760 283192 79828 283248
rect 79884 283192 79952 283248
rect 80008 283192 590970 283248
rect 591026 283192 591094 283248
rect 591150 283192 591218 283248
rect 591274 283192 591342 283248
rect 591398 283192 591466 283248
rect 591522 283192 591590 283248
rect 591646 283192 591714 283248
rect 591770 283192 591840 283248
rect 79078 283188 591840 283192
rect 79078 283132 99294 283188
rect 99350 283132 99418 283188
rect 99474 283132 109294 283188
rect 109350 283132 109418 283188
rect 109474 283132 119294 283188
rect 119350 283132 119418 283188
rect 119474 283132 129294 283188
rect 129350 283132 129418 283188
rect 129474 283132 139294 283188
rect 139350 283132 139418 283188
rect 139474 283132 149294 283188
rect 149350 283132 149418 283188
rect 149474 283132 159294 283188
rect 159350 283132 159418 283188
rect 159474 283132 169294 283188
rect 169350 283132 169418 283188
rect 169474 283132 179294 283188
rect 179350 283132 179418 283188
rect 179474 283132 189294 283188
rect 189350 283132 189418 283188
rect 189474 283132 199294 283188
rect 199350 283132 199418 283188
rect 199474 283132 209294 283188
rect 209350 283132 209418 283188
rect 209474 283132 219294 283188
rect 219350 283132 219418 283188
rect 219474 283132 229294 283188
rect 229350 283132 229418 283188
rect 229474 283132 239294 283188
rect 239350 283132 239418 283188
rect 239474 283132 249294 283188
rect 249350 283132 249418 283188
rect 249474 283132 259294 283188
rect 259350 283132 259418 283188
rect 259474 283132 269294 283188
rect 269350 283132 269418 283188
rect 269474 283132 279294 283188
rect 279350 283132 279418 283188
rect 279474 283132 289294 283188
rect 289350 283132 289418 283188
rect 289474 283132 299294 283188
rect 299350 283132 299418 283188
rect 299474 283132 309294 283188
rect 309350 283132 309418 283188
rect 309474 283132 319294 283188
rect 319350 283132 319418 283188
rect 319474 283132 329294 283188
rect 329350 283132 329418 283188
rect 329474 283132 339294 283188
rect 339350 283132 339418 283188
rect 339474 283132 349294 283188
rect 349350 283132 349418 283188
rect 349474 283132 359294 283188
rect 359350 283132 359418 283188
rect 359474 283132 369294 283188
rect 369350 283132 369418 283188
rect 369474 283132 379294 283188
rect 379350 283132 379418 283188
rect 379474 283132 389294 283188
rect 389350 283132 389418 283188
rect 389474 283132 399294 283188
rect 399350 283132 399418 283188
rect 399474 283132 409294 283188
rect 409350 283132 409418 283188
rect 409474 283132 419294 283188
rect 419350 283132 419418 283188
rect 419474 283132 429294 283188
rect 429350 283132 429418 283188
rect 429474 283132 439294 283188
rect 439350 283132 439418 283188
rect 439474 283132 449294 283188
rect 449350 283132 449418 283188
rect 449474 283132 459294 283188
rect 459350 283132 459418 283188
rect 459474 283132 469294 283188
rect 469350 283132 469418 283188
rect 469474 283132 479294 283188
rect 479350 283132 479418 283188
rect 479474 283132 489294 283188
rect 489350 283132 489418 283188
rect 489474 283132 499294 283188
rect 499350 283132 499418 283188
rect 499474 283132 509294 283188
rect 509350 283132 509418 283188
rect 509474 283132 519294 283188
rect 519350 283132 519418 283188
rect 519474 283132 529294 283188
rect 529350 283132 529418 283188
rect 529474 283132 539294 283188
rect 539350 283132 539418 283188
rect 539474 283132 549294 283188
rect 549350 283132 549418 283188
rect 549474 283132 591840 283188
rect 79078 283124 591840 283132
rect 79078 283068 79208 283124
rect 79264 283068 79332 283124
rect 79388 283068 79456 283124
rect 79512 283068 79580 283124
rect 79636 283068 79704 283124
rect 79760 283068 79828 283124
rect 79884 283068 79952 283124
rect 80008 283068 590970 283124
rect 591026 283068 591094 283124
rect 591150 283068 591218 283124
rect 591274 283068 591342 283124
rect 591398 283068 591466 283124
rect 591522 283068 591590 283124
rect 591646 283068 591714 283124
rect 591770 283068 591840 283124
rect 79078 283064 591840 283068
rect 79078 283008 99294 283064
rect 99350 283008 99418 283064
rect 99474 283008 109294 283064
rect 109350 283008 109418 283064
rect 109474 283008 119294 283064
rect 119350 283008 119418 283064
rect 119474 283008 129294 283064
rect 129350 283008 129418 283064
rect 129474 283008 139294 283064
rect 139350 283008 139418 283064
rect 139474 283008 149294 283064
rect 149350 283008 149418 283064
rect 149474 283008 159294 283064
rect 159350 283008 159418 283064
rect 159474 283008 169294 283064
rect 169350 283008 169418 283064
rect 169474 283008 179294 283064
rect 179350 283008 179418 283064
rect 179474 283008 189294 283064
rect 189350 283008 189418 283064
rect 189474 283008 199294 283064
rect 199350 283008 199418 283064
rect 199474 283008 209294 283064
rect 209350 283008 209418 283064
rect 209474 283008 219294 283064
rect 219350 283008 219418 283064
rect 219474 283008 229294 283064
rect 229350 283008 229418 283064
rect 229474 283008 239294 283064
rect 239350 283008 239418 283064
rect 239474 283008 249294 283064
rect 249350 283008 249418 283064
rect 249474 283008 259294 283064
rect 259350 283008 259418 283064
rect 259474 283008 269294 283064
rect 269350 283008 269418 283064
rect 269474 283008 279294 283064
rect 279350 283008 279418 283064
rect 279474 283008 289294 283064
rect 289350 283008 289418 283064
rect 289474 283008 299294 283064
rect 299350 283008 299418 283064
rect 299474 283008 309294 283064
rect 309350 283008 309418 283064
rect 309474 283008 319294 283064
rect 319350 283008 319418 283064
rect 319474 283008 329294 283064
rect 329350 283008 329418 283064
rect 329474 283008 339294 283064
rect 339350 283008 339418 283064
rect 339474 283008 349294 283064
rect 349350 283008 349418 283064
rect 349474 283008 359294 283064
rect 359350 283008 359418 283064
rect 359474 283008 369294 283064
rect 369350 283008 369418 283064
rect 369474 283008 379294 283064
rect 379350 283008 379418 283064
rect 379474 283008 389294 283064
rect 389350 283008 389418 283064
rect 389474 283008 399294 283064
rect 399350 283008 399418 283064
rect 399474 283008 409294 283064
rect 409350 283008 409418 283064
rect 409474 283008 419294 283064
rect 419350 283008 419418 283064
rect 419474 283008 429294 283064
rect 429350 283008 429418 283064
rect 429474 283008 439294 283064
rect 439350 283008 439418 283064
rect 439474 283008 449294 283064
rect 449350 283008 449418 283064
rect 449474 283008 459294 283064
rect 459350 283008 459418 283064
rect 459474 283008 469294 283064
rect 469350 283008 469418 283064
rect 469474 283008 479294 283064
rect 479350 283008 479418 283064
rect 479474 283008 489294 283064
rect 489350 283008 489418 283064
rect 489474 283008 499294 283064
rect 499350 283008 499418 283064
rect 499474 283008 509294 283064
rect 509350 283008 509418 283064
rect 509474 283008 519294 283064
rect 519350 283008 519418 283064
rect 519474 283008 529294 283064
rect 529350 283008 529418 283064
rect 529474 283008 539294 283064
rect 539350 283008 539418 283064
rect 539474 283008 549294 283064
rect 549350 283008 549418 283064
rect 549474 283008 591840 283064
rect 79078 283000 591840 283008
rect 79078 282944 79208 283000
rect 79264 282944 79332 283000
rect 79388 282944 79456 283000
rect 79512 282944 79580 283000
rect 79636 282944 79704 283000
rect 79760 282944 79828 283000
rect 79884 282944 79952 283000
rect 80008 282944 590970 283000
rect 591026 282944 591094 283000
rect 591150 282944 591218 283000
rect 591274 282944 591342 283000
rect 591398 282944 591466 283000
rect 591522 282944 591590 283000
rect 591646 282944 591714 283000
rect 591770 282944 591840 283000
rect 79078 282940 591840 282944
rect 79078 282884 99294 282940
rect 99350 282884 99418 282940
rect 99474 282884 109294 282940
rect 109350 282884 109418 282940
rect 109474 282884 119294 282940
rect 119350 282884 119418 282940
rect 119474 282884 129294 282940
rect 129350 282884 129418 282940
rect 129474 282884 139294 282940
rect 139350 282884 139418 282940
rect 139474 282884 149294 282940
rect 149350 282884 149418 282940
rect 149474 282884 159294 282940
rect 159350 282884 159418 282940
rect 159474 282884 169294 282940
rect 169350 282884 169418 282940
rect 169474 282884 179294 282940
rect 179350 282884 179418 282940
rect 179474 282884 189294 282940
rect 189350 282884 189418 282940
rect 189474 282884 199294 282940
rect 199350 282884 199418 282940
rect 199474 282884 209294 282940
rect 209350 282884 209418 282940
rect 209474 282884 219294 282940
rect 219350 282884 219418 282940
rect 219474 282884 229294 282940
rect 229350 282884 229418 282940
rect 229474 282884 239294 282940
rect 239350 282884 239418 282940
rect 239474 282884 249294 282940
rect 249350 282884 249418 282940
rect 249474 282884 259294 282940
rect 259350 282884 259418 282940
rect 259474 282884 269294 282940
rect 269350 282884 269418 282940
rect 269474 282884 279294 282940
rect 279350 282884 279418 282940
rect 279474 282884 289294 282940
rect 289350 282884 289418 282940
rect 289474 282884 299294 282940
rect 299350 282884 299418 282940
rect 299474 282884 309294 282940
rect 309350 282884 309418 282940
rect 309474 282884 319294 282940
rect 319350 282884 319418 282940
rect 319474 282884 329294 282940
rect 329350 282884 329418 282940
rect 329474 282884 339294 282940
rect 339350 282884 339418 282940
rect 339474 282884 349294 282940
rect 349350 282884 349418 282940
rect 349474 282884 359294 282940
rect 359350 282884 359418 282940
rect 359474 282884 369294 282940
rect 369350 282884 369418 282940
rect 369474 282884 379294 282940
rect 379350 282884 379418 282940
rect 379474 282884 389294 282940
rect 389350 282884 389418 282940
rect 389474 282884 399294 282940
rect 399350 282884 399418 282940
rect 399474 282884 409294 282940
rect 409350 282884 409418 282940
rect 409474 282884 419294 282940
rect 419350 282884 419418 282940
rect 419474 282884 429294 282940
rect 429350 282884 429418 282940
rect 429474 282884 439294 282940
rect 439350 282884 439418 282940
rect 439474 282884 449294 282940
rect 449350 282884 449418 282940
rect 449474 282884 459294 282940
rect 459350 282884 459418 282940
rect 459474 282884 469294 282940
rect 469350 282884 469418 282940
rect 469474 282884 479294 282940
rect 479350 282884 479418 282940
rect 479474 282884 489294 282940
rect 489350 282884 489418 282940
rect 489474 282884 499294 282940
rect 499350 282884 499418 282940
rect 499474 282884 509294 282940
rect 509350 282884 509418 282940
rect 509474 282884 519294 282940
rect 519350 282884 519418 282940
rect 519474 282884 529294 282940
rect 529350 282884 529418 282940
rect 529474 282884 539294 282940
rect 539350 282884 539418 282940
rect 539474 282884 549294 282940
rect 549350 282884 549418 282940
rect 549474 282884 591840 282940
rect 79078 282876 591840 282884
rect 79078 282820 79208 282876
rect 79264 282820 79332 282876
rect 79388 282820 79456 282876
rect 79512 282820 79580 282876
rect 79636 282820 79704 282876
rect 79760 282820 79828 282876
rect 79884 282820 79952 282876
rect 80008 282820 590970 282876
rect 591026 282820 591094 282876
rect 591150 282820 591218 282876
rect 591274 282820 591342 282876
rect 591398 282820 591466 282876
rect 591522 282820 591590 282876
rect 591646 282820 591714 282876
rect 591770 282820 591840 282876
rect 79078 282816 591840 282820
rect 79078 282760 99294 282816
rect 99350 282760 99418 282816
rect 99474 282760 109294 282816
rect 109350 282760 109418 282816
rect 109474 282760 119294 282816
rect 119350 282760 119418 282816
rect 119474 282760 129294 282816
rect 129350 282760 129418 282816
rect 129474 282760 139294 282816
rect 139350 282760 139418 282816
rect 139474 282760 149294 282816
rect 149350 282760 149418 282816
rect 149474 282760 159294 282816
rect 159350 282760 159418 282816
rect 159474 282760 169294 282816
rect 169350 282760 169418 282816
rect 169474 282760 179294 282816
rect 179350 282760 179418 282816
rect 179474 282760 189294 282816
rect 189350 282760 189418 282816
rect 189474 282760 199294 282816
rect 199350 282760 199418 282816
rect 199474 282760 209294 282816
rect 209350 282760 209418 282816
rect 209474 282760 219294 282816
rect 219350 282760 219418 282816
rect 219474 282760 229294 282816
rect 229350 282760 229418 282816
rect 229474 282760 239294 282816
rect 239350 282760 239418 282816
rect 239474 282760 249294 282816
rect 249350 282760 249418 282816
rect 249474 282760 259294 282816
rect 259350 282760 259418 282816
rect 259474 282760 269294 282816
rect 269350 282760 269418 282816
rect 269474 282760 279294 282816
rect 279350 282760 279418 282816
rect 279474 282760 289294 282816
rect 289350 282760 289418 282816
rect 289474 282760 299294 282816
rect 299350 282760 299418 282816
rect 299474 282760 309294 282816
rect 309350 282760 309418 282816
rect 309474 282760 319294 282816
rect 319350 282760 319418 282816
rect 319474 282760 329294 282816
rect 329350 282760 329418 282816
rect 329474 282760 339294 282816
rect 339350 282760 339418 282816
rect 339474 282760 349294 282816
rect 349350 282760 349418 282816
rect 349474 282760 359294 282816
rect 359350 282760 359418 282816
rect 359474 282760 369294 282816
rect 369350 282760 369418 282816
rect 369474 282760 379294 282816
rect 379350 282760 379418 282816
rect 379474 282760 389294 282816
rect 389350 282760 389418 282816
rect 389474 282760 399294 282816
rect 399350 282760 399418 282816
rect 399474 282760 409294 282816
rect 409350 282760 409418 282816
rect 409474 282760 419294 282816
rect 419350 282760 419418 282816
rect 419474 282760 429294 282816
rect 429350 282760 429418 282816
rect 429474 282760 439294 282816
rect 439350 282760 439418 282816
rect 439474 282760 449294 282816
rect 449350 282760 449418 282816
rect 449474 282760 459294 282816
rect 459350 282760 459418 282816
rect 459474 282760 469294 282816
rect 469350 282760 469418 282816
rect 469474 282760 479294 282816
rect 479350 282760 479418 282816
rect 479474 282760 489294 282816
rect 489350 282760 489418 282816
rect 489474 282760 499294 282816
rect 499350 282760 499418 282816
rect 499474 282760 509294 282816
rect 509350 282760 509418 282816
rect 509474 282760 519294 282816
rect 519350 282760 519418 282816
rect 519474 282760 529294 282816
rect 529350 282760 529418 282816
rect 529474 282760 539294 282816
rect 539350 282760 539418 282816
rect 539474 282760 549294 282816
rect 549350 282760 549418 282816
rect 549474 282760 591840 282816
rect 79078 282752 591840 282760
rect 79078 282696 79208 282752
rect 79264 282696 79332 282752
rect 79388 282696 79456 282752
rect 79512 282696 79580 282752
rect 79636 282696 79704 282752
rect 79760 282696 79828 282752
rect 79884 282696 79952 282752
rect 80008 282696 590970 282752
rect 591026 282696 591094 282752
rect 591150 282696 591218 282752
rect 591274 282696 591342 282752
rect 591398 282696 591466 282752
rect 591522 282696 591590 282752
rect 591646 282696 591714 282752
rect 591770 282696 591840 282752
rect 79078 282692 591840 282696
rect 79078 282636 99294 282692
rect 99350 282636 99418 282692
rect 99474 282636 109294 282692
rect 109350 282636 109418 282692
rect 109474 282636 119294 282692
rect 119350 282636 119418 282692
rect 119474 282636 129294 282692
rect 129350 282636 129418 282692
rect 129474 282636 139294 282692
rect 139350 282636 139418 282692
rect 139474 282636 149294 282692
rect 149350 282636 149418 282692
rect 149474 282636 159294 282692
rect 159350 282636 159418 282692
rect 159474 282636 169294 282692
rect 169350 282636 169418 282692
rect 169474 282636 179294 282692
rect 179350 282636 179418 282692
rect 179474 282636 189294 282692
rect 189350 282636 189418 282692
rect 189474 282636 199294 282692
rect 199350 282636 199418 282692
rect 199474 282636 209294 282692
rect 209350 282636 209418 282692
rect 209474 282636 219294 282692
rect 219350 282636 219418 282692
rect 219474 282636 229294 282692
rect 229350 282636 229418 282692
rect 229474 282636 239294 282692
rect 239350 282636 239418 282692
rect 239474 282636 249294 282692
rect 249350 282636 249418 282692
rect 249474 282636 259294 282692
rect 259350 282636 259418 282692
rect 259474 282636 269294 282692
rect 269350 282636 269418 282692
rect 269474 282636 279294 282692
rect 279350 282636 279418 282692
rect 279474 282636 289294 282692
rect 289350 282636 289418 282692
rect 289474 282636 299294 282692
rect 299350 282636 299418 282692
rect 299474 282636 309294 282692
rect 309350 282636 309418 282692
rect 309474 282636 319294 282692
rect 319350 282636 319418 282692
rect 319474 282636 329294 282692
rect 329350 282636 329418 282692
rect 329474 282636 339294 282692
rect 339350 282636 339418 282692
rect 339474 282636 349294 282692
rect 349350 282636 349418 282692
rect 349474 282636 359294 282692
rect 359350 282636 359418 282692
rect 359474 282636 369294 282692
rect 369350 282636 369418 282692
rect 369474 282636 379294 282692
rect 379350 282636 379418 282692
rect 379474 282636 389294 282692
rect 389350 282636 389418 282692
rect 389474 282636 399294 282692
rect 399350 282636 399418 282692
rect 399474 282636 409294 282692
rect 409350 282636 409418 282692
rect 409474 282636 419294 282692
rect 419350 282636 419418 282692
rect 419474 282636 429294 282692
rect 429350 282636 429418 282692
rect 429474 282636 439294 282692
rect 439350 282636 439418 282692
rect 439474 282636 449294 282692
rect 449350 282636 449418 282692
rect 449474 282636 459294 282692
rect 459350 282636 459418 282692
rect 459474 282636 469294 282692
rect 469350 282636 469418 282692
rect 469474 282636 479294 282692
rect 479350 282636 479418 282692
rect 479474 282636 489294 282692
rect 489350 282636 489418 282692
rect 489474 282636 499294 282692
rect 499350 282636 499418 282692
rect 499474 282636 509294 282692
rect 509350 282636 509418 282692
rect 509474 282636 519294 282692
rect 519350 282636 519418 282692
rect 519474 282636 529294 282692
rect 529350 282636 529418 282692
rect 529474 282636 539294 282692
rect 539350 282636 539418 282692
rect 539474 282636 549294 282692
rect 549350 282636 549418 282692
rect 549474 282636 591840 282692
rect 79078 282628 591840 282636
rect 79078 282572 79208 282628
rect 79264 282572 79332 282628
rect 79388 282572 79456 282628
rect 79512 282572 79580 282628
rect 79636 282572 79704 282628
rect 79760 282572 79828 282628
rect 79884 282572 79952 282628
rect 80008 282572 590970 282628
rect 591026 282572 591094 282628
rect 591150 282572 591218 282628
rect 591274 282572 591342 282628
rect 591398 282572 591466 282628
rect 591522 282572 591590 282628
rect 591646 282572 591714 282628
rect 591770 282572 591840 282628
rect 79078 282568 591840 282572
rect 79078 282512 99294 282568
rect 99350 282512 99418 282568
rect 99474 282512 109294 282568
rect 109350 282512 109418 282568
rect 109474 282512 119294 282568
rect 119350 282512 119418 282568
rect 119474 282512 129294 282568
rect 129350 282512 129418 282568
rect 129474 282512 139294 282568
rect 139350 282512 139418 282568
rect 139474 282512 149294 282568
rect 149350 282512 149418 282568
rect 149474 282512 159294 282568
rect 159350 282512 159418 282568
rect 159474 282512 169294 282568
rect 169350 282512 169418 282568
rect 169474 282512 179294 282568
rect 179350 282512 179418 282568
rect 179474 282512 189294 282568
rect 189350 282512 189418 282568
rect 189474 282512 199294 282568
rect 199350 282512 199418 282568
rect 199474 282512 209294 282568
rect 209350 282512 209418 282568
rect 209474 282512 219294 282568
rect 219350 282512 219418 282568
rect 219474 282512 229294 282568
rect 229350 282512 229418 282568
rect 229474 282512 239294 282568
rect 239350 282512 239418 282568
rect 239474 282512 249294 282568
rect 249350 282512 249418 282568
rect 249474 282512 259294 282568
rect 259350 282512 259418 282568
rect 259474 282512 269294 282568
rect 269350 282512 269418 282568
rect 269474 282512 279294 282568
rect 279350 282512 279418 282568
rect 279474 282512 289294 282568
rect 289350 282512 289418 282568
rect 289474 282512 299294 282568
rect 299350 282512 299418 282568
rect 299474 282512 309294 282568
rect 309350 282512 309418 282568
rect 309474 282512 319294 282568
rect 319350 282512 319418 282568
rect 319474 282512 329294 282568
rect 329350 282512 329418 282568
rect 329474 282512 339294 282568
rect 339350 282512 339418 282568
rect 339474 282512 349294 282568
rect 349350 282512 349418 282568
rect 349474 282512 359294 282568
rect 359350 282512 359418 282568
rect 359474 282512 369294 282568
rect 369350 282512 369418 282568
rect 369474 282512 379294 282568
rect 379350 282512 379418 282568
rect 379474 282512 389294 282568
rect 389350 282512 389418 282568
rect 389474 282512 399294 282568
rect 399350 282512 399418 282568
rect 399474 282512 409294 282568
rect 409350 282512 409418 282568
rect 409474 282512 419294 282568
rect 419350 282512 419418 282568
rect 419474 282512 429294 282568
rect 429350 282512 429418 282568
rect 429474 282512 439294 282568
rect 439350 282512 439418 282568
rect 439474 282512 449294 282568
rect 449350 282512 449418 282568
rect 449474 282512 459294 282568
rect 459350 282512 459418 282568
rect 459474 282512 469294 282568
rect 469350 282512 469418 282568
rect 469474 282512 479294 282568
rect 479350 282512 479418 282568
rect 479474 282512 489294 282568
rect 489350 282512 489418 282568
rect 489474 282512 499294 282568
rect 499350 282512 499418 282568
rect 499474 282512 509294 282568
rect 509350 282512 509418 282568
rect 509474 282512 519294 282568
rect 519350 282512 519418 282568
rect 519474 282512 529294 282568
rect 529350 282512 529418 282568
rect 529474 282512 539294 282568
rect 539350 282512 539418 282568
rect 539474 282512 549294 282568
rect 549350 282512 549418 282568
rect 549474 282512 591840 282568
rect 79078 282442 591840 282512
rect 77678 281972 593240 282042
rect 77678 281916 77808 281972
rect 77864 281916 77932 281972
rect 77988 281916 78056 281972
rect 78112 281916 78180 281972
rect 78236 281916 78304 281972
rect 78360 281916 78428 281972
rect 78484 281916 78552 281972
rect 78608 281916 592370 281972
rect 592426 281916 592494 281972
rect 592550 281916 592618 281972
rect 592674 281916 592742 281972
rect 592798 281916 592866 281972
rect 592922 281916 592990 281972
rect 593046 281916 593114 281972
rect 593170 281916 593240 281972
rect 77678 281912 593240 281916
rect 77678 281856 94294 281912
rect 94350 281856 94418 281912
rect 94474 281856 104294 281912
rect 104350 281856 104418 281912
rect 104474 281856 114294 281912
rect 114350 281856 114418 281912
rect 114474 281856 124294 281912
rect 124350 281856 124418 281912
rect 124474 281856 134294 281912
rect 134350 281856 134418 281912
rect 134474 281856 144294 281912
rect 144350 281856 144418 281912
rect 144474 281856 154294 281912
rect 154350 281856 154418 281912
rect 154474 281856 164294 281912
rect 164350 281856 164418 281912
rect 164474 281856 174294 281912
rect 174350 281856 174418 281912
rect 174474 281856 184294 281912
rect 184350 281856 184418 281912
rect 184474 281856 194294 281912
rect 194350 281856 194418 281912
rect 194474 281856 204294 281912
rect 204350 281856 204418 281912
rect 204474 281856 214294 281912
rect 214350 281856 214418 281912
rect 214474 281856 224294 281912
rect 224350 281856 224418 281912
rect 224474 281856 234294 281912
rect 234350 281856 234418 281912
rect 234474 281856 244294 281912
rect 244350 281856 244418 281912
rect 244474 281856 254294 281912
rect 254350 281856 254418 281912
rect 254474 281856 264294 281912
rect 264350 281856 264418 281912
rect 264474 281856 274294 281912
rect 274350 281856 274418 281912
rect 274474 281856 284294 281912
rect 284350 281856 284418 281912
rect 284474 281856 294294 281912
rect 294350 281856 294418 281912
rect 294474 281856 304294 281912
rect 304350 281856 304418 281912
rect 304474 281856 314294 281912
rect 314350 281856 314418 281912
rect 314474 281856 324294 281912
rect 324350 281856 324418 281912
rect 324474 281856 334294 281912
rect 334350 281856 334418 281912
rect 334474 281856 344294 281912
rect 344350 281856 344418 281912
rect 344474 281856 354294 281912
rect 354350 281856 354418 281912
rect 354474 281856 364294 281912
rect 364350 281856 364418 281912
rect 364474 281856 374294 281912
rect 374350 281856 374418 281912
rect 374474 281856 384294 281912
rect 384350 281856 384418 281912
rect 384474 281856 394294 281912
rect 394350 281856 394418 281912
rect 394474 281856 404294 281912
rect 404350 281856 404418 281912
rect 404474 281856 414294 281912
rect 414350 281856 414418 281912
rect 414474 281856 424294 281912
rect 424350 281856 424418 281912
rect 424474 281856 434294 281912
rect 434350 281856 434418 281912
rect 434474 281856 444294 281912
rect 444350 281856 444418 281912
rect 444474 281856 454294 281912
rect 454350 281856 454418 281912
rect 454474 281856 464294 281912
rect 464350 281856 464418 281912
rect 464474 281856 474294 281912
rect 474350 281856 474418 281912
rect 474474 281856 484294 281912
rect 484350 281856 484418 281912
rect 484474 281856 494294 281912
rect 494350 281856 494418 281912
rect 494474 281856 504294 281912
rect 504350 281856 504418 281912
rect 504474 281856 514294 281912
rect 514350 281856 514418 281912
rect 514474 281856 524294 281912
rect 524350 281856 524418 281912
rect 524474 281856 534294 281912
rect 534350 281856 534418 281912
rect 534474 281856 544294 281912
rect 544350 281856 544418 281912
rect 544474 281856 554294 281912
rect 554350 281856 554418 281912
rect 554474 281856 593240 281912
rect 77678 281848 593240 281856
rect 77678 281792 77808 281848
rect 77864 281792 77932 281848
rect 77988 281792 78056 281848
rect 78112 281792 78180 281848
rect 78236 281792 78304 281848
rect 78360 281792 78428 281848
rect 78484 281792 78552 281848
rect 78608 281792 592370 281848
rect 592426 281792 592494 281848
rect 592550 281792 592618 281848
rect 592674 281792 592742 281848
rect 592798 281792 592866 281848
rect 592922 281792 592990 281848
rect 593046 281792 593114 281848
rect 593170 281792 593240 281848
rect 77678 281788 593240 281792
rect 77678 281732 94294 281788
rect 94350 281732 94418 281788
rect 94474 281732 104294 281788
rect 104350 281732 104418 281788
rect 104474 281732 114294 281788
rect 114350 281732 114418 281788
rect 114474 281732 124294 281788
rect 124350 281732 124418 281788
rect 124474 281732 134294 281788
rect 134350 281732 134418 281788
rect 134474 281732 144294 281788
rect 144350 281732 144418 281788
rect 144474 281732 154294 281788
rect 154350 281732 154418 281788
rect 154474 281732 164294 281788
rect 164350 281732 164418 281788
rect 164474 281732 174294 281788
rect 174350 281732 174418 281788
rect 174474 281732 184294 281788
rect 184350 281732 184418 281788
rect 184474 281732 194294 281788
rect 194350 281732 194418 281788
rect 194474 281732 204294 281788
rect 204350 281732 204418 281788
rect 204474 281732 214294 281788
rect 214350 281732 214418 281788
rect 214474 281732 224294 281788
rect 224350 281732 224418 281788
rect 224474 281732 234294 281788
rect 234350 281732 234418 281788
rect 234474 281732 244294 281788
rect 244350 281732 244418 281788
rect 244474 281732 254294 281788
rect 254350 281732 254418 281788
rect 254474 281732 264294 281788
rect 264350 281732 264418 281788
rect 264474 281732 274294 281788
rect 274350 281732 274418 281788
rect 274474 281732 284294 281788
rect 284350 281732 284418 281788
rect 284474 281732 294294 281788
rect 294350 281732 294418 281788
rect 294474 281732 304294 281788
rect 304350 281732 304418 281788
rect 304474 281732 314294 281788
rect 314350 281732 314418 281788
rect 314474 281732 324294 281788
rect 324350 281732 324418 281788
rect 324474 281732 334294 281788
rect 334350 281732 334418 281788
rect 334474 281732 344294 281788
rect 344350 281732 344418 281788
rect 344474 281732 354294 281788
rect 354350 281732 354418 281788
rect 354474 281732 364294 281788
rect 364350 281732 364418 281788
rect 364474 281732 374294 281788
rect 374350 281732 374418 281788
rect 374474 281732 384294 281788
rect 384350 281732 384418 281788
rect 384474 281732 394294 281788
rect 394350 281732 394418 281788
rect 394474 281732 404294 281788
rect 404350 281732 404418 281788
rect 404474 281732 414294 281788
rect 414350 281732 414418 281788
rect 414474 281732 424294 281788
rect 424350 281732 424418 281788
rect 424474 281732 434294 281788
rect 434350 281732 434418 281788
rect 434474 281732 444294 281788
rect 444350 281732 444418 281788
rect 444474 281732 454294 281788
rect 454350 281732 454418 281788
rect 454474 281732 464294 281788
rect 464350 281732 464418 281788
rect 464474 281732 474294 281788
rect 474350 281732 474418 281788
rect 474474 281732 484294 281788
rect 484350 281732 484418 281788
rect 484474 281732 494294 281788
rect 494350 281732 494418 281788
rect 494474 281732 504294 281788
rect 504350 281732 504418 281788
rect 504474 281732 514294 281788
rect 514350 281732 514418 281788
rect 514474 281732 524294 281788
rect 524350 281732 524418 281788
rect 524474 281732 534294 281788
rect 534350 281732 534418 281788
rect 534474 281732 544294 281788
rect 544350 281732 544418 281788
rect 544474 281732 554294 281788
rect 554350 281732 554418 281788
rect 554474 281732 593240 281788
rect 77678 281724 593240 281732
rect 77678 281668 77808 281724
rect 77864 281668 77932 281724
rect 77988 281668 78056 281724
rect 78112 281668 78180 281724
rect 78236 281668 78304 281724
rect 78360 281668 78428 281724
rect 78484 281668 78552 281724
rect 78608 281668 592370 281724
rect 592426 281668 592494 281724
rect 592550 281668 592618 281724
rect 592674 281668 592742 281724
rect 592798 281668 592866 281724
rect 592922 281668 592990 281724
rect 593046 281668 593114 281724
rect 593170 281668 593240 281724
rect 77678 281664 593240 281668
rect 77678 281608 94294 281664
rect 94350 281608 94418 281664
rect 94474 281608 104294 281664
rect 104350 281608 104418 281664
rect 104474 281608 114294 281664
rect 114350 281608 114418 281664
rect 114474 281608 124294 281664
rect 124350 281608 124418 281664
rect 124474 281608 134294 281664
rect 134350 281608 134418 281664
rect 134474 281608 144294 281664
rect 144350 281608 144418 281664
rect 144474 281608 154294 281664
rect 154350 281608 154418 281664
rect 154474 281608 164294 281664
rect 164350 281608 164418 281664
rect 164474 281608 174294 281664
rect 174350 281608 174418 281664
rect 174474 281608 184294 281664
rect 184350 281608 184418 281664
rect 184474 281608 194294 281664
rect 194350 281608 194418 281664
rect 194474 281608 204294 281664
rect 204350 281608 204418 281664
rect 204474 281608 214294 281664
rect 214350 281608 214418 281664
rect 214474 281608 224294 281664
rect 224350 281608 224418 281664
rect 224474 281608 234294 281664
rect 234350 281608 234418 281664
rect 234474 281608 244294 281664
rect 244350 281608 244418 281664
rect 244474 281608 254294 281664
rect 254350 281608 254418 281664
rect 254474 281608 264294 281664
rect 264350 281608 264418 281664
rect 264474 281608 274294 281664
rect 274350 281608 274418 281664
rect 274474 281608 284294 281664
rect 284350 281608 284418 281664
rect 284474 281608 294294 281664
rect 294350 281608 294418 281664
rect 294474 281608 304294 281664
rect 304350 281608 304418 281664
rect 304474 281608 314294 281664
rect 314350 281608 314418 281664
rect 314474 281608 324294 281664
rect 324350 281608 324418 281664
rect 324474 281608 334294 281664
rect 334350 281608 334418 281664
rect 334474 281608 344294 281664
rect 344350 281608 344418 281664
rect 344474 281608 354294 281664
rect 354350 281608 354418 281664
rect 354474 281608 364294 281664
rect 364350 281608 364418 281664
rect 364474 281608 374294 281664
rect 374350 281608 374418 281664
rect 374474 281608 384294 281664
rect 384350 281608 384418 281664
rect 384474 281608 394294 281664
rect 394350 281608 394418 281664
rect 394474 281608 404294 281664
rect 404350 281608 404418 281664
rect 404474 281608 414294 281664
rect 414350 281608 414418 281664
rect 414474 281608 424294 281664
rect 424350 281608 424418 281664
rect 424474 281608 434294 281664
rect 434350 281608 434418 281664
rect 434474 281608 444294 281664
rect 444350 281608 444418 281664
rect 444474 281608 454294 281664
rect 454350 281608 454418 281664
rect 454474 281608 464294 281664
rect 464350 281608 464418 281664
rect 464474 281608 474294 281664
rect 474350 281608 474418 281664
rect 474474 281608 484294 281664
rect 484350 281608 484418 281664
rect 484474 281608 494294 281664
rect 494350 281608 494418 281664
rect 494474 281608 504294 281664
rect 504350 281608 504418 281664
rect 504474 281608 514294 281664
rect 514350 281608 514418 281664
rect 514474 281608 524294 281664
rect 524350 281608 524418 281664
rect 524474 281608 534294 281664
rect 534350 281608 534418 281664
rect 534474 281608 544294 281664
rect 544350 281608 544418 281664
rect 544474 281608 554294 281664
rect 554350 281608 554418 281664
rect 554474 281608 593240 281664
rect 77678 281600 593240 281608
rect 77678 281544 77808 281600
rect 77864 281544 77932 281600
rect 77988 281544 78056 281600
rect 78112 281544 78180 281600
rect 78236 281544 78304 281600
rect 78360 281544 78428 281600
rect 78484 281544 78552 281600
rect 78608 281544 592370 281600
rect 592426 281544 592494 281600
rect 592550 281544 592618 281600
rect 592674 281544 592742 281600
rect 592798 281544 592866 281600
rect 592922 281544 592990 281600
rect 593046 281544 593114 281600
rect 593170 281544 593240 281600
rect 77678 281540 593240 281544
rect 77678 281484 94294 281540
rect 94350 281484 94418 281540
rect 94474 281484 104294 281540
rect 104350 281484 104418 281540
rect 104474 281484 114294 281540
rect 114350 281484 114418 281540
rect 114474 281484 124294 281540
rect 124350 281484 124418 281540
rect 124474 281484 134294 281540
rect 134350 281484 134418 281540
rect 134474 281484 144294 281540
rect 144350 281484 144418 281540
rect 144474 281484 154294 281540
rect 154350 281484 154418 281540
rect 154474 281484 164294 281540
rect 164350 281484 164418 281540
rect 164474 281484 174294 281540
rect 174350 281484 174418 281540
rect 174474 281484 184294 281540
rect 184350 281484 184418 281540
rect 184474 281484 194294 281540
rect 194350 281484 194418 281540
rect 194474 281484 204294 281540
rect 204350 281484 204418 281540
rect 204474 281484 214294 281540
rect 214350 281484 214418 281540
rect 214474 281484 224294 281540
rect 224350 281484 224418 281540
rect 224474 281484 234294 281540
rect 234350 281484 234418 281540
rect 234474 281484 244294 281540
rect 244350 281484 244418 281540
rect 244474 281484 254294 281540
rect 254350 281484 254418 281540
rect 254474 281484 264294 281540
rect 264350 281484 264418 281540
rect 264474 281484 274294 281540
rect 274350 281484 274418 281540
rect 274474 281484 284294 281540
rect 284350 281484 284418 281540
rect 284474 281484 294294 281540
rect 294350 281484 294418 281540
rect 294474 281484 304294 281540
rect 304350 281484 304418 281540
rect 304474 281484 314294 281540
rect 314350 281484 314418 281540
rect 314474 281484 324294 281540
rect 324350 281484 324418 281540
rect 324474 281484 334294 281540
rect 334350 281484 334418 281540
rect 334474 281484 344294 281540
rect 344350 281484 344418 281540
rect 344474 281484 354294 281540
rect 354350 281484 354418 281540
rect 354474 281484 364294 281540
rect 364350 281484 364418 281540
rect 364474 281484 374294 281540
rect 374350 281484 374418 281540
rect 374474 281484 384294 281540
rect 384350 281484 384418 281540
rect 384474 281484 394294 281540
rect 394350 281484 394418 281540
rect 394474 281484 404294 281540
rect 404350 281484 404418 281540
rect 404474 281484 414294 281540
rect 414350 281484 414418 281540
rect 414474 281484 424294 281540
rect 424350 281484 424418 281540
rect 424474 281484 434294 281540
rect 434350 281484 434418 281540
rect 434474 281484 444294 281540
rect 444350 281484 444418 281540
rect 444474 281484 454294 281540
rect 454350 281484 454418 281540
rect 454474 281484 464294 281540
rect 464350 281484 464418 281540
rect 464474 281484 474294 281540
rect 474350 281484 474418 281540
rect 474474 281484 484294 281540
rect 484350 281484 484418 281540
rect 484474 281484 494294 281540
rect 494350 281484 494418 281540
rect 494474 281484 504294 281540
rect 504350 281484 504418 281540
rect 504474 281484 514294 281540
rect 514350 281484 514418 281540
rect 514474 281484 524294 281540
rect 524350 281484 524418 281540
rect 524474 281484 534294 281540
rect 534350 281484 534418 281540
rect 534474 281484 544294 281540
rect 544350 281484 544418 281540
rect 544474 281484 554294 281540
rect 554350 281484 554418 281540
rect 554474 281484 593240 281540
rect 77678 281476 593240 281484
rect 77678 281420 77808 281476
rect 77864 281420 77932 281476
rect 77988 281420 78056 281476
rect 78112 281420 78180 281476
rect 78236 281420 78304 281476
rect 78360 281420 78428 281476
rect 78484 281420 78552 281476
rect 78608 281420 592370 281476
rect 592426 281420 592494 281476
rect 592550 281420 592618 281476
rect 592674 281420 592742 281476
rect 592798 281420 592866 281476
rect 592922 281420 592990 281476
rect 593046 281420 593114 281476
rect 593170 281420 593240 281476
rect 77678 281416 593240 281420
rect 77678 281360 94294 281416
rect 94350 281360 94418 281416
rect 94474 281360 104294 281416
rect 104350 281360 104418 281416
rect 104474 281360 114294 281416
rect 114350 281360 114418 281416
rect 114474 281360 124294 281416
rect 124350 281360 124418 281416
rect 124474 281360 134294 281416
rect 134350 281360 134418 281416
rect 134474 281360 144294 281416
rect 144350 281360 144418 281416
rect 144474 281360 154294 281416
rect 154350 281360 154418 281416
rect 154474 281360 164294 281416
rect 164350 281360 164418 281416
rect 164474 281360 174294 281416
rect 174350 281360 174418 281416
rect 174474 281360 184294 281416
rect 184350 281360 184418 281416
rect 184474 281360 194294 281416
rect 194350 281360 194418 281416
rect 194474 281360 204294 281416
rect 204350 281360 204418 281416
rect 204474 281360 214294 281416
rect 214350 281360 214418 281416
rect 214474 281360 224294 281416
rect 224350 281360 224418 281416
rect 224474 281360 234294 281416
rect 234350 281360 234418 281416
rect 234474 281360 244294 281416
rect 244350 281360 244418 281416
rect 244474 281360 254294 281416
rect 254350 281360 254418 281416
rect 254474 281360 264294 281416
rect 264350 281360 264418 281416
rect 264474 281360 274294 281416
rect 274350 281360 274418 281416
rect 274474 281360 284294 281416
rect 284350 281360 284418 281416
rect 284474 281360 294294 281416
rect 294350 281360 294418 281416
rect 294474 281360 304294 281416
rect 304350 281360 304418 281416
rect 304474 281360 314294 281416
rect 314350 281360 314418 281416
rect 314474 281360 324294 281416
rect 324350 281360 324418 281416
rect 324474 281360 334294 281416
rect 334350 281360 334418 281416
rect 334474 281360 344294 281416
rect 344350 281360 344418 281416
rect 344474 281360 354294 281416
rect 354350 281360 354418 281416
rect 354474 281360 364294 281416
rect 364350 281360 364418 281416
rect 364474 281360 374294 281416
rect 374350 281360 374418 281416
rect 374474 281360 384294 281416
rect 384350 281360 384418 281416
rect 384474 281360 394294 281416
rect 394350 281360 394418 281416
rect 394474 281360 404294 281416
rect 404350 281360 404418 281416
rect 404474 281360 414294 281416
rect 414350 281360 414418 281416
rect 414474 281360 424294 281416
rect 424350 281360 424418 281416
rect 424474 281360 434294 281416
rect 434350 281360 434418 281416
rect 434474 281360 444294 281416
rect 444350 281360 444418 281416
rect 444474 281360 454294 281416
rect 454350 281360 454418 281416
rect 454474 281360 464294 281416
rect 464350 281360 464418 281416
rect 464474 281360 474294 281416
rect 474350 281360 474418 281416
rect 474474 281360 484294 281416
rect 484350 281360 484418 281416
rect 484474 281360 494294 281416
rect 494350 281360 494418 281416
rect 494474 281360 504294 281416
rect 504350 281360 504418 281416
rect 504474 281360 514294 281416
rect 514350 281360 514418 281416
rect 514474 281360 524294 281416
rect 524350 281360 524418 281416
rect 524474 281360 534294 281416
rect 534350 281360 534418 281416
rect 534474 281360 544294 281416
rect 544350 281360 544418 281416
rect 544474 281360 554294 281416
rect 554350 281360 554418 281416
rect 554474 281360 593240 281416
rect 77678 281352 593240 281360
rect 77678 281296 77808 281352
rect 77864 281296 77932 281352
rect 77988 281296 78056 281352
rect 78112 281296 78180 281352
rect 78236 281296 78304 281352
rect 78360 281296 78428 281352
rect 78484 281296 78552 281352
rect 78608 281296 592370 281352
rect 592426 281296 592494 281352
rect 592550 281296 592618 281352
rect 592674 281296 592742 281352
rect 592798 281296 592866 281352
rect 592922 281296 592990 281352
rect 593046 281296 593114 281352
rect 593170 281296 593240 281352
rect 77678 281292 593240 281296
rect 77678 281236 94294 281292
rect 94350 281236 94418 281292
rect 94474 281236 104294 281292
rect 104350 281236 104418 281292
rect 104474 281236 114294 281292
rect 114350 281236 114418 281292
rect 114474 281236 124294 281292
rect 124350 281236 124418 281292
rect 124474 281236 134294 281292
rect 134350 281236 134418 281292
rect 134474 281236 144294 281292
rect 144350 281236 144418 281292
rect 144474 281236 154294 281292
rect 154350 281236 154418 281292
rect 154474 281236 164294 281292
rect 164350 281236 164418 281292
rect 164474 281236 174294 281292
rect 174350 281236 174418 281292
rect 174474 281236 184294 281292
rect 184350 281236 184418 281292
rect 184474 281236 194294 281292
rect 194350 281236 194418 281292
rect 194474 281236 204294 281292
rect 204350 281236 204418 281292
rect 204474 281236 214294 281292
rect 214350 281236 214418 281292
rect 214474 281236 224294 281292
rect 224350 281236 224418 281292
rect 224474 281236 234294 281292
rect 234350 281236 234418 281292
rect 234474 281236 244294 281292
rect 244350 281236 244418 281292
rect 244474 281236 254294 281292
rect 254350 281236 254418 281292
rect 254474 281236 264294 281292
rect 264350 281236 264418 281292
rect 264474 281236 274294 281292
rect 274350 281236 274418 281292
rect 274474 281236 284294 281292
rect 284350 281236 284418 281292
rect 284474 281236 294294 281292
rect 294350 281236 294418 281292
rect 294474 281236 304294 281292
rect 304350 281236 304418 281292
rect 304474 281236 314294 281292
rect 314350 281236 314418 281292
rect 314474 281236 324294 281292
rect 324350 281236 324418 281292
rect 324474 281236 334294 281292
rect 334350 281236 334418 281292
rect 334474 281236 344294 281292
rect 344350 281236 344418 281292
rect 344474 281236 354294 281292
rect 354350 281236 354418 281292
rect 354474 281236 364294 281292
rect 364350 281236 364418 281292
rect 364474 281236 374294 281292
rect 374350 281236 374418 281292
rect 374474 281236 384294 281292
rect 384350 281236 384418 281292
rect 384474 281236 394294 281292
rect 394350 281236 394418 281292
rect 394474 281236 404294 281292
rect 404350 281236 404418 281292
rect 404474 281236 414294 281292
rect 414350 281236 414418 281292
rect 414474 281236 424294 281292
rect 424350 281236 424418 281292
rect 424474 281236 434294 281292
rect 434350 281236 434418 281292
rect 434474 281236 444294 281292
rect 444350 281236 444418 281292
rect 444474 281236 454294 281292
rect 454350 281236 454418 281292
rect 454474 281236 464294 281292
rect 464350 281236 464418 281292
rect 464474 281236 474294 281292
rect 474350 281236 474418 281292
rect 474474 281236 484294 281292
rect 484350 281236 484418 281292
rect 484474 281236 494294 281292
rect 494350 281236 494418 281292
rect 494474 281236 504294 281292
rect 504350 281236 504418 281292
rect 504474 281236 514294 281292
rect 514350 281236 514418 281292
rect 514474 281236 524294 281292
rect 524350 281236 524418 281292
rect 524474 281236 534294 281292
rect 534350 281236 534418 281292
rect 534474 281236 544294 281292
rect 544350 281236 544418 281292
rect 544474 281236 554294 281292
rect 554350 281236 554418 281292
rect 554474 281236 593240 281292
rect 77678 281228 593240 281236
rect 77678 281172 77808 281228
rect 77864 281172 77932 281228
rect 77988 281172 78056 281228
rect 78112 281172 78180 281228
rect 78236 281172 78304 281228
rect 78360 281172 78428 281228
rect 78484 281172 78552 281228
rect 78608 281172 592370 281228
rect 592426 281172 592494 281228
rect 592550 281172 592618 281228
rect 592674 281172 592742 281228
rect 592798 281172 592866 281228
rect 592922 281172 592990 281228
rect 593046 281172 593114 281228
rect 593170 281172 593240 281228
rect 77678 281168 593240 281172
rect 77678 281112 94294 281168
rect 94350 281112 94418 281168
rect 94474 281112 104294 281168
rect 104350 281112 104418 281168
rect 104474 281112 114294 281168
rect 114350 281112 114418 281168
rect 114474 281112 124294 281168
rect 124350 281112 124418 281168
rect 124474 281112 134294 281168
rect 134350 281112 134418 281168
rect 134474 281112 144294 281168
rect 144350 281112 144418 281168
rect 144474 281112 154294 281168
rect 154350 281112 154418 281168
rect 154474 281112 164294 281168
rect 164350 281112 164418 281168
rect 164474 281112 174294 281168
rect 174350 281112 174418 281168
rect 174474 281112 184294 281168
rect 184350 281112 184418 281168
rect 184474 281112 194294 281168
rect 194350 281112 194418 281168
rect 194474 281112 204294 281168
rect 204350 281112 204418 281168
rect 204474 281112 214294 281168
rect 214350 281112 214418 281168
rect 214474 281112 224294 281168
rect 224350 281112 224418 281168
rect 224474 281112 234294 281168
rect 234350 281112 234418 281168
rect 234474 281112 244294 281168
rect 244350 281112 244418 281168
rect 244474 281112 254294 281168
rect 254350 281112 254418 281168
rect 254474 281112 264294 281168
rect 264350 281112 264418 281168
rect 264474 281112 274294 281168
rect 274350 281112 274418 281168
rect 274474 281112 284294 281168
rect 284350 281112 284418 281168
rect 284474 281112 294294 281168
rect 294350 281112 294418 281168
rect 294474 281112 304294 281168
rect 304350 281112 304418 281168
rect 304474 281112 314294 281168
rect 314350 281112 314418 281168
rect 314474 281112 324294 281168
rect 324350 281112 324418 281168
rect 324474 281112 334294 281168
rect 334350 281112 334418 281168
rect 334474 281112 344294 281168
rect 344350 281112 344418 281168
rect 344474 281112 354294 281168
rect 354350 281112 354418 281168
rect 354474 281112 364294 281168
rect 364350 281112 364418 281168
rect 364474 281112 374294 281168
rect 374350 281112 374418 281168
rect 374474 281112 384294 281168
rect 384350 281112 384418 281168
rect 384474 281112 394294 281168
rect 394350 281112 394418 281168
rect 394474 281112 404294 281168
rect 404350 281112 404418 281168
rect 404474 281112 414294 281168
rect 414350 281112 414418 281168
rect 414474 281112 424294 281168
rect 424350 281112 424418 281168
rect 424474 281112 434294 281168
rect 434350 281112 434418 281168
rect 434474 281112 444294 281168
rect 444350 281112 444418 281168
rect 444474 281112 454294 281168
rect 454350 281112 454418 281168
rect 454474 281112 464294 281168
rect 464350 281112 464418 281168
rect 464474 281112 474294 281168
rect 474350 281112 474418 281168
rect 474474 281112 484294 281168
rect 484350 281112 484418 281168
rect 484474 281112 494294 281168
rect 494350 281112 494418 281168
rect 494474 281112 504294 281168
rect 504350 281112 504418 281168
rect 504474 281112 514294 281168
rect 514350 281112 514418 281168
rect 514474 281112 524294 281168
rect 524350 281112 524418 281168
rect 524474 281112 534294 281168
rect 534350 281112 534418 281168
rect 534474 281112 544294 281168
rect 544350 281112 544418 281168
rect 544474 281112 554294 281168
rect 554350 281112 554418 281168
rect 554474 281112 593240 281168
rect 77678 281042 593240 281112
rect 699322 280954 702688 281076
rect 699322 280898 699444 280954
rect 699500 280898 699744 280954
rect 699800 280898 700044 280954
rect 700100 280898 702688 280954
rect 699322 280756 702688 280898
rect 697922 277434 702624 277576
rect 697922 277378 698044 277434
rect 698100 277378 698344 277434
rect 698400 277378 698644 277434
rect 698700 277378 702624 277434
rect 697922 277256 702624 277378
rect 699322 273954 702688 274076
rect 699322 273898 699444 273954
rect 699500 273898 699744 273954
rect 699800 273898 700044 273954
rect 700100 273898 702688 273954
rect 699322 273756 702688 273898
rect 75376 273622 80078 273744
rect 75376 273566 79300 273622
rect 79356 273566 79600 273622
rect 79656 273566 79900 273622
rect 79956 273566 80078 273622
rect 75376 273424 80078 273566
rect 697922 270434 702624 270576
rect 697922 270378 698044 270434
rect 698100 270378 698344 270434
rect 698400 270378 698644 270434
rect 698700 270378 702624 270434
rect 697922 270256 702624 270378
rect 75312 270102 78678 270244
rect 75312 270046 77900 270102
rect 77956 270046 78200 270102
rect 78256 270046 78500 270102
rect 78556 270046 78678 270102
rect 75312 269924 78678 270046
rect 666132 268607 700322 268749
rect 666132 268551 699444 268607
rect 699500 268551 699744 268607
rect 699800 268551 700044 268607
rect 700100 268551 700322 268607
rect 77678 268372 89920 268442
rect 77678 268316 77748 268372
rect 77804 268316 77872 268372
rect 77928 268316 77996 268372
rect 78052 268316 78120 268372
rect 78176 268316 78244 268372
rect 78300 268316 78368 268372
rect 78424 268316 78492 268372
rect 78548 268316 89920 268372
rect 77678 268248 89920 268316
rect 77678 268192 77748 268248
rect 77804 268192 77872 268248
rect 77928 268192 77996 268248
rect 78052 268192 78120 268248
rect 78176 268192 78244 268248
rect 78300 268192 78368 268248
rect 78424 268192 78492 268248
rect 78548 268192 89920 268248
rect 77678 268122 89920 268192
rect 560032 268372 593240 268442
rect 666132 268429 700322 268551
rect 560032 268316 592370 268372
rect 592426 268316 592494 268372
rect 592550 268316 592618 268372
rect 592674 268316 592742 268372
rect 592798 268316 592866 268372
rect 592922 268316 592990 268372
rect 593046 268316 593114 268372
rect 593170 268316 593240 268372
rect 560032 268248 593240 268316
rect 560032 268192 592370 268248
rect 592426 268192 592494 268248
rect 592550 268192 592618 268248
rect 592674 268192 592742 268248
rect 592798 268192 592866 268248
rect 592922 268192 592990 268248
rect 593046 268192 593114 268248
rect 593170 268192 593240 268248
rect 560032 268122 593240 268192
rect 699322 266954 702688 267076
rect 699322 266898 699444 266954
rect 699500 266898 699744 266954
rect 699800 266898 700044 266954
rect 700100 266898 702688 266954
rect 699322 266756 702688 266898
rect 75376 266622 80078 266744
rect 75376 266566 79300 266622
rect 79356 266566 79600 266622
rect 79656 266566 79900 266622
rect 79956 266566 80078 266622
rect 75376 266424 80078 266566
rect 697922 263434 702624 263576
rect 697922 263378 698044 263434
rect 698100 263378 698344 263434
rect 698400 263378 698644 263434
rect 698700 263378 702624 263434
rect 697922 263256 702624 263378
rect 75312 263102 78678 263244
rect 75312 263046 77900 263102
rect 77956 263046 78200 263102
rect 78256 263046 78500 263102
rect 78556 263046 78678 263102
rect 75312 262924 78678 263046
rect 75376 259622 80078 259744
rect 75376 259566 79300 259622
rect 79356 259566 79600 259622
rect 79656 259566 79900 259622
rect 79956 259566 80078 259622
rect 75376 259424 80078 259566
rect 75312 256102 78678 256244
rect 75312 256046 77900 256102
rect 77956 256046 78200 256102
rect 78256 256046 78500 256102
rect 78556 256046 78678 256102
rect 75312 255924 78678 256046
rect 79078 255372 89920 255442
rect 79078 255316 79148 255372
rect 79204 255316 79272 255372
rect 79328 255316 79396 255372
rect 79452 255316 79520 255372
rect 79576 255316 79644 255372
rect 79700 255316 79768 255372
rect 79824 255316 79892 255372
rect 79948 255316 89920 255372
rect 79078 255248 89920 255316
rect 79078 255192 79148 255248
rect 79204 255192 79272 255248
rect 79328 255192 79396 255248
rect 79452 255192 79520 255248
rect 79576 255192 79644 255248
rect 79700 255192 79768 255248
rect 79824 255192 79892 255248
rect 79948 255192 89920 255248
rect 79078 255122 89920 255192
rect 560032 255372 591840 255442
rect 560032 255316 590970 255372
rect 591026 255316 591094 255372
rect 591150 255316 591218 255372
rect 591274 255316 591342 255372
rect 591398 255316 591466 255372
rect 591522 255316 591590 255372
rect 591646 255316 591714 255372
rect 591770 255316 591840 255372
rect 560032 255248 591840 255316
rect 560032 255192 590970 255248
rect 591026 255192 591094 255248
rect 591150 255192 591218 255248
rect 591274 255192 591342 255248
rect 591398 255192 591466 255248
rect 591522 255192 591590 255248
rect 591646 255192 591714 255248
rect 591770 255192 591840 255248
rect 560032 255122 591840 255192
rect 666132 253289 698922 253431
rect 666132 253233 698044 253289
rect 698100 253233 698344 253289
rect 698400 253233 698644 253289
rect 698700 253233 698922 253289
rect 666132 253111 698922 253233
rect 76115 249048 80078 249110
rect 76115 248992 79284 249048
rect 79340 248992 79584 249048
rect 79640 248992 79884 249048
rect 79940 248992 80078 249048
rect 76115 248910 80078 248992
rect 76115 248510 76435 248910
rect 76915 248633 78678 248710
rect 76915 248577 77847 248633
rect 77903 248577 78147 248633
rect 78203 248577 78447 248633
rect 78503 248577 78678 248633
rect 76915 248510 78678 248577
rect 699322 247423 701085 247490
rect 699322 247367 699497 247423
rect 699553 247367 699797 247423
rect 699853 247367 700097 247423
rect 700153 247367 701085 247423
rect 699322 247290 701085 247367
rect 701565 247090 701885 247490
rect 697922 247008 701885 247090
rect 697922 246952 698060 247008
rect 698116 246952 698360 247008
rect 698416 246952 698660 247008
rect 698716 246952 701885 247008
rect 697922 246890 701885 246952
rect 77678 242372 89920 242442
rect 77678 242316 77748 242372
rect 77804 242316 77872 242372
rect 77928 242316 77996 242372
rect 78052 242316 78120 242372
rect 78176 242316 78244 242372
rect 78300 242316 78368 242372
rect 78424 242316 78492 242372
rect 78548 242316 89920 242372
rect 77678 242248 89920 242316
rect 77678 242192 77748 242248
rect 77804 242192 77872 242248
rect 77928 242192 77996 242248
rect 78052 242192 78120 242248
rect 78176 242192 78244 242248
rect 78300 242192 78368 242248
rect 78424 242192 78492 242248
rect 78548 242192 89920 242248
rect 77678 242122 89920 242192
rect 560032 242372 593240 242442
rect 560032 242316 592370 242372
rect 592426 242316 592494 242372
rect 592550 242316 592618 242372
rect 592674 242316 592742 242372
rect 592798 242316 592866 242372
rect 592922 242316 592990 242372
rect 593046 242316 593114 242372
rect 593170 242316 593240 242372
rect 560032 242248 593240 242316
rect 560032 242192 592370 242248
rect 592426 242192 592494 242248
rect 592550 242192 592618 242248
rect 592674 242192 592742 242248
rect 592798 242192 592866 242248
rect 592922 242192 592990 242248
rect 593046 242192 593114 242248
rect 593170 242192 593240 242248
rect 560032 242122 593240 242192
rect 699322 237971 702688 238076
rect 699322 237915 699444 237971
rect 699500 237915 699744 237971
rect 699800 237915 700044 237971
rect 700100 237915 702688 237971
rect 699322 237756 702688 237915
rect 697922 234434 702624 234576
rect 697922 234378 698044 234434
rect 698100 234378 698344 234434
rect 698400 234378 698644 234434
rect 698700 234378 702624 234434
rect 697922 234256 702624 234378
rect 75376 232622 80078 232744
rect 75376 232566 79300 232622
rect 79356 232566 79600 232622
rect 79656 232566 79900 232622
rect 79956 232566 80078 232622
rect 75376 232424 80078 232566
rect 699322 230954 702688 231076
rect 699322 230898 699444 230954
rect 699500 230898 699744 230954
rect 699800 230898 700044 230954
rect 700100 230898 702688 230954
rect 699322 230756 702688 230898
rect 79078 229372 89920 229442
rect 79078 229316 79148 229372
rect 79204 229316 79272 229372
rect 79328 229316 79396 229372
rect 79452 229316 79520 229372
rect 79576 229316 79644 229372
rect 79700 229316 79768 229372
rect 79824 229316 79892 229372
rect 79948 229316 89920 229372
rect 79078 229248 89920 229316
rect 75312 229102 78678 229244
rect 79078 229192 79148 229248
rect 79204 229192 79272 229248
rect 79328 229192 79396 229248
rect 79452 229192 79520 229248
rect 79576 229192 79644 229248
rect 79700 229192 79768 229248
rect 79824 229192 79892 229248
rect 79948 229192 89920 229248
rect 79078 229122 89920 229192
rect 560032 229372 591840 229442
rect 560032 229316 590970 229372
rect 591026 229316 591094 229372
rect 591150 229316 591218 229372
rect 591274 229316 591342 229372
rect 591398 229316 591466 229372
rect 591522 229316 591590 229372
rect 591646 229316 591714 229372
rect 591770 229316 591840 229372
rect 560032 229248 591840 229316
rect 560032 229192 590970 229248
rect 591026 229192 591094 229248
rect 591150 229192 591218 229248
rect 591274 229192 591342 229248
rect 591398 229192 591466 229248
rect 591522 229192 591590 229248
rect 591646 229192 591714 229248
rect 591770 229192 591840 229248
rect 560032 229122 591840 229192
rect 75312 229046 77900 229102
rect 77956 229046 78200 229102
rect 78256 229046 78500 229102
rect 78556 229046 78678 229102
rect 75312 228924 78678 229046
rect 697922 227434 702624 227576
rect 697922 227378 698044 227434
rect 698100 227378 698344 227434
rect 698400 227378 698644 227434
rect 698700 227378 702624 227434
rect 697922 227256 702624 227378
rect 75376 225622 80078 225744
rect 75376 225566 79300 225622
rect 79356 225566 79600 225622
rect 79656 225566 79900 225622
rect 79956 225566 80078 225622
rect 75376 225424 80078 225566
rect 699322 223954 702688 224076
rect 699322 223898 699444 223954
rect 699500 223898 699744 223954
rect 699800 223898 700044 223954
rect 700100 223898 702688 223954
rect 699322 223756 702688 223898
rect 666132 222653 698922 222795
rect 666132 222597 698044 222653
rect 698100 222597 698344 222653
rect 698400 222597 698644 222653
rect 698700 222597 698922 222653
rect 666132 222475 698922 222597
rect 75312 222102 78678 222244
rect 75312 222046 77900 222102
rect 77956 222046 78200 222102
rect 78256 222046 78500 222102
rect 78556 222046 78678 222102
rect 75312 221924 78678 222046
rect 697922 220434 702624 220576
rect 697922 220378 698044 220434
rect 698100 220378 698344 220434
rect 698400 220378 698644 220434
rect 698700 220378 702624 220434
rect 697922 220256 702624 220378
rect 75376 218622 80078 218744
rect 75376 218566 79300 218622
rect 79356 218566 79600 218622
rect 79656 218566 79900 218622
rect 79956 218566 80078 218622
rect 75376 218424 80078 218566
rect 77678 216372 89920 216442
rect 77678 216316 77748 216372
rect 77804 216316 77872 216372
rect 77928 216316 77996 216372
rect 78052 216316 78120 216372
rect 78176 216316 78244 216372
rect 78300 216316 78368 216372
rect 78424 216316 78492 216372
rect 78548 216316 89920 216372
rect 77678 216248 89920 216316
rect 77678 216192 77748 216248
rect 77804 216192 77872 216248
rect 77928 216192 77996 216248
rect 78052 216192 78120 216248
rect 78176 216192 78244 216248
rect 78300 216192 78368 216248
rect 78424 216192 78492 216248
rect 78548 216192 89920 216248
rect 77678 216122 89920 216192
rect 560032 216372 593240 216442
rect 560032 216316 592370 216372
rect 592426 216316 592494 216372
rect 592550 216316 592618 216372
rect 592674 216316 592742 216372
rect 592798 216316 592866 216372
rect 592922 216316 592990 216372
rect 593046 216316 593114 216372
rect 593170 216316 593240 216372
rect 560032 216248 593240 216316
rect 560032 216192 592370 216248
rect 592426 216192 592494 216248
rect 592550 216192 592618 216248
rect 592674 216192 592742 216248
rect 592798 216192 592866 216248
rect 592922 216192 592990 216248
rect 593046 216192 593114 216248
rect 593170 216192 593240 216248
rect 560032 216122 593240 216192
rect 75312 215102 78678 215244
rect 75312 215046 77900 215102
rect 77956 215046 78200 215102
rect 78256 215046 78500 215102
rect 78556 215046 78678 215102
rect 75312 214924 78678 215046
rect 76115 208048 80078 208110
rect 76115 207992 79284 208048
rect 79340 207992 79584 208048
rect 79640 207992 79884 208048
rect 79940 207992 80078 208048
rect 76115 207910 80078 207992
rect 76115 207510 76435 207910
rect 76915 207633 78678 207710
rect 76915 207577 77847 207633
rect 77903 207577 78147 207633
rect 78203 207577 78447 207633
rect 78503 207577 78678 207633
rect 76915 207510 78678 207577
rect 666132 207335 700322 207477
rect 666132 207279 699444 207335
rect 699500 207279 699744 207335
rect 699800 207279 700044 207335
rect 700100 207279 700322 207335
rect 666132 207157 700322 207279
rect 699322 204423 701085 204490
rect 699322 204367 699497 204423
rect 699553 204367 699797 204423
rect 699853 204367 700097 204423
rect 700153 204367 701085 204423
rect 699322 204290 701085 204367
rect 701565 204090 701885 204490
rect 697922 204008 701885 204090
rect 697922 203952 698060 204008
rect 698116 203952 698360 204008
rect 698416 203952 698660 204008
rect 698716 203952 701885 204008
rect 697922 203890 701885 203952
rect 79078 203372 89920 203442
rect 79078 203316 79148 203372
rect 79204 203316 79272 203372
rect 79328 203316 79396 203372
rect 79452 203316 79520 203372
rect 79576 203316 79644 203372
rect 79700 203316 79768 203372
rect 79824 203316 79892 203372
rect 79948 203316 89920 203372
rect 79078 203248 89920 203316
rect 79078 203192 79148 203248
rect 79204 203192 79272 203248
rect 79328 203192 79396 203248
rect 79452 203192 79520 203248
rect 79576 203192 79644 203248
rect 79700 203192 79768 203248
rect 79824 203192 79892 203248
rect 79948 203192 89920 203248
rect 79078 203122 89920 203192
rect 560032 203372 591840 203442
rect 560032 203316 590970 203372
rect 591026 203316 591094 203372
rect 591150 203316 591218 203372
rect 591274 203316 591342 203372
rect 591398 203316 591466 203372
rect 591522 203316 591590 203372
rect 591646 203316 591714 203372
rect 591770 203316 591840 203372
rect 560032 203248 591840 203316
rect 560032 203192 590970 203248
rect 591026 203192 591094 203248
rect 591150 203192 591218 203248
rect 591274 203192 591342 203248
rect 591398 203192 591466 203248
rect 591522 203192 591590 203248
rect 591646 203192 591714 203248
rect 591770 203192 591840 203248
rect 560032 203122 591840 203192
rect 699322 194954 702688 195076
rect 699322 194898 699444 194954
rect 699500 194898 699744 194954
rect 699800 194898 700044 194954
rect 700100 194898 702688 194954
rect 699322 194756 702688 194898
rect 666132 192017 698922 192159
rect 666132 191961 698044 192017
rect 698100 191961 698344 192017
rect 698400 191961 698644 192017
rect 698700 191961 698922 192017
rect 666132 191839 698922 191961
rect 75376 191622 80078 191744
rect 75376 191566 79300 191622
rect 79356 191566 79600 191622
rect 79656 191566 79900 191622
rect 79956 191566 80078 191622
rect 75376 191424 80078 191566
rect 697922 191434 702624 191576
rect 697922 191378 698044 191434
rect 698100 191378 698344 191434
rect 698400 191378 698644 191434
rect 698700 191378 702624 191434
rect 697922 191256 702624 191378
rect 77678 190372 89920 190442
rect 77678 190316 77748 190372
rect 77804 190316 77872 190372
rect 77928 190316 77996 190372
rect 78052 190316 78120 190372
rect 78176 190316 78244 190372
rect 78300 190316 78368 190372
rect 78424 190316 78492 190372
rect 78548 190316 89920 190372
rect 77678 190248 89920 190316
rect 77678 190192 77748 190248
rect 77804 190192 77872 190248
rect 77928 190192 77996 190248
rect 78052 190192 78120 190248
rect 78176 190192 78244 190248
rect 78300 190192 78368 190248
rect 78424 190192 78492 190248
rect 78548 190192 89920 190248
rect 77678 190122 89920 190192
rect 560032 190372 593240 190442
rect 560032 190316 592370 190372
rect 592426 190316 592494 190372
rect 592550 190316 592618 190372
rect 592674 190316 592742 190372
rect 592798 190316 592866 190372
rect 592922 190316 592990 190372
rect 593046 190316 593114 190372
rect 593170 190316 593240 190372
rect 560032 190248 593240 190316
rect 560032 190192 592370 190248
rect 592426 190192 592494 190248
rect 592550 190192 592618 190248
rect 592674 190192 592742 190248
rect 592798 190192 592866 190248
rect 592922 190192 592990 190248
rect 593046 190192 593114 190248
rect 593170 190192 593240 190248
rect 560032 190122 593240 190192
rect 75312 188102 78678 188244
rect 75312 188046 77900 188102
rect 77956 188046 78200 188102
rect 78256 188046 78500 188102
rect 78556 188046 78678 188102
rect 75312 187924 78678 188046
rect 699322 187954 702688 188076
rect 699322 187898 699444 187954
rect 699500 187898 699744 187954
rect 699800 187898 700044 187954
rect 700100 187898 702688 187954
rect 699322 187756 702688 187898
rect 75376 184622 80078 184744
rect 75376 184566 79300 184622
rect 79356 184566 79600 184622
rect 79656 184566 79900 184622
rect 79956 184566 80078 184622
rect 75376 184424 80078 184566
rect 697922 184434 702624 184576
rect 697922 184378 698044 184434
rect 698100 184378 698344 184434
rect 698400 184378 698644 184434
rect 698700 184378 702624 184434
rect 697922 184256 702624 184378
rect 75312 181102 78678 181244
rect 75312 181046 77900 181102
rect 77956 181046 78200 181102
rect 78256 181046 78500 181102
rect 78556 181046 78678 181102
rect 75312 180924 78678 181046
rect 699322 180954 702688 181076
rect 699322 180898 699444 180954
rect 699500 180898 699744 180954
rect 699800 180898 700044 180954
rect 700100 180898 702688 180954
rect 699322 180756 702688 180898
rect 75376 177622 80078 177744
rect 75376 177566 79300 177622
rect 79356 177566 79600 177622
rect 79656 177566 79900 177622
rect 79956 177566 80078 177622
rect 75376 177442 80078 177566
rect 75376 177424 89920 177442
rect 79078 177372 89920 177424
rect 79078 177316 79148 177372
rect 79204 177316 79272 177372
rect 79328 177316 79396 177372
rect 79452 177316 79520 177372
rect 79576 177316 79644 177372
rect 79700 177316 79768 177372
rect 79824 177316 79892 177372
rect 79948 177316 89920 177372
rect 79078 177248 89920 177316
rect 79078 177192 79148 177248
rect 79204 177192 79272 177248
rect 79328 177192 79396 177248
rect 79452 177192 79520 177248
rect 79576 177192 79644 177248
rect 79700 177192 79768 177248
rect 79824 177192 79892 177248
rect 79948 177192 89920 177248
rect 79078 177122 89920 177192
rect 560032 177372 591840 177442
rect 560032 177316 590970 177372
rect 591026 177316 591094 177372
rect 591150 177316 591218 177372
rect 591274 177316 591342 177372
rect 591398 177316 591466 177372
rect 591522 177316 591590 177372
rect 591646 177316 591714 177372
rect 591770 177316 591840 177372
rect 560032 177248 591840 177316
rect 697922 177434 702624 177576
rect 697922 177378 698044 177434
rect 698100 177378 698344 177434
rect 698400 177378 698644 177434
rect 698700 177378 702624 177434
rect 697922 177256 702624 177378
rect 560032 177192 590970 177248
rect 591026 177192 591094 177248
rect 591150 177192 591218 177248
rect 591274 177192 591342 177248
rect 591398 177192 591466 177248
rect 591522 177192 591590 177248
rect 591646 177192 591714 177248
rect 591770 177192 591840 177248
rect 560032 177122 591840 177192
rect 666132 176699 700322 176841
rect 666132 176643 699444 176699
rect 699500 176643 699744 176699
rect 699800 176643 700044 176699
rect 700100 176643 700322 176699
rect 666132 176521 700322 176643
rect 75312 174102 78678 174244
rect 75312 174046 77900 174102
rect 77956 174046 78200 174102
rect 78256 174046 78500 174102
rect 78556 174046 78678 174102
rect 75312 173924 78678 174046
rect 77678 164372 89920 164442
rect 77678 164316 77748 164372
rect 77804 164316 77872 164372
rect 77928 164316 77996 164372
rect 78052 164316 78120 164372
rect 78176 164316 78244 164372
rect 78300 164316 78368 164372
rect 78424 164316 78492 164372
rect 78548 164316 89920 164372
rect 77678 164248 89920 164316
rect 77678 164192 77748 164248
rect 77804 164192 77872 164248
rect 77928 164192 77996 164248
rect 78052 164192 78120 164248
rect 78176 164192 78244 164248
rect 78300 164192 78368 164248
rect 78424 164192 78492 164248
rect 78548 164192 89920 164248
rect 77678 164122 89920 164192
rect 560032 164372 593240 164442
rect 560032 164316 592370 164372
rect 592426 164316 592494 164372
rect 592550 164316 592618 164372
rect 592674 164316 592742 164372
rect 592798 164316 592866 164372
rect 592922 164316 592990 164372
rect 593046 164316 593114 164372
rect 593170 164316 593240 164372
rect 560032 164248 593240 164316
rect 560032 164192 592370 164248
rect 592426 164192 592494 164248
rect 592550 164192 592618 164248
rect 592674 164192 592742 164248
rect 592798 164192 592866 164248
rect 592922 164192 592990 164248
rect 593046 164192 593114 164248
rect 593170 164192 593240 164248
rect 560032 164122 593240 164192
rect 666132 161381 698922 161523
rect 666132 161325 698044 161381
rect 698100 161325 698344 161381
rect 698400 161325 698644 161381
rect 698700 161325 698922 161381
rect 666132 161203 698922 161325
rect 699322 161423 701085 161490
rect 699322 161367 699497 161423
rect 699553 161367 699797 161423
rect 699853 161367 700097 161423
rect 700153 161367 701085 161423
rect 699322 161290 701085 161367
rect 701565 161090 701885 161490
rect 697922 161008 701885 161090
rect 697922 160952 698060 161008
rect 698116 160952 698360 161008
rect 698416 160952 698660 161008
rect 698716 160952 701885 161008
rect 697922 160890 701885 160952
rect 699322 151954 702688 152076
rect 699322 151898 699444 151954
rect 699500 151898 699744 151954
rect 699800 151898 700044 151954
rect 700100 151898 702688 151954
rect 699322 151756 702688 151898
rect 79078 151372 89920 151442
rect 79078 151316 79148 151372
rect 79204 151316 79272 151372
rect 79328 151316 79396 151372
rect 79452 151316 79520 151372
rect 79576 151316 79644 151372
rect 79700 151316 79768 151372
rect 79824 151316 79892 151372
rect 79948 151316 89920 151372
rect 79078 151248 89920 151316
rect 79078 151192 79148 151248
rect 79204 151192 79272 151248
rect 79328 151192 79396 151248
rect 79452 151192 79520 151248
rect 79576 151192 79644 151248
rect 79700 151192 79768 151248
rect 79824 151192 79892 151248
rect 79948 151192 89920 151248
rect 79078 151122 89920 151192
rect 560032 151372 591840 151442
rect 560032 151316 590970 151372
rect 591026 151316 591094 151372
rect 591150 151316 591218 151372
rect 591274 151316 591342 151372
rect 591398 151316 591466 151372
rect 591522 151316 591590 151372
rect 591646 151316 591714 151372
rect 591770 151316 591840 151372
rect 560032 151248 591840 151316
rect 560032 151192 590970 151248
rect 591026 151192 591094 151248
rect 591150 151192 591218 151248
rect 591274 151192 591342 151248
rect 591398 151192 591466 151248
rect 591522 151192 591590 151248
rect 591646 151192 591714 151248
rect 591770 151192 591840 151248
rect 560032 151122 591840 151192
rect 697922 148434 702624 148576
rect 697922 148378 698044 148434
rect 698100 148378 698344 148434
rect 698400 148378 698644 148434
rect 698700 148378 702624 148434
rect 697922 148256 702624 148378
rect 70000 146670 78678 146728
rect 70000 146658 77808 146670
rect 70000 146602 70074 146658
rect 70130 146614 77808 146658
rect 77864 146614 77932 146670
rect 77988 146614 78056 146670
rect 78112 146614 78180 146670
rect 78236 146614 78304 146670
rect 78360 146614 78428 146670
rect 78484 146614 78552 146670
rect 78608 146614 78678 146670
rect 70130 146602 78678 146614
rect 70000 146546 78678 146602
rect 70000 146534 77808 146546
rect 70000 146478 70074 146534
rect 70130 146490 77808 146534
rect 77864 146490 77932 146546
rect 77988 146490 78056 146546
rect 78112 146490 78180 146546
rect 78236 146490 78304 146546
rect 78360 146490 78428 146546
rect 78484 146490 78552 146546
rect 78608 146490 78678 146546
rect 70130 146478 78678 146490
rect 70000 146422 78678 146478
rect 70000 146410 77808 146422
rect 70000 146354 70074 146410
rect 70130 146366 77808 146410
rect 77864 146366 77932 146422
rect 77988 146366 78056 146422
rect 78112 146366 78180 146422
rect 78236 146366 78304 146422
rect 78360 146366 78428 146422
rect 78484 146366 78552 146422
rect 78608 146366 78678 146422
rect 70130 146354 78678 146366
rect 70000 146298 78678 146354
rect 70000 146286 77808 146298
rect 70000 146230 70074 146286
rect 70130 146242 77808 146286
rect 77864 146242 77932 146298
rect 77988 146242 78056 146298
rect 78112 146242 78180 146298
rect 78236 146242 78304 146298
rect 78360 146242 78428 146298
rect 78484 146242 78552 146298
rect 78608 146242 78678 146298
rect 70130 146230 78678 146242
rect 70000 146174 78678 146230
rect 70000 146162 77808 146174
rect 70000 146106 70074 146162
rect 70130 146118 77808 146162
rect 77864 146118 77932 146174
rect 77988 146118 78056 146174
rect 78112 146118 78180 146174
rect 78236 146118 78304 146174
rect 78360 146118 78428 146174
rect 78484 146118 78552 146174
rect 78608 146118 78678 146174
rect 70130 146106 78678 146118
rect 70000 146050 78678 146106
rect 70000 146038 77808 146050
rect 70000 145982 70074 146038
rect 70130 145994 77808 146038
rect 77864 145994 77932 146050
rect 77988 145994 78056 146050
rect 78112 145994 78180 146050
rect 78236 145994 78304 146050
rect 78360 145994 78428 146050
rect 78484 145994 78552 146050
rect 78608 145994 78678 146050
rect 70130 145982 78678 145994
rect 70000 145926 78678 145982
rect 70000 145914 77808 145926
rect 70000 145858 70074 145914
rect 70130 145870 77808 145914
rect 77864 145870 77932 145926
rect 77988 145870 78056 145926
rect 78112 145870 78180 145926
rect 78236 145870 78304 145926
rect 78360 145870 78428 145926
rect 78484 145870 78552 145926
rect 78608 145870 78678 145926
rect 666132 146063 700322 146205
rect 666132 146007 699444 146063
rect 699500 146007 699744 146063
rect 699800 146007 700044 146063
rect 700100 146007 700322 146063
rect 666132 145885 700322 146007
rect 70130 145858 78678 145870
rect 70000 145802 78678 145858
rect 70000 145790 77808 145802
rect 70000 145734 70074 145790
rect 70130 145746 77808 145790
rect 77864 145746 77932 145802
rect 77988 145746 78056 145802
rect 78112 145746 78180 145802
rect 78236 145746 78304 145802
rect 78360 145746 78428 145802
rect 78484 145746 78552 145802
rect 78608 145746 78678 145802
rect 70130 145734 78678 145746
rect 70000 145678 78678 145734
rect 70000 145666 77808 145678
rect 70000 145610 70074 145666
rect 70130 145622 77808 145666
rect 77864 145622 77932 145678
rect 77988 145622 78056 145678
rect 78112 145622 78180 145678
rect 78236 145622 78304 145678
rect 78360 145622 78428 145678
rect 78484 145622 78552 145678
rect 78608 145622 78678 145678
rect 70130 145610 78678 145622
rect 70000 145554 78678 145610
rect 70000 145542 77808 145554
rect 70000 145486 70074 145542
rect 70130 145498 77808 145542
rect 77864 145498 77932 145554
rect 77988 145498 78056 145554
rect 78112 145498 78180 145554
rect 78236 145498 78304 145554
rect 78360 145498 78428 145554
rect 78484 145498 78552 145554
rect 78608 145498 78678 145554
rect 70130 145486 78678 145498
rect 70000 145430 78678 145486
rect 70000 145418 77808 145430
rect 70000 145362 70074 145418
rect 70130 145374 77808 145418
rect 77864 145374 77932 145430
rect 77988 145374 78056 145430
rect 78112 145374 78180 145430
rect 78236 145374 78304 145430
rect 78360 145374 78428 145430
rect 78484 145374 78552 145430
rect 78608 145374 78678 145430
rect 70130 145362 78678 145374
rect 70000 145306 78678 145362
rect 70000 145294 77808 145306
rect 70000 145238 70074 145294
rect 70130 145250 77808 145294
rect 77864 145250 77932 145306
rect 77988 145250 78056 145306
rect 78112 145250 78180 145306
rect 78236 145250 78304 145306
rect 78360 145250 78428 145306
rect 78484 145250 78552 145306
rect 78608 145250 78678 145306
rect 70130 145238 78678 145250
rect 70000 145182 78678 145238
rect 70000 145170 77808 145182
rect 70000 145114 70074 145170
rect 70130 145126 77808 145170
rect 77864 145126 77932 145182
rect 77988 145126 78056 145182
rect 78112 145126 78180 145182
rect 78236 145126 78304 145182
rect 78360 145126 78428 145182
rect 78484 145126 78552 145182
rect 78608 145126 78678 145182
rect 70130 145114 78678 145126
rect 70000 145058 78678 145114
rect 70000 145046 77808 145058
rect 70000 144990 70074 145046
rect 70130 145002 77808 145046
rect 77864 145002 77932 145058
rect 77988 145002 78056 145058
rect 78112 145002 78180 145058
rect 78236 145002 78304 145058
rect 78360 145002 78428 145058
rect 78484 145002 78552 145058
rect 78608 145002 78678 145058
rect 70130 144990 78678 145002
rect 70000 144934 78678 144990
rect 70000 144922 77808 144934
rect 70000 144866 70074 144922
rect 70130 144878 77808 144922
rect 77864 144878 77932 144934
rect 77988 144878 78056 144934
rect 78112 144878 78180 144934
rect 78236 144878 78304 144934
rect 78360 144878 78428 144934
rect 78484 144878 78552 144934
rect 78608 144878 78678 144934
rect 70130 144866 78678 144878
rect 70000 144828 78678 144866
rect 699322 144954 702688 145076
rect 699322 144898 699444 144954
rect 699500 144898 699744 144954
rect 699800 144898 700044 144954
rect 700100 144898 702688 144954
rect 699322 144756 702688 144898
rect 70000 144190 78678 144248
rect 70000 144184 77808 144190
rect 70000 144128 70074 144184
rect 70130 144134 77808 144184
rect 77864 144134 77932 144190
rect 77988 144134 78056 144190
rect 78112 144134 78180 144190
rect 78236 144134 78304 144190
rect 78360 144134 78428 144190
rect 78484 144134 78552 144190
rect 78608 144134 78678 144190
rect 70130 144128 78678 144134
rect 70000 144066 78678 144128
rect 70000 144060 77808 144066
rect 70000 144004 70074 144060
rect 70130 144010 77808 144060
rect 77864 144010 77932 144066
rect 77988 144010 78056 144066
rect 78112 144010 78180 144066
rect 78236 144010 78304 144066
rect 78360 144010 78428 144066
rect 78484 144010 78552 144066
rect 78608 144010 78678 144066
rect 70130 144004 78678 144010
rect 70000 143942 78678 144004
rect 70000 143936 77808 143942
rect 70000 143880 70074 143936
rect 70130 143886 77808 143936
rect 77864 143886 77932 143942
rect 77988 143886 78056 143942
rect 78112 143886 78180 143942
rect 78236 143886 78304 143942
rect 78360 143886 78428 143942
rect 78484 143886 78552 143942
rect 78608 143886 78678 143942
rect 70130 143880 78678 143886
rect 70000 143818 78678 143880
rect 70000 143812 77808 143818
rect 70000 143756 70074 143812
rect 70130 143762 77808 143812
rect 77864 143762 77932 143818
rect 77988 143762 78056 143818
rect 78112 143762 78180 143818
rect 78236 143762 78304 143818
rect 78360 143762 78428 143818
rect 78484 143762 78552 143818
rect 78608 143762 78678 143818
rect 70130 143756 78678 143762
rect 70000 143694 78678 143756
rect 70000 143688 77808 143694
rect 70000 143632 70074 143688
rect 70130 143638 77808 143688
rect 77864 143638 77932 143694
rect 77988 143638 78056 143694
rect 78112 143638 78180 143694
rect 78236 143638 78304 143694
rect 78360 143638 78428 143694
rect 78484 143638 78552 143694
rect 78608 143638 78678 143694
rect 70130 143632 78678 143638
rect 70000 143570 78678 143632
rect 70000 143564 77808 143570
rect 70000 143508 70074 143564
rect 70130 143514 77808 143564
rect 77864 143514 77932 143570
rect 77988 143514 78056 143570
rect 78112 143514 78180 143570
rect 78236 143514 78304 143570
rect 78360 143514 78428 143570
rect 78484 143514 78552 143570
rect 78608 143514 78678 143570
rect 70130 143508 78678 143514
rect 70000 143446 78678 143508
rect 70000 143440 77808 143446
rect 70000 143384 70074 143440
rect 70130 143390 77808 143440
rect 77864 143390 77932 143446
rect 77988 143390 78056 143446
rect 78112 143390 78180 143446
rect 78236 143390 78304 143446
rect 78360 143390 78428 143446
rect 78484 143390 78552 143446
rect 78608 143390 78678 143446
rect 70130 143384 78678 143390
rect 70000 143322 78678 143384
rect 70000 143316 77808 143322
rect 70000 143260 70074 143316
rect 70130 143266 77808 143316
rect 77864 143266 77932 143322
rect 77988 143266 78056 143322
rect 78112 143266 78180 143322
rect 78236 143266 78304 143322
rect 78360 143266 78428 143322
rect 78484 143266 78552 143322
rect 78608 143266 78678 143322
rect 70130 143260 78678 143266
rect 70000 143198 78678 143260
rect 70000 143192 77808 143198
rect 70000 143136 70074 143192
rect 70130 143142 77808 143192
rect 77864 143142 77932 143198
rect 77988 143142 78056 143198
rect 78112 143142 78180 143198
rect 78236 143142 78304 143198
rect 78360 143142 78428 143198
rect 78484 143142 78552 143198
rect 78608 143142 78678 143198
rect 70130 143136 78678 143142
rect 70000 143074 78678 143136
rect 70000 143068 77808 143074
rect 70000 143012 70074 143068
rect 70130 143018 77808 143068
rect 77864 143018 77932 143074
rect 77988 143018 78056 143074
rect 78112 143018 78180 143074
rect 78236 143018 78304 143074
rect 78360 143018 78428 143074
rect 78484 143018 78552 143074
rect 78608 143018 78678 143074
rect 70130 143012 78678 143018
rect 70000 142950 78678 143012
rect 70000 142944 77808 142950
rect 70000 142888 70074 142944
rect 70130 142894 77808 142944
rect 77864 142894 77932 142950
rect 77988 142894 78056 142950
rect 78112 142894 78180 142950
rect 78236 142894 78304 142950
rect 78360 142894 78428 142950
rect 78484 142894 78552 142950
rect 78608 142894 78678 142950
rect 70130 142888 78678 142894
rect 70000 142826 78678 142888
rect 70000 142820 77808 142826
rect 70000 142764 70074 142820
rect 70130 142770 77808 142820
rect 77864 142770 77932 142826
rect 77988 142770 78056 142826
rect 78112 142770 78180 142826
rect 78236 142770 78304 142826
rect 78360 142770 78428 142826
rect 78484 142770 78552 142826
rect 78608 142770 78678 142826
rect 70130 142764 78678 142770
rect 70000 142702 78678 142764
rect 70000 142696 77808 142702
rect 70000 142640 70074 142696
rect 70130 142646 77808 142696
rect 77864 142646 77932 142702
rect 77988 142646 78056 142702
rect 78112 142646 78180 142702
rect 78236 142646 78304 142702
rect 78360 142646 78428 142702
rect 78484 142646 78552 142702
rect 78608 142646 78678 142702
rect 70130 142640 78678 142646
rect 70000 142578 78678 142640
rect 70000 142572 77808 142578
rect 70000 142516 70074 142572
rect 70130 142522 77808 142572
rect 77864 142522 77932 142578
rect 77988 142522 78056 142578
rect 78112 142522 78180 142578
rect 78236 142522 78304 142578
rect 78360 142522 78428 142578
rect 78484 142522 78552 142578
rect 78608 142522 78678 142578
rect 70130 142516 78678 142522
rect 70000 142454 78678 142516
rect 70000 142448 77808 142454
rect 70000 142392 70074 142448
rect 70130 142398 77808 142448
rect 77864 142398 77932 142454
rect 77988 142398 78056 142454
rect 78112 142398 78180 142454
rect 78236 142398 78304 142454
rect 78360 142398 78428 142454
rect 78484 142398 78552 142454
rect 78608 142398 78678 142454
rect 70130 142392 78678 142398
rect 70000 142330 78678 142392
rect 70000 142324 77808 142330
rect 70000 142268 70074 142324
rect 70130 142274 77808 142324
rect 77864 142274 77932 142330
rect 77988 142274 78056 142330
rect 78112 142274 78180 142330
rect 78236 142274 78304 142330
rect 78360 142274 78428 142330
rect 78484 142274 78552 142330
rect 78608 142274 78678 142330
rect 70130 142268 78678 142274
rect 70000 142198 78678 142268
rect 70000 141820 78678 141878
rect 70000 141814 77808 141820
rect 70000 141758 70074 141814
rect 70130 141764 77808 141814
rect 77864 141764 77932 141820
rect 77988 141764 78056 141820
rect 78112 141764 78180 141820
rect 78236 141764 78304 141820
rect 78360 141764 78428 141820
rect 78484 141764 78552 141820
rect 78608 141764 78678 141820
rect 70130 141758 78678 141764
rect 70000 141696 78678 141758
rect 70000 141690 77808 141696
rect 70000 141634 70074 141690
rect 70130 141640 77808 141690
rect 77864 141640 77932 141696
rect 77988 141640 78056 141696
rect 78112 141640 78180 141696
rect 78236 141640 78304 141696
rect 78360 141640 78428 141696
rect 78484 141640 78552 141696
rect 78608 141640 78678 141696
rect 70130 141634 78678 141640
rect 70000 141572 78678 141634
rect 70000 141566 77808 141572
rect 70000 141510 70074 141566
rect 70130 141516 77808 141566
rect 77864 141516 77932 141572
rect 77988 141516 78056 141572
rect 78112 141516 78180 141572
rect 78236 141516 78304 141572
rect 78360 141516 78428 141572
rect 78484 141516 78552 141572
rect 78608 141516 78678 141572
rect 70130 141510 78678 141516
rect 70000 141448 78678 141510
rect 70000 141442 77808 141448
rect 70000 141386 70074 141442
rect 70130 141392 77808 141442
rect 77864 141392 77932 141448
rect 77988 141392 78056 141448
rect 78112 141392 78180 141448
rect 78236 141392 78304 141448
rect 78360 141392 78428 141448
rect 78484 141392 78552 141448
rect 78608 141392 78678 141448
rect 70130 141386 78678 141392
rect 70000 141324 78678 141386
rect 70000 141318 77808 141324
rect 70000 141262 70074 141318
rect 70130 141268 77808 141318
rect 77864 141268 77932 141324
rect 77988 141268 78056 141324
rect 78112 141268 78180 141324
rect 78236 141268 78304 141324
rect 78360 141268 78428 141324
rect 78484 141268 78552 141324
rect 78608 141268 78678 141324
rect 70130 141262 78678 141268
rect 70000 141200 78678 141262
rect 697922 141434 702624 141576
rect 697922 141378 698044 141434
rect 698100 141378 698344 141434
rect 698400 141378 698644 141434
rect 698700 141378 702624 141434
rect 697922 141256 702624 141378
rect 70000 141194 77808 141200
rect 70000 141138 70074 141194
rect 70130 141144 77808 141194
rect 77864 141144 77932 141200
rect 77988 141144 78056 141200
rect 78112 141144 78180 141200
rect 78236 141144 78304 141200
rect 78360 141144 78428 141200
rect 78484 141144 78552 141200
rect 78608 141144 78678 141200
rect 70130 141138 78678 141144
rect 70000 141076 78678 141138
rect 70000 141070 77808 141076
rect 70000 141014 70074 141070
rect 70130 141020 77808 141070
rect 77864 141020 77932 141076
rect 77988 141020 78056 141076
rect 78112 141020 78180 141076
rect 78236 141020 78304 141076
rect 78360 141020 78428 141076
rect 78484 141020 78552 141076
rect 78608 141020 78678 141076
rect 70130 141014 78678 141020
rect 70000 140952 78678 141014
rect 70000 140946 77808 140952
rect 70000 140890 70074 140946
rect 70130 140896 77808 140946
rect 77864 140896 77932 140952
rect 77988 140896 78056 140952
rect 78112 140896 78180 140952
rect 78236 140896 78304 140952
rect 78360 140896 78428 140952
rect 78484 140896 78552 140952
rect 78608 140896 78678 140952
rect 70130 140890 78678 140896
rect 70000 140828 78678 140890
rect 70000 140822 77808 140828
rect 70000 140766 70074 140822
rect 70130 140772 77808 140822
rect 77864 140772 77932 140828
rect 77988 140772 78056 140828
rect 78112 140772 78180 140828
rect 78236 140772 78304 140828
rect 78360 140772 78428 140828
rect 78484 140772 78552 140828
rect 78608 140772 78678 140828
rect 70130 140766 78678 140772
rect 70000 140704 78678 140766
rect 70000 140698 77808 140704
rect 70000 140642 70074 140698
rect 70130 140648 77808 140698
rect 77864 140648 77932 140704
rect 77988 140648 78056 140704
rect 78112 140648 78180 140704
rect 78236 140648 78304 140704
rect 78360 140648 78428 140704
rect 78484 140648 78552 140704
rect 78608 140648 78678 140704
rect 70130 140642 78678 140648
rect 70000 140580 78678 140642
rect 70000 140574 77808 140580
rect 70000 140518 70074 140574
rect 70130 140524 77808 140574
rect 77864 140524 77932 140580
rect 77988 140524 78056 140580
rect 78112 140524 78180 140580
rect 78236 140524 78304 140580
rect 78360 140524 78428 140580
rect 78484 140524 78552 140580
rect 78608 140524 78678 140580
rect 70130 140518 78678 140524
rect 70000 140456 78678 140518
rect 70000 140450 77808 140456
rect 70000 140394 70074 140450
rect 70130 140400 77808 140450
rect 77864 140400 77932 140456
rect 77988 140400 78056 140456
rect 78112 140400 78180 140456
rect 78236 140400 78304 140456
rect 78360 140400 78428 140456
rect 78484 140400 78552 140456
rect 78608 140400 78678 140456
rect 70130 140394 78678 140400
rect 70000 140332 78678 140394
rect 70000 140326 77808 140332
rect 70000 140270 70074 140326
rect 70130 140276 77808 140326
rect 77864 140276 77932 140332
rect 77988 140276 78056 140332
rect 78112 140276 78180 140332
rect 78236 140276 78304 140332
rect 78360 140276 78428 140332
rect 78484 140276 78552 140332
rect 78608 140276 78678 140332
rect 70130 140270 78678 140276
rect 70000 140208 78678 140270
rect 70000 140202 77808 140208
rect 70000 140146 70074 140202
rect 70130 140152 77808 140202
rect 77864 140152 77932 140208
rect 77988 140152 78056 140208
rect 78112 140152 78180 140208
rect 78236 140152 78304 140208
rect 78360 140152 78428 140208
rect 78484 140152 78552 140208
rect 78608 140152 78678 140208
rect 70130 140146 78678 140152
rect 70000 140084 78678 140146
rect 70000 140078 77808 140084
rect 70000 140022 70074 140078
rect 70130 140028 77808 140078
rect 77864 140028 77932 140084
rect 77988 140028 78056 140084
rect 78112 140028 78180 140084
rect 78236 140028 78304 140084
rect 78360 140028 78428 140084
rect 78484 140028 78552 140084
rect 78608 140028 78678 140084
rect 70130 140022 78678 140028
rect 70000 139960 78678 140022
rect 70000 139954 77808 139960
rect 70000 139898 70074 139954
rect 70130 139904 77808 139954
rect 77864 139904 77932 139960
rect 77988 139904 78056 139960
rect 78112 139904 78180 139960
rect 78236 139904 78304 139960
rect 78360 139904 78428 139960
rect 78484 139904 78552 139960
rect 78608 139904 78678 139960
rect 70130 139898 78678 139904
rect 70000 139828 78678 139898
rect 70000 139114 78678 139172
rect 70000 139108 77808 139114
rect 70000 139052 70074 139108
rect 70130 139058 77808 139108
rect 77864 139058 77932 139114
rect 77988 139058 78056 139114
rect 78112 139058 78180 139114
rect 78236 139058 78304 139114
rect 78360 139058 78428 139114
rect 78484 139058 78552 139114
rect 78608 139058 78678 139114
rect 70130 139052 78678 139058
rect 70000 138990 78678 139052
rect 70000 138984 77808 138990
rect 70000 138928 70074 138984
rect 70130 138934 77808 138984
rect 77864 138934 77932 138990
rect 77988 138934 78056 138990
rect 78112 138934 78180 138990
rect 78236 138934 78304 138990
rect 78360 138934 78428 138990
rect 78484 138934 78552 138990
rect 78608 138934 78678 138990
rect 70130 138928 78678 138934
rect 70000 138866 78678 138928
rect 70000 138860 77808 138866
rect 70000 138804 70074 138860
rect 70130 138810 77808 138860
rect 77864 138810 77932 138866
rect 77988 138810 78056 138866
rect 78112 138810 78180 138866
rect 78236 138810 78304 138866
rect 78360 138810 78428 138866
rect 78484 138810 78552 138866
rect 78608 138810 78678 138866
rect 70130 138804 78678 138810
rect 70000 138742 78678 138804
rect 70000 138736 77808 138742
rect 70000 138680 70074 138736
rect 70130 138686 77808 138736
rect 77864 138686 77932 138742
rect 77988 138686 78056 138742
rect 78112 138686 78180 138742
rect 78236 138686 78304 138742
rect 78360 138686 78428 138742
rect 78484 138686 78552 138742
rect 78608 138686 78678 138742
rect 70130 138680 78678 138686
rect 70000 138618 78678 138680
rect 70000 138612 77808 138618
rect 70000 138556 70074 138612
rect 70130 138562 77808 138612
rect 77864 138562 77932 138618
rect 77988 138562 78056 138618
rect 78112 138562 78180 138618
rect 78236 138562 78304 138618
rect 78360 138562 78428 138618
rect 78484 138562 78552 138618
rect 78608 138562 78678 138618
rect 70130 138556 78678 138562
rect 70000 138494 78678 138556
rect 70000 138488 77808 138494
rect 70000 138432 70074 138488
rect 70130 138438 77808 138488
rect 77864 138438 77932 138494
rect 77988 138438 78056 138494
rect 78112 138438 78180 138494
rect 78236 138438 78304 138494
rect 78360 138438 78428 138494
rect 78484 138438 78552 138494
rect 78608 138438 78678 138494
rect 70130 138432 78678 138438
rect 70000 138370 78678 138432
rect 70000 138364 77808 138370
rect 70000 138308 70074 138364
rect 70130 138314 77808 138364
rect 77864 138314 77932 138370
rect 77988 138314 78056 138370
rect 78112 138314 78180 138370
rect 78236 138314 78304 138370
rect 78360 138314 78428 138370
rect 78484 138314 78552 138370
rect 78608 138314 78678 138370
rect 70130 138308 78678 138314
rect 70000 138246 78678 138308
rect 70000 138240 77808 138246
rect 70000 138184 70074 138240
rect 70130 138190 77808 138240
rect 77864 138190 77932 138246
rect 77988 138190 78056 138246
rect 78112 138190 78180 138246
rect 78236 138190 78304 138246
rect 78360 138190 78428 138246
rect 78484 138190 78552 138246
rect 78608 138190 78678 138246
rect 70130 138184 78678 138190
rect 70000 138122 78678 138184
rect 560032 138372 593240 138442
rect 560032 138316 592370 138372
rect 592426 138316 592494 138372
rect 592550 138316 592618 138372
rect 592674 138316 592742 138372
rect 592798 138316 592866 138372
rect 592922 138316 592990 138372
rect 593046 138316 593114 138372
rect 593170 138316 593240 138372
rect 560032 138248 593240 138316
rect 560032 138192 592370 138248
rect 592426 138192 592494 138248
rect 592550 138192 592618 138248
rect 592674 138192 592742 138248
rect 592798 138192 592866 138248
rect 592922 138192 592990 138248
rect 593046 138192 593114 138248
rect 593170 138192 593240 138248
rect 560032 138122 593240 138192
rect 70000 138116 77808 138122
rect 70000 138060 70074 138116
rect 70130 138066 77808 138116
rect 77864 138066 77932 138122
rect 77988 138066 78056 138122
rect 78112 138066 78180 138122
rect 78236 138066 78304 138122
rect 78360 138066 78428 138122
rect 78484 138066 78552 138122
rect 78608 138066 78678 138122
rect 70130 138060 78678 138066
rect 70000 137998 78678 138060
rect 70000 137992 77808 137998
rect 70000 137936 70074 137992
rect 70130 137942 77808 137992
rect 77864 137942 77932 137998
rect 77988 137942 78056 137998
rect 78112 137942 78180 137998
rect 78236 137942 78304 137998
rect 78360 137942 78428 137998
rect 78484 137942 78552 137998
rect 78608 137942 78678 137998
rect 70130 137936 78678 137942
rect 70000 137874 78678 137936
rect 70000 137868 77808 137874
rect 70000 137812 70074 137868
rect 70130 137818 77808 137868
rect 77864 137818 77932 137874
rect 77988 137818 78056 137874
rect 78112 137818 78180 137874
rect 78236 137818 78304 137874
rect 78360 137818 78428 137874
rect 78484 137818 78552 137874
rect 78608 137818 78678 137874
rect 70130 137812 78678 137818
rect 70000 137750 78678 137812
rect 699322 137954 702688 138076
rect 699322 137898 699444 137954
rect 699500 137898 699744 137954
rect 699800 137898 700044 137954
rect 700100 137898 702688 137954
rect 699322 137756 702688 137898
rect 70000 137744 77808 137750
rect 70000 137688 70074 137744
rect 70130 137694 77808 137744
rect 77864 137694 77932 137750
rect 77988 137694 78056 137750
rect 78112 137694 78180 137750
rect 78236 137694 78304 137750
rect 78360 137694 78428 137750
rect 78484 137694 78552 137750
rect 78608 137694 78678 137750
rect 70130 137688 78678 137694
rect 70000 137626 78678 137688
rect 70000 137620 77808 137626
rect 70000 137564 70074 137620
rect 70130 137570 77808 137620
rect 77864 137570 77932 137626
rect 77988 137570 78056 137626
rect 78112 137570 78180 137626
rect 78236 137570 78304 137626
rect 78360 137570 78428 137626
rect 78484 137570 78552 137626
rect 78608 137570 78678 137626
rect 70130 137564 78678 137570
rect 70000 137502 78678 137564
rect 70000 137496 77808 137502
rect 70000 137440 70074 137496
rect 70130 137446 77808 137496
rect 77864 137446 77932 137502
rect 77988 137446 78056 137502
rect 78112 137446 78180 137502
rect 78236 137446 78304 137502
rect 78360 137446 78428 137502
rect 78484 137446 78552 137502
rect 78608 137446 78678 137502
rect 70130 137440 78678 137446
rect 70000 137378 78678 137440
rect 70000 137372 77808 137378
rect 70000 137316 70074 137372
rect 70130 137322 77808 137372
rect 77864 137322 77932 137378
rect 77988 137322 78056 137378
rect 78112 137322 78180 137378
rect 78236 137322 78304 137378
rect 78360 137322 78428 137378
rect 78484 137322 78552 137378
rect 78608 137322 78678 137378
rect 70130 137316 78678 137322
rect 70000 137254 78678 137316
rect 70000 137248 77808 137254
rect 70000 137192 70074 137248
rect 70130 137198 77808 137248
rect 77864 137198 77932 137254
rect 77988 137198 78056 137254
rect 78112 137198 78180 137254
rect 78236 137198 78304 137254
rect 78360 137198 78428 137254
rect 78484 137198 78552 137254
rect 78608 137198 78678 137254
rect 70130 137192 78678 137198
rect 70000 137122 78678 137192
rect 70000 136744 78678 136802
rect 70000 136738 77808 136744
rect 70000 136682 70074 136738
rect 70130 136688 77808 136738
rect 77864 136688 77932 136744
rect 77988 136688 78056 136744
rect 78112 136688 78180 136744
rect 78236 136688 78304 136744
rect 78360 136688 78428 136744
rect 78484 136688 78552 136744
rect 78608 136688 78678 136744
rect 70130 136682 78678 136688
rect 70000 136620 78678 136682
rect 70000 136614 77808 136620
rect 70000 136558 70074 136614
rect 70130 136564 77808 136614
rect 77864 136564 77932 136620
rect 77988 136564 78056 136620
rect 78112 136564 78180 136620
rect 78236 136564 78304 136620
rect 78360 136564 78428 136620
rect 78484 136564 78552 136620
rect 78608 136564 78678 136620
rect 70130 136558 78678 136564
rect 70000 136496 78678 136558
rect 70000 136490 77808 136496
rect 70000 136434 70074 136490
rect 70130 136440 77808 136490
rect 77864 136440 77932 136496
rect 77988 136440 78056 136496
rect 78112 136440 78180 136496
rect 78236 136440 78304 136496
rect 78360 136440 78428 136496
rect 78484 136440 78552 136496
rect 78608 136440 78678 136496
rect 70130 136434 78678 136440
rect 70000 136372 78678 136434
rect 70000 136366 77808 136372
rect 70000 136310 70074 136366
rect 70130 136316 77808 136366
rect 77864 136316 77932 136372
rect 77988 136316 78056 136372
rect 78112 136316 78180 136372
rect 78236 136316 78304 136372
rect 78360 136316 78428 136372
rect 78484 136316 78552 136372
rect 78608 136316 78678 136372
rect 70130 136310 78678 136316
rect 70000 136248 78678 136310
rect 70000 136242 77808 136248
rect 70000 136186 70074 136242
rect 70130 136192 77808 136242
rect 77864 136192 77932 136248
rect 77988 136192 78056 136248
rect 78112 136192 78180 136248
rect 78236 136192 78304 136248
rect 78360 136192 78428 136248
rect 78484 136192 78552 136248
rect 78608 136192 78678 136248
rect 70130 136186 78678 136192
rect 70000 136124 78678 136186
rect 70000 136118 77808 136124
rect 70000 136062 70074 136118
rect 70130 136068 77808 136118
rect 77864 136068 77932 136124
rect 77988 136068 78056 136124
rect 78112 136068 78180 136124
rect 78236 136068 78304 136124
rect 78360 136068 78428 136124
rect 78484 136068 78552 136124
rect 78608 136068 78678 136124
rect 70130 136062 78678 136068
rect 70000 136000 78678 136062
rect 70000 135994 77808 136000
rect 70000 135938 70074 135994
rect 70130 135944 77808 135994
rect 77864 135944 77932 136000
rect 77988 135944 78056 136000
rect 78112 135944 78180 136000
rect 78236 135944 78304 136000
rect 78360 135944 78428 136000
rect 78484 135944 78552 136000
rect 78608 135944 78678 136000
rect 70130 135938 78678 135944
rect 70000 135876 78678 135938
rect 70000 135870 77808 135876
rect 70000 135814 70074 135870
rect 70130 135820 77808 135870
rect 77864 135820 77932 135876
rect 77988 135820 78056 135876
rect 78112 135820 78180 135876
rect 78236 135820 78304 135876
rect 78360 135820 78428 135876
rect 78484 135820 78552 135876
rect 78608 135820 78678 135876
rect 70130 135814 78678 135820
rect 70000 135752 78678 135814
rect 70000 135746 77808 135752
rect 70000 135690 70074 135746
rect 70130 135696 77808 135746
rect 77864 135696 77932 135752
rect 77988 135696 78056 135752
rect 78112 135696 78180 135752
rect 78236 135696 78304 135752
rect 78360 135696 78428 135752
rect 78484 135696 78552 135752
rect 78608 135696 78678 135752
rect 70130 135690 78678 135696
rect 70000 135628 78678 135690
rect 70000 135622 77808 135628
rect 70000 135566 70074 135622
rect 70130 135572 77808 135622
rect 77864 135572 77932 135628
rect 77988 135572 78056 135628
rect 78112 135572 78180 135628
rect 78236 135572 78304 135628
rect 78360 135572 78428 135628
rect 78484 135572 78552 135628
rect 78608 135572 78678 135628
rect 70130 135566 78678 135572
rect 70000 135504 78678 135566
rect 70000 135498 77808 135504
rect 70000 135442 70074 135498
rect 70130 135448 77808 135498
rect 77864 135448 77932 135504
rect 77988 135448 78056 135504
rect 78112 135448 78180 135504
rect 78236 135448 78304 135504
rect 78360 135448 78428 135504
rect 78484 135448 78552 135504
rect 78608 135448 78678 135504
rect 70130 135442 78678 135448
rect 70000 135380 78678 135442
rect 70000 135374 77808 135380
rect 70000 135318 70074 135374
rect 70130 135324 77808 135374
rect 77864 135324 77932 135380
rect 77988 135324 78056 135380
rect 78112 135324 78180 135380
rect 78236 135324 78304 135380
rect 78360 135324 78428 135380
rect 78484 135324 78552 135380
rect 78608 135324 78678 135380
rect 70130 135318 78678 135324
rect 70000 135256 78678 135318
rect 70000 135250 77808 135256
rect 70000 135194 70074 135250
rect 70130 135200 77808 135250
rect 77864 135200 77932 135256
rect 77988 135200 78056 135256
rect 78112 135200 78180 135256
rect 78236 135200 78304 135256
rect 78360 135200 78428 135256
rect 78484 135200 78552 135256
rect 78608 135200 78678 135256
rect 70130 135194 78678 135200
rect 70000 135132 78678 135194
rect 70000 135126 77808 135132
rect 70000 135070 70074 135126
rect 70130 135076 77808 135126
rect 77864 135076 77932 135132
rect 77988 135076 78056 135132
rect 78112 135076 78180 135132
rect 78236 135076 78304 135132
rect 78360 135076 78428 135132
rect 78484 135076 78552 135132
rect 78608 135076 78678 135132
rect 70130 135070 78678 135076
rect 70000 135008 78678 135070
rect 70000 135002 77808 135008
rect 70000 134946 70074 135002
rect 70130 134952 77808 135002
rect 77864 134952 77932 135008
rect 77988 134952 78056 135008
rect 78112 134952 78180 135008
rect 78236 134952 78304 135008
rect 78360 134952 78428 135008
rect 78484 134952 78552 135008
rect 78608 134952 78678 135008
rect 70130 134946 78678 134952
rect 70000 134884 78678 134946
rect 70000 134878 77808 134884
rect 70000 134822 70074 134878
rect 70130 134828 77808 134878
rect 77864 134828 77932 134884
rect 77988 134828 78056 134884
rect 78112 134828 78180 134884
rect 78236 134828 78304 134884
rect 78360 134828 78428 134884
rect 78484 134828 78552 134884
rect 78608 134828 78678 134884
rect 70130 134822 78678 134828
rect 70000 134752 78678 134822
rect 697922 134418 702624 134576
rect 697922 134362 698044 134418
rect 698100 134362 698344 134418
rect 698400 134362 698644 134418
rect 698700 134362 702624 134418
rect 697922 134256 702624 134362
rect 70000 134140 78678 134172
rect 70000 134134 77808 134140
rect 70000 134078 70074 134134
rect 70130 134084 77808 134134
rect 77864 134084 77932 134140
rect 77988 134084 78056 134140
rect 78112 134084 78180 134140
rect 78236 134084 78304 134140
rect 78360 134084 78428 134140
rect 78484 134084 78552 134140
rect 78608 134084 78678 134140
rect 70130 134078 78678 134084
rect 70000 134016 78678 134078
rect 70000 134010 77808 134016
rect 70000 133954 70074 134010
rect 70130 133960 77808 134010
rect 77864 133960 77932 134016
rect 77988 133960 78056 134016
rect 78112 133960 78180 134016
rect 78236 133960 78304 134016
rect 78360 133960 78428 134016
rect 78484 133960 78552 134016
rect 78608 133960 78678 134016
rect 70130 133954 78678 133960
rect 70000 133892 78678 133954
rect 70000 133886 77808 133892
rect 70000 133830 70074 133886
rect 70130 133836 77808 133886
rect 77864 133836 77932 133892
rect 77988 133836 78056 133892
rect 78112 133836 78180 133892
rect 78236 133836 78304 133892
rect 78360 133836 78428 133892
rect 78484 133836 78552 133892
rect 78608 133836 78678 133892
rect 70130 133830 78678 133836
rect 70000 133768 78678 133830
rect 70000 133762 77808 133768
rect 70000 133706 70074 133762
rect 70130 133712 77808 133762
rect 77864 133712 77932 133768
rect 77988 133712 78056 133768
rect 78112 133712 78180 133768
rect 78236 133712 78304 133768
rect 78360 133712 78428 133768
rect 78484 133712 78552 133768
rect 78608 133712 78678 133768
rect 70130 133706 78678 133712
rect 70000 133644 78678 133706
rect 70000 133638 77808 133644
rect 70000 133582 70074 133638
rect 70130 133588 77808 133638
rect 77864 133588 77932 133644
rect 77988 133588 78056 133644
rect 78112 133588 78180 133644
rect 78236 133588 78304 133644
rect 78360 133588 78428 133644
rect 78484 133588 78552 133644
rect 78608 133588 78678 133644
rect 670161 133803 700322 133945
rect 670161 133747 699444 133803
rect 699500 133747 699744 133803
rect 699800 133747 700044 133803
rect 700100 133747 700322 133803
rect 670161 133625 700322 133747
rect 70130 133582 78678 133588
rect 70000 133520 78678 133582
rect 70000 133514 77808 133520
rect 70000 133458 70074 133514
rect 70130 133464 77808 133514
rect 77864 133464 77932 133520
rect 77988 133464 78056 133520
rect 78112 133464 78180 133520
rect 78236 133464 78304 133520
rect 78360 133464 78428 133520
rect 78484 133464 78552 133520
rect 78608 133464 78678 133520
rect 70130 133458 78678 133464
rect 70000 133396 78678 133458
rect 70000 133390 77808 133396
rect 70000 133334 70074 133390
rect 70130 133340 77808 133390
rect 77864 133340 77932 133396
rect 77988 133340 78056 133396
rect 78112 133340 78180 133396
rect 78236 133340 78304 133396
rect 78360 133340 78428 133396
rect 78484 133340 78552 133396
rect 78608 133340 78678 133396
rect 70130 133334 78678 133340
rect 70000 133272 78678 133334
rect 70000 133266 77808 133272
rect 70000 133210 70074 133266
rect 70130 133216 77808 133266
rect 77864 133216 77932 133272
rect 77988 133216 78056 133272
rect 78112 133216 78180 133272
rect 78236 133216 78304 133272
rect 78360 133216 78428 133272
rect 78484 133216 78552 133272
rect 78608 133216 78678 133272
rect 70130 133210 78678 133216
rect 70000 133148 78678 133210
rect 70000 133142 77808 133148
rect 70000 133086 70074 133142
rect 70130 133092 77808 133142
rect 77864 133092 77932 133148
rect 77988 133092 78056 133148
rect 78112 133092 78180 133148
rect 78236 133092 78304 133148
rect 78360 133092 78428 133148
rect 78484 133092 78552 133148
rect 78608 133092 78678 133148
rect 70130 133086 78678 133092
rect 70000 133024 78678 133086
rect 70000 133018 77808 133024
rect 70000 132962 70074 133018
rect 70130 132968 77808 133018
rect 77864 132968 77932 133024
rect 77988 132968 78056 133024
rect 78112 132968 78180 133024
rect 78236 132968 78304 133024
rect 78360 132968 78428 133024
rect 78484 132968 78552 133024
rect 78608 132968 78678 133024
rect 70130 132962 78678 132968
rect 70000 132900 78678 132962
rect 70000 132894 77808 132900
rect 70000 132838 70074 132894
rect 70130 132844 77808 132894
rect 77864 132844 77932 132900
rect 77988 132844 78056 132900
rect 78112 132844 78180 132900
rect 78236 132844 78304 132900
rect 78360 132844 78428 132900
rect 78484 132844 78552 132900
rect 78608 132844 78678 132900
rect 70130 132838 78678 132844
rect 70000 132776 78678 132838
rect 670161 133003 698922 133145
rect 670161 132947 698044 133003
rect 698100 132947 698344 133003
rect 698400 132947 698644 133003
rect 698700 132947 698922 133003
rect 670161 132825 698922 132947
rect 70000 132770 77808 132776
rect 70000 132714 70074 132770
rect 70130 132720 77808 132770
rect 77864 132720 77932 132776
rect 77988 132720 78056 132776
rect 78112 132720 78180 132776
rect 78236 132720 78304 132776
rect 78360 132720 78428 132776
rect 78484 132720 78552 132776
rect 78608 132720 78678 132776
rect 70130 132714 78678 132720
rect 70000 132652 78678 132714
rect 70000 132646 77808 132652
rect 70000 132590 70074 132646
rect 70130 132596 77808 132646
rect 77864 132596 77932 132652
rect 77988 132596 78056 132652
rect 78112 132596 78180 132652
rect 78236 132596 78304 132652
rect 78360 132596 78428 132652
rect 78484 132596 78552 132652
rect 78608 132596 78678 132652
rect 70130 132590 78678 132596
rect 70000 132528 78678 132590
rect 70000 132522 77808 132528
rect 70000 132466 70074 132522
rect 70130 132472 77808 132522
rect 77864 132472 77932 132528
rect 77988 132472 78056 132528
rect 78112 132472 78180 132528
rect 78236 132472 78304 132528
rect 78360 132472 78428 132528
rect 78484 132472 78552 132528
rect 78608 132472 78678 132528
rect 70130 132466 78678 132472
rect 70000 132404 78678 132466
rect 70000 132398 77808 132404
rect 70000 132342 70074 132398
rect 70130 132348 77808 132398
rect 77864 132348 77932 132404
rect 77988 132348 78056 132404
rect 78112 132348 78180 132404
rect 78236 132348 78304 132404
rect 78360 132348 78428 132404
rect 78484 132348 78552 132404
rect 78608 132348 78678 132404
rect 70130 132342 78678 132348
rect 70000 132272 78678 132342
rect 79078 125372 89920 125442
rect 79078 125316 79148 125372
rect 79204 125316 79272 125372
rect 79328 125316 79396 125372
rect 79452 125316 79520 125372
rect 79576 125316 79644 125372
rect 79700 125316 79768 125372
rect 79824 125316 79892 125372
rect 79948 125316 89920 125372
rect 79078 125248 89920 125316
rect 79078 125192 79148 125248
rect 79204 125192 79272 125248
rect 79328 125192 79396 125248
rect 79452 125192 79520 125248
rect 79576 125192 79644 125248
rect 79700 125192 79768 125248
rect 79824 125192 79892 125248
rect 79948 125192 89920 125248
rect 79078 125122 89920 125192
rect 560032 125372 591840 125442
rect 560032 125316 590970 125372
rect 591026 125316 591094 125372
rect 591150 125316 591218 125372
rect 591274 125316 591342 125372
rect 591398 125316 591466 125372
rect 591522 125316 591590 125372
rect 591646 125316 591714 125372
rect 591770 125316 591840 125372
rect 560032 125248 591840 125316
rect 560032 125192 590970 125248
rect 591026 125192 591094 125248
rect 591150 125192 591218 125248
rect 591274 125192 591342 125248
rect 591398 125192 591466 125248
rect 591522 125192 591590 125248
rect 591646 125192 591714 125248
rect 591770 125192 591840 125248
rect 560032 125122 591840 125192
rect 592240 121691 620622 121822
rect 592240 121635 592359 121691
rect 592415 121635 592659 121691
rect 592715 121635 592959 121691
rect 593015 121635 620622 121691
rect 592240 121502 620622 121635
rect 590840 120137 620622 120268
rect 590840 120081 590959 120137
rect 591015 120081 591259 120137
rect 591315 120081 591559 120137
rect 591615 120081 620622 120137
rect 590840 119948 620622 120081
rect 592240 118583 620622 118714
rect 592240 118527 592359 118583
rect 592415 118527 592659 118583
rect 592715 118527 592959 118583
rect 593015 118527 620622 118583
rect 592240 118394 620622 118527
rect 699322 118423 701085 118490
rect 699322 118367 699497 118423
rect 699553 118367 699797 118423
rect 699853 118367 700097 118423
rect 700153 118367 701085 118423
rect 699322 118290 701085 118367
rect 701565 118090 701885 118490
rect 697922 118008 701885 118090
rect 697922 117952 698060 118008
rect 698116 117952 698360 118008
rect 698416 117952 698660 118008
rect 698716 117952 701885 118008
rect 697922 117890 701885 117952
rect 590840 117029 620622 117160
rect 590840 116973 590959 117029
rect 591015 116973 591259 117029
rect 591315 116973 591559 117029
rect 591615 116973 620622 117029
rect 590840 116840 620622 116973
rect 592240 115475 620622 115606
rect 592240 115419 592359 115475
rect 592415 115419 592659 115475
rect 592715 115419 592959 115475
rect 593015 115419 620622 115475
rect 592240 115286 620622 115419
rect 590840 113921 620622 114052
rect 590840 113865 590959 113921
rect 591015 113865 591259 113921
rect 591315 113865 591559 113921
rect 591615 113865 620622 113921
rect 590840 113732 620622 113865
rect 592240 112442 620622 112498
rect 77678 112372 89920 112442
rect 77678 112316 77748 112372
rect 77804 112316 77872 112372
rect 77928 112316 77996 112372
rect 78052 112316 78120 112372
rect 78176 112316 78244 112372
rect 78300 112316 78368 112372
rect 78424 112316 78492 112372
rect 78548 112316 89920 112372
rect 77678 112248 89920 112316
rect 77678 112192 77748 112248
rect 77804 112192 77872 112248
rect 77928 112192 77996 112248
rect 78052 112192 78120 112248
rect 78176 112192 78244 112248
rect 78300 112192 78368 112248
rect 78424 112192 78492 112248
rect 78548 112192 89920 112248
rect 77678 112122 89920 112192
rect 560032 112372 620622 112442
rect 560032 112316 592370 112372
rect 592426 112316 592494 112372
rect 592550 112316 592618 112372
rect 592674 112316 592742 112372
rect 592798 112316 592866 112372
rect 592922 112316 592990 112372
rect 593046 112316 593114 112372
rect 593170 112316 620622 112372
rect 560032 112248 620622 112316
rect 560032 112192 592370 112248
rect 592426 112192 592494 112248
rect 592550 112192 592618 112248
rect 592674 112192 592742 112248
rect 592798 112192 592866 112248
rect 592922 112192 592990 112248
rect 593046 112192 593114 112248
rect 593170 112192 620622 112248
rect 560032 112178 620622 112192
rect 560032 112122 593240 112178
rect 699322 108954 702688 109076
rect 699322 108898 699444 108954
rect 699500 108898 699744 108954
rect 699800 108898 700044 108954
rect 700100 108898 702688 108954
rect 699322 108756 702688 108898
rect 70000 105670 78678 105728
rect 70000 105658 77808 105670
rect 70000 105602 70074 105658
rect 70130 105614 77808 105658
rect 77864 105614 77932 105670
rect 77988 105614 78056 105670
rect 78112 105614 78180 105670
rect 78236 105614 78304 105670
rect 78360 105614 78428 105670
rect 78484 105614 78552 105670
rect 78608 105614 78678 105670
rect 70130 105602 78678 105614
rect 70000 105546 78678 105602
rect 70000 105534 77808 105546
rect 70000 105478 70074 105534
rect 70130 105490 77808 105534
rect 77864 105490 77932 105546
rect 77988 105490 78056 105546
rect 78112 105490 78180 105546
rect 78236 105490 78304 105546
rect 78360 105490 78428 105546
rect 78484 105490 78552 105546
rect 78608 105490 78678 105546
rect 70130 105478 78678 105490
rect 70000 105422 78678 105478
rect 70000 105410 77808 105422
rect 70000 105354 70074 105410
rect 70130 105366 77808 105410
rect 77864 105366 77932 105422
rect 77988 105366 78056 105422
rect 78112 105366 78180 105422
rect 78236 105366 78304 105422
rect 78360 105366 78428 105422
rect 78484 105366 78552 105422
rect 78608 105366 78678 105422
rect 70130 105354 78678 105366
rect 70000 105298 78678 105354
rect 70000 105286 77808 105298
rect 70000 105230 70074 105286
rect 70130 105242 77808 105286
rect 77864 105242 77932 105298
rect 77988 105242 78056 105298
rect 78112 105242 78180 105298
rect 78236 105242 78304 105298
rect 78360 105242 78428 105298
rect 78484 105242 78552 105298
rect 78608 105242 78678 105298
rect 697922 105434 702624 105576
rect 697922 105378 698044 105434
rect 698100 105378 698344 105434
rect 698400 105378 698644 105434
rect 698700 105378 702624 105434
rect 697922 105256 702624 105378
rect 70130 105230 78678 105242
rect 70000 105174 78678 105230
rect 70000 105162 77808 105174
rect 70000 105106 70074 105162
rect 70130 105118 77808 105162
rect 77864 105118 77932 105174
rect 77988 105118 78056 105174
rect 78112 105118 78180 105174
rect 78236 105118 78304 105174
rect 78360 105118 78428 105174
rect 78484 105118 78552 105174
rect 78608 105118 78678 105174
rect 70130 105106 78678 105118
rect 70000 105050 78678 105106
rect 70000 105038 77808 105050
rect 70000 104982 70074 105038
rect 70130 104994 77808 105038
rect 77864 104994 77932 105050
rect 77988 104994 78056 105050
rect 78112 104994 78180 105050
rect 78236 104994 78304 105050
rect 78360 104994 78428 105050
rect 78484 104994 78552 105050
rect 78608 104994 78678 105050
rect 70130 104982 78678 104994
rect 70000 104926 78678 104982
rect 70000 104914 77808 104926
rect 70000 104858 70074 104914
rect 70130 104870 77808 104914
rect 77864 104870 77932 104926
rect 77988 104870 78056 104926
rect 78112 104870 78180 104926
rect 78236 104870 78304 104926
rect 78360 104870 78428 104926
rect 78484 104870 78552 104926
rect 78608 104870 78678 104926
rect 70130 104858 78678 104870
rect 70000 104802 78678 104858
rect 70000 104790 77808 104802
rect 70000 104734 70074 104790
rect 70130 104746 77808 104790
rect 77864 104746 77932 104802
rect 77988 104746 78056 104802
rect 78112 104746 78180 104802
rect 78236 104746 78304 104802
rect 78360 104746 78428 104802
rect 78484 104746 78552 104802
rect 78608 104746 78678 104802
rect 70130 104734 78678 104746
rect 70000 104678 78678 104734
rect 70000 104666 77808 104678
rect 70000 104610 70074 104666
rect 70130 104622 77808 104666
rect 77864 104622 77932 104678
rect 77988 104622 78056 104678
rect 78112 104622 78180 104678
rect 78236 104622 78304 104678
rect 78360 104622 78428 104678
rect 78484 104622 78552 104678
rect 78608 104622 78678 104678
rect 70130 104610 78678 104622
rect 70000 104554 78678 104610
rect 70000 104542 77808 104554
rect 70000 104486 70074 104542
rect 70130 104498 77808 104542
rect 77864 104498 77932 104554
rect 77988 104498 78056 104554
rect 78112 104498 78180 104554
rect 78236 104498 78304 104554
rect 78360 104498 78428 104554
rect 78484 104498 78552 104554
rect 78608 104498 78678 104554
rect 70130 104486 78678 104498
rect 70000 104430 78678 104486
rect 70000 104418 77808 104430
rect 70000 104362 70074 104418
rect 70130 104374 77808 104418
rect 77864 104374 77932 104430
rect 77988 104374 78056 104430
rect 78112 104374 78180 104430
rect 78236 104374 78304 104430
rect 78360 104374 78428 104430
rect 78484 104374 78552 104430
rect 78608 104374 78678 104430
rect 70130 104362 78678 104374
rect 70000 104306 78678 104362
rect 70000 104294 77808 104306
rect 70000 104238 70074 104294
rect 70130 104250 77808 104294
rect 77864 104250 77932 104306
rect 77988 104250 78056 104306
rect 78112 104250 78180 104306
rect 78236 104250 78304 104306
rect 78360 104250 78428 104306
rect 78484 104250 78552 104306
rect 78608 104250 78678 104306
rect 70130 104238 78678 104250
rect 70000 104182 78678 104238
rect 70000 104170 77808 104182
rect 70000 104114 70074 104170
rect 70130 104126 77808 104170
rect 77864 104126 77932 104182
rect 77988 104126 78056 104182
rect 78112 104126 78180 104182
rect 78236 104126 78304 104182
rect 78360 104126 78428 104182
rect 78484 104126 78552 104182
rect 78608 104126 78678 104182
rect 70130 104114 78678 104126
rect 70000 104058 78678 104114
rect 70000 104046 77808 104058
rect 70000 103990 70074 104046
rect 70130 104002 77808 104046
rect 77864 104002 77932 104058
rect 77988 104002 78056 104058
rect 78112 104002 78180 104058
rect 78236 104002 78304 104058
rect 78360 104002 78428 104058
rect 78484 104002 78552 104058
rect 78608 104002 78678 104058
rect 70130 103990 78678 104002
rect 70000 103934 78678 103990
rect 70000 103922 77808 103934
rect 70000 103866 70074 103922
rect 70130 103878 77808 103922
rect 77864 103878 77932 103934
rect 77988 103878 78056 103934
rect 78112 103878 78180 103934
rect 78236 103878 78304 103934
rect 78360 103878 78428 103934
rect 78484 103878 78552 103934
rect 78608 103878 78678 103934
rect 70130 103866 78678 103878
rect 70000 103828 78678 103866
rect 70000 103190 78678 103248
rect 70000 103184 77808 103190
rect 70000 103128 70074 103184
rect 70130 103134 77808 103184
rect 77864 103134 77932 103190
rect 77988 103134 78056 103190
rect 78112 103134 78180 103190
rect 78236 103134 78304 103190
rect 78360 103134 78428 103190
rect 78484 103134 78552 103190
rect 78608 103134 78678 103190
rect 70130 103128 78678 103134
rect 70000 103066 78678 103128
rect 70000 103060 77808 103066
rect 70000 103004 70074 103060
rect 70130 103010 77808 103060
rect 77864 103010 77932 103066
rect 77988 103010 78056 103066
rect 78112 103010 78180 103066
rect 78236 103010 78304 103066
rect 78360 103010 78428 103066
rect 78484 103010 78552 103066
rect 78608 103010 78678 103066
rect 70130 103004 78678 103010
rect 70000 102942 78678 103004
rect 70000 102936 77808 102942
rect 70000 102880 70074 102936
rect 70130 102886 77808 102936
rect 77864 102886 77932 102942
rect 77988 102886 78056 102942
rect 78112 102886 78180 102942
rect 78236 102886 78304 102942
rect 78360 102886 78428 102942
rect 78484 102886 78552 102942
rect 78608 102886 78678 102942
rect 70130 102880 78678 102886
rect 70000 102818 78678 102880
rect 70000 102812 77808 102818
rect 70000 102756 70074 102812
rect 70130 102762 77808 102812
rect 77864 102762 77932 102818
rect 77988 102762 78056 102818
rect 78112 102762 78180 102818
rect 78236 102762 78304 102818
rect 78360 102762 78428 102818
rect 78484 102762 78552 102818
rect 78608 102762 78678 102818
rect 70130 102756 78678 102762
rect 70000 102694 78678 102756
rect 70000 102688 77808 102694
rect 70000 102632 70074 102688
rect 70130 102638 77808 102688
rect 77864 102638 77932 102694
rect 77988 102638 78056 102694
rect 78112 102638 78180 102694
rect 78236 102638 78304 102694
rect 78360 102638 78428 102694
rect 78484 102638 78552 102694
rect 78608 102638 78678 102694
rect 70130 102632 78678 102638
rect 70000 102570 78678 102632
rect 70000 102564 77808 102570
rect 70000 102508 70074 102564
rect 70130 102514 77808 102564
rect 77864 102514 77932 102570
rect 77988 102514 78056 102570
rect 78112 102514 78180 102570
rect 78236 102514 78304 102570
rect 78360 102514 78428 102570
rect 78484 102514 78552 102570
rect 78608 102514 78678 102570
rect 70130 102508 78678 102514
rect 70000 102446 78678 102508
rect 70000 102440 77808 102446
rect 70000 102384 70074 102440
rect 70130 102390 77808 102440
rect 77864 102390 77932 102446
rect 77988 102390 78056 102446
rect 78112 102390 78180 102446
rect 78236 102390 78304 102446
rect 78360 102390 78428 102446
rect 78484 102390 78552 102446
rect 78608 102390 78678 102446
rect 70130 102384 78678 102390
rect 70000 102322 78678 102384
rect 70000 102316 77808 102322
rect 70000 102260 70074 102316
rect 70130 102266 77808 102316
rect 77864 102266 77932 102322
rect 77988 102266 78056 102322
rect 78112 102266 78180 102322
rect 78236 102266 78304 102322
rect 78360 102266 78428 102322
rect 78484 102266 78552 102322
rect 78608 102266 78678 102322
rect 70130 102260 78678 102266
rect 70000 102198 78678 102260
rect 70000 102192 77808 102198
rect 70000 102136 70074 102192
rect 70130 102142 77808 102192
rect 77864 102142 77932 102198
rect 77988 102142 78056 102198
rect 78112 102142 78180 102198
rect 78236 102142 78304 102198
rect 78360 102142 78428 102198
rect 78484 102142 78552 102198
rect 78608 102142 78678 102198
rect 70130 102136 78678 102142
rect 70000 102074 78678 102136
rect 70000 102068 77808 102074
rect 70000 102012 70074 102068
rect 70130 102018 77808 102068
rect 77864 102018 77932 102074
rect 77988 102018 78056 102074
rect 78112 102018 78180 102074
rect 78236 102018 78304 102074
rect 78360 102018 78428 102074
rect 78484 102018 78552 102074
rect 78608 102018 78678 102074
rect 70130 102012 78678 102018
rect 70000 101950 78678 102012
rect 70000 101944 77808 101950
rect 70000 101888 70074 101944
rect 70130 101894 77808 101944
rect 77864 101894 77932 101950
rect 77988 101894 78056 101950
rect 78112 101894 78180 101950
rect 78236 101894 78304 101950
rect 78360 101894 78428 101950
rect 78484 101894 78552 101950
rect 78608 101894 78678 101950
rect 70130 101888 78678 101894
rect 70000 101826 78678 101888
rect 70000 101820 77808 101826
rect 70000 101764 70074 101820
rect 70130 101770 77808 101820
rect 77864 101770 77932 101826
rect 77988 101770 78056 101826
rect 78112 101770 78180 101826
rect 78236 101770 78304 101826
rect 78360 101770 78428 101826
rect 78484 101770 78552 101826
rect 78608 101770 78678 101826
rect 70130 101764 78678 101770
rect 70000 101702 78678 101764
rect 699322 101954 702688 102076
rect 699322 101898 699444 101954
rect 699500 101898 699744 101954
rect 699800 101898 700044 101954
rect 700100 101898 702688 101954
rect 699322 101756 702688 101898
rect 70000 101696 77808 101702
rect 70000 101640 70074 101696
rect 70130 101646 77808 101696
rect 77864 101646 77932 101702
rect 77988 101646 78056 101702
rect 78112 101646 78180 101702
rect 78236 101646 78304 101702
rect 78360 101646 78428 101702
rect 78484 101646 78552 101702
rect 78608 101646 78678 101702
rect 70130 101640 78678 101646
rect 70000 101578 78678 101640
rect 70000 101572 77808 101578
rect 70000 101516 70074 101572
rect 70130 101522 77808 101572
rect 77864 101522 77932 101578
rect 77988 101522 78056 101578
rect 78112 101522 78180 101578
rect 78236 101522 78304 101578
rect 78360 101522 78428 101578
rect 78484 101522 78552 101578
rect 78608 101522 78678 101578
rect 70130 101516 78678 101522
rect 70000 101454 78678 101516
rect 70000 101448 77808 101454
rect 70000 101392 70074 101448
rect 70130 101398 77808 101448
rect 77864 101398 77932 101454
rect 77988 101398 78056 101454
rect 78112 101398 78180 101454
rect 78236 101398 78304 101454
rect 78360 101398 78428 101454
rect 78484 101398 78552 101454
rect 78608 101398 78678 101454
rect 70130 101392 78678 101398
rect 70000 101330 78678 101392
rect 70000 101324 77808 101330
rect 70000 101268 70074 101324
rect 70130 101274 77808 101324
rect 77864 101274 77932 101330
rect 77988 101274 78056 101330
rect 78112 101274 78180 101330
rect 78236 101274 78304 101330
rect 78360 101274 78428 101330
rect 78484 101274 78552 101330
rect 78608 101274 78678 101330
rect 70130 101268 78678 101274
rect 70000 101198 78678 101268
rect 70000 100820 78678 100878
rect 70000 100814 77808 100820
rect 70000 100758 70074 100814
rect 70130 100764 77808 100814
rect 77864 100764 77932 100820
rect 77988 100764 78056 100820
rect 78112 100764 78180 100820
rect 78236 100764 78304 100820
rect 78360 100764 78428 100820
rect 78484 100764 78552 100820
rect 78608 100764 78678 100820
rect 70130 100758 78678 100764
rect 70000 100696 78678 100758
rect 70000 100690 77808 100696
rect 70000 100634 70074 100690
rect 70130 100640 77808 100690
rect 77864 100640 77932 100696
rect 77988 100640 78056 100696
rect 78112 100640 78180 100696
rect 78236 100640 78304 100696
rect 78360 100640 78428 100696
rect 78484 100640 78552 100696
rect 78608 100640 78678 100696
rect 70130 100634 78678 100640
rect 70000 100572 78678 100634
rect 70000 100566 77808 100572
rect 70000 100510 70074 100566
rect 70130 100516 77808 100566
rect 77864 100516 77932 100572
rect 77988 100516 78056 100572
rect 78112 100516 78180 100572
rect 78236 100516 78304 100572
rect 78360 100516 78428 100572
rect 78484 100516 78552 100572
rect 78608 100516 78678 100572
rect 70130 100510 78678 100516
rect 70000 100448 78678 100510
rect 70000 100442 77808 100448
rect 70000 100386 70074 100442
rect 70130 100392 77808 100442
rect 77864 100392 77932 100448
rect 77988 100392 78056 100448
rect 78112 100392 78180 100448
rect 78236 100392 78304 100448
rect 78360 100392 78428 100448
rect 78484 100392 78552 100448
rect 78608 100392 78678 100448
rect 70130 100386 78678 100392
rect 70000 100324 78678 100386
rect 70000 100318 77808 100324
rect 70000 100262 70074 100318
rect 70130 100268 77808 100318
rect 77864 100268 77932 100324
rect 77988 100268 78056 100324
rect 78112 100268 78180 100324
rect 78236 100268 78304 100324
rect 78360 100268 78428 100324
rect 78484 100268 78552 100324
rect 78608 100268 78678 100324
rect 70130 100262 78678 100268
rect 70000 100200 78678 100262
rect 70000 100194 77808 100200
rect 70000 100138 70074 100194
rect 70130 100144 77808 100194
rect 77864 100144 77932 100200
rect 77988 100144 78056 100200
rect 78112 100144 78180 100200
rect 78236 100144 78304 100200
rect 78360 100144 78428 100200
rect 78484 100144 78552 100200
rect 78608 100144 78678 100200
rect 70130 100138 78678 100144
rect 70000 100076 78678 100138
rect 70000 100070 77808 100076
rect 70000 100014 70074 100070
rect 70130 100020 77808 100070
rect 77864 100020 77932 100076
rect 77988 100020 78056 100076
rect 78112 100020 78180 100076
rect 78236 100020 78304 100076
rect 78360 100020 78428 100076
rect 78484 100020 78552 100076
rect 78608 100020 78678 100076
rect 70130 100014 78678 100020
rect 70000 99952 78678 100014
rect 70000 99946 77808 99952
rect 70000 99890 70074 99946
rect 70130 99896 77808 99946
rect 77864 99896 77932 99952
rect 77988 99896 78056 99952
rect 78112 99896 78180 99952
rect 78236 99896 78304 99952
rect 78360 99896 78428 99952
rect 78484 99896 78552 99952
rect 78608 99896 78678 99952
rect 70130 99890 78678 99896
rect 70000 99828 78678 99890
rect 70000 99822 77808 99828
rect 70000 99766 70074 99822
rect 70130 99772 77808 99822
rect 77864 99772 77932 99828
rect 77988 99772 78056 99828
rect 78112 99772 78180 99828
rect 78236 99772 78304 99828
rect 78360 99772 78428 99828
rect 78484 99772 78552 99828
rect 78608 99772 78678 99828
rect 70130 99766 78678 99772
rect 70000 99704 78678 99766
rect 70000 99698 77808 99704
rect 70000 99642 70074 99698
rect 70130 99648 77808 99698
rect 77864 99648 77932 99704
rect 77988 99648 78056 99704
rect 78112 99648 78180 99704
rect 78236 99648 78304 99704
rect 78360 99648 78428 99704
rect 78484 99648 78552 99704
rect 78608 99648 78678 99704
rect 70130 99642 78678 99648
rect 70000 99580 78678 99642
rect 70000 99574 77808 99580
rect 70000 99518 70074 99574
rect 70130 99524 77808 99574
rect 77864 99524 77932 99580
rect 77988 99524 78056 99580
rect 78112 99524 78180 99580
rect 78236 99524 78304 99580
rect 78360 99524 78428 99580
rect 78484 99524 78552 99580
rect 78608 99524 78678 99580
rect 70130 99518 78678 99524
rect 70000 99456 78678 99518
rect 70000 99450 77808 99456
rect 70000 99394 70074 99450
rect 70130 99400 77808 99450
rect 77864 99400 77932 99456
rect 77988 99400 78056 99456
rect 78112 99400 78180 99456
rect 78236 99400 78304 99456
rect 78360 99400 78428 99456
rect 78484 99400 78552 99456
rect 78608 99400 78678 99456
rect 70130 99394 78678 99400
rect 70000 99332 78678 99394
rect 70000 99326 77808 99332
rect 70000 99270 70074 99326
rect 70130 99276 77808 99326
rect 77864 99276 77932 99332
rect 77988 99276 78056 99332
rect 78112 99276 78180 99332
rect 78236 99276 78304 99332
rect 78360 99276 78428 99332
rect 78484 99276 78552 99332
rect 78608 99276 78678 99332
rect 70130 99270 78678 99276
rect 70000 99208 78678 99270
rect 70000 99202 77808 99208
rect 70000 99146 70074 99202
rect 70130 99152 77808 99202
rect 77864 99152 77932 99208
rect 77988 99152 78056 99208
rect 78112 99152 78180 99208
rect 78236 99152 78304 99208
rect 78360 99152 78428 99208
rect 78484 99152 78552 99208
rect 78608 99152 78678 99208
rect 70130 99146 78678 99152
rect 70000 99084 78678 99146
rect 79078 99372 89920 99442
rect 79078 99316 79148 99372
rect 79204 99316 79272 99372
rect 79328 99316 79396 99372
rect 79452 99316 79520 99372
rect 79576 99316 79644 99372
rect 79700 99316 79768 99372
rect 79824 99316 79892 99372
rect 79948 99316 89920 99372
rect 79078 99248 89920 99316
rect 79078 99192 79148 99248
rect 79204 99192 79272 99248
rect 79328 99192 79396 99248
rect 79452 99192 79520 99248
rect 79576 99192 79644 99248
rect 79700 99192 79768 99248
rect 79824 99192 79892 99248
rect 79948 99192 89920 99248
rect 79078 99122 89920 99192
rect 560032 99372 591840 99442
rect 560032 99316 590970 99372
rect 591026 99316 591094 99372
rect 591150 99316 591218 99372
rect 591274 99316 591342 99372
rect 591398 99316 591466 99372
rect 591522 99316 591590 99372
rect 591646 99316 591714 99372
rect 591770 99316 591840 99372
rect 560032 99248 591840 99316
rect 560032 99192 590970 99248
rect 591026 99192 591094 99248
rect 591150 99192 591218 99248
rect 591274 99192 591342 99248
rect 591398 99192 591466 99248
rect 591522 99192 591590 99248
rect 591646 99192 591714 99248
rect 591770 99192 591840 99248
rect 560032 99122 591840 99192
rect 70000 99078 77808 99084
rect 70000 99022 70074 99078
rect 70130 99028 77808 99078
rect 77864 99028 77932 99084
rect 77988 99028 78056 99084
rect 78112 99028 78180 99084
rect 78236 99028 78304 99084
rect 78360 99028 78428 99084
rect 78484 99028 78552 99084
rect 78608 99028 78678 99084
rect 70130 99022 78678 99028
rect 70000 98960 78678 99022
rect 70000 98954 77808 98960
rect 70000 98898 70074 98954
rect 70130 98904 77808 98954
rect 77864 98904 77932 98960
rect 77988 98904 78056 98960
rect 78112 98904 78180 98960
rect 78236 98904 78304 98960
rect 78360 98904 78428 98960
rect 78484 98904 78552 98960
rect 78608 98904 78678 98960
rect 70130 98898 78678 98904
rect 70000 98828 78678 98898
rect 697922 98434 702624 98576
rect 697922 98378 698044 98434
rect 698100 98378 698344 98434
rect 698400 98378 698644 98434
rect 698700 98378 702624 98434
rect 697922 98256 702624 98378
rect 70000 98114 78678 98172
rect 70000 98108 77808 98114
rect 70000 98052 70074 98108
rect 70130 98058 77808 98108
rect 77864 98058 77932 98114
rect 77988 98058 78056 98114
rect 78112 98058 78180 98114
rect 78236 98058 78304 98114
rect 78360 98058 78428 98114
rect 78484 98058 78552 98114
rect 78608 98058 78678 98114
rect 70130 98052 78678 98058
rect 70000 97990 78678 98052
rect 70000 97984 77808 97990
rect 70000 97928 70074 97984
rect 70130 97934 77808 97984
rect 77864 97934 77932 97990
rect 77988 97934 78056 97990
rect 78112 97934 78180 97990
rect 78236 97934 78304 97990
rect 78360 97934 78428 97990
rect 78484 97934 78552 97990
rect 78608 97934 78678 97990
rect 70130 97928 78678 97934
rect 70000 97866 78678 97928
rect 70000 97860 77808 97866
rect 70000 97804 70074 97860
rect 70130 97810 77808 97860
rect 77864 97810 77932 97866
rect 77988 97810 78056 97866
rect 78112 97810 78180 97866
rect 78236 97810 78304 97866
rect 78360 97810 78428 97866
rect 78484 97810 78552 97866
rect 78608 97810 78678 97866
rect 70130 97804 78678 97810
rect 70000 97742 78678 97804
rect 70000 97736 77808 97742
rect 70000 97680 70074 97736
rect 70130 97686 77808 97736
rect 77864 97686 77932 97742
rect 77988 97686 78056 97742
rect 78112 97686 78180 97742
rect 78236 97686 78304 97742
rect 78360 97686 78428 97742
rect 78484 97686 78552 97742
rect 78608 97686 78678 97742
rect 70130 97680 78678 97686
rect 70000 97618 78678 97680
rect 70000 97612 77808 97618
rect 70000 97556 70074 97612
rect 70130 97562 77808 97612
rect 77864 97562 77932 97618
rect 77988 97562 78056 97618
rect 78112 97562 78180 97618
rect 78236 97562 78304 97618
rect 78360 97562 78428 97618
rect 78484 97562 78552 97618
rect 78608 97562 78678 97618
rect 70130 97556 78678 97562
rect 70000 97494 78678 97556
rect 70000 97488 77808 97494
rect 70000 97432 70074 97488
rect 70130 97438 77808 97488
rect 77864 97438 77932 97494
rect 77988 97438 78056 97494
rect 78112 97438 78180 97494
rect 78236 97438 78304 97494
rect 78360 97438 78428 97494
rect 78484 97438 78552 97494
rect 78608 97438 78678 97494
rect 70130 97432 78678 97438
rect 70000 97370 78678 97432
rect 70000 97364 77808 97370
rect 70000 97308 70074 97364
rect 70130 97314 77808 97364
rect 77864 97314 77932 97370
rect 77988 97314 78056 97370
rect 78112 97314 78180 97370
rect 78236 97314 78304 97370
rect 78360 97314 78428 97370
rect 78484 97314 78552 97370
rect 78608 97314 78678 97370
rect 70130 97308 78678 97314
rect 70000 97246 78678 97308
rect 70000 97240 77808 97246
rect 70000 97184 70074 97240
rect 70130 97190 77808 97240
rect 77864 97190 77932 97246
rect 77988 97190 78056 97246
rect 78112 97190 78180 97246
rect 78236 97190 78304 97246
rect 78360 97190 78428 97246
rect 78484 97190 78552 97246
rect 78608 97190 78678 97246
rect 70130 97184 78678 97190
rect 70000 97122 78678 97184
rect 70000 97116 77808 97122
rect 70000 97060 70074 97116
rect 70130 97066 77808 97116
rect 77864 97066 77932 97122
rect 77988 97066 78056 97122
rect 78112 97066 78180 97122
rect 78236 97066 78304 97122
rect 78360 97066 78428 97122
rect 78484 97066 78552 97122
rect 78608 97066 78678 97122
rect 70130 97060 78678 97066
rect 70000 96998 78678 97060
rect 70000 96992 77808 96998
rect 70000 96936 70074 96992
rect 70130 96942 77808 96992
rect 77864 96942 77932 96998
rect 77988 96942 78056 96998
rect 78112 96942 78180 96998
rect 78236 96942 78304 96998
rect 78360 96942 78428 96998
rect 78484 96942 78552 96998
rect 78608 96942 78678 96998
rect 70130 96936 78678 96942
rect 70000 96874 78678 96936
rect 70000 96868 77808 96874
rect 70000 96812 70074 96868
rect 70130 96818 77808 96868
rect 77864 96818 77932 96874
rect 77988 96818 78056 96874
rect 78112 96818 78180 96874
rect 78236 96818 78304 96874
rect 78360 96818 78428 96874
rect 78484 96818 78552 96874
rect 78608 96818 78678 96874
rect 70130 96812 78678 96818
rect 70000 96750 78678 96812
rect 70000 96744 77808 96750
rect 70000 96688 70074 96744
rect 70130 96694 77808 96744
rect 77864 96694 77932 96750
rect 77988 96694 78056 96750
rect 78112 96694 78180 96750
rect 78236 96694 78304 96750
rect 78360 96694 78428 96750
rect 78484 96694 78552 96750
rect 78608 96694 78678 96750
rect 70130 96688 78678 96694
rect 70000 96626 78678 96688
rect 70000 96620 77808 96626
rect 70000 96564 70074 96620
rect 70130 96570 77808 96620
rect 77864 96570 77932 96626
rect 77988 96570 78056 96626
rect 78112 96570 78180 96626
rect 78236 96570 78304 96626
rect 78360 96570 78428 96626
rect 78484 96570 78552 96626
rect 78608 96570 78678 96626
rect 70130 96564 78678 96570
rect 70000 96502 78678 96564
rect 70000 96496 77808 96502
rect 70000 96440 70074 96496
rect 70130 96446 77808 96496
rect 77864 96446 77932 96502
rect 77988 96446 78056 96502
rect 78112 96446 78180 96502
rect 78236 96446 78304 96502
rect 78360 96446 78428 96502
rect 78484 96446 78552 96502
rect 78608 96446 78678 96502
rect 70130 96440 78678 96446
rect 70000 96378 78678 96440
rect 70000 96372 77808 96378
rect 70000 96316 70074 96372
rect 70130 96322 77808 96372
rect 77864 96322 77932 96378
rect 77988 96322 78056 96378
rect 78112 96322 78180 96378
rect 78236 96322 78304 96378
rect 78360 96322 78428 96378
rect 78484 96322 78552 96378
rect 78608 96322 78678 96378
rect 70130 96316 78678 96322
rect 70000 96254 78678 96316
rect 70000 96248 77808 96254
rect 70000 96192 70074 96248
rect 70130 96198 77808 96248
rect 77864 96198 77932 96254
rect 77988 96198 78056 96254
rect 78112 96198 78180 96254
rect 78236 96198 78304 96254
rect 78360 96198 78428 96254
rect 78484 96198 78552 96254
rect 78608 96198 78678 96254
rect 70130 96192 78678 96198
rect 70000 96122 78678 96192
rect 70000 95744 78678 95802
rect 70000 95738 77808 95744
rect 70000 95682 70074 95738
rect 70130 95688 77808 95738
rect 77864 95688 77932 95744
rect 77988 95688 78056 95744
rect 78112 95688 78180 95744
rect 78236 95688 78304 95744
rect 78360 95688 78428 95744
rect 78484 95688 78552 95744
rect 78608 95688 78678 95744
rect 70130 95682 78678 95688
rect 70000 95620 78678 95682
rect 70000 95614 77808 95620
rect 70000 95558 70074 95614
rect 70130 95564 77808 95614
rect 77864 95564 77932 95620
rect 77988 95564 78056 95620
rect 78112 95564 78180 95620
rect 78236 95564 78304 95620
rect 78360 95564 78428 95620
rect 78484 95564 78552 95620
rect 78608 95564 78678 95620
rect 70130 95558 78678 95564
rect 70000 95496 78678 95558
rect 70000 95490 77808 95496
rect 70000 95434 70074 95490
rect 70130 95440 77808 95490
rect 77864 95440 77932 95496
rect 77988 95440 78056 95496
rect 78112 95440 78180 95496
rect 78236 95440 78304 95496
rect 78360 95440 78428 95496
rect 78484 95440 78552 95496
rect 78608 95440 78678 95496
rect 70130 95434 78678 95440
rect 70000 95372 78678 95434
rect 70000 95366 77808 95372
rect 70000 95310 70074 95366
rect 70130 95316 77808 95366
rect 77864 95316 77932 95372
rect 77988 95316 78056 95372
rect 78112 95316 78180 95372
rect 78236 95316 78304 95372
rect 78360 95316 78428 95372
rect 78484 95316 78552 95372
rect 78608 95316 78678 95372
rect 70130 95310 78678 95316
rect 70000 95248 78678 95310
rect 70000 95242 77808 95248
rect 70000 95186 70074 95242
rect 70130 95192 77808 95242
rect 77864 95192 77932 95248
rect 77988 95192 78056 95248
rect 78112 95192 78180 95248
rect 78236 95192 78304 95248
rect 78360 95192 78428 95248
rect 78484 95192 78552 95248
rect 78608 95192 78678 95248
rect 70130 95186 78678 95192
rect 70000 95124 78678 95186
rect 70000 95118 77808 95124
rect 70000 95062 70074 95118
rect 70130 95068 77808 95118
rect 77864 95068 77932 95124
rect 77988 95068 78056 95124
rect 78112 95068 78180 95124
rect 78236 95068 78304 95124
rect 78360 95068 78428 95124
rect 78484 95068 78552 95124
rect 78608 95068 78678 95124
rect 70130 95062 78678 95068
rect 70000 95000 78678 95062
rect 70000 94994 77808 95000
rect 70000 94938 70074 94994
rect 70130 94944 77808 94994
rect 77864 94944 77932 95000
rect 77988 94944 78056 95000
rect 78112 94944 78180 95000
rect 78236 94944 78304 95000
rect 78360 94944 78428 95000
rect 78484 94944 78552 95000
rect 78608 94944 78678 95000
rect 70130 94938 78678 94944
rect 70000 94876 78678 94938
rect 70000 94870 77808 94876
rect 70000 94814 70074 94870
rect 70130 94820 77808 94870
rect 77864 94820 77932 94876
rect 77988 94820 78056 94876
rect 78112 94820 78180 94876
rect 78236 94820 78304 94876
rect 78360 94820 78428 94876
rect 78484 94820 78552 94876
rect 78608 94820 78678 94876
rect 70130 94814 78678 94820
rect 70000 94752 78678 94814
rect 699322 94954 702688 95076
rect 699322 94898 699444 94954
rect 699500 94898 699744 94954
rect 699800 94898 700044 94954
rect 700100 94898 702688 94954
rect 699322 94756 702688 94898
rect 70000 94746 77808 94752
rect 70000 94690 70074 94746
rect 70130 94696 77808 94746
rect 77864 94696 77932 94752
rect 77988 94696 78056 94752
rect 78112 94696 78180 94752
rect 78236 94696 78304 94752
rect 78360 94696 78428 94752
rect 78484 94696 78552 94752
rect 78608 94696 78678 94752
rect 70130 94690 78678 94696
rect 70000 94628 78678 94690
rect 70000 94622 77808 94628
rect 70000 94566 70074 94622
rect 70130 94572 77808 94622
rect 77864 94572 77932 94628
rect 77988 94572 78056 94628
rect 78112 94572 78180 94628
rect 78236 94572 78304 94628
rect 78360 94572 78428 94628
rect 78484 94572 78552 94628
rect 78608 94572 78678 94628
rect 70130 94566 78678 94572
rect 70000 94504 78678 94566
rect 70000 94498 77808 94504
rect 70000 94442 70074 94498
rect 70130 94448 77808 94498
rect 77864 94448 77932 94504
rect 77988 94448 78056 94504
rect 78112 94448 78180 94504
rect 78236 94448 78304 94504
rect 78360 94448 78428 94504
rect 78484 94448 78552 94504
rect 78608 94448 78678 94504
rect 70130 94442 78678 94448
rect 70000 94380 78678 94442
rect 70000 94374 77808 94380
rect 70000 94318 70074 94374
rect 70130 94324 77808 94374
rect 77864 94324 77932 94380
rect 77988 94324 78056 94380
rect 78112 94324 78180 94380
rect 78236 94324 78304 94380
rect 78360 94324 78428 94380
rect 78484 94324 78552 94380
rect 78608 94324 78678 94380
rect 70130 94318 78678 94324
rect 70000 94256 78678 94318
rect 70000 94250 77808 94256
rect 70000 94194 70074 94250
rect 70130 94200 77808 94250
rect 77864 94200 77932 94256
rect 77988 94200 78056 94256
rect 78112 94200 78180 94256
rect 78236 94200 78304 94256
rect 78360 94200 78428 94256
rect 78484 94200 78552 94256
rect 78608 94200 78678 94256
rect 70130 94194 78678 94200
rect 70000 94132 78678 94194
rect 70000 94126 77808 94132
rect 70000 94070 70074 94126
rect 70130 94076 77808 94126
rect 77864 94076 77932 94132
rect 77988 94076 78056 94132
rect 78112 94076 78180 94132
rect 78236 94076 78304 94132
rect 78360 94076 78428 94132
rect 78484 94076 78552 94132
rect 78608 94076 78678 94132
rect 70130 94070 78678 94076
rect 70000 94008 78678 94070
rect 70000 94002 77808 94008
rect 70000 93946 70074 94002
rect 70130 93952 77808 94002
rect 77864 93952 77932 94008
rect 77988 93952 78056 94008
rect 78112 93952 78180 94008
rect 78236 93952 78304 94008
rect 78360 93952 78428 94008
rect 78484 93952 78552 94008
rect 78608 93952 78678 94008
rect 70130 93946 78678 93952
rect 70000 93884 78678 93946
rect 70000 93878 77808 93884
rect 70000 93822 70074 93878
rect 70130 93828 77808 93878
rect 77864 93828 77932 93884
rect 77988 93828 78056 93884
rect 78112 93828 78180 93884
rect 78236 93828 78304 93884
rect 78360 93828 78428 93884
rect 78484 93828 78552 93884
rect 78608 93828 78678 93884
rect 70130 93822 78678 93828
rect 70000 93752 78678 93822
rect 70000 93140 78678 93172
rect 70000 93134 77808 93140
rect 70000 93078 70074 93134
rect 70130 93084 77808 93134
rect 77864 93084 77932 93140
rect 77988 93084 78056 93140
rect 78112 93084 78180 93140
rect 78236 93084 78304 93140
rect 78360 93084 78428 93140
rect 78484 93084 78552 93140
rect 78608 93084 78678 93140
rect 70130 93078 78678 93084
rect 70000 93016 78678 93078
rect 70000 93010 77808 93016
rect 70000 92954 70074 93010
rect 70130 92960 77808 93010
rect 77864 92960 77932 93016
rect 77988 92960 78056 93016
rect 78112 92960 78180 93016
rect 78236 92960 78304 93016
rect 78360 92960 78428 93016
rect 78484 92960 78552 93016
rect 78608 92960 78678 93016
rect 70130 92954 78678 92960
rect 70000 92892 78678 92954
rect 70000 92886 77808 92892
rect 70000 92830 70074 92886
rect 70130 92836 77808 92886
rect 77864 92836 77932 92892
rect 77988 92836 78056 92892
rect 78112 92836 78180 92892
rect 78236 92836 78304 92892
rect 78360 92836 78428 92892
rect 78484 92836 78552 92892
rect 78608 92836 78678 92892
rect 70130 92830 78678 92836
rect 70000 92768 78678 92830
rect 70000 92762 77808 92768
rect 70000 92706 70074 92762
rect 70130 92712 77808 92762
rect 77864 92712 77932 92768
rect 77988 92712 78056 92768
rect 78112 92712 78180 92768
rect 78236 92712 78304 92768
rect 78360 92712 78428 92768
rect 78484 92712 78552 92768
rect 78608 92712 78678 92768
rect 70130 92706 78678 92712
rect 70000 92644 78678 92706
rect 70000 92638 77808 92644
rect 70000 92582 70074 92638
rect 70130 92588 77808 92638
rect 77864 92588 77932 92644
rect 77988 92588 78056 92644
rect 78112 92588 78180 92644
rect 78236 92588 78304 92644
rect 78360 92588 78428 92644
rect 78484 92588 78552 92644
rect 78608 92588 78678 92644
rect 70130 92582 78678 92588
rect 70000 92520 78678 92582
rect 70000 92514 77808 92520
rect 70000 92458 70074 92514
rect 70130 92464 77808 92514
rect 77864 92464 77932 92520
rect 77988 92464 78056 92520
rect 78112 92464 78180 92520
rect 78236 92464 78304 92520
rect 78360 92464 78428 92520
rect 78484 92464 78552 92520
rect 78608 92464 78678 92520
rect 70130 92458 78678 92464
rect 70000 92396 78678 92458
rect 70000 92390 77808 92396
rect 70000 92334 70074 92390
rect 70130 92340 77808 92390
rect 77864 92340 77932 92396
rect 77988 92340 78056 92396
rect 78112 92340 78180 92396
rect 78236 92340 78304 92396
rect 78360 92340 78428 92396
rect 78484 92340 78552 92396
rect 78608 92340 78678 92396
rect 70130 92334 78678 92340
rect 70000 92272 78678 92334
rect 70000 92266 77808 92272
rect 70000 92210 70074 92266
rect 70130 92216 77808 92266
rect 77864 92216 77932 92272
rect 77988 92216 78056 92272
rect 78112 92216 78180 92272
rect 78236 92216 78304 92272
rect 78360 92216 78428 92272
rect 78484 92216 78552 92272
rect 78608 92216 78678 92272
rect 70130 92210 78678 92216
rect 70000 92148 78678 92210
rect 70000 92142 77808 92148
rect 70000 92086 70074 92142
rect 70130 92092 77808 92142
rect 77864 92092 77932 92148
rect 77988 92092 78056 92148
rect 78112 92092 78180 92148
rect 78236 92092 78304 92148
rect 78360 92092 78428 92148
rect 78484 92092 78552 92148
rect 78608 92092 78678 92148
rect 70130 92086 78678 92092
rect 70000 92024 78678 92086
rect 70000 92018 77808 92024
rect 70000 91962 70074 92018
rect 70130 91968 77808 92018
rect 77864 91968 77932 92024
rect 77988 91968 78056 92024
rect 78112 91968 78180 92024
rect 78236 91968 78304 92024
rect 78360 91968 78428 92024
rect 78484 91968 78552 92024
rect 78608 91968 78678 92024
rect 70130 91962 78678 91968
rect 70000 91900 78678 91962
rect 70000 91894 77808 91900
rect 70000 91838 70074 91894
rect 70130 91844 77808 91894
rect 77864 91844 77932 91900
rect 77988 91844 78056 91900
rect 78112 91844 78180 91900
rect 78236 91844 78304 91900
rect 78360 91844 78428 91900
rect 78484 91844 78552 91900
rect 78608 91844 78678 91900
rect 70130 91838 78678 91844
rect 70000 91776 78678 91838
rect 70000 91770 77808 91776
rect 70000 91714 70074 91770
rect 70130 91720 77808 91770
rect 77864 91720 77932 91776
rect 77988 91720 78056 91776
rect 78112 91720 78180 91776
rect 78236 91720 78304 91776
rect 78360 91720 78428 91776
rect 78484 91720 78552 91776
rect 78608 91720 78678 91776
rect 70130 91714 78678 91720
rect 70000 91652 78678 91714
rect 70000 91646 77808 91652
rect 70000 91590 70074 91646
rect 70130 91596 77808 91646
rect 77864 91596 77932 91652
rect 77988 91596 78056 91652
rect 78112 91596 78180 91652
rect 78236 91596 78304 91652
rect 78360 91596 78428 91652
rect 78484 91596 78552 91652
rect 78608 91596 78678 91652
rect 70130 91590 78678 91596
rect 70000 91528 78678 91590
rect 70000 91522 77808 91528
rect 70000 91466 70074 91522
rect 70130 91472 77808 91522
rect 77864 91472 77932 91528
rect 77988 91472 78056 91528
rect 78112 91472 78180 91528
rect 78236 91472 78304 91528
rect 78360 91472 78428 91528
rect 78484 91472 78552 91528
rect 78608 91472 78678 91528
rect 70130 91466 78678 91472
rect 70000 91404 78678 91466
rect 70000 91398 77808 91404
rect 70000 91342 70074 91398
rect 70130 91348 77808 91398
rect 77864 91348 77932 91404
rect 77988 91348 78056 91404
rect 78112 91348 78180 91404
rect 78236 91348 78304 91404
rect 78360 91348 78428 91404
rect 78484 91348 78552 91404
rect 78608 91348 78678 91404
rect 70130 91342 78678 91348
rect 70000 91272 78678 91342
rect 697922 91434 702624 91576
rect 697922 91378 698044 91434
rect 698100 91378 698344 91434
rect 698400 91378 698644 91434
rect 698700 91378 702624 91434
rect 697922 91256 702624 91378
rect 77678 86372 89920 86442
rect 77678 86316 77748 86372
rect 77804 86316 77872 86372
rect 77928 86316 77996 86372
rect 78052 86316 78120 86372
rect 78176 86316 78244 86372
rect 78300 86316 78368 86372
rect 78424 86316 78492 86372
rect 78548 86316 89920 86372
rect 77678 86248 89920 86316
rect 77678 86192 77748 86248
rect 77804 86192 77872 86248
rect 77928 86192 77996 86248
rect 78052 86192 78120 86248
rect 78176 86192 78244 86248
rect 78300 86192 78368 86248
rect 78424 86192 78492 86248
rect 78548 86192 89920 86248
rect 77678 86122 89920 86192
rect 560032 86372 593240 86442
rect 560032 86316 592370 86372
rect 592426 86316 592494 86372
rect 592550 86316 592618 86372
rect 592674 86316 592742 86372
rect 592798 86316 592866 86372
rect 592922 86316 592990 86372
rect 593046 86316 593114 86372
rect 593170 86316 593240 86372
rect 560032 86248 593240 86316
rect 560032 86192 592370 86248
rect 592426 86192 592494 86248
rect 592550 86192 592618 86248
rect 592674 86192 592742 86248
rect 592798 86192 592866 86248
rect 592922 86192 592990 86248
rect 593046 86192 593114 86248
rect 593170 86192 593240 86248
rect 560032 86122 593240 86192
rect 79078 80008 698922 80078
rect 79078 79952 79208 80008
rect 79264 79952 79332 80008
rect 79388 79952 79456 80008
rect 79512 79952 79580 80008
rect 79636 79952 79704 80008
rect 79760 79952 79828 80008
rect 79884 79952 79952 80008
rect 80008 79952 99294 80008
rect 99350 79952 99418 80008
rect 99474 79952 107330 80008
rect 107386 79952 107454 80008
rect 107510 79952 107578 80008
rect 107634 79952 107702 80008
rect 107758 79952 107826 80008
rect 107882 79952 107950 80008
rect 108006 79952 108074 80008
rect 108130 79952 108198 80008
rect 108254 79952 108322 80008
rect 108378 79952 108446 80008
rect 108502 79952 108570 80008
rect 108626 79952 108694 80008
rect 108750 79952 108818 80008
rect 108874 79952 108942 80008
rect 108998 79952 109066 80008
rect 109122 79952 109810 80008
rect 109866 79952 109934 80008
rect 109990 79952 110058 80008
rect 110114 79952 110182 80008
rect 110238 79952 110306 80008
rect 110362 79952 110430 80008
rect 110486 79952 110554 80008
rect 110610 79952 110678 80008
rect 110734 79952 110802 80008
rect 110858 79952 110926 80008
rect 110982 79952 111050 80008
rect 111106 79952 111174 80008
rect 111230 79952 111298 80008
rect 111354 79952 111422 80008
rect 111478 79952 111546 80008
rect 111602 79952 111670 80008
rect 111726 79952 112180 80008
rect 112236 79952 112304 80008
rect 112360 79952 112428 80008
rect 112484 79952 112552 80008
rect 112608 79952 112676 80008
rect 112732 79952 112800 80008
rect 112856 79952 112924 80008
rect 112980 79952 113048 80008
rect 113104 79952 113172 80008
rect 113228 79952 113296 80008
rect 113352 79952 113420 80008
rect 113476 79952 113544 80008
rect 113600 79952 113668 80008
rect 113724 79952 113792 80008
rect 113848 79952 113916 80008
rect 113972 79952 114040 80008
rect 114096 79952 114886 80008
rect 114942 79952 115010 80008
rect 115066 79952 115134 80008
rect 115190 79952 115258 80008
rect 115314 79952 115382 80008
rect 115438 79952 115506 80008
rect 115562 79952 115630 80008
rect 115686 79952 115754 80008
rect 115810 79952 115878 80008
rect 115934 79952 116002 80008
rect 116058 79952 116126 80008
rect 116182 79952 116250 80008
rect 116306 79952 116374 80008
rect 116430 79952 116498 80008
rect 116554 79952 116622 80008
rect 116678 79952 116746 80008
rect 116802 79952 117256 80008
rect 117312 79952 117380 80008
rect 117436 79952 117504 80008
rect 117560 79952 117628 80008
rect 117684 79952 117752 80008
rect 117808 79952 117876 80008
rect 117932 79952 118000 80008
rect 118056 79952 118124 80008
rect 118180 79952 118248 80008
rect 118304 79952 118372 80008
rect 118428 79952 118496 80008
rect 118552 79952 118620 80008
rect 118676 79952 118744 80008
rect 118800 79952 118868 80008
rect 118924 79952 118992 80008
rect 119048 79952 119116 80008
rect 119172 79952 119860 80008
rect 119916 79952 119984 80008
rect 120040 79952 120108 80008
rect 120164 79952 120232 80008
rect 120288 79952 120356 80008
rect 120412 79952 120480 80008
rect 120536 79952 120604 80008
rect 120660 79952 120728 80008
rect 120784 79952 120852 80008
rect 120908 79952 120976 80008
rect 121032 79952 121100 80008
rect 121156 79952 121224 80008
rect 121280 79952 121348 80008
rect 121404 79952 121472 80008
rect 121528 79952 121596 80008
rect 121652 79952 129294 80008
rect 129350 79952 129418 80008
rect 129474 79952 139294 80008
rect 139350 79952 139418 80008
rect 139474 79952 149294 80008
rect 149350 79952 149418 80008
rect 149474 79952 159294 80008
rect 159350 79952 159418 80008
rect 159474 79952 169294 80008
rect 169350 79952 169418 80008
rect 169474 79952 179294 80008
rect 179350 79952 179418 80008
rect 179474 79952 189294 80008
rect 189350 79952 189418 80008
rect 189474 79952 199294 80008
rect 199350 79952 199418 80008
rect 199474 79952 209294 80008
rect 209350 79952 209418 80008
rect 209474 79952 219294 80008
rect 219350 79952 219418 80008
rect 219474 79952 229294 80008
rect 229350 79952 229418 80008
rect 229474 79952 239294 80008
rect 239350 79952 239418 80008
rect 239474 79952 249294 80008
rect 249350 79952 249418 80008
rect 249474 79952 259294 80008
rect 259350 79952 259418 80008
rect 259474 79952 269294 80008
rect 269350 79952 269418 80008
rect 269474 79952 272330 80008
rect 272386 79952 272454 80008
rect 272510 79952 272578 80008
rect 272634 79952 272702 80008
rect 272758 79952 272826 80008
rect 272882 79952 272950 80008
rect 273006 79952 273074 80008
rect 273130 79952 273198 80008
rect 273254 79952 273322 80008
rect 273378 79952 273446 80008
rect 273502 79952 273570 80008
rect 273626 79952 273694 80008
rect 273750 79952 273818 80008
rect 273874 79952 273942 80008
rect 273998 79952 274066 80008
rect 274122 79952 274810 80008
rect 274866 79952 274934 80008
rect 274990 79952 275058 80008
rect 275114 79952 275182 80008
rect 275238 79952 275306 80008
rect 275362 79952 275430 80008
rect 275486 79952 275554 80008
rect 275610 79952 275678 80008
rect 275734 79952 275802 80008
rect 275858 79952 275926 80008
rect 275982 79952 276050 80008
rect 276106 79952 276174 80008
rect 276230 79952 276298 80008
rect 276354 79952 276422 80008
rect 276478 79952 276546 80008
rect 276602 79952 276670 80008
rect 276726 79952 277180 80008
rect 277236 79952 277304 80008
rect 277360 79952 277428 80008
rect 277484 79952 277552 80008
rect 277608 79952 277676 80008
rect 277732 79952 277800 80008
rect 277856 79952 277924 80008
rect 277980 79952 278048 80008
rect 278104 79952 278172 80008
rect 278228 79952 278296 80008
rect 278352 79952 278420 80008
rect 278476 79952 278544 80008
rect 278600 79952 278668 80008
rect 278724 79952 278792 80008
rect 278848 79952 278916 80008
rect 278972 79952 279040 80008
rect 279096 79952 279886 80008
rect 279942 79952 280010 80008
rect 280066 79952 280134 80008
rect 280190 79952 280258 80008
rect 280314 79952 280382 80008
rect 280438 79952 280506 80008
rect 280562 79952 280630 80008
rect 280686 79952 280754 80008
rect 280810 79952 280878 80008
rect 280934 79952 281002 80008
rect 281058 79952 281126 80008
rect 281182 79952 281250 80008
rect 281306 79952 281374 80008
rect 281430 79952 281498 80008
rect 281554 79952 281622 80008
rect 281678 79952 281746 80008
rect 281802 79952 282256 80008
rect 282312 79952 282380 80008
rect 282436 79952 282504 80008
rect 282560 79952 282628 80008
rect 282684 79952 282752 80008
rect 282808 79952 282876 80008
rect 282932 79952 283000 80008
rect 283056 79952 283124 80008
rect 283180 79952 283248 80008
rect 283304 79952 283372 80008
rect 283428 79952 283496 80008
rect 283552 79952 283620 80008
rect 283676 79952 283744 80008
rect 283800 79952 283868 80008
rect 283924 79952 283992 80008
rect 284048 79952 284116 80008
rect 284172 79952 284860 80008
rect 284916 79952 284984 80008
rect 285040 79952 285108 80008
rect 285164 79952 285232 80008
rect 285288 79952 285356 80008
rect 285412 79952 285480 80008
rect 285536 79952 285604 80008
rect 285660 79952 285728 80008
rect 285784 79952 285852 80008
rect 285908 79952 285976 80008
rect 286032 79952 286100 80008
rect 286156 79952 286224 80008
rect 286280 79952 286348 80008
rect 286404 79952 286472 80008
rect 286528 79952 286596 80008
rect 286652 79952 289294 80008
rect 289350 79952 289418 80008
rect 289474 79952 299294 80008
rect 299350 79952 299418 80008
rect 299474 79952 309294 80008
rect 309350 79952 309418 80008
rect 309474 79952 319294 80008
rect 319350 79952 319418 80008
rect 319474 79952 329294 80008
rect 329350 79952 329418 80008
rect 329474 79952 339294 80008
rect 339350 79952 339418 80008
rect 339474 79952 349294 80008
rect 349350 79952 349418 80008
rect 349474 79952 359294 80008
rect 359350 79952 359418 80008
rect 359474 79952 369294 80008
rect 369350 79952 369418 80008
rect 369474 79952 379294 80008
rect 379350 79952 379418 80008
rect 379474 79952 389294 80008
rect 389350 79952 389418 80008
rect 389474 79952 399294 80008
rect 399350 79952 399418 80008
rect 399474 79952 409294 80008
rect 409350 79952 409418 80008
rect 409474 79952 419294 80008
rect 419350 79952 419418 80008
rect 419474 79952 429294 80008
rect 429350 79952 429418 80008
rect 429474 79952 439294 80008
rect 439350 79952 439418 80008
rect 439474 79952 449294 80008
rect 449350 79952 449418 80008
rect 449474 79952 459294 80008
rect 459350 79952 459418 80008
rect 459474 79952 469294 80008
rect 469350 79952 469418 80008
rect 469474 79952 479294 80008
rect 479350 79952 479418 80008
rect 479474 79952 489294 80008
rect 489350 79952 489418 80008
rect 489474 79952 499294 80008
rect 499350 79952 499418 80008
rect 499474 79952 509294 80008
rect 509350 79952 509418 80008
rect 509474 79952 519294 80008
rect 519350 79952 519418 80008
rect 519474 79952 529294 80008
rect 529350 79952 529418 80008
rect 529474 79952 539294 80008
rect 539350 79952 539418 80008
rect 539474 79952 549294 80008
rect 549350 79952 549418 80008
rect 549474 79952 590970 80008
rect 591026 79952 591094 80008
rect 591150 79952 591218 80008
rect 591274 79952 591342 80008
rect 591398 79952 591466 80008
rect 591522 79952 591590 80008
rect 591646 79952 591714 80008
rect 591770 79952 602330 80008
rect 602386 79952 602454 80008
rect 602510 79952 602578 80008
rect 602634 79952 602702 80008
rect 602758 79952 602826 80008
rect 602882 79952 602950 80008
rect 603006 79952 603074 80008
rect 603130 79952 603198 80008
rect 603254 79952 603322 80008
rect 603378 79952 603446 80008
rect 603502 79952 603570 80008
rect 603626 79952 603694 80008
rect 603750 79952 603818 80008
rect 603874 79952 603942 80008
rect 603998 79952 604066 80008
rect 604122 79952 604810 80008
rect 604866 79952 604934 80008
rect 604990 79952 605058 80008
rect 605114 79952 605182 80008
rect 605238 79952 605306 80008
rect 605362 79952 605430 80008
rect 605486 79952 605554 80008
rect 605610 79952 605678 80008
rect 605734 79952 605802 80008
rect 605858 79952 605926 80008
rect 605982 79952 606050 80008
rect 606106 79952 606174 80008
rect 606230 79952 606298 80008
rect 606354 79952 606422 80008
rect 606478 79952 606546 80008
rect 606602 79952 606670 80008
rect 606726 79952 607180 80008
rect 607236 79952 607304 80008
rect 607360 79952 607428 80008
rect 607484 79952 607552 80008
rect 607608 79952 607676 80008
rect 607732 79952 607800 80008
rect 607856 79952 607924 80008
rect 607980 79952 608048 80008
rect 608104 79952 608172 80008
rect 608228 79952 608296 80008
rect 608352 79952 608420 80008
rect 608476 79952 608544 80008
rect 608600 79952 608668 80008
rect 608724 79952 608792 80008
rect 608848 79952 608916 80008
rect 608972 79952 609040 80008
rect 609096 79952 609886 80008
rect 609942 79952 610010 80008
rect 610066 79952 610134 80008
rect 610190 79952 610258 80008
rect 610314 79952 610382 80008
rect 610438 79952 610506 80008
rect 610562 79952 610630 80008
rect 610686 79952 610754 80008
rect 610810 79952 610878 80008
rect 610934 79952 611002 80008
rect 611058 79952 611126 80008
rect 611182 79952 611250 80008
rect 611306 79952 611374 80008
rect 611430 79952 611498 80008
rect 611554 79952 611622 80008
rect 611678 79952 611746 80008
rect 611802 79952 612256 80008
rect 612312 79952 612380 80008
rect 612436 79952 612504 80008
rect 612560 79952 612628 80008
rect 612684 79952 612752 80008
rect 612808 79952 612876 80008
rect 612932 79952 613000 80008
rect 613056 79952 613124 80008
rect 613180 79952 613248 80008
rect 613304 79952 613372 80008
rect 613428 79952 613496 80008
rect 613552 79952 613620 80008
rect 613676 79952 613744 80008
rect 613800 79952 613868 80008
rect 613924 79952 613992 80008
rect 614048 79952 614116 80008
rect 614172 79952 614860 80008
rect 614916 79952 614984 80008
rect 615040 79952 615108 80008
rect 615164 79952 615232 80008
rect 615288 79952 615356 80008
rect 615412 79952 615480 80008
rect 615536 79952 615604 80008
rect 615660 79952 615728 80008
rect 615784 79952 615852 80008
rect 615908 79952 615976 80008
rect 616032 79952 616100 80008
rect 616156 79952 616224 80008
rect 616280 79952 616348 80008
rect 616404 79952 616472 80008
rect 616528 79952 616596 80008
rect 616652 79952 628697 80008
rect 628753 79952 628821 80008
rect 628877 79952 636637 80008
rect 636693 79952 636761 80008
rect 636817 79952 644577 80008
rect 644633 79952 644701 80008
rect 644757 79952 670090 80008
rect 670146 79952 670214 80008
rect 670270 79952 670338 80008
rect 670394 79952 670462 80008
rect 670518 79952 670586 80008
rect 670642 79952 670710 80008
rect 670766 79952 698052 80008
rect 698108 79952 698176 80008
rect 698232 79952 698300 80008
rect 698356 79952 698424 80008
rect 698480 79952 698548 80008
rect 698604 79952 698672 80008
rect 698728 79952 698796 80008
rect 698852 79952 698922 80008
rect 79078 79884 698922 79952
rect 79078 79828 79208 79884
rect 79264 79828 79332 79884
rect 79388 79828 79456 79884
rect 79512 79828 79580 79884
rect 79636 79828 79704 79884
rect 79760 79828 79828 79884
rect 79884 79828 79952 79884
rect 80008 79828 99294 79884
rect 99350 79828 99418 79884
rect 99474 79828 107330 79884
rect 107386 79828 107454 79884
rect 107510 79828 107578 79884
rect 107634 79828 107702 79884
rect 107758 79828 107826 79884
rect 107882 79828 107950 79884
rect 108006 79828 108074 79884
rect 108130 79828 108198 79884
rect 108254 79828 108322 79884
rect 108378 79828 108446 79884
rect 108502 79828 108570 79884
rect 108626 79828 108694 79884
rect 108750 79828 108818 79884
rect 108874 79828 108942 79884
rect 108998 79828 109066 79884
rect 109122 79828 109810 79884
rect 109866 79828 109934 79884
rect 109990 79828 110058 79884
rect 110114 79828 110182 79884
rect 110238 79828 110306 79884
rect 110362 79828 110430 79884
rect 110486 79828 110554 79884
rect 110610 79828 110678 79884
rect 110734 79828 110802 79884
rect 110858 79828 110926 79884
rect 110982 79828 111050 79884
rect 111106 79828 111174 79884
rect 111230 79828 111298 79884
rect 111354 79828 111422 79884
rect 111478 79828 111546 79884
rect 111602 79828 111670 79884
rect 111726 79828 112180 79884
rect 112236 79828 112304 79884
rect 112360 79828 112428 79884
rect 112484 79828 112552 79884
rect 112608 79828 112676 79884
rect 112732 79828 112800 79884
rect 112856 79828 112924 79884
rect 112980 79828 113048 79884
rect 113104 79828 113172 79884
rect 113228 79828 113296 79884
rect 113352 79828 113420 79884
rect 113476 79828 113544 79884
rect 113600 79828 113668 79884
rect 113724 79828 113792 79884
rect 113848 79828 113916 79884
rect 113972 79828 114040 79884
rect 114096 79828 114886 79884
rect 114942 79828 115010 79884
rect 115066 79828 115134 79884
rect 115190 79828 115258 79884
rect 115314 79828 115382 79884
rect 115438 79828 115506 79884
rect 115562 79828 115630 79884
rect 115686 79828 115754 79884
rect 115810 79828 115878 79884
rect 115934 79828 116002 79884
rect 116058 79828 116126 79884
rect 116182 79828 116250 79884
rect 116306 79828 116374 79884
rect 116430 79828 116498 79884
rect 116554 79828 116622 79884
rect 116678 79828 116746 79884
rect 116802 79828 117256 79884
rect 117312 79828 117380 79884
rect 117436 79828 117504 79884
rect 117560 79828 117628 79884
rect 117684 79828 117752 79884
rect 117808 79828 117876 79884
rect 117932 79828 118000 79884
rect 118056 79828 118124 79884
rect 118180 79828 118248 79884
rect 118304 79828 118372 79884
rect 118428 79828 118496 79884
rect 118552 79828 118620 79884
rect 118676 79828 118744 79884
rect 118800 79828 118868 79884
rect 118924 79828 118992 79884
rect 119048 79828 119116 79884
rect 119172 79828 119860 79884
rect 119916 79828 119984 79884
rect 120040 79828 120108 79884
rect 120164 79828 120232 79884
rect 120288 79828 120356 79884
rect 120412 79828 120480 79884
rect 120536 79828 120604 79884
rect 120660 79828 120728 79884
rect 120784 79828 120852 79884
rect 120908 79828 120976 79884
rect 121032 79828 121100 79884
rect 121156 79828 121224 79884
rect 121280 79828 121348 79884
rect 121404 79828 121472 79884
rect 121528 79828 121596 79884
rect 121652 79828 129294 79884
rect 129350 79828 129418 79884
rect 129474 79828 139294 79884
rect 139350 79828 139418 79884
rect 139474 79828 149294 79884
rect 149350 79828 149418 79884
rect 149474 79828 159294 79884
rect 159350 79828 159418 79884
rect 159474 79828 169294 79884
rect 169350 79828 169418 79884
rect 169474 79828 179294 79884
rect 179350 79828 179418 79884
rect 179474 79828 189294 79884
rect 189350 79828 189418 79884
rect 189474 79828 199294 79884
rect 199350 79828 199418 79884
rect 199474 79828 209294 79884
rect 209350 79828 209418 79884
rect 209474 79828 219294 79884
rect 219350 79828 219418 79884
rect 219474 79828 229294 79884
rect 229350 79828 229418 79884
rect 229474 79828 239294 79884
rect 239350 79828 239418 79884
rect 239474 79828 249294 79884
rect 249350 79828 249418 79884
rect 249474 79828 259294 79884
rect 259350 79828 259418 79884
rect 259474 79828 269294 79884
rect 269350 79828 269418 79884
rect 269474 79828 272330 79884
rect 272386 79828 272454 79884
rect 272510 79828 272578 79884
rect 272634 79828 272702 79884
rect 272758 79828 272826 79884
rect 272882 79828 272950 79884
rect 273006 79828 273074 79884
rect 273130 79828 273198 79884
rect 273254 79828 273322 79884
rect 273378 79828 273446 79884
rect 273502 79828 273570 79884
rect 273626 79828 273694 79884
rect 273750 79828 273818 79884
rect 273874 79828 273942 79884
rect 273998 79828 274066 79884
rect 274122 79828 274810 79884
rect 274866 79828 274934 79884
rect 274990 79828 275058 79884
rect 275114 79828 275182 79884
rect 275238 79828 275306 79884
rect 275362 79828 275430 79884
rect 275486 79828 275554 79884
rect 275610 79828 275678 79884
rect 275734 79828 275802 79884
rect 275858 79828 275926 79884
rect 275982 79828 276050 79884
rect 276106 79828 276174 79884
rect 276230 79828 276298 79884
rect 276354 79828 276422 79884
rect 276478 79828 276546 79884
rect 276602 79828 276670 79884
rect 276726 79828 277180 79884
rect 277236 79828 277304 79884
rect 277360 79828 277428 79884
rect 277484 79828 277552 79884
rect 277608 79828 277676 79884
rect 277732 79828 277800 79884
rect 277856 79828 277924 79884
rect 277980 79828 278048 79884
rect 278104 79828 278172 79884
rect 278228 79828 278296 79884
rect 278352 79828 278420 79884
rect 278476 79828 278544 79884
rect 278600 79828 278668 79884
rect 278724 79828 278792 79884
rect 278848 79828 278916 79884
rect 278972 79828 279040 79884
rect 279096 79828 279886 79884
rect 279942 79828 280010 79884
rect 280066 79828 280134 79884
rect 280190 79828 280258 79884
rect 280314 79828 280382 79884
rect 280438 79828 280506 79884
rect 280562 79828 280630 79884
rect 280686 79828 280754 79884
rect 280810 79828 280878 79884
rect 280934 79828 281002 79884
rect 281058 79828 281126 79884
rect 281182 79828 281250 79884
rect 281306 79828 281374 79884
rect 281430 79828 281498 79884
rect 281554 79828 281622 79884
rect 281678 79828 281746 79884
rect 281802 79828 282256 79884
rect 282312 79828 282380 79884
rect 282436 79828 282504 79884
rect 282560 79828 282628 79884
rect 282684 79828 282752 79884
rect 282808 79828 282876 79884
rect 282932 79828 283000 79884
rect 283056 79828 283124 79884
rect 283180 79828 283248 79884
rect 283304 79828 283372 79884
rect 283428 79828 283496 79884
rect 283552 79828 283620 79884
rect 283676 79828 283744 79884
rect 283800 79828 283868 79884
rect 283924 79828 283992 79884
rect 284048 79828 284116 79884
rect 284172 79828 284860 79884
rect 284916 79828 284984 79884
rect 285040 79828 285108 79884
rect 285164 79828 285232 79884
rect 285288 79828 285356 79884
rect 285412 79828 285480 79884
rect 285536 79828 285604 79884
rect 285660 79828 285728 79884
rect 285784 79828 285852 79884
rect 285908 79828 285976 79884
rect 286032 79828 286100 79884
rect 286156 79828 286224 79884
rect 286280 79828 286348 79884
rect 286404 79828 286472 79884
rect 286528 79828 286596 79884
rect 286652 79828 289294 79884
rect 289350 79828 289418 79884
rect 289474 79828 299294 79884
rect 299350 79828 299418 79884
rect 299474 79828 309294 79884
rect 309350 79828 309418 79884
rect 309474 79828 319294 79884
rect 319350 79828 319418 79884
rect 319474 79828 329294 79884
rect 329350 79828 329418 79884
rect 329474 79828 339294 79884
rect 339350 79828 339418 79884
rect 339474 79828 349294 79884
rect 349350 79828 349418 79884
rect 349474 79828 359294 79884
rect 359350 79828 359418 79884
rect 359474 79828 369294 79884
rect 369350 79828 369418 79884
rect 369474 79828 379294 79884
rect 379350 79828 379418 79884
rect 379474 79828 389294 79884
rect 389350 79828 389418 79884
rect 389474 79828 399294 79884
rect 399350 79828 399418 79884
rect 399474 79828 409294 79884
rect 409350 79828 409418 79884
rect 409474 79828 419294 79884
rect 419350 79828 419418 79884
rect 419474 79828 429294 79884
rect 429350 79828 429418 79884
rect 429474 79828 439294 79884
rect 439350 79828 439418 79884
rect 439474 79828 449294 79884
rect 449350 79828 449418 79884
rect 449474 79828 459294 79884
rect 459350 79828 459418 79884
rect 459474 79828 469294 79884
rect 469350 79828 469418 79884
rect 469474 79828 479294 79884
rect 479350 79828 479418 79884
rect 479474 79828 489294 79884
rect 489350 79828 489418 79884
rect 489474 79828 499294 79884
rect 499350 79828 499418 79884
rect 499474 79828 509294 79884
rect 509350 79828 509418 79884
rect 509474 79828 519294 79884
rect 519350 79828 519418 79884
rect 519474 79828 529294 79884
rect 529350 79828 529418 79884
rect 529474 79828 539294 79884
rect 539350 79828 539418 79884
rect 539474 79828 549294 79884
rect 549350 79828 549418 79884
rect 549474 79828 590970 79884
rect 591026 79828 591094 79884
rect 591150 79828 591218 79884
rect 591274 79828 591342 79884
rect 591398 79828 591466 79884
rect 591522 79828 591590 79884
rect 591646 79828 591714 79884
rect 591770 79828 602330 79884
rect 602386 79828 602454 79884
rect 602510 79828 602578 79884
rect 602634 79828 602702 79884
rect 602758 79828 602826 79884
rect 602882 79828 602950 79884
rect 603006 79828 603074 79884
rect 603130 79828 603198 79884
rect 603254 79828 603322 79884
rect 603378 79828 603446 79884
rect 603502 79828 603570 79884
rect 603626 79828 603694 79884
rect 603750 79828 603818 79884
rect 603874 79828 603942 79884
rect 603998 79828 604066 79884
rect 604122 79828 604810 79884
rect 604866 79828 604934 79884
rect 604990 79828 605058 79884
rect 605114 79828 605182 79884
rect 605238 79828 605306 79884
rect 605362 79828 605430 79884
rect 605486 79828 605554 79884
rect 605610 79828 605678 79884
rect 605734 79828 605802 79884
rect 605858 79828 605926 79884
rect 605982 79828 606050 79884
rect 606106 79828 606174 79884
rect 606230 79828 606298 79884
rect 606354 79828 606422 79884
rect 606478 79828 606546 79884
rect 606602 79828 606670 79884
rect 606726 79828 607180 79884
rect 607236 79828 607304 79884
rect 607360 79828 607428 79884
rect 607484 79828 607552 79884
rect 607608 79828 607676 79884
rect 607732 79828 607800 79884
rect 607856 79828 607924 79884
rect 607980 79828 608048 79884
rect 608104 79828 608172 79884
rect 608228 79828 608296 79884
rect 608352 79828 608420 79884
rect 608476 79828 608544 79884
rect 608600 79828 608668 79884
rect 608724 79828 608792 79884
rect 608848 79828 608916 79884
rect 608972 79828 609040 79884
rect 609096 79828 609886 79884
rect 609942 79828 610010 79884
rect 610066 79828 610134 79884
rect 610190 79828 610258 79884
rect 610314 79828 610382 79884
rect 610438 79828 610506 79884
rect 610562 79828 610630 79884
rect 610686 79828 610754 79884
rect 610810 79828 610878 79884
rect 610934 79828 611002 79884
rect 611058 79828 611126 79884
rect 611182 79828 611250 79884
rect 611306 79828 611374 79884
rect 611430 79828 611498 79884
rect 611554 79828 611622 79884
rect 611678 79828 611746 79884
rect 611802 79828 612256 79884
rect 612312 79828 612380 79884
rect 612436 79828 612504 79884
rect 612560 79828 612628 79884
rect 612684 79828 612752 79884
rect 612808 79828 612876 79884
rect 612932 79828 613000 79884
rect 613056 79828 613124 79884
rect 613180 79828 613248 79884
rect 613304 79828 613372 79884
rect 613428 79828 613496 79884
rect 613552 79828 613620 79884
rect 613676 79828 613744 79884
rect 613800 79828 613868 79884
rect 613924 79828 613992 79884
rect 614048 79828 614116 79884
rect 614172 79828 614860 79884
rect 614916 79828 614984 79884
rect 615040 79828 615108 79884
rect 615164 79828 615232 79884
rect 615288 79828 615356 79884
rect 615412 79828 615480 79884
rect 615536 79828 615604 79884
rect 615660 79828 615728 79884
rect 615784 79828 615852 79884
rect 615908 79828 615976 79884
rect 616032 79828 616100 79884
rect 616156 79828 616224 79884
rect 616280 79828 616348 79884
rect 616404 79828 616472 79884
rect 616528 79828 616596 79884
rect 616652 79828 628697 79884
rect 628753 79828 628821 79884
rect 628877 79828 636637 79884
rect 636693 79828 636761 79884
rect 636817 79828 644577 79884
rect 644633 79828 644701 79884
rect 644757 79828 670090 79884
rect 670146 79828 670214 79884
rect 670270 79828 670338 79884
rect 670394 79828 670462 79884
rect 670518 79828 670586 79884
rect 670642 79828 670710 79884
rect 670766 79828 698052 79884
rect 698108 79828 698176 79884
rect 698232 79828 698300 79884
rect 698356 79828 698424 79884
rect 698480 79828 698548 79884
rect 698604 79828 698672 79884
rect 698728 79828 698796 79884
rect 698852 79828 698922 79884
rect 79078 79760 698922 79828
rect 79078 79704 79208 79760
rect 79264 79704 79332 79760
rect 79388 79704 79456 79760
rect 79512 79704 79580 79760
rect 79636 79704 79704 79760
rect 79760 79704 79828 79760
rect 79884 79704 79952 79760
rect 80008 79704 99294 79760
rect 99350 79704 99418 79760
rect 99474 79704 107330 79760
rect 107386 79704 107454 79760
rect 107510 79704 107578 79760
rect 107634 79704 107702 79760
rect 107758 79704 107826 79760
rect 107882 79704 107950 79760
rect 108006 79704 108074 79760
rect 108130 79704 108198 79760
rect 108254 79704 108322 79760
rect 108378 79704 108446 79760
rect 108502 79704 108570 79760
rect 108626 79704 108694 79760
rect 108750 79704 108818 79760
rect 108874 79704 108942 79760
rect 108998 79704 109066 79760
rect 109122 79704 109810 79760
rect 109866 79704 109934 79760
rect 109990 79704 110058 79760
rect 110114 79704 110182 79760
rect 110238 79704 110306 79760
rect 110362 79704 110430 79760
rect 110486 79704 110554 79760
rect 110610 79704 110678 79760
rect 110734 79704 110802 79760
rect 110858 79704 110926 79760
rect 110982 79704 111050 79760
rect 111106 79704 111174 79760
rect 111230 79704 111298 79760
rect 111354 79704 111422 79760
rect 111478 79704 111546 79760
rect 111602 79704 111670 79760
rect 111726 79704 112180 79760
rect 112236 79704 112304 79760
rect 112360 79704 112428 79760
rect 112484 79704 112552 79760
rect 112608 79704 112676 79760
rect 112732 79704 112800 79760
rect 112856 79704 112924 79760
rect 112980 79704 113048 79760
rect 113104 79704 113172 79760
rect 113228 79704 113296 79760
rect 113352 79704 113420 79760
rect 113476 79704 113544 79760
rect 113600 79704 113668 79760
rect 113724 79704 113792 79760
rect 113848 79704 113916 79760
rect 113972 79704 114040 79760
rect 114096 79704 114886 79760
rect 114942 79704 115010 79760
rect 115066 79704 115134 79760
rect 115190 79704 115258 79760
rect 115314 79704 115382 79760
rect 115438 79704 115506 79760
rect 115562 79704 115630 79760
rect 115686 79704 115754 79760
rect 115810 79704 115878 79760
rect 115934 79704 116002 79760
rect 116058 79704 116126 79760
rect 116182 79704 116250 79760
rect 116306 79704 116374 79760
rect 116430 79704 116498 79760
rect 116554 79704 116622 79760
rect 116678 79704 116746 79760
rect 116802 79704 117256 79760
rect 117312 79704 117380 79760
rect 117436 79704 117504 79760
rect 117560 79704 117628 79760
rect 117684 79704 117752 79760
rect 117808 79704 117876 79760
rect 117932 79704 118000 79760
rect 118056 79704 118124 79760
rect 118180 79704 118248 79760
rect 118304 79704 118372 79760
rect 118428 79704 118496 79760
rect 118552 79704 118620 79760
rect 118676 79704 118744 79760
rect 118800 79704 118868 79760
rect 118924 79704 118992 79760
rect 119048 79704 119116 79760
rect 119172 79704 119860 79760
rect 119916 79704 119984 79760
rect 120040 79704 120108 79760
rect 120164 79704 120232 79760
rect 120288 79704 120356 79760
rect 120412 79704 120480 79760
rect 120536 79704 120604 79760
rect 120660 79704 120728 79760
rect 120784 79704 120852 79760
rect 120908 79704 120976 79760
rect 121032 79704 121100 79760
rect 121156 79704 121224 79760
rect 121280 79704 121348 79760
rect 121404 79704 121472 79760
rect 121528 79704 121596 79760
rect 121652 79704 129294 79760
rect 129350 79704 129418 79760
rect 129474 79704 139294 79760
rect 139350 79704 139418 79760
rect 139474 79704 149294 79760
rect 149350 79704 149418 79760
rect 149474 79704 159294 79760
rect 159350 79704 159418 79760
rect 159474 79704 169294 79760
rect 169350 79704 169418 79760
rect 169474 79704 179294 79760
rect 179350 79704 179418 79760
rect 179474 79704 189294 79760
rect 189350 79704 189418 79760
rect 189474 79704 199294 79760
rect 199350 79704 199418 79760
rect 199474 79704 209294 79760
rect 209350 79704 209418 79760
rect 209474 79704 219294 79760
rect 219350 79704 219418 79760
rect 219474 79704 229294 79760
rect 229350 79704 229418 79760
rect 229474 79704 239294 79760
rect 239350 79704 239418 79760
rect 239474 79704 249294 79760
rect 249350 79704 249418 79760
rect 249474 79704 259294 79760
rect 259350 79704 259418 79760
rect 259474 79704 269294 79760
rect 269350 79704 269418 79760
rect 269474 79704 272330 79760
rect 272386 79704 272454 79760
rect 272510 79704 272578 79760
rect 272634 79704 272702 79760
rect 272758 79704 272826 79760
rect 272882 79704 272950 79760
rect 273006 79704 273074 79760
rect 273130 79704 273198 79760
rect 273254 79704 273322 79760
rect 273378 79704 273446 79760
rect 273502 79704 273570 79760
rect 273626 79704 273694 79760
rect 273750 79704 273818 79760
rect 273874 79704 273942 79760
rect 273998 79704 274066 79760
rect 274122 79704 274810 79760
rect 274866 79704 274934 79760
rect 274990 79704 275058 79760
rect 275114 79704 275182 79760
rect 275238 79704 275306 79760
rect 275362 79704 275430 79760
rect 275486 79704 275554 79760
rect 275610 79704 275678 79760
rect 275734 79704 275802 79760
rect 275858 79704 275926 79760
rect 275982 79704 276050 79760
rect 276106 79704 276174 79760
rect 276230 79704 276298 79760
rect 276354 79704 276422 79760
rect 276478 79704 276546 79760
rect 276602 79704 276670 79760
rect 276726 79704 277180 79760
rect 277236 79704 277304 79760
rect 277360 79704 277428 79760
rect 277484 79704 277552 79760
rect 277608 79704 277676 79760
rect 277732 79704 277800 79760
rect 277856 79704 277924 79760
rect 277980 79704 278048 79760
rect 278104 79704 278172 79760
rect 278228 79704 278296 79760
rect 278352 79704 278420 79760
rect 278476 79704 278544 79760
rect 278600 79704 278668 79760
rect 278724 79704 278792 79760
rect 278848 79704 278916 79760
rect 278972 79704 279040 79760
rect 279096 79704 279886 79760
rect 279942 79704 280010 79760
rect 280066 79704 280134 79760
rect 280190 79704 280258 79760
rect 280314 79704 280382 79760
rect 280438 79704 280506 79760
rect 280562 79704 280630 79760
rect 280686 79704 280754 79760
rect 280810 79704 280878 79760
rect 280934 79704 281002 79760
rect 281058 79704 281126 79760
rect 281182 79704 281250 79760
rect 281306 79704 281374 79760
rect 281430 79704 281498 79760
rect 281554 79704 281622 79760
rect 281678 79704 281746 79760
rect 281802 79704 282256 79760
rect 282312 79704 282380 79760
rect 282436 79704 282504 79760
rect 282560 79704 282628 79760
rect 282684 79704 282752 79760
rect 282808 79704 282876 79760
rect 282932 79704 283000 79760
rect 283056 79704 283124 79760
rect 283180 79704 283248 79760
rect 283304 79704 283372 79760
rect 283428 79704 283496 79760
rect 283552 79704 283620 79760
rect 283676 79704 283744 79760
rect 283800 79704 283868 79760
rect 283924 79704 283992 79760
rect 284048 79704 284116 79760
rect 284172 79704 284860 79760
rect 284916 79704 284984 79760
rect 285040 79704 285108 79760
rect 285164 79704 285232 79760
rect 285288 79704 285356 79760
rect 285412 79704 285480 79760
rect 285536 79704 285604 79760
rect 285660 79704 285728 79760
rect 285784 79704 285852 79760
rect 285908 79704 285976 79760
rect 286032 79704 286100 79760
rect 286156 79704 286224 79760
rect 286280 79704 286348 79760
rect 286404 79704 286472 79760
rect 286528 79704 286596 79760
rect 286652 79704 289294 79760
rect 289350 79704 289418 79760
rect 289474 79704 299294 79760
rect 299350 79704 299418 79760
rect 299474 79704 309294 79760
rect 309350 79704 309418 79760
rect 309474 79704 319294 79760
rect 319350 79704 319418 79760
rect 319474 79704 329294 79760
rect 329350 79704 329418 79760
rect 329474 79704 339294 79760
rect 339350 79704 339418 79760
rect 339474 79704 349294 79760
rect 349350 79704 349418 79760
rect 349474 79704 359294 79760
rect 359350 79704 359418 79760
rect 359474 79704 369294 79760
rect 369350 79704 369418 79760
rect 369474 79704 379294 79760
rect 379350 79704 379418 79760
rect 379474 79704 389294 79760
rect 389350 79704 389418 79760
rect 389474 79704 399294 79760
rect 399350 79704 399418 79760
rect 399474 79704 409294 79760
rect 409350 79704 409418 79760
rect 409474 79704 419294 79760
rect 419350 79704 419418 79760
rect 419474 79704 429294 79760
rect 429350 79704 429418 79760
rect 429474 79704 439294 79760
rect 439350 79704 439418 79760
rect 439474 79704 449294 79760
rect 449350 79704 449418 79760
rect 449474 79704 459294 79760
rect 459350 79704 459418 79760
rect 459474 79704 469294 79760
rect 469350 79704 469418 79760
rect 469474 79704 479294 79760
rect 479350 79704 479418 79760
rect 479474 79704 489294 79760
rect 489350 79704 489418 79760
rect 489474 79704 499294 79760
rect 499350 79704 499418 79760
rect 499474 79704 509294 79760
rect 509350 79704 509418 79760
rect 509474 79704 519294 79760
rect 519350 79704 519418 79760
rect 519474 79704 529294 79760
rect 529350 79704 529418 79760
rect 529474 79704 539294 79760
rect 539350 79704 539418 79760
rect 539474 79704 549294 79760
rect 549350 79704 549418 79760
rect 549474 79704 590970 79760
rect 591026 79704 591094 79760
rect 591150 79704 591218 79760
rect 591274 79704 591342 79760
rect 591398 79704 591466 79760
rect 591522 79704 591590 79760
rect 591646 79704 591714 79760
rect 591770 79704 602330 79760
rect 602386 79704 602454 79760
rect 602510 79704 602578 79760
rect 602634 79704 602702 79760
rect 602758 79704 602826 79760
rect 602882 79704 602950 79760
rect 603006 79704 603074 79760
rect 603130 79704 603198 79760
rect 603254 79704 603322 79760
rect 603378 79704 603446 79760
rect 603502 79704 603570 79760
rect 603626 79704 603694 79760
rect 603750 79704 603818 79760
rect 603874 79704 603942 79760
rect 603998 79704 604066 79760
rect 604122 79704 604810 79760
rect 604866 79704 604934 79760
rect 604990 79704 605058 79760
rect 605114 79704 605182 79760
rect 605238 79704 605306 79760
rect 605362 79704 605430 79760
rect 605486 79704 605554 79760
rect 605610 79704 605678 79760
rect 605734 79704 605802 79760
rect 605858 79704 605926 79760
rect 605982 79704 606050 79760
rect 606106 79704 606174 79760
rect 606230 79704 606298 79760
rect 606354 79704 606422 79760
rect 606478 79704 606546 79760
rect 606602 79704 606670 79760
rect 606726 79704 607180 79760
rect 607236 79704 607304 79760
rect 607360 79704 607428 79760
rect 607484 79704 607552 79760
rect 607608 79704 607676 79760
rect 607732 79704 607800 79760
rect 607856 79704 607924 79760
rect 607980 79704 608048 79760
rect 608104 79704 608172 79760
rect 608228 79704 608296 79760
rect 608352 79704 608420 79760
rect 608476 79704 608544 79760
rect 608600 79704 608668 79760
rect 608724 79704 608792 79760
rect 608848 79704 608916 79760
rect 608972 79704 609040 79760
rect 609096 79704 609886 79760
rect 609942 79704 610010 79760
rect 610066 79704 610134 79760
rect 610190 79704 610258 79760
rect 610314 79704 610382 79760
rect 610438 79704 610506 79760
rect 610562 79704 610630 79760
rect 610686 79704 610754 79760
rect 610810 79704 610878 79760
rect 610934 79704 611002 79760
rect 611058 79704 611126 79760
rect 611182 79704 611250 79760
rect 611306 79704 611374 79760
rect 611430 79704 611498 79760
rect 611554 79704 611622 79760
rect 611678 79704 611746 79760
rect 611802 79704 612256 79760
rect 612312 79704 612380 79760
rect 612436 79704 612504 79760
rect 612560 79704 612628 79760
rect 612684 79704 612752 79760
rect 612808 79704 612876 79760
rect 612932 79704 613000 79760
rect 613056 79704 613124 79760
rect 613180 79704 613248 79760
rect 613304 79704 613372 79760
rect 613428 79704 613496 79760
rect 613552 79704 613620 79760
rect 613676 79704 613744 79760
rect 613800 79704 613868 79760
rect 613924 79704 613992 79760
rect 614048 79704 614116 79760
rect 614172 79704 614860 79760
rect 614916 79704 614984 79760
rect 615040 79704 615108 79760
rect 615164 79704 615232 79760
rect 615288 79704 615356 79760
rect 615412 79704 615480 79760
rect 615536 79704 615604 79760
rect 615660 79704 615728 79760
rect 615784 79704 615852 79760
rect 615908 79704 615976 79760
rect 616032 79704 616100 79760
rect 616156 79704 616224 79760
rect 616280 79704 616348 79760
rect 616404 79704 616472 79760
rect 616528 79704 616596 79760
rect 616652 79704 628697 79760
rect 628753 79704 628821 79760
rect 628877 79704 636637 79760
rect 636693 79704 636761 79760
rect 636817 79704 644577 79760
rect 644633 79704 644701 79760
rect 644757 79704 670090 79760
rect 670146 79704 670214 79760
rect 670270 79704 670338 79760
rect 670394 79704 670462 79760
rect 670518 79704 670586 79760
rect 670642 79704 670710 79760
rect 670766 79704 698052 79760
rect 698108 79704 698176 79760
rect 698232 79704 698300 79760
rect 698356 79704 698424 79760
rect 698480 79704 698548 79760
rect 698604 79704 698672 79760
rect 698728 79704 698796 79760
rect 698852 79704 698922 79760
rect 79078 79636 698922 79704
rect 79078 79580 79208 79636
rect 79264 79580 79332 79636
rect 79388 79580 79456 79636
rect 79512 79580 79580 79636
rect 79636 79580 79704 79636
rect 79760 79580 79828 79636
rect 79884 79580 79952 79636
rect 80008 79580 99294 79636
rect 99350 79580 99418 79636
rect 99474 79580 107330 79636
rect 107386 79580 107454 79636
rect 107510 79580 107578 79636
rect 107634 79580 107702 79636
rect 107758 79580 107826 79636
rect 107882 79580 107950 79636
rect 108006 79580 108074 79636
rect 108130 79580 108198 79636
rect 108254 79580 108322 79636
rect 108378 79580 108446 79636
rect 108502 79580 108570 79636
rect 108626 79580 108694 79636
rect 108750 79580 108818 79636
rect 108874 79580 108942 79636
rect 108998 79580 109066 79636
rect 109122 79580 109810 79636
rect 109866 79580 109934 79636
rect 109990 79580 110058 79636
rect 110114 79580 110182 79636
rect 110238 79580 110306 79636
rect 110362 79580 110430 79636
rect 110486 79580 110554 79636
rect 110610 79580 110678 79636
rect 110734 79580 110802 79636
rect 110858 79580 110926 79636
rect 110982 79580 111050 79636
rect 111106 79580 111174 79636
rect 111230 79580 111298 79636
rect 111354 79580 111422 79636
rect 111478 79580 111546 79636
rect 111602 79580 111670 79636
rect 111726 79580 112180 79636
rect 112236 79580 112304 79636
rect 112360 79580 112428 79636
rect 112484 79580 112552 79636
rect 112608 79580 112676 79636
rect 112732 79580 112800 79636
rect 112856 79580 112924 79636
rect 112980 79580 113048 79636
rect 113104 79580 113172 79636
rect 113228 79580 113296 79636
rect 113352 79580 113420 79636
rect 113476 79580 113544 79636
rect 113600 79580 113668 79636
rect 113724 79580 113792 79636
rect 113848 79580 113916 79636
rect 113972 79580 114040 79636
rect 114096 79580 114886 79636
rect 114942 79580 115010 79636
rect 115066 79580 115134 79636
rect 115190 79580 115258 79636
rect 115314 79580 115382 79636
rect 115438 79580 115506 79636
rect 115562 79580 115630 79636
rect 115686 79580 115754 79636
rect 115810 79580 115878 79636
rect 115934 79580 116002 79636
rect 116058 79580 116126 79636
rect 116182 79580 116250 79636
rect 116306 79580 116374 79636
rect 116430 79580 116498 79636
rect 116554 79580 116622 79636
rect 116678 79580 116746 79636
rect 116802 79580 117256 79636
rect 117312 79580 117380 79636
rect 117436 79580 117504 79636
rect 117560 79580 117628 79636
rect 117684 79580 117752 79636
rect 117808 79580 117876 79636
rect 117932 79580 118000 79636
rect 118056 79580 118124 79636
rect 118180 79580 118248 79636
rect 118304 79580 118372 79636
rect 118428 79580 118496 79636
rect 118552 79580 118620 79636
rect 118676 79580 118744 79636
rect 118800 79580 118868 79636
rect 118924 79580 118992 79636
rect 119048 79580 119116 79636
rect 119172 79580 119860 79636
rect 119916 79580 119984 79636
rect 120040 79580 120108 79636
rect 120164 79580 120232 79636
rect 120288 79580 120356 79636
rect 120412 79580 120480 79636
rect 120536 79580 120604 79636
rect 120660 79580 120728 79636
rect 120784 79580 120852 79636
rect 120908 79580 120976 79636
rect 121032 79580 121100 79636
rect 121156 79580 121224 79636
rect 121280 79580 121348 79636
rect 121404 79580 121472 79636
rect 121528 79580 121596 79636
rect 121652 79580 129294 79636
rect 129350 79580 129418 79636
rect 129474 79580 139294 79636
rect 139350 79580 139418 79636
rect 139474 79580 149294 79636
rect 149350 79580 149418 79636
rect 149474 79580 159294 79636
rect 159350 79580 159418 79636
rect 159474 79580 169294 79636
rect 169350 79580 169418 79636
rect 169474 79580 179294 79636
rect 179350 79580 179418 79636
rect 179474 79580 189294 79636
rect 189350 79580 189418 79636
rect 189474 79580 199294 79636
rect 199350 79580 199418 79636
rect 199474 79580 209294 79636
rect 209350 79580 209418 79636
rect 209474 79580 219294 79636
rect 219350 79580 219418 79636
rect 219474 79580 229294 79636
rect 229350 79580 229418 79636
rect 229474 79580 239294 79636
rect 239350 79580 239418 79636
rect 239474 79580 249294 79636
rect 249350 79580 249418 79636
rect 249474 79580 259294 79636
rect 259350 79580 259418 79636
rect 259474 79580 269294 79636
rect 269350 79580 269418 79636
rect 269474 79580 272330 79636
rect 272386 79580 272454 79636
rect 272510 79580 272578 79636
rect 272634 79580 272702 79636
rect 272758 79580 272826 79636
rect 272882 79580 272950 79636
rect 273006 79580 273074 79636
rect 273130 79580 273198 79636
rect 273254 79580 273322 79636
rect 273378 79580 273446 79636
rect 273502 79580 273570 79636
rect 273626 79580 273694 79636
rect 273750 79580 273818 79636
rect 273874 79580 273942 79636
rect 273998 79580 274066 79636
rect 274122 79580 274810 79636
rect 274866 79580 274934 79636
rect 274990 79580 275058 79636
rect 275114 79580 275182 79636
rect 275238 79580 275306 79636
rect 275362 79580 275430 79636
rect 275486 79580 275554 79636
rect 275610 79580 275678 79636
rect 275734 79580 275802 79636
rect 275858 79580 275926 79636
rect 275982 79580 276050 79636
rect 276106 79580 276174 79636
rect 276230 79580 276298 79636
rect 276354 79580 276422 79636
rect 276478 79580 276546 79636
rect 276602 79580 276670 79636
rect 276726 79580 277180 79636
rect 277236 79580 277304 79636
rect 277360 79580 277428 79636
rect 277484 79580 277552 79636
rect 277608 79580 277676 79636
rect 277732 79580 277800 79636
rect 277856 79580 277924 79636
rect 277980 79580 278048 79636
rect 278104 79580 278172 79636
rect 278228 79580 278296 79636
rect 278352 79580 278420 79636
rect 278476 79580 278544 79636
rect 278600 79580 278668 79636
rect 278724 79580 278792 79636
rect 278848 79580 278916 79636
rect 278972 79580 279040 79636
rect 279096 79580 279886 79636
rect 279942 79580 280010 79636
rect 280066 79580 280134 79636
rect 280190 79580 280258 79636
rect 280314 79580 280382 79636
rect 280438 79580 280506 79636
rect 280562 79580 280630 79636
rect 280686 79580 280754 79636
rect 280810 79580 280878 79636
rect 280934 79580 281002 79636
rect 281058 79580 281126 79636
rect 281182 79580 281250 79636
rect 281306 79580 281374 79636
rect 281430 79580 281498 79636
rect 281554 79580 281622 79636
rect 281678 79580 281746 79636
rect 281802 79580 282256 79636
rect 282312 79580 282380 79636
rect 282436 79580 282504 79636
rect 282560 79580 282628 79636
rect 282684 79580 282752 79636
rect 282808 79580 282876 79636
rect 282932 79580 283000 79636
rect 283056 79580 283124 79636
rect 283180 79580 283248 79636
rect 283304 79580 283372 79636
rect 283428 79580 283496 79636
rect 283552 79580 283620 79636
rect 283676 79580 283744 79636
rect 283800 79580 283868 79636
rect 283924 79580 283992 79636
rect 284048 79580 284116 79636
rect 284172 79580 284860 79636
rect 284916 79580 284984 79636
rect 285040 79580 285108 79636
rect 285164 79580 285232 79636
rect 285288 79580 285356 79636
rect 285412 79580 285480 79636
rect 285536 79580 285604 79636
rect 285660 79580 285728 79636
rect 285784 79580 285852 79636
rect 285908 79580 285976 79636
rect 286032 79580 286100 79636
rect 286156 79580 286224 79636
rect 286280 79580 286348 79636
rect 286404 79580 286472 79636
rect 286528 79580 286596 79636
rect 286652 79580 289294 79636
rect 289350 79580 289418 79636
rect 289474 79580 299294 79636
rect 299350 79580 299418 79636
rect 299474 79580 309294 79636
rect 309350 79580 309418 79636
rect 309474 79580 319294 79636
rect 319350 79580 319418 79636
rect 319474 79580 329294 79636
rect 329350 79580 329418 79636
rect 329474 79580 339294 79636
rect 339350 79580 339418 79636
rect 339474 79580 349294 79636
rect 349350 79580 349418 79636
rect 349474 79580 359294 79636
rect 359350 79580 359418 79636
rect 359474 79580 369294 79636
rect 369350 79580 369418 79636
rect 369474 79580 379294 79636
rect 379350 79580 379418 79636
rect 379474 79580 389294 79636
rect 389350 79580 389418 79636
rect 389474 79580 399294 79636
rect 399350 79580 399418 79636
rect 399474 79580 409294 79636
rect 409350 79580 409418 79636
rect 409474 79580 419294 79636
rect 419350 79580 419418 79636
rect 419474 79580 429294 79636
rect 429350 79580 429418 79636
rect 429474 79580 439294 79636
rect 439350 79580 439418 79636
rect 439474 79580 449294 79636
rect 449350 79580 449418 79636
rect 449474 79580 459294 79636
rect 459350 79580 459418 79636
rect 459474 79580 469294 79636
rect 469350 79580 469418 79636
rect 469474 79580 479294 79636
rect 479350 79580 479418 79636
rect 479474 79580 489294 79636
rect 489350 79580 489418 79636
rect 489474 79580 499294 79636
rect 499350 79580 499418 79636
rect 499474 79580 509294 79636
rect 509350 79580 509418 79636
rect 509474 79580 519294 79636
rect 519350 79580 519418 79636
rect 519474 79580 529294 79636
rect 529350 79580 529418 79636
rect 529474 79580 539294 79636
rect 539350 79580 539418 79636
rect 539474 79580 549294 79636
rect 549350 79580 549418 79636
rect 549474 79580 590970 79636
rect 591026 79580 591094 79636
rect 591150 79580 591218 79636
rect 591274 79580 591342 79636
rect 591398 79580 591466 79636
rect 591522 79580 591590 79636
rect 591646 79580 591714 79636
rect 591770 79580 602330 79636
rect 602386 79580 602454 79636
rect 602510 79580 602578 79636
rect 602634 79580 602702 79636
rect 602758 79580 602826 79636
rect 602882 79580 602950 79636
rect 603006 79580 603074 79636
rect 603130 79580 603198 79636
rect 603254 79580 603322 79636
rect 603378 79580 603446 79636
rect 603502 79580 603570 79636
rect 603626 79580 603694 79636
rect 603750 79580 603818 79636
rect 603874 79580 603942 79636
rect 603998 79580 604066 79636
rect 604122 79580 604810 79636
rect 604866 79580 604934 79636
rect 604990 79580 605058 79636
rect 605114 79580 605182 79636
rect 605238 79580 605306 79636
rect 605362 79580 605430 79636
rect 605486 79580 605554 79636
rect 605610 79580 605678 79636
rect 605734 79580 605802 79636
rect 605858 79580 605926 79636
rect 605982 79580 606050 79636
rect 606106 79580 606174 79636
rect 606230 79580 606298 79636
rect 606354 79580 606422 79636
rect 606478 79580 606546 79636
rect 606602 79580 606670 79636
rect 606726 79580 607180 79636
rect 607236 79580 607304 79636
rect 607360 79580 607428 79636
rect 607484 79580 607552 79636
rect 607608 79580 607676 79636
rect 607732 79580 607800 79636
rect 607856 79580 607924 79636
rect 607980 79580 608048 79636
rect 608104 79580 608172 79636
rect 608228 79580 608296 79636
rect 608352 79580 608420 79636
rect 608476 79580 608544 79636
rect 608600 79580 608668 79636
rect 608724 79580 608792 79636
rect 608848 79580 608916 79636
rect 608972 79580 609040 79636
rect 609096 79580 609886 79636
rect 609942 79580 610010 79636
rect 610066 79580 610134 79636
rect 610190 79580 610258 79636
rect 610314 79580 610382 79636
rect 610438 79580 610506 79636
rect 610562 79580 610630 79636
rect 610686 79580 610754 79636
rect 610810 79580 610878 79636
rect 610934 79580 611002 79636
rect 611058 79580 611126 79636
rect 611182 79580 611250 79636
rect 611306 79580 611374 79636
rect 611430 79580 611498 79636
rect 611554 79580 611622 79636
rect 611678 79580 611746 79636
rect 611802 79580 612256 79636
rect 612312 79580 612380 79636
rect 612436 79580 612504 79636
rect 612560 79580 612628 79636
rect 612684 79580 612752 79636
rect 612808 79580 612876 79636
rect 612932 79580 613000 79636
rect 613056 79580 613124 79636
rect 613180 79580 613248 79636
rect 613304 79580 613372 79636
rect 613428 79580 613496 79636
rect 613552 79580 613620 79636
rect 613676 79580 613744 79636
rect 613800 79580 613868 79636
rect 613924 79580 613992 79636
rect 614048 79580 614116 79636
rect 614172 79580 614860 79636
rect 614916 79580 614984 79636
rect 615040 79580 615108 79636
rect 615164 79580 615232 79636
rect 615288 79580 615356 79636
rect 615412 79580 615480 79636
rect 615536 79580 615604 79636
rect 615660 79580 615728 79636
rect 615784 79580 615852 79636
rect 615908 79580 615976 79636
rect 616032 79580 616100 79636
rect 616156 79580 616224 79636
rect 616280 79580 616348 79636
rect 616404 79580 616472 79636
rect 616528 79580 616596 79636
rect 616652 79580 628697 79636
rect 628753 79580 628821 79636
rect 628877 79580 636637 79636
rect 636693 79580 636761 79636
rect 636817 79580 644577 79636
rect 644633 79580 644701 79636
rect 644757 79580 670090 79636
rect 670146 79580 670214 79636
rect 670270 79580 670338 79636
rect 670394 79580 670462 79636
rect 670518 79580 670586 79636
rect 670642 79580 670710 79636
rect 670766 79580 698052 79636
rect 698108 79580 698176 79636
rect 698232 79580 698300 79636
rect 698356 79580 698424 79636
rect 698480 79580 698548 79636
rect 698604 79580 698672 79636
rect 698728 79580 698796 79636
rect 698852 79580 698922 79636
rect 79078 79512 698922 79580
rect 79078 79456 79208 79512
rect 79264 79456 79332 79512
rect 79388 79456 79456 79512
rect 79512 79456 79580 79512
rect 79636 79456 79704 79512
rect 79760 79456 79828 79512
rect 79884 79456 79952 79512
rect 80008 79456 99294 79512
rect 99350 79456 99418 79512
rect 99474 79456 107330 79512
rect 107386 79456 107454 79512
rect 107510 79456 107578 79512
rect 107634 79456 107702 79512
rect 107758 79456 107826 79512
rect 107882 79456 107950 79512
rect 108006 79456 108074 79512
rect 108130 79456 108198 79512
rect 108254 79456 108322 79512
rect 108378 79456 108446 79512
rect 108502 79456 108570 79512
rect 108626 79456 108694 79512
rect 108750 79456 108818 79512
rect 108874 79456 108942 79512
rect 108998 79456 109066 79512
rect 109122 79456 109810 79512
rect 109866 79456 109934 79512
rect 109990 79456 110058 79512
rect 110114 79456 110182 79512
rect 110238 79456 110306 79512
rect 110362 79456 110430 79512
rect 110486 79456 110554 79512
rect 110610 79456 110678 79512
rect 110734 79456 110802 79512
rect 110858 79456 110926 79512
rect 110982 79456 111050 79512
rect 111106 79456 111174 79512
rect 111230 79456 111298 79512
rect 111354 79456 111422 79512
rect 111478 79456 111546 79512
rect 111602 79456 111670 79512
rect 111726 79456 112180 79512
rect 112236 79456 112304 79512
rect 112360 79456 112428 79512
rect 112484 79456 112552 79512
rect 112608 79456 112676 79512
rect 112732 79456 112800 79512
rect 112856 79456 112924 79512
rect 112980 79456 113048 79512
rect 113104 79456 113172 79512
rect 113228 79456 113296 79512
rect 113352 79456 113420 79512
rect 113476 79456 113544 79512
rect 113600 79456 113668 79512
rect 113724 79456 113792 79512
rect 113848 79456 113916 79512
rect 113972 79456 114040 79512
rect 114096 79456 114886 79512
rect 114942 79456 115010 79512
rect 115066 79456 115134 79512
rect 115190 79456 115258 79512
rect 115314 79456 115382 79512
rect 115438 79456 115506 79512
rect 115562 79456 115630 79512
rect 115686 79456 115754 79512
rect 115810 79456 115878 79512
rect 115934 79456 116002 79512
rect 116058 79456 116126 79512
rect 116182 79456 116250 79512
rect 116306 79456 116374 79512
rect 116430 79456 116498 79512
rect 116554 79456 116622 79512
rect 116678 79456 116746 79512
rect 116802 79456 117256 79512
rect 117312 79456 117380 79512
rect 117436 79456 117504 79512
rect 117560 79456 117628 79512
rect 117684 79456 117752 79512
rect 117808 79456 117876 79512
rect 117932 79456 118000 79512
rect 118056 79456 118124 79512
rect 118180 79456 118248 79512
rect 118304 79456 118372 79512
rect 118428 79456 118496 79512
rect 118552 79456 118620 79512
rect 118676 79456 118744 79512
rect 118800 79456 118868 79512
rect 118924 79456 118992 79512
rect 119048 79456 119116 79512
rect 119172 79456 119860 79512
rect 119916 79456 119984 79512
rect 120040 79456 120108 79512
rect 120164 79456 120232 79512
rect 120288 79456 120356 79512
rect 120412 79456 120480 79512
rect 120536 79456 120604 79512
rect 120660 79456 120728 79512
rect 120784 79456 120852 79512
rect 120908 79456 120976 79512
rect 121032 79456 121100 79512
rect 121156 79456 121224 79512
rect 121280 79456 121348 79512
rect 121404 79456 121472 79512
rect 121528 79456 121596 79512
rect 121652 79456 129294 79512
rect 129350 79456 129418 79512
rect 129474 79456 139294 79512
rect 139350 79456 139418 79512
rect 139474 79456 149294 79512
rect 149350 79456 149418 79512
rect 149474 79456 159294 79512
rect 159350 79456 159418 79512
rect 159474 79456 169294 79512
rect 169350 79456 169418 79512
rect 169474 79456 179294 79512
rect 179350 79456 179418 79512
rect 179474 79456 189294 79512
rect 189350 79456 189418 79512
rect 189474 79456 199294 79512
rect 199350 79456 199418 79512
rect 199474 79456 209294 79512
rect 209350 79456 209418 79512
rect 209474 79456 219294 79512
rect 219350 79456 219418 79512
rect 219474 79456 229294 79512
rect 229350 79456 229418 79512
rect 229474 79456 239294 79512
rect 239350 79456 239418 79512
rect 239474 79456 249294 79512
rect 249350 79456 249418 79512
rect 249474 79456 259294 79512
rect 259350 79456 259418 79512
rect 259474 79456 269294 79512
rect 269350 79456 269418 79512
rect 269474 79456 272330 79512
rect 272386 79456 272454 79512
rect 272510 79456 272578 79512
rect 272634 79456 272702 79512
rect 272758 79456 272826 79512
rect 272882 79456 272950 79512
rect 273006 79456 273074 79512
rect 273130 79456 273198 79512
rect 273254 79456 273322 79512
rect 273378 79456 273446 79512
rect 273502 79456 273570 79512
rect 273626 79456 273694 79512
rect 273750 79456 273818 79512
rect 273874 79456 273942 79512
rect 273998 79456 274066 79512
rect 274122 79456 274810 79512
rect 274866 79456 274934 79512
rect 274990 79456 275058 79512
rect 275114 79456 275182 79512
rect 275238 79456 275306 79512
rect 275362 79456 275430 79512
rect 275486 79456 275554 79512
rect 275610 79456 275678 79512
rect 275734 79456 275802 79512
rect 275858 79456 275926 79512
rect 275982 79456 276050 79512
rect 276106 79456 276174 79512
rect 276230 79456 276298 79512
rect 276354 79456 276422 79512
rect 276478 79456 276546 79512
rect 276602 79456 276670 79512
rect 276726 79456 277180 79512
rect 277236 79456 277304 79512
rect 277360 79456 277428 79512
rect 277484 79456 277552 79512
rect 277608 79456 277676 79512
rect 277732 79456 277800 79512
rect 277856 79456 277924 79512
rect 277980 79456 278048 79512
rect 278104 79456 278172 79512
rect 278228 79456 278296 79512
rect 278352 79456 278420 79512
rect 278476 79456 278544 79512
rect 278600 79456 278668 79512
rect 278724 79456 278792 79512
rect 278848 79456 278916 79512
rect 278972 79456 279040 79512
rect 279096 79456 279886 79512
rect 279942 79456 280010 79512
rect 280066 79456 280134 79512
rect 280190 79456 280258 79512
rect 280314 79456 280382 79512
rect 280438 79456 280506 79512
rect 280562 79456 280630 79512
rect 280686 79456 280754 79512
rect 280810 79456 280878 79512
rect 280934 79456 281002 79512
rect 281058 79456 281126 79512
rect 281182 79456 281250 79512
rect 281306 79456 281374 79512
rect 281430 79456 281498 79512
rect 281554 79456 281622 79512
rect 281678 79456 281746 79512
rect 281802 79456 282256 79512
rect 282312 79456 282380 79512
rect 282436 79456 282504 79512
rect 282560 79456 282628 79512
rect 282684 79456 282752 79512
rect 282808 79456 282876 79512
rect 282932 79456 283000 79512
rect 283056 79456 283124 79512
rect 283180 79456 283248 79512
rect 283304 79456 283372 79512
rect 283428 79456 283496 79512
rect 283552 79456 283620 79512
rect 283676 79456 283744 79512
rect 283800 79456 283868 79512
rect 283924 79456 283992 79512
rect 284048 79456 284116 79512
rect 284172 79456 284860 79512
rect 284916 79456 284984 79512
rect 285040 79456 285108 79512
rect 285164 79456 285232 79512
rect 285288 79456 285356 79512
rect 285412 79456 285480 79512
rect 285536 79456 285604 79512
rect 285660 79456 285728 79512
rect 285784 79456 285852 79512
rect 285908 79456 285976 79512
rect 286032 79456 286100 79512
rect 286156 79456 286224 79512
rect 286280 79456 286348 79512
rect 286404 79456 286472 79512
rect 286528 79456 286596 79512
rect 286652 79456 289294 79512
rect 289350 79456 289418 79512
rect 289474 79456 299294 79512
rect 299350 79456 299418 79512
rect 299474 79456 309294 79512
rect 309350 79456 309418 79512
rect 309474 79456 319294 79512
rect 319350 79456 319418 79512
rect 319474 79456 329294 79512
rect 329350 79456 329418 79512
rect 329474 79456 339294 79512
rect 339350 79456 339418 79512
rect 339474 79456 349294 79512
rect 349350 79456 349418 79512
rect 349474 79456 359294 79512
rect 359350 79456 359418 79512
rect 359474 79456 369294 79512
rect 369350 79456 369418 79512
rect 369474 79456 379294 79512
rect 379350 79456 379418 79512
rect 379474 79456 389294 79512
rect 389350 79456 389418 79512
rect 389474 79456 399294 79512
rect 399350 79456 399418 79512
rect 399474 79456 409294 79512
rect 409350 79456 409418 79512
rect 409474 79456 419294 79512
rect 419350 79456 419418 79512
rect 419474 79456 429294 79512
rect 429350 79456 429418 79512
rect 429474 79456 439294 79512
rect 439350 79456 439418 79512
rect 439474 79456 449294 79512
rect 449350 79456 449418 79512
rect 449474 79456 459294 79512
rect 459350 79456 459418 79512
rect 459474 79456 469294 79512
rect 469350 79456 469418 79512
rect 469474 79456 479294 79512
rect 479350 79456 479418 79512
rect 479474 79456 489294 79512
rect 489350 79456 489418 79512
rect 489474 79456 499294 79512
rect 499350 79456 499418 79512
rect 499474 79456 509294 79512
rect 509350 79456 509418 79512
rect 509474 79456 519294 79512
rect 519350 79456 519418 79512
rect 519474 79456 529294 79512
rect 529350 79456 529418 79512
rect 529474 79456 539294 79512
rect 539350 79456 539418 79512
rect 539474 79456 549294 79512
rect 549350 79456 549418 79512
rect 549474 79456 590970 79512
rect 591026 79456 591094 79512
rect 591150 79456 591218 79512
rect 591274 79456 591342 79512
rect 591398 79456 591466 79512
rect 591522 79456 591590 79512
rect 591646 79456 591714 79512
rect 591770 79456 602330 79512
rect 602386 79456 602454 79512
rect 602510 79456 602578 79512
rect 602634 79456 602702 79512
rect 602758 79456 602826 79512
rect 602882 79456 602950 79512
rect 603006 79456 603074 79512
rect 603130 79456 603198 79512
rect 603254 79456 603322 79512
rect 603378 79456 603446 79512
rect 603502 79456 603570 79512
rect 603626 79456 603694 79512
rect 603750 79456 603818 79512
rect 603874 79456 603942 79512
rect 603998 79456 604066 79512
rect 604122 79456 604810 79512
rect 604866 79456 604934 79512
rect 604990 79456 605058 79512
rect 605114 79456 605182 79512
rect 605238 79456 605306 79512
rect 605362 79456 605430 79512
rect 605486 79456 605554 79512
rect 605610 79456 605678 79512
rect 605734 79456 605802 79512
rect 605858 79456 605926 79512
rect 605982 79456 606050 79512
rect 606106 79456 606174 79512
rect 606230 79456 606298 79512
rect 606354 79456 606422 79512
rect 606478 79456 606546 79512
rect 606602 79456 606670 79512
rect 606726 79456 607180 79512
rect 607236 79456 607304 79512
rect 607360 79456 607428 79512
rect 607484 79456 607552 79512
rect 607608 79456 607676 79512
rect 607732 79456 607800 79512
rect 607856 79456 607924 79512
rect 607980 79456 608048 79512
rect 608104 79456 608172 79512
rect 608228 79456 608296 79512
rect 608352 79456 608420 79512
rect 608476 79456 608544 79512
rect 608600 79456 608668 79512
rect 608724 79456 608792 79512
rect 608848 79456 608916 79512
rect 608972 79456 609040 79512
rect 609096 79456 609886 79512
rect 609942 79456 610010 79512
rect 610066 79456 610134 79512
rect 610190 79456 610258 79512
rect 610314 79456 610382 79512
rect 610438 79456 610506 79512
rect 610562 79456 610630 79512
rect 610686 79456 610754 79512
rect 610810 79456 610878 79512
rect 610934 79456 611002 79512
rect 611058 79456 611126 79512
rect 611182 79456 611250 79512
rect 611306 79456 611374 79512
rect 611430 79456 611498 79512
rect 611554 79456 611622 79512
rect 611678 79456 611746 79512
rect 611802 79456 612256 79512
rect 612312 79456 612380 79512
rect 612436 79456 612504 79512
rect 612560 79456 612628 79512
rect 612684 79456 612752 79512
rect 612808 79456 612876 79512
rect 612932 79456 613000 79512
rect 613056 79456 613124 79512
rect 613180 79456 613248 79512
rect 613304 79456 613372 79512
rect 613428 79456 613496 79512
rect 613552 79456 613620 79512
rect 613676 79456 613744 79512
rect 613800 79456 613868 79512
rect 613924 79456 613992 79512
rect 614048 79456 614116 79512
rect 614172 79456 614860 79512
rect 614916 79456 614984 79512
rect 615040 79456 615108 79512
rect 615164 79456 615232 79512
rect 615288 79456 615356 79512
rect 615412 79456 615480 79512
rect 615536 79456 615604 79512
rect 615660 79456 615728 79512
rect 615784 79456 615852 79512
rect 615908 79456 615976 79512
rect 616032 79456 616100 79512
rect 616156 79456 616224 79512
rect 616280 79456 616348 79512
rect 616404 79456 616472 79512
rect 616528 79456 616596 79512
rect 616652 79456 628697 79512
rect 628753 79456 628821 79512
rect 628877 79456 636637 79512
rect 636693 79456 636761 79512
rect 636817 79456 644577 79512
rect 644633 79456 644701 79512
rect 644757 79456 670090 79512
rect 670146 79456 670214 79512
rect 670270 79456 670338 79512
rect 670394 79456 670462 79512
rect 670518 79456 670586 79512
rect 670642 79456 670710 79512
rect 670766 79456 698052 79512
rect 698108 79456 698176 79512
rect 698232 79456 698300 79512
rect 698356 79456 698424 79512
rect 698480 79456 698548 79512
rect 698604 79456 698672 79512
rect 698728 79456 698796 79512
rect 698852 79456 698922 79512
rect 79078 79388 698922 79456
rect 79078 79332 79208 79388
rect 79264 79332 79332 79388
rect 79388 79332 79456 79388
rect 79512 79332 79580 79388
rect 79636 79332 79704 79388
rect 79760 79332 79828 79388
rect 79884 79332 79952 79388
rect 80008 79332 99294 79388
rect 99350 79332 99418 79388
rect 99474 79332 107330 79388
rect 107386 79332 107454 79388
rect 107510 79332 107578 79388
rect 107634 79332 107702 79388
rect 107758 79332 107826 79388
rect 107882 79332 107950 79388
rect 108006 79332 108074 79388
rect 108130 79332 108198 79388
rect 108254 79332 108322 79388
rect 108378 79332 108446 79388
rect 108502 79332 108570 79388
rect 108626 79332 108694 79388
rect 108750 79332 108818 79388
rect 108874 79332 108942 79388
rect 108998 79332 109066 79388
rect 109122 79332 109810 79388
rect 109866 79332 109934 79388
rect 109990 79332 110058 79388
rect 110114 79332 110182 79388
rect 110238 79332 110306 79388
rect 110362 79332 110430 79388
rect 110486 79332 110554 79388
rect 110610 79332 110678 79388
rect 110734 79332 110802 79388
rect 110858 79332 110926 79388
rect 110982 79332 111050 79388
rect 111106 79332 111174 79388
rect 111230 79332 111298 79388
rect 111354 79332 111422 79388
rect 111478 79332 111546 79388
rect 111602 79332 111670 79388
rect 111726 79332 112180 79388
rect 112236 79332 112304 79388
rect 112360 79332 112428 79388
rect 112484 79332 112552 79388
rect 112608 79332 112676 79388
rect 112732 79332 112800 79388
rect 112856 79332 112924 79388
rect 112980 79332 113048 79388
rect 113104 79332 113172 79388
rect 113228 79332 113296 79388
rect 113352 79332 113420 79388
rect 113476 79332 113544 79388
rect 113600 79332 113668 79388
rect 113724 79332 113792 79388
rect 113848 79332 113916 79388
rect 113972 79332 114040 79388
rect 114096 79332 114886 79388
rect 114942 79332 115010 79388
rect 115066 79332 115134 79388
rect 115190 79332 115258 79388
rect 115314 79332 115382 79388
rect 115438 79332 115506 79388
rect 115562 79332 115630 79388
rect 115686 79332 115754 79388
rect 115810 79332 115878 79388
rect 115934 79332 116002 79388
rect 116058 79332 116126 79388
rect 116182 79332 116250 79388
rect 116306 79332 116374 79388
rect 116430 79332 116498 79388
rect 116554 79332 116622 79388
rect 116678 79332 116746 79388
rect 116802 79332 117256 79388
rect 117312 79332 117380 79388
rect 117436 79332 117504 79388
rect 117560 79332 117628 79388
rect 117684 79332 117752 79388
rect 117808 79332 117876 79388
rect 117932 79332 118000 79388
rect 118056 79332 118124 79388
rect 118180 79332 118248 79388
rect 118304 79332 118372 79388
rect 118428 79332 118496 79388
rect 118552 79332 118620 79388
rect 118676 79332 118744 79388
rect 118800 79332 118868 79388
rect 118924 79332 118992 79388
rect 119048 79332 119116 79388
rect 119172 79332 119860 79388
rect 119916 79332 119984 79388
rect 120040 79332 120108 79388
rect 120164 79332 120232 79388
rect 120288 79332 120356 79388
rect 120412 79332 120480 79388
rect 120536 79332 120604 79388
rect 120660 79332 120728 79388
rect 120784 79332 120852 79388
rect 120908 79332 120976 79388
rect 121032 79332 121100 79388
rect 121156 79332 121224 79388
rect 121280 79332 121348 79388
rect 121404 79332 121472 79388
rect 121528 79332 121596 79388
rect 121652 79332 129294 79388
rect 129350 79332 129418 79388
rect 129474 79332 139294 79388
rect 139350 79332 139418 79388
rect 139474 79332 149294 79388
rect 149350 79332 149418 79388
rect 149474 79332 159294 79388
rect 159350 79332 159418 79388
rect 159474 79332 169294 79388
rect 169350 79332 169418 79388
rect 169474 79332 179294 79388
rect 179350 79332 179418 79388
rect 179474 79332 189294 79388
rect 189350 79332 189418 79388
rect 189474 79332 199294 79388
rect 199350 79332 199418 79388
rect 199474 79332 209294 79388
rect 209350 79332 209418 79388
rect 209474 79332 219294 79388
rect 219350 79332 219418 79388
rect 219474 79332 229294 79388
rect 229350 79332 229418 79388
rect 229474 79332 239294 79388
rect 239350 79332 239418 79388
rect 239474 79332 249294 79388
rect 249350 79332 249418 79388
rect 249474 79332 259294 79388
rect 259350 79332 259418 79388
rect 259474 79332 269294 79388
rect 269350 79332 269418 79388
rect 269474 79332 272330 79388
rect 272386 79332 272454 79388
rect 272510 79332 272578 79388
rect 272634 79332 272702 79388
rect 272758 79332 272826 79388
rect 272882 79332 272950 79388
rect 273006 79332 273074 79388
rect 273130 79332 273198 79388
rect 273254 79332 273322 79388
rect 273378 79332 273446 79388
rect 273502 79332 273570 79388
rect 273626 79332 273694 79388
rect 273750 79332 273818 79388
rect 273874 79332 273942 79388
rect 273998 79332 274066 79388
rect 274122 79332 274810 79388
rect 274866 79332 274934 79388
rect 274990 79332 275058 79388
rect 275114 79332 275182 79388
rect 275238 79332 275306 79388
rect 275362 79332 275430 79388
rect 275486 79332 275554 79388
rect 275610 79332 275678 79388
rect 275734 79332 275802 79388
rect 275858 79332 275926 79388
rect 275982 79332 276050 79388
rect 276106 79332 276174 79388
rect 276230 79332 276298 79388
rect 276354 79332 276422 79388
rect 276478 79332 276546 79388
rect 276602 79332 276670 79388
rect 276726 79332 277180 79388
rect 277236 79332 277304 79388
rect 277360 79332 277428 79388
rect 277484 79332 277552 79388
rect 277608 79332 277676 79388
rect 277732 79332 277800 79388
rect 277856 79332 277924 79388
rect 277980 79332 278048 79388
rect 278104 79332 278172 79388
rect 278228 79332 278296 79388
rect 278352 79332 278420 79388
rect 278476 79332 278544 79388
rect 278600 79332 278668 79388
rect 278724 79332 278792 79388
rect 278848 79332 278916 79388
rect 278972 79332 279040 79388
rect 279096 79332 279886 79388
rect 279942 79332 280010 79388
rect 280066 79332 280134 79388
rect 280190 79332 280258 79388
rect 280314 79332 280382 79388
rect 280438 79332 280506 79388
rect 280562 79332 280630 79388
rect 280686 79332 280754 79388
rect 280810 79332 280878 79388
rect 280934 79332 281002 79388
rect 281058 79332 281126 79388
rect 281182 79332 281250 79388
rect 281306 79332 281374 79388
rect 281430 79332 281498 79388
rect 281554 79332 281622 79388
rect 281678 79332 281746 79388
rect 281802 79332 282256 79388
rect 282312 79332 282380 79388
rect 282436 79332 282504 79388
rect 282560 79332 282628 79388
rect 282684 79332 282752 79388
rect 282808 79332 282876 79388
rect 282932 79332 283000 79388
rect 283056 79332 283124 79388
rect 283180 79332 283248 79388
rect 283304 79332 283372 79388
rect 283428 79332 283496 79388
rect 283552 79332 283620 79388
rect 283676 79332 283744 79388
rect 283800 79332 283868 79388
rect 283924 79332 283992 79388
rect 284048 79332 284116 79388
rect 284172 79332 284860 79388
rect 284916 79332 284984 79388
rect 285040 79332 285108 79388
rect 285164 79332 285232 79388
rect 285288 79332 285356 79388
rect 285412 79332 285480 79388
rect 285536 79332 285604 79388
rect 285660 79332 285728 79388
rect 285784 79332 285852 79388
rect 285908 79332 285976 79388
rect 286032 79332 286100 79388
rect 286156 79332 286224 79388
rect 286280 79332 286348 79388
rect 286404 79332 286472 79388
rect 286528 79332 286596 79388
rect 286652 79332 289294 79388
rect 289350 79332 289418 79388
rect 289474 79332 299294 79388
rect 299350 79332 299418 79388
rect 299474 79332 309294 79388
rect 309350 79332 309418 79388
rect 309474 79332 319294 79388
rect 319350 79332 319418 79388
rect 319474 79332 329294 79388
rect 329350 79332 329418 79388
rect 329474 79332 339294 79388
rect 339350 79332 339418 79388
rect 339474 79332 349294 79388
rect 349350 79332 349418 79388
rect 349474 79332 359294 79388
rect 359350 79332 359418 79388
rect 359474 79332 369294 79388
rect 369350 79332 369418 79388
rect 369474 79332 379294 79388
rect 379350 79332 379418 79388
rect 379474 79332 389294 79388
rect 389350 79332 389418 79388
rect 389474 79332 399294 79388
rect 399350 79332 399418 79388
rect 399474 79332 409294 79388
rect 409350 79332 409418 79388
rect 409474 79332 419294 79388
rect 419350 79332 419418 79388
rect 419474 79332 429294 79388
rect 429350 79332 429418 79388
rect 429474 79332 439294 79388
rect 439350 79332 439418 79388
rect 439474 79332 449294 79388
rect 449350 79332 449418 79388
rect 449474 79332 459294 79388
rect 459350 79332 459418 79388
rect 459474 79332 469294 79388
rect 469350 79332 469418 79388
rect 469474 79332 479294 79388
rect 479350 79332 479418 79388
rect 479474 79332 489294 79388
rect 489350 79332 489418 79388
rect 489474 79332 499294 79388
rect 499350 79332 499418 79388
rect 499474 79332 509294 79388
rect 509350 79332 509418 79388
rect 509474 79332 519294 79388
rect 519350 79332 519418 79388
rect 519474 79332 529294 79388
rect 529350 79332 529418 79388
rect 529474 79332 539294 79388
rect 539350 79332 539418 79388
rect 539474 79332 549294 79388
rect 549350 79332 549418 79388
rect 549474 79332 590970 79388
rect 591026 79332 591094 79388
rect 591150 79332 591218 79388
rect 591274 79332 591342 79388
rect 591398 79332 591466 79388
rect 591522 79332 591590 79388
rect 591646 79332 591714 79388
rect 591770 79332 602330 79388
rect 602386 79332 602454 79388
rect 602510 79332 602578 79388
rect 602634 79332 602702 79388
rect 602758 79332 602826 79388
rect 602882 79332 602950 79388
rect 603006 79332 603074 79388
rect 603130 79332 603198 79388
rect 603254 79332 603322 79388
rect 603378 79332 603446 79388
rect 603502 79332 603570 79388
rect 603626 79332 603694 79388
rect 603750 79332 603818 79388
rect 603874 79332 603942 79388
rect 603998 79332 604066 79388
rect 604122 79332 604810 79388
rect 604866 79332 604934 79388
rect 604990 79332 605058 79388
rect 605114 79332 605182 79388
rect 605238 79332 605306 79388
rect 605362 79332 605430 79388
rect 605486 79332 605554 79388
rect 605610 79332 605678 79388
rect 605734 79332 605802 79388
rect 605858 79332 605926 79388
rect 605982 79332 606050 79388
rect 606106 79332 606174 79388
rect 606230 79332 606298 79388
rect 606354 79332 606422 79388
rect 606478 79332 606546 79388
rect 606602 79332 606670 79388
rect 606726 79332 607180 79388
rect 607236 79332 607304 79388
rect 607360 79332 607428 79388
rect 607484 79332 607552 79388
rect 607608 79332 607676 79388
rect 607732 79332 607800 79388
rect 607856 79332 607924 79388
rect 607980 79332 608048 79388
rect 608104 79332 608172 79388
rect 608228 79332 608296 79388
rect 608352 79332 608420 79388
rect 608476 79332 608544 79388
rect 608600 79332 608668 79388
rect 608724 79332 608792 79388
rect 608848 79332 608916 79388
rect 608972 79332 609040 79388
rect 609096 79332 609886 79388
rect 609942 79332 610010 79388
rect 610066 79332 610134 79388
rect 610190 79332 610258 79388
rect 610314 79332 610382 79388
rect 610438 79332 610506 79388
rect 610562 79332 610630 79388
rect 610686 79332 610754 79388
rect 610810 79332 610878 79388
rect 610934 79332 611002 79388
rect 611058 79332 611126 79388
rect 611182 79332 611250 79388
rect 611306 79332 611374 79388
rect 611430 79332 611498 79388
rect 611554 79332 611622 79388
rect 611678 79332 611746 79388
rect 611802 79332 612256 79388
rect 612312 79332 612380 79388
rect 612436 79332 612504 79388
rect 612560 79332 612628 79388
rect 612684 79332 612752 79388
rect 612808 79332 612876 79388
rect 612932 79332 613000 79388
rect 613056 79332 613124 79388
rect 613180 79332 613248 79388
rect 613304 79332 613372 79388
rect 613428 79332 613496 79388
rect 613552 79332 613620 79388
rect 613676 79332 613744 79388
rect 613800 79332 613868 79388
rect 613924 79332 613992 79388
rect 614048 79332 614116 79388
rect 614172 79332 614860 79388
rect 614916 79332 614984 79388
rect 615040 79332 615108 79388
rect 615164 79332 615232 79388
rect 615288 79332 615356 79388
rect 615412 79332 615480 79388
rect 615536 79332 615604 79388
rect 615660 79332 615728 79388
rect 615784 79332 615852 79388
rect 615908 79332 615976 79388
rect 616032 79332 616100 79388
rect 616156 79332 616224 79388
rect 616280 79332 616348 79388
rect 616404 79332 616472 79388
rect 616528 79332 616596 79388
rect 616652 79332 628697 79388
rect 628753 79332 628821 79388
rect 628877 79332 636637 79388
rect 636693 79332 636761 79388
rect 636817 79332 644577 79388
rect 644633 79332 644701 79388
rect 644757 79332 670090 79388
rect 670146 79332 670214 79388
rect 670270 79332 670338 79388
rect 670394 79332 670462 79388
rect 670518 79332 670586 79388
rect 670642 79332 670710 79388
rect 670766 79332 698052 79388
rect 698108 79332 698176 79388
rect 698232 79332 698300 79388
rect 698356 79332 698424 79388
rect 698480 79332 698548 79388
rect 698604 79332 698672 79388
rect 698728 79332 698796 79388
rect 698852 79332 698922 79388
rect 79078 79264 698922 79332
rect 79078 79208 79208 79264
rect 79264 79208 79332 79264
rect 79388 79208 79456 79264
rect 79512 79208 79580 79264
rect 79636 79208 79704 79264
rect 79760 79208 79828 79264
rect 79884 79208 79952 79264
rect 80008 79208 99294 79264
rect 99350 79208 99418 79264
rect 99474 79208 107330 79264
rect 107386 79208 107454 79264
rect 107510 79208 107578 79264
rect 107634 79208 107702 79264
rect 107758 79208 107826 79264
rect 107882 79208 107950 79264
rect 108006 79208 108074 79264
rect 108130 79208 108198 79264
rect 108254 79208 108322 79264
rect 108378 79208 108446 79264
rect 108502 79208 108570 79264
rect 108626 79208 108694 79264
rect 108750 79208 108818 79264
rect 108874 79208 108942 79264
rect 108998 79208 109066 79264
rect 109122 79208 109810 79264
rect 109866 79208 109934 79264
rect 109990 79208 110058 79264
rect 110114 79208 110182 79264
rect 110238 79208 110306 79264
rect 110362 79208 110430 79264
rect 110486 79208 110554 79264
rect 110610 79208 110678 79264
rect 110734 79208 110802 79264
rect 110858 79208 110926 79264
rect 110982 79208 111050 79264
rect 111106 79208 111174 79264
rect 111230 79208 111298 79264
rect 111354 79208 111422 79264
rect 111478 79208 111546 79264
rect 111602 79208 111670 79264
rect 111726 79208 112180 79264
rect 112236 79208 112304 79264
rect 112360 79208 112428 79264
rect 112484 79208 112552 79264
rect 112608 79208 112676 79264
rect 112732 79208 112800 79264
rect 112856 79208 112924 79264
rect 112980 79208 113048 79264
rect 113104 79208 113172 79264
rect 113228 79208 113296 79264
rect 113352 79208 113420 79264
rect 113476 79208 113544 79264
rect 113600 79208 113668 79264
rect 113724 79208 113792 79264
rect 113848 79208 113916 79264
rect 113972 79208 114040 79264
rect 114096 79208 114886 79264
rect 114942 79208 115010 79264
rect 115066 79208 115134 79264
rect 115190 79208 115258 79264
rect 115314 79208 115382 79264
rect 115438 79208 115506 79264
rect 115562 79208 115630 79264
rect 115686 79208 115754 79264
rect 115810 79208 115878 79264
rect 115934 79208 116002 79264
rect 116058 79208 116126 79264
rect 116182 79208 116250 79264
rect 116306 79208 116374 79264
rect 116430 79208 116498 79264
rect 116554 79208 116622 79264
rect 116678 79208 116746 79264
rect 116802 79208 117256 79264
rect 117312 79208 117380 79264
rect 117436 79208 117504 79264
rect 117560 79208 117628 79264
rect 117684 79208 117752 79264
rect 117808 79208 117876 79264
rect 117932 79208 118000 79264
rect 118056 79208 118124 79264
rect 118180 79208 118248 79264
rect 118304 79208 118372 79264
rect 118428 79208 118496 79264
rect 118552 79208 118620 79264
rect 118676 79208 118744 79264
rect 118800 79208 118868 79264
rect 118924 79208 118992 79264
rect 119048 79208 119116 79264
rect 119172 79208 119860 79264
rect 119916 79208 119984 79264
rect 120040 79208 120108 79264
rect 120164 79208 120232 79264
rect 120288 79208 120356 79264
rect 120412 79208 120480 79264
rect 120536 79208 120604 79264
rect 120660 79208 120728 79264
rect 120784 79208 120852 79264
rect 120908 79208 120976 79264
rect 121032 79208 121100 79264
rect 121156 79208 121224 79264
rect 121280 79208 121348 79264
rect 121404 79208 121472 79264
rect 121528 79208 121596 79264
rect 121652 79208 129294 79264
rect 129350 79208 129418 79264
rect 129474 79208 139294 79264
rect 139350 79208 139418 79264
rect 139474 79208 149294 79264
rect 149350 79208 149418 79264
rect 149474 79208 159294 79264
rect 159350 79208 159418 79264
rect 159474 79208 169294 79264
rect 169350 79208 169418 79264
rect 169474 79208 179294 79264
rect 179350 79208 179418 79264
rect 179474 79208 189294 79264
rect 189350 79208 189418 79264
rect 189474 79208 199294 79264
rect 199350 79208 199418 79264
rect 199474 79208 209294 79264
rect 209350 79208 209418 79264
rect 209474 79208 219294 79264
rect 219350 79208 219418 79264
rect 219474 79208 229294 79264
rect 229350 79208 229418 79264
rect 229474 79208 239294 79264
rect 239350 79208 239418 79264
rect 239474 79208 249294 79264
rect 249350 79208 249418 79264
rect 249474 79208 259294 79264
rect 259350 79208 259418 79264
rect 259474 79208 269294 79264
rect 269350 79208 269418 79264
rect 269474 79208 272330 79264
rect 272386 79208 272454 79264
rect 272510 79208 272578 79264
rect 272634 79208 272702 79264
rect 272758 79208 272826 79264
rect 272882 79208 272950 79264
rect 273006 79208 273074 79264
rect 273130 79208 273198 79264
rect 273254 79208 273322 79264
rect 273378 79208 273446 79264
rect 273502 79208 273570 79264
rect 273626 79208 273694 79264
rect 273750 79208 273818 79264
rect 273874 79208 273942 79264
rect 273998 79208 274066 79264
rect 274122 79208 274810 79264
rect 274866 79208 274934 79264
rect 274990 79208 275058 79264
rect 275114 79208 275182 79264
rect 275238 79208 275306 79264
rect 275362 79208 275430 79264
rect 275486 79208 275554 79264
rect 275610 79208 275678 79264
rect 275734 79208 275802 79264
rect 275858 79208 275926 79264
rect 275982 79208 276050 79264
rect 276106 79208 276174 79264
rect 276230 79208 276298 79264
rect 276354 79208 276422 79264
rect 276478 79208 276546 79264
rect 276602 79208 276670 79264
rect 276726 79208 277180 79264
rect 277236 79208 277304 79264
rect 277360 79208 277428 79264
rect 277484 79208 277552 79264
rect 277608 79208 277676 79264
rect 277732 79208 277800 79264
rect 277856 79208 277924 79264
rect 277980 79208 278048 79264
rect 278104 79208 278172 79264
rect 278228 79208 278296 79264
rect 278352 79208 278420 79264
rect 278476 79208 278544 79264
rect 278600 79208 278668 79264
rect 278724 79208 278792 79264
rect 278848 79208 278916 79264
rect 278972 79208 279040 79264
rect 279096 79208 279886 79264
rect 279942 79208 280010 79264
rect 280066 79208 280134 79264
rect 280190 79208 280258 79264
rect 280314 79208 280382 79264
rect 280438 79208 280506 79264
rect 280562 79208 280630 79264
rect 280686 79208 280754 79264
rect 280810 79208 280878 79264
rect 280934 79208 281002 79264
rect 281058 79208 281126 79264
rect 281182 79208 281250 79264
rect 281306 79208 281374 79264
rect 281430 79208 281498 79264
rect 281554 79208 281622 79264
rect 281678 79208 281746 79264
rect 281802 79208 282256 79264
rect 282312 79208 282380 79264
rect 282436 79208 282504 79264
rect 282560 79208 282628 79264
rect 282684 79208 282752 79264
rect 282808 79208 282876 79264
rect 282932 79208 283000 79264
rect 283056 79208 283124 79264
rect 283180 79208 283248 79264
rect 283304 79208 283372 79264
rect 283428 79208 283496 79264
rect 283552 79208 283620 79264
rect 283676 79208 283744 79264
rect 283800 79208 283868 79264
rect 283924 79208 283992 79264
rect 284048 79208 284116 79264
rect 284172 79208 284860 79264
rect 284916 79208 284984 79264
rect 285040 79208 285108 79264
rect 285164 79208 285232 79264
rect 285288 79208 285356 79264
rect 285412 79208 285480 79264
rect 285536 79208 285604 79264
rect 285660 79208 285728 79264
rect 285784 79208 285852 79264
rect 285908 79208 285976 79264
rect 286032 79208 286100 79264
rect 286156 79208 286224 79264
rect 286280 79208 286348 79264
rect 286404 79208 286472 79264
rect 286528 79208 286596 79264
rect 286652 79208 289294 79264
rect 289350 79208 289418 79264
rect 289474 79208 299294 79264
rect 299350 79208 299418 79264
rect 299474 79208 309294 79264
rect 309350 79208 309418 79264
rect 309474 79208 319294 79264
rect 319350 79208 319418 79264
rect 319474 79208 329294 79264
rect 329350 79208 329418 79264
rect 329474 79208 339294 79264
rect 339350 79208 339418 79264
rect 339474 79208 349294 79264
rect 349350 79208 349418 79264
rect 349474 79208 359294 79264
rect 359350 79208 359418 79264
rect 359474 79208 369294 79264
rect 369350 79208 369418 79264
rect 369474 79208 379294 79264
rect 379350 79208 379418 79264
rect 379474 79208 389294 79264
rect 389350 79208 389418 79264
rect 389474 79208 399294 79264
rect 399350 79208 399418 79264
rect 399474 79208 409294 79264
rect 409350 79208 409418 79264
rect 409474 79208 419294 79264
rect 419350 79208 419418 79264
rect 419474 79208 429294 79264
rect 429350 79208 429418 79264
rect 429474 79208 439294 79264
rect 439350 79208 439418 79264
rect 439474 79208 449294 79264
rect 449350 79208 449418 79264
rect 449474 79208 459294 79264
rect 459350 79208 459418 79264
rect 459474 79208 469294 79264
rect 469350 79208 469418 79264
rect 469474 79208 479294 79264
rect 479350 79208 479418 79264
rect 479474 79208 489294 79264
rect 489350 79208 489418 79264
rect 489474 79208 499294 79264
rect 499350 79208 499418 79264
rect 499474 79208 509294 79264
rect 509350 79208 509418 79264
rect 509474 79208 519294 79264
rect 519350 79208 519418 79264
rect 519474 79208 529294 79264
rect 529350 79208 529418 79264
rect 529474 79208 539294 79264
rect 539350 79208 539418 79264
rect 539474 79208 549294 79264
rect 549350 79208 549418 79264
rect 549474 79208 590970 79264
rect 591026 79208 591094 79264
rect 591150 79208 591218 79264
rect 591274 79208 591342 79264
rect 591398 79208 591466 79264
rect 591522 79208 591590 79264
rect 591646 79208 591714 79264
rect 591770 79208 602330 79264
rect 602386 79208 602454 79264
rect 602510 79208 602578 79264
rect 602634 79208 602702 79264
rect 602758 79208 602826 79264
rect 602882 79208 602950 79264
rect 603006 79208 603074 79264
rect 603130 79208 603198 79264
rect 603254 79208 603322 79264
rect 603378 79208 603446 79264
rect 603502 79208 603570 79264
rect 603626 79208 603694 79264
rect 603750 79208 603818 79264
rect 603874 79208 603942 79264
rect 603998 79208 604066 79264
rect 604122 79208 604810 79264
rect 604866 79208 604934 79264
rect 604990 79208 605058 79264
rect 605114 79208 605182 79264
rect 605238 79208 605306 79264
rect 605362 79208 605430 79264
rect 605486 79208 605554 79264
rect 605610 79208 605678 79264
rect 605734 79208 605802 79264
rect 605858 79208 605926 79264
rect 605982 79208 606050 79264
rect 606106 79208 606174 79264
rect 606230 79208 606298 79264
rect 606354 79208 606422 79264
rect 606478 79208 606546 79264
rect 606602 79208 606670 79264
rect 606726 79208 607180 79264
rect 607236 79208 607304 79264
rect 607360 79208 607428 79264
rect 607484 79208 607552 79264
rect 607608 79208 607676 79264
rect 607732 79208 607800 79264
rect 607856 79208 607924 79264
rect 607980 79208 608048 79264
rect 608104 79208 608172 79264
rect 608228 79208 608296 79264
rect 608352 79208 608420 79264
rect 608476 79208 608544 79264
rect 608600 79208 608668 79264
rect 608724 79208 608792 79264
rect 608848 79208 608916 79264
rect 608972 79208 609040 79264
rect 609096 79208 609886 79264
rect 609942 79208 610010 79264
rect 610066 79208 610134 79264
rect 610190 79208 610258 79264
rect 610314 79208 610382 79264
rect 610438 79208 610506 79264
rect 610562 79208 610630 79264
rect 610686 79208 610754 79264
rect 610810 79208 610878 79264
rect 610934 79208 611002 79264
rect 611058 79208 611126 79264
rect 611182 79208 611250 79264
rect 611306 79208 611374 79264
rect 611430 79208 611498 79264
rect 611554 79208 611622 79264
rect 611678 79208 611746 79264
rect 611802 79208 612256 79264
rect 612312 79208 612380 79264
rect 612436 79208 612504 79264
rect 612560 79208 612628 79264
rect 612684 79208 612752 79264
rect 612808 79208 612876 79264
rect 612932 79208 613000 79264
rect 613056 79208 613124 79264
rect 613180 79208 613248 79264
rect 613304 79208 613372 79264
rect 613428 79208 613496 79264
rect 613552 79208 613620 79264
rect 613676 79208 613744 79264
rect 613800 79208 613868 79264
rect 613924 79208 613992 79264
rect 614048 79208 614116 79264
rect 614172 79208 614860 79264
rect 614916 79208 614984 79264
rect 615040 79208 615108 79264
rect 615164 79208 615232 79264
rect 615288 79208 615356 79264
rect 615412 79208 615480 79264
rect 615536 79208 615604 79264
rect 615660 79208 615728 79264
rect 615784 79208 615852 79264
rect 615908 79208 615976 79264
rect 616032 79208 616100 79264
rect 616156 79208 616224 79264
rect 616280 79208 616348 79264
rect 616404 79208 616472 79264
rect 616528 79208 616596 79264
rect 616652 79208 628697 79264
rect 628753 79208 628821 79264
rect 628877 79208 636637 79264
rect 636693 79208 636761 79264
rect 636817 79208 644577 79264
rect 644633 79208 644701 79264
rect 644757 79208 670090 79264
rect 670146 79208 670214 79264
rect 670270 79208 670338 79264
rect 670394 79208 670462 79264
rect 670518 79208 670586 79264
rect 670642 79208 670710 79264
rect 670766 79208 698052 79264
rect 698108 79208 698176 79264
rect 698232 79208 698300 79264
rect 698356 79208 698424 79264
rect 698480 79208 698548 79264
rect 698604 79208 698672 79264
rect 698728 79208 698796 79264
rect 698852 79208 698922 79264
rect 79078 79078 698922 79208
rect 77678 78608 700322 78678
rect 77678 78552 77808 78608
rect 77864 78552 77932 78608
rect 77988 78552 78056 78608
rect 78112 78552 78180 78608
rect 78236 78552 78304 78608
rect 78360 78552 78428 78608
rect 78484 78552 78552 78608
rect 78608 78552 94294 78608
rect 94350 78552 94418 78608
rect 94474 78552 104294 78608
rect 104350 78552 104418 78608
rect 104474 78552 124294 78608
rect 124350 78552 124418 78608
rect 124474 78552 134294 78608
rect 134350 78552 134418 78608
rect 134474 78552 144294 78608
rect 144350 78552 144418 78608
rect 144474 78552 154294 78608
rect 154350 78552 154418 78608
rect 154474 78552 164294 78608
rect 164350 78552 164418 78608
rect 164474 78552 174294 78608
rect 174350 78552 174418 78608
rect 174474 78552 184294 78608
rect 184350 78552 184418 78608
rect 184474 78552 194294 78608
rect 194350 78552 194418 78608
rect 194474 78552 204294 78608
rect 204350 78552 204418 78608
rect 204474 78552 214294 78608
rect 214350 78552 214418 78608
rect 214474 78552 224294 78608
rect 224350 78552 224418 78608
rect 224474 78552 234294 78608
rect 234350 78552 234418 78608
rect 234474 78552 244294 78608
rect 244350 78552 244418 78608
rect 244474 78552 254294 78608
rect 254350 78552 254418 78608
rect 254474 78552 264294 78608
rect 264350 78552 264418 78608
rect 264474 78552 294294 78608
rect 294350 78552 294418 78608
rect 294474 78552 304294 78608
rect 304350 78552 304418 78608
rect 304474 78552 314294 78608
rect 314350 78552 314418 78608
rect 314474 78552 324294 78608
rect 324350 78552 324418 78608
rect 324474 78552 334294 78608
rect 334350 78552 334418 78608
rect 334474 78552 344294 78608
rect 344350 78552 344418 78608
rect 344474 78552 354294 78608
rect 354350 78552 354418 78608
rect 354474 78552 364294 78608
rect 364350 78552 364418 78608
rect 364474 78552 374294 78608
rect 374350 78552 374418 78608
rect 374474 78552 384294 78608
rect 384350 78552 384418 78608
rect 384474 78552 394294 78608
rect 394350 78552 394418 78608
rect 394474 78552 404294 78608
rect 404350 78552 404418 78608
rect 404474 78552 414294 78608
rect 414350 78552 414418 78608
rect 414474 78552 424294 78608
rect 424350 78552 424418 78608
rect 424474 78552 434294 78608
rect 434350 78552 434418 78608
rect 434474 78552 444294 78608
rect 444350 78552 444418 78608
rect 444474 78552 454294 78608
rect 454350 78552 454418 78608
rect 454474 78552 464294 78608
rect 464350 78552 464418 78608
rect 464474 78552 474294 78608
rect 474350 78552 474418 78608
rect 474474 78552 484294 78608
rect 484350 78552 484418 78608
rect 484474 78552 494294 78608
rect 494350 78552 494418 78608
rect 494474 78552 504294 78608
rect 504350 78552 504418 78608
rect 504474 78552 514294 78608
rect 514350 78552 514418 78608
rect 514474 78552 524294 78608
rect 524350 78552 524418 78608
rect 524474 78552 534294 78608
rect 534350 78552 534418 78608
rect 534474 78552 544294 78608
rect 544350 78552 544418 78608
rect 544474 78552 554294 78608
rect 554350 78552 554418 78608
rect 554474 78552 592370 78608
rect 592426 78552 592494 78608
rect 592550 78552 592618 78608
rect 592674 78552 592742 78608
rect 592798 78552 592866 78608
rect 592922 78552 592990 78608
rect 593046 78552 593114 78608
rect 593170 78552 624727 78608
rect 624783 78552 624851 78608
rect 624907 78552 632667 78608
rect 632723 78552 632791 78608
rect 632847 78552 640607 78608
rect 640663 78552 640731 78608
rect 640787 78552 648547 78608
rect 648603 78552 648671 78608
rect 648727 78552 657330 78608
rect 657386 78552 657454 78608
rect 657510 78552 657578 78608
rect 657634 78552 657702 78608
rect 657758 78552 657826 78608
rect 657882 78552 657950 78608
rect 658006 78552 658074 78608
rect 658130 78552 658198 78608
rect 658254 78552 658322 78608
rect 658378 78552 658446 78608
rect 658502 78552 658570 78608
rect 658626 78552 658694 78608
rect 658750 78552 658818 78608
rect 658874 78552 658942 78608
rect 658998 78552 659066 78608
rect 659122 78552 659810 78608
rect 659866 78552 659934 78608
rect 659990 78552 660058 78608
rect 660114 78552 660182 78608
rect 660238 78552 660306 78608
rect 660362 78552 660430 78608
rect 660486 78552 660554 78608
rect 660610 78552 660678 78608
rect 660734 78552 660802 78608
rect 660858 78552 660926 78608
rect 660982 78552 661050 78608
rect 661106 78552 661174 78608
rect 661230 78552 661298 78608
rect 661354 78552 661422 78608
rect 661478 78552 661546 78608
rect 661602 78552 661670 78608
rect 661726 78552 662180 78608
rect 662236 78552 662304 78608
rect 662360 78552 662428 78608
rect 662484 78552 662552 78608
rect 662608 78552 662676 78608
rect 662732 78552 662800 78608
rect 662856 78552 662924 78608
rect 662980 78552 663048 78608
rect 663104 78552 663172 78608
rect 663228 78552 663296 78608
rect 663352 78552 663420 78608
rect 663476 78552 663544 78608
rect 663600 78552 663668 78608
rect 663724 78552 663792 78608
rect 663848 78552 663916 78608
rect 663972 78552 664040 78608
rect 664096 78552 664886 78608
rect 664942 78552 665010 78608
rect 665066 78552 665134 78608
rect 665190 78552 665258 78608
rect 665314 78552 665382 78608
rect 665438 78552 665506 78608
rect 665562 78552 665630 78608
rect 665686 78552 665754 78608
rect 665810 78552 665878 78608
rect 665934 78552 666002 78608
rect 666058 78552 666126 78608
rect 666182 78552 666250 78608
rect 666306 78552 666374 78608
rect 666430 78552 666498 78608
rect 666554 78552 666622 78608
rect 666678 78552 666746 78608
rect 666802 78552 667256 78608
rect 667312 78552 667380 78608
rect 667436 78552 667504 78608
rect 667560 78552 667628 78608
rect 667684 78552 667752 78608
rect 667808 78552 667876 78608
rect 667932 78552 668000 78608
rect 668056 78552 668124 78608
rect 668180 78552 668248 78608
rect 668304 78552 668372 78608
rect 668428 78552 668496 78608
rect 668552 78552 668620 78608
rect 668676 78552 668744 78608
rect 668800 78552 668868 78608
rect 668924 78552 668992 78608
rect 669048 78552 669116 78608
rect 669172 78552 669860 78608
rect 669916 78552 669984 78608
rect 670040 78552 670108 78608
rect 670164 78552 670232 78608
rect 670288 78552 670356 78608
rect 670412 78552 670480 78608
rect 670536 78552 670604 78608
rect 670660 78552 670728 78608
rect 670784 78552 670852 78608
rect 670908 78552 670976 78608
rect 671032 78552 671100 78608
rect 671156 78552 671224 78608
rect 671280 78552 671348 78608
rect 671404 78552 671472 78608
rect 671528 78552 671596 78608
rect 671652 78552 699452 78608
rect 699508 78552 699576 78608
rect 699632 78552 699700 78608
rect 699756 78552 699824 78608
rect 699880 78552 699948 78608
rect 700004 78552 700072 78608
rect 700128 78552 700196 78608
rect 700252 78552 700322 78608
rect 77678 78484 700322 78552
rect 77678 78428 77808 78484
rect 77864 78428 77932 78484
rect 77988 78428 78056 78484
rect 78112 78428 78180 78484
rect 78236 78428 78304 78484
rect 78360 78428 78428 78484
rect 78484 78428 78552 78484
rect 78608 78428 94294 78484
rect 94350 78428 94418 78484
rect 94474 78428 104294 78484
rect 104350 78428 104418 78484
rect 104474 78428 124294 78484
rect 124350 78428 124418 78484
rect 124474 78428 134294 78484
rect 134350 78428 134418 78484
rect 134474 78428 144294 78484
rect 144350 78428 144418 78484
rect 144474 78428 154294 78484
rect 154350 78428 154418 78484
rect 154474 78428 164294 78484
rect 164350 78428 164418 78484
rect 164474 78428 174294 78484
rect 174350 78428 174418 78484
rect 174474 78428 184294 78484
rect 184350 78428 184418 78484
rect 184474 78428 194294 78484
rect 194350 78428 194418 78484
rect 194474 78428 204294 78484
rect 204350 78428 204418 78484
rect 204474 78428 214294 78484
rect 214350 78428 214418 78484
rect 214474 78428 224294 78484
rect 224350 78428 224418 78484
rect 224474 78428 234294 78484
rect 234350 78428 234418 78484
rect 234474 78428 244294 78484
rect 244350 78428 244418 78484
rect 244474 78428 254294 78484
rect 254350 78428 254418 78484
rect 254474 78428 264294 78484
rect 264350 78428 264418 78484
rect 264474 78428 294294 78484
rect 294350 78428 294418 78484
rect 294474 78428 304294 78484
rect 304350 78428 304418 78484
rect 304474 78428 314294 78484
rect 314350 78428 314418 78484
rect 314474 78428 324294 78484
rect 324350 78428 324418 78484
rect 324474 78428 334294 78484
rect 334350 78428 334418 78484
rect 334474 78428 344294 78484
rect 344350 78428 344418 78484
rect 344474 78428 354294 78484
rect 354350 78428 354418 78484
rect 354474 78428 364294 78484
rect 364350 78428 364418 78484
rect 364474 78428 374294 78484
rect 374350 78428 374418 78484
rect 374474 78428 384294 78484
rect 384350 78428 384418 78484
rect 384474 78428 394294 78484
rect 394350 78428 394418 78484
rect 394474 78428 404294 78484
rect 404350 78428 404418 78484
rect 404474 78428 414294 78484
rect 414350 78428 414418 78484
rect 414474 78428 424294 78484
rect 424350 78428 424418 78484
rect 424474 78428 434294 78484
rect 434350 78428 434418 78484
rect 434474 78428 444294 78484
rect 444350 78428 444418 78484
rect 444474 78428 454294 78484
rect 454350 78428 454418 78484
rect 454474 78428 464294 78484
rect 464350 78428 464418 78484
rect 464474 78428 474294 78484
rect 474350 78428 474418 78484
rect 474474 78428 484294 78484
rect 484350 78428 484418 78484
rect 484474 78428 494294 78484
rect 494350 78428 494418 78484
rect 494474 78428 504294 78484
rect 504350 78428 504418 78484
rect 504474 78428 514294 78484
rect 514350 78428 514418 78484
rect 514474 78428 524294 78484
rect 524350 78428 524418 78484
rect 524474 78428 534294 78484
rect 534350 78428 534418 78484
rect 534474 78428 544294 78484
rect 544350 78428 544418 78484
rect 544474 78428 554294 78484
rect 554350 78428 554418 78484
rect 554474 78428 592370 78484
rect 592426 78428 592494 78484
rect 592550 78428 592618 78484
rect 592674 78428 592742 78484
rect 592798 78428 592866 78484
rect 592922 78428 592990 78484
rect 593046 78428 593114 78484
rect 593170 78428 624727 78484
rect 624783 78428 624851 78484
rect 624907 78428 632667 78484
rect 632723 78428 632791 78484
rect 632847 78428 640607 78484
rect 640663 78428 640731 78484
rect 640787 78428 648547 78484
rect 648603 78428 648671 78484
rect 648727 78428 657330 78484
rect 657386 78428 657454 78484
rect 657510 78428 657578 78484
rect 657634 78428 657702 78484
rect 657758 78428 657826 78484
rect 657882 78428 657950 78484
rect 658006 78428 658074 78484
rect 658130 78428 658198 78484
rect 658254 78428 658322 78484
rect 658378 78428 658446 78484
rect 658502 78428 658570 78484
rect 658626 78428 658694 78484
rect 658750 78428 658818 78484
rect 658874 78428 658942 78484
rect 658998 78428 659066 78484
rect 659122 78428 659810 78484
rect 659866 78428 659934 78484
rect 659990 78428 660058 78484
rect 660114 78428 660182 78484
rect 660238 78428 660306 78484
rect 660362 78428 660430 78484
rect 660486 78428 660554 78484
rect 660610 78428 660678 78484
rect 660734 78428 660802 78484
rect 660858 78428 660926 78484
rect 660982 78428 661050 78484
rect 661106 78428 661174 78484
rect 661230 78428 661298 78484
rect 661354 78428 661422 78484
rect 661478 78428 661546 78484
rect 661602 78428 661670 78484
rect 661726 78428 662180 78484
rect 662236 78428 662304 78484
rect 662360 78428 662428 78484
rect 662484 78428 662552 78484
rect 662608 78428 662676 78484
rect 662732 78428 662800 78484
rect 662856 78428 662924 78484
rect 662980 78428 663048 78484
rect 663104 78428 663172 78484
rect 663228 78428 663296 78484
rect 663352 78428 663420 78484
rect 663476 78428 663544 78484
rect 663600 78428 663668 78484
rect 663724 78428 663792 78484
rect 663848 78428 663916 78484
rect 663972 78428 664040 78484
rect 664096 78428 664886 78484
rect 664942 78428 665010 78484
rect 665066 78428 665134 78484
rect 665190 78428 665258 78484
rect 665314 78428 665382 78484
rect 665438 78428 665506 78484
rect 665562 78428 665630 78484
rect 665686 78428 665754 78484
rect 665810 78428 665878 78484
rect 665934 78428 666002 78484
rect 666058 78428 666126 78484
rect 666182 78428 666250 78484
rect 666306 78428 666374 78484
rect 666430 78428 666498 78484
rect 666554 78428 666622 78484
rect 666678 78428 666746 78484
rect 666802 78428 667256 78484
rect 667312 78428 667380 78484
rect 667436 78428 667504 78484
rect 667560 78428 667628 78484
rect 667684 78428 667752 78484
rect 667808 78428 667876 78484
rect 667932 78428 668000 78484
rect 668056 78428 668124 78484
rect 668180 78428 668248 78484
rect 668304 78428 668372 78484
rect 668428 78428 668496 78484
rect 668552 78428 668620 78484
rect 668676 78428 668744 78484
rect 668800 78428 668868 78484
rect 668924 78428 668992 78484
rect 669048 78428 669116 78484
rect 669172 78428 669860 78484
rect 669916 78428 669984 78484
rect 670040 78428 670108 78484
rect 670164 78428 670232 78484
rect 670288 78428 670356 78484
rect 670412 78428 670480 78484
rect 670536 78428 670604 78484
rect 670660 78428 670728 78484
rect 670784 78428 670852 78484
rect 670908 78428 670976 78484
rect 671032 78428 671100 78484
rect 671156 78428 671224 78484
rect 671280 78428 671348 78484
rect 671404 78428 671472 78484
rect 671528 78428 671596 78484
rect 671652 78428 699452 78484
rect 699508 78428 699576 78484
rect 699632 78428 699700 78484
rect 699756 78428 699824 78484
rect 699880 78428 699948 78484
rect 700004 78428 700072 78484
rect 700128 78428 700196 78484
rect 700252 78428 700322 78484
rect 77678 78360 700322 78428
rect 77678 78304 77808 78360
rect 77864 78304 77932 78360
rect 77988 78304 78056 78360
rect 78112 78304 78180 78360
rect 78236 78304 78304 78360
rect 78360 78304 78428 78360
rect 78484 78304 78552 78360
rect 78608 78304 94294 78360
rect 94350 78304 94418 78360
rect 94474 78304 104294 78360
rect 104350 78304 104418 78360
rect 104474 78304 124294 78360
rect 124350 78304 124418 78360
rect 124474 78304 134294 78360
rect 134350 78304 134418 78360
rect 134474 78304 144294 78360
rect 144350 78304 144418 78360
rect 144474 78304 154294 78360
rect 154350 78304 154418 78360
rect 154474 78304 164294 78360
rect 164350 78304 164418 78360
rect 164474 78304 174294 78360
rect 174350 78304 174418 78360
rect 174474 78304 184294 78360
rect 184350 78304 184418 78360
rect 184474 78304 194294 78360
rect 194350 78304 194418 78360
rect 194474 78304 204294 78360
rect 204350 78304 204418 78360
rect 204474 78304 214294 78360
rect 214350 78304 214418 78360
rect 214474 78304 224294 78360
rect 224350 78304 224418 78360
rect 224474 78304 234294 78360
rect 234350 78304 234418 78360
rect 234474 78304 244294 78360
rect 244350 78304 244418 78360
rect 244474 78304 254294 78360
rect 254350 78304 254418 78360
rect 254474 78304 264294 78360
rect 264350 78304 264418 78360
rect 264474 78304 294294 78360
rect 294350 78304 294418 78360
rect 294474 78304 304294 78360
rect 304350 78304 304418 78360
rect 304474 78304 314294 78360
rect 314350 78304 314418 78360
rect 314474 78304 324294 78360
rect 324350 78304 324418 78360
rect 324474 78304 334294 78360
rect 334350 78304 334418 78360
rect 334474 78304 344294 78360
rect 344350 78304 344418 78360
rect 344474 78304 354294 78360
rect 354350 78304 354418 78360
rect 354474 78304 364294 78360
rect 364350 78304 364418 78360
rect 364474 78304 374294 78360
rect 374350 78304 374418 78360
rect 374474 78304 384294 78360
rect 384350 78304 384418 78360
rect 384474 78304 394294 78360
rect 394350 78304 394418 78360
rect 394474 78304 404294 78360
rect 404350 78304 404418 78360
rect 404474 78304 414294 78360
rect 414350 78304 414418 78360
rect 414474 78304 424294 78360
rect 424350 78304 424418 78360
rect 424474 78304 434294 78360
rect 434350 78304 434418 78360
rect 434474 78304 444294 78360
rect 444350 78304 444418 78360
rect 444474 78304 454294 78360
rect 454350 78304 454418 78360
rect 454474 78304 464294 78360
rect 464350 78304 464418 78360
rect 464474 78304 474294 78360
rect 474350 78304 474418 78360
rect 474474 78304 484294 78360
rect 484350 78304 484418 78360
rect 484474 78304 494294 78360
rect 494350 78304 494418 78360
rect 494474 78304 504294 78360
rect 504350 78304 504418 78360
rect 504474 78304 514294 78360
rect 514350 78304 514418 78360
rect 514474 78304 524294 78360
rect 524350 78304 524418 78360
rect 524474 78304 534294 78360
rect 534350 78304 534418 78360
rect 534474 78304 544294 78360
rect 544350 78304 544418 78360
rect 544474 78304 554294 78360
rect 554350 78304 554418 78360
rect 554474 78304 592370 78360
rect 592426 78304 592494 78360
rect 592550 78304 592618 78360
rect 592674 78304 592742 78360
rect 592798 78304 592866 78360
rect 592922 78304 592990 78360
rect 593046 78304 593114 78360
rect 593170 78304 624727 78360
rect 624783 78304 624851 78360
rect 624907 78304 632667 78360
rect 632723 78304 632791 78360
rect 632847 78304 640607 78360
rect 640663 78304 640731 78360
rect 640787 78304 648547 78360
rect 648603 78304 648671 78360
rect 648727 78304 657330 78360
rect 657386 78304 657454 78360
rect 657510 78304 657578 78360
rect 657634 78304 657702 78360
rect 657758 78304 657826 78360
rect 657882 78304 657950 78360
rect 658006 78304 658074 78360
rect 658130 78304 658198 78360
rect 658254 78304 658322 78360
rect 658378 78304 658446 78360
rect 658502 78304 658570 78360
rect 658626 78304 658694 78360
rect 658750 78304 658818 78360
rect 658874 78304 658942 78360
rect 658998 78304 659066 78360
rect 659122 78304 659810 78360
rect 659866 78304 659934 78360
rect 659990 78304 660058 78360
rect 660114 78304 660182 78360
rect 660238 78304 660306 78360
rect 660362 78304 660430 78360
rect 660486 78304 660554 78360
rect 660610 78304 660678 78360
rect 660734 78304 660802 78360
rect 660858 78304 660926 78360
rect 660982 78304 661050 78360
rect 661106 78304 661174 78360
rect 661230 78304 661298 78360
rect 661354 78304 661422 78360
rect 661478 78304 661546 78360
rect 661602 78304 661670 78360
rect 661726 78304 662180 78360
rect 662236 78304 662304 78360
rect 662360 78304 662428 78360
rect 662484 78304 662552 78360
rect 662608 78304 662676 78360
rect 662732 78304 662800 78360
rect 662856 78304 662924 78360
rect 662980 78304 663048 78360
rect 663104 78304 663172 78360
rect 663228 78304 663296 78360
rect 663352 78304 663420 78360
rect 663476 78304 663544 78360
rect 663600 78304 663668 78360
rect 663724 78304 663792 78360
rect 663848 78304 663916 78360
rect 663972 78304 664040 78360
rect 664096 78304 664886 78360
rect 664942 78304 665010 78360
rect 665066 78304 665134 78360
rect 665190 78304 665258 78360
rect 665314 78304 665382 78360
rect 665438 78304 665506 78360
rect 665562 78304 665630 78360
rect 665686 78304 665754 78360
rect 665810 78304 665878 78360
rect 665934 78304 666002 78360
rect 666058 78304 666126 78360
rect 666182 78304 666250 78360
rect 666306 78304 666374 78360
rect 666430 78304 666498 78360
rect 666554 78304 666622 78360
rect 666678 78304 666746 78360
rect 666802 78304 667256 78360
rect 667312 78304 667380 78360
rect 667436 78304 667504 78360
rect 667560 78304 667628 78360
rect 667684 78304 667752 78360
rect 667808 78304 667876 78360
rect 667932 78304 668000 78360
rect 668056 78304 668124 78360
rect 668180 78304 668248 78360
rect 668304 78304 668372 78360
rect 668428 78304 668496 78360
rect 668552 78304 668620 78360
rect 668676 78304 668744 78360
rect 668800 78304 668868 78360
rect 668924 78304 668992 78360
rect 669048 78304 669116 78360
rect 669172 78304 669860 78360
rect 669916 78304 669984 78360
rect 670040 78304 670108 78360
rect 670164 78304 670232 78360
rect 670288 78304 670356 78360
rect 670412 78304 670480 78360
rect 670536 78304 670604 78360
rect 670660 78304 670728 78360
rect 670784 78304 670852 78360
rect 670908 78304 670976 78360
rect 671032 78304 671100 78360
rect 671156 78304 671224 78360
rect 671280 78304 671348 78360
rect 671404 78304 671472 78360
rect 671528 78304 671596 78360
rect 671652 78304 699452 78360
rect 699508 78304 699576 78360
rect 699632 78304 699700 78360
rect 699756 78304 699824 78360
rect 699880 78304 699948 78360
rect 700004 78304 700072 78360
rect 700128 78304 700196 78360
rect 700252 78304 700322 78360
rect 77678 78236 700322 78304
rect 77678 78180 77808 78236
rect 77864 78180 77932 78236
rect 77988 78180 78056 78236
rect 78112 78180 78180 78236
rect 78236 78180 78304 78236
rect 78360 78180 78428 78236
rect 78484 78180 78552 78236
rect 78608 78180 94294 78236
rect 94350 78180 94418 78236
rect 94474 78180 104294 78236
rect 104350 78180 104418 78236
rect 104474 78180 124294 78236
rect 124350 78180 124418 78236
rect 124474 78180 134294 78236
rect 134350 78180 134418 78236
rect 134474 78180 144294 78236
rect 144350 78180 144418 78236
rect 144474 78180 154294 78236
rect 154350 78180 154418 78236
rect 154474 78180 164294 78236
rect 164350 78180 164418 78236
rect 164474 78180 174294 78236
rect 174350 78180 174418 78236
rect 174474 78180 184294 78236
rect 184350 78180 184418 78236
rect 184474 78180 194294 78236
rect 194350 78180 194418 78236
rect 194474 78180 204294 78236
rect 204350 78180 204418 78236
rect 204474 78180 214294 78236
rect 214350 78180 214418 78236
rect 214474 78180 224294 78236
rect 224350 78180 224418 78236
rect 224474 78180 234294 78236
rect 234350 78180 234418 78236
rect 234474 78180 244294 78236
rect 244350 78180 244418 78236
rect 244474 78180 254294 78236
rect 254350 78180 254418 78236
rect 254474 78180 264294 78236
rect 264350 78180 264418 78236
rect 264474 78180 294294 78236
rect 294350 78180 294418 78236
rect 294474 78180 304294 78236
rect 304350 78180 304418 78236
rect 304474 78180 314294 78236
rect 314350 78180 314418 78236
rect 314474 78180 324294 78236
rect 324350 78180 324418 78236
rect 324474 78180 334294 78236
rect 334350 78180 334418 78236
rect 334474 78180 344294 78236
rect 344350 78180 344418 78236
rect 344474 78180 354294 78236
rect 354350 78180 354418 78236
rect 354474 78180 364294 78236
rect 364350 78180 364418 78236
rect 364474 78180 374294 78236
rect 374350 78180 374418 78236
rect 374474 78180 384294 78236
rect 384350 78180 384418 78236
rect 384474 78180 394294 78236
rect 394350 78180 394418 78236
rect 394474 78180 404294 78236
rect 404350 78180 404418 78236
rect 404474 78180 414294 78236
rect 414350 78180 414418 78236
rect 414474 78180 424294 78236
rect 424350 78180 424418 78236
rect 424474 78180 434294 78236
rect 434350 78180 434418 78236
rect 434474 78180 444294 78236
rect 444350 78180 444418 78236
rect 444474 78180 454294 78236
rect 454350 78180 454418 78236
rect 454474 78180 464294 78236
rect 464350 78180 464418 78236
rect 464474 78180 474294 78236
rect 474350 78180 474418 78236
rect 474474 78180 484294 78236
rect 484350 78180 484418 78236
rect 484474 78180 494294 78236
rect 494350 78180 494418 78236
rect 494474 78180 504294 78236
rect 504350 78180 504418 78236
rect 504474 78180 514294 78236
rect 514350 78180 514418 78236
rect 514474 78180 524294 78236
rect 524350 78180 524418 78236
rect 524474 78180 534294 78236
rect 534350 78180 534418 78236
rect 534474 78180 544294 78236
rect 544350 78180 544418 78236
rect 544474 78180 554294 78236
rect 554350 78180 554418 78236
rect 554474 78180 592370 78236
rect 592426 78180 592494 78236
rect 592550 78180 592618 78236
rect 592674 78180 592742 78236
rect 592798 78180 592866 78236
rect 592922 78180 592990 78236
rect 593046 78180 593114 78236
rect 593170 78180 624727 78236
rect 624783 78180 624851 78236
rect 624907 78180 632667 78236
rect 632723 78180 632791 78236
rect 632847 78180 640607 78236
rect 640663 78180 640731 78236
rect 640787 78180 648547 78236
rect 648603 78180 648671 78236
rect 648727 78180 657330 78236
rect 657386 78180 657454 78236
rect 657510 78180 657578 78236
rect 657634 78180 657702 78236
rect 657758 78180 657826 78236
rect 657882 78180 657950 78236
rect 658006 78180 658074 78236
rect 658130 78180 658198 78236
rect 658254 78180 658322 78236
rect 658378 78180 658446 78236
rect 658502 78180 658570 78236
rect 658626 78180 658694 78236
rect 658750 78180 658818 78236
rect 658874 78180 658942 78236
rect 658998 78180 659066 78236
rect 659122 78180 659810 78236
rect 659866 78180 659934 78236
rect 659990 78180 660058 78236
rect 660114 78180 660182 78236
rect 660238 78180 660306 78236
rect 660362 78180 660430 78236
rect 660486 78180 660554 78236
rect 660610 78180 660678 78236
rect 660734 78180 660802 78236
rect 660858 78180 660926 78236
rect 660982 78180 661050 78236
rect 661106 78180 661174 78236
rect 661230 78180 661298 78236
rect 661354 78180 661422 78236
rect 661478 78180 661546 78236
rect 661602 78180 661670 78236
rect 661726 78180 662180 78236
rect 662236 78180 662304 78236
rect 662360 78180 662428 78236
rect 662484 78180 662552 78236
rect 662608 78180 662676 78236
rect 662732 78180 662800 78236
rect 662856 78180 662924 78236
rect 662980 78180 663048 78236
rect 663104 78180 663172 78236
rect 663228 78180 663296 78236
rect 663352 78180 663420 78236
rect 663476 78180 663544 78236
rect 663600 78180 663668 78236
rect 663724 78180 663792 78236
rect 663848 78180 663916 78236
rect 663972 78180 664040 78236
rect 664096 78180 664886 78236
rect 664942 78180 665010 78236
rect 665066 78180 665134 78236
rect 665190 78180 665258 78236
rect 665314 78180 665382 78236
rect 665438 78180 665506 78236
rect 665562 78180 665630 78236
rect 665686 78180 665754 78236
rect 665810 78180 665878 78236
rect 665934 78180 666002 78236
rect 666058 78180 666126 78236
rect 666182 78180 666250 78236
rect 666306 78180 666374 78236
rect 666430 78180 666498 78236
rect 666554 78180 666622 78236
rect 666678 78180 666746 78236
rect 666802 78180 667256 78236
rect 667312 78180 667380 78236
rect 667436 78180 667504 78236
rect 667560 78180 667628 78236
rect 667684 78180 667752 78236
rect 667808 78180 667876 78236
rect 667932 78180 668000 78236
rect 668056 78180 668124 78236
rect 668180 78180 668248 78236
rect 668304 78180 668372 78236
rect 668428 78180 668496 78236
rect 668552 78180 668620 78236
rect 668676 78180 668744 78236
rect 668800 78180 668868 78236
rect 668924 78180 668992 78236
rect 669048 78180 669116 78236
rect 669172 78180 669860 78236
rect 669916 78180 669984 78236
rect 670040 78180 670108 78236
rect 670164 78180 670232 78236
rect 670288 78180 670356 78236
rect 670412 78180 670480 78236
rect 670536 78180 670604 78236
rect 670660 78180 670728 78236
rect 670784 78180 670852 78236
rect 670908 78180 670976 78236
rect 671032 78180 671100 78236
rect 671156 78180 671224 78236
rect 671280 78180 671348 78236
rect 671404 78180 671472 78236
rect 671528 78180 671596 78236
rect 671652 78180 699452 78236
rect 699508 78180 699576 78236
rect 699632 78180 699700 78236
rect 699756 78180 699824 78236
rect 699880 78180 699948 78236
rect 700004 78180 700072 78236
rect 700128 78180 700196 78236
rect 700252 78180 700322 78236
rect 77678 78112 700322 78180
rect 77678 78056 77808 78112
rect 77864 78056 77932 78112
rect 77988 78056 78056 78112
rect 78112 78056 78180 78112
rect 78236 78056 78304 78112
rect 78360 78056 78428 78112
rect 78484 78056 78552 78112
rect 78608 78056 94294 78112
rect 94350 78056 94418 78112
rect 94474 78056 104294 78112
rect 104350 78056 104418 78112
rect 104474 78056 124294 78112
rect 124350 78056 124418 78112
rect 124474 78056 134294 78112
rect 134350 78056 134418 78112
rect 134474 78056 144294 78112
rect 144350 78056 144418 78112
rect 144474 78056 154294 78112
rect 154350 78056 154418 78112
rect 154474 78056 164294 78112
rect 164350 78056 164418 78112
rect 164474 78056 174294 78112
rect 174350 78056 174418 78112
rect 174474 78056 184294 78112
rect 184350 78056 184418 78112
rect 184474 78056 194294 78112
rect 194350 78056 194418 78112
rect 194474 78056 204294 78112
rect 204350 78056 204418 78112
rect 204474 78056 214294 78112
rect 214350 78056 214418 78112
rect 214474 78056 224294 78112
rect 224350 78056 224418 78112
rect 224474 78056 234294 78112
rect 234350 78056 234418 78112
rect 234474 78056 244294 78112
rect 244350 78056 244418 78112
rect 244474 78056 254294 78112
rect 254350 78056 254418 78112
rect 254474 78056 264294 78112
rect 264350 78056 264418 78112
rect 264474 78056 294294 78112
rect 294350 78056 294418 78112
rect 294474 78056 304294 78112
rect 304350 78056 304418 78112
rect 304474 78056 314294 78112
rect 314350 78056 314418 78112
rect 314474 78056 324294 78112
rect 324350 78056 324418 78112
rect 324474 78056 334294 78112
rect 334350 78056 334418 78112
rect 334474 78056 344294 78112
rect 344350 78056 344418 78112
rect 344474 78056 354294 78112
rect 354350 78056 354418 78112
rect 354474 78056 364294 78112
rect 364350 78056 364418 78112
rect 364474 78056 374294 78112
rect 374350 78056 374418 78112
rect 374474 78056 384294 78112
rect 384350 78056 384418 78112
rect 384474 78056 394294 78112
rect 394350 78056 394418 78112
rect 394474 78056 404294 78112
rect 404350 78056 404418 78112
rect 404474 78056 414294 78112
rect 414350 78056 414418 78112
rect 414474 78056 424294 78112
rect 424350 78056 424418 78112
rect 424474 78056 434294 78112
rect 434350 78056 434418 78112
rect 434474 78056 444294 78112
rect 444350 78056 444418 78112
rect 444474 78056 454294 78112
rect 454350 78056 454418 78112
rect 454474 78056 464294 78112
rect 464350 78056 464418 78112
rect 464474 78056 474294 78112
rect 474350 78056 474418 78112
rect 474474 78056 484294 78112
rect 484350 78056 484418 78112
rect 484474 78056 494294 78112
rect 494350 78056 494418 78112
rect 494474 78056 504294 78112
rect 504350 78056 504418 78112
rect 504474 78056 514294 78112
rect 514350 78056 514418 78112
rect 514474 78056 524294 78112
rect 524350 78056 524418 78112
rect 524474 78056 534294 78112
rect 534350 78056 534418 78112
rect 534474 78056 544294 78112
rect 544350 78056 544418 78112
rect 544474 78056 554294 78112
rect 554350 78056 554418 78112
rect 554474 78056 592370 78112
rect 592426 78056 592494 78112
rect 592550 78056 592618 78112
rect 592674 78056 592742 78112
rect 592798 78056 592866 78112
rect 592922 78056 592990 78112
rect 593046 78056 593114 78112
rect 593170 78056 624727 78112
rect 624783 78056 624851 78112
rect 624907 78056 632667 78112
rect 632723 78056 632791 78112
rect 632847 78056 640607 78112
rect 640663 78056 640731 78112
rect 640787 78056 648547 78112
rect 648603 78056 648671 78112
rect 648727 78056 657330 78112
rect 657386 78056 657454 78112
rect 657510 78056 657578 78112
rect 657634 78056 657702 78112
rect 657758 78056 657826 78112
rect 657882 78056 657950 78112
rect 658006 78056 658074 78112
rect 658130 78056 658198 78112
rect 658254 78056 658322 78112
rect 658378 78056 658446 78112
rect 658502 78056 658570 78112
rect 658626 78056 658694 78112
rect 658750 78056 658818 78112
rect 658874 78056 658942 78112
rect 658998 78056 659066 78112
rect 659122 78056 659810 78112
rect 659866 78056 659934 78112
rect 659990 78056 660058 78112
rect 660114 78056 660182 78112
rect 660238 78056 660306 78112
rect 660362 78056 660430 78112
rect 660486 78056 660554 78112
rect 660610 78056 660678 78112
rect 660734 78056 660802 78112
rect 660858 78056 660926 78112
rect 660982 78056 661050 78112
rect 661106 78056 661174 78112
rect 661230 78056 661298 78112
rect 661354 78056 661422 78112
rect 661478 78056 661546 78112
rect 661602 78056 661670 78112
rect 661726 78056 662180 78112
rect 662236 78056 662304 78112
rect 662360 78056 662428 78112
rect 662484 78056 662552 78112
rect 662608 78056 662676 78112
rect 662732 78056 662800 78112
rect 662856 78056 662924 78112
rect 662980 78056 663048 78112
rect 663104 78056 663172 78112
rect 663228 78056 663296 78112
rect 663352 78056 663420 78112
rect 663476 78056 663544 78112
rect 663600 78056 663668 78112
rect 663724 78056 663792 78112
rect 663848 78056 663916 78112
rect 663972 78056 664040 78112
rect 664096 78056 664886 78112
rect 664942 78056 665010 78112
rect 665066 78056 665134 78112
rect 665190 78056 665258 78112
rect 665314 78056 665382 78112
rect 665438 78056 665506 78112
rect 665562 78056 665630 78112
rect 665686 78056 665754 78112
rect 665810 78056 665878 78112
rect 665934 78056 666002 78112
rect 666058 78056 666126 78112
rect 666182 78056 666250 78112
rect 666306 78056 666374 78112
rect 666430 78056 666498 78112
rect 666554 78056 666622 78112
rect 666678 78056 666746 78112
rect 666802 78056 667256 78112
rect 667312 78056 667380 78112
rect 667436 78056 667504 78112
rect 667560 78056 667628 78112
rect 667684 78056 667752 78112
rect 667808 78056 667876 78112
rect 667932 78056 668000 78112
rect 668056 78056 668124 78112
rect 668180 78056 668248 78112
rect 668304 78056 668372 78112
rect 668428 78056 668496 78112
rect 668552 78056 668620 78112
rect 668676 78056 668744 78112
rect 668800 78056 668868 78112
rect 668924 78056 668992 78112
rect 669048 78056 669116 78112
rect 669172 78056 669860 78112
rect 669916 78056 669984 78112
rect 670040 78056 670108 78112
rect 670164 78056 670232 78112
rect 670288 78056 670356 78112
rect 670412 78056 670480 78112
rect 670536 78056 670604 78112
rect 670660 78056 670728 78112
rect 670784 78056 670852 78112
rect 670908 78056 670976 78112
rect 671032 78056 671100 78112
rect 671156 78056 671224 78112
rect 671280 78056 671348 78112
rect 671404 78056 671472 78112
rect 671528 78056 671596 78112
rect 671652 78056 699452 78112
rect 699508 78056 699576 78112
rect 699632 78056 699700 78112
rect 699756 78056 699824 78112
rect 699880 78056 699948 78112
rect 700004 78056 700072 78112
rect 700128 78056 700196 78112
rect 700252 78056 700322 78112
rect 77678 77988 700322 78056
rect 77678 77932 77808 77988
rect 77864 77932 77932 77988
rect 77988 77932 78056 77988
rect 78112 77932 78180 77988
rect 78236 77932 78304 77988
rect 78360 77932 78428 77988
rect 78484 77932 78552 77988
rect 78608 77932 94294 77988
rect 94350 77932 94418 77988
rect 94474 77932 104294 77988
rect 104350 77932 104418 77988
rect 104474 77932 124294 77988
rect 124350 77932 124418 77988
rect 124474 77932 134294 77988
rect 134350 77932 134418 77988
rect 134474 77932 144294 77988
rect 144350 77932 144418 77988
rect 144474 77932 154294 77988
rect 154350 77932 154418 77988
rect 154474 77932 164294 77988
rect 164350 77932 164418 77988
rect 164474 77932 174294 77988
rect 174350 77932 174418 77988
rect 174474 77932 184294 77988
rect 184350 77932 184418 77988
rect 184474 77932 194294 77988
rect 194350 77932 194418 77988
rect 194474 77932 204294 77988
rect 204350 77932 204418 77988
rect 204474 77932 214294 77988
rect 214350 77932 214418 77988
rect 214474 77932 224294 77988
rect 224350 77932 224418 77988
rect 224474 77932 234294 77988
rect 234350 77932 234418 77988
rect 234474 77932 244294 77988
rect 244350 77932 244418 77988
rect 244474 77932 254294 77988
rect 254350 77932 254418 77988
rect 254474 77932 264294 77988
rect 264350 77932 264418 77988
rect 264474 77932 294294 77988
rect 294350 77932 294418 77988
rect 294474 77932 304294 77988
rect 304350 77932 304418 77988
rect 304474 77932 314294 77988
rect 314350 77932 314418 77988
rect 314474 77932 324294 77988
rect 324350 77932 324418 77988
rect 324474 77932 334294 77988
rect 334350 77932 334418 77988
rect 334474 77932 344294 77988
rect 344350 77932 344418 77988
rect 344474 77932 354294 77988
rect 354350 77932 354418 77988
rect 354474 77932 364294 77988
rect 364350 77932 364418 77988
rect 364474 77932 374294 77988
rect 374350 77932 374418 77988
rect 374474 77932 384294 77988
rect 384350 77932 384418 77988
rect 384474 77932 394294 77988
rect 394350 77932 394418 77988
rect 394474 77932 404294 77988
rect 404350 77932 404418 77988
rect 404474 77932 414294 77988
rect 414350 77932 414418 77988
rect 414474 77932 424294 77988
rect 424350 77932 424418 77988
rect 424474 77932 434294 77988
rect 434350 77932 434418 77988
rect 434474 77932 444294 77988
rect 444350 77932 444418 77988
rect 444474 77932 454294 77988
rect 454350 77932 454418 77988
rect 454474 77932 464294 77988
rect 464350 77932 464418 77988
rect 464474 77932 474294 77988
rect 474350 77932 474418 77988
rect 474474 77932 484294 77988
rect 484350 77932 484418 77988
rect 484474 77932 494294 77988
rect 494350 77932 494418 77988
rect 494474 77932 504294 77988
rect 504350 77932 504418 77988
rect 504474 77932 514294 77988
rect 514350 77932 514418 77988
rect 514474 77932 524294 77988
rect 524350 77932 524418 77988
rect 524474 77932 534294 77988
rect 534350 77932 534418 77988
rect 534474 77932 544294 77988
rect 544350 77932 544418 77988
rect 544474 77932 554294 77988
rect 554350 77932 554418 77988
rect 554474 77932 592370 77988
rect 592426 77932 592494 77988
rect 592550 77932 592618 77988
rect 592674 77932 592742 77988
rect 592798 77932 592866 77988
rect 592922 77932 592990 77988
rect 593046 77932 593114 77988
rect 593170 77932 624727 77988
rect 624783 77932 624851 77988
rect 624907 77932 632667 77988
rect 632723 77932 632791 77988
rect 632847 77932 640607 77988
rect 640663 77932 640731 77988
rect 640787 77932 648547 77988
rect 648603 77932 648671 77988
rect 648727 77932 657330 77988
rect 657386 77932 657454 77988
rect 657510 77932 657578 77988
rect 657634 77932 657702 77988
rect 657758 77932 657826 77988
rect 657882 77932 657950 77988
rect 658006 77932 658074 77988
rect 658130 77932 658198 77988
rect 658254 77932 658322 77988
rect 658378 77932 658446 77988
rect 658502 77932 658570 77988
rect 658626 77932 658694 77988
rect 658750 77932 658818 77988
rect 658874 77932 658942 77988
rect 658998 77932 659066 77988
rect 659122 77932 659810 77988
rect 659866 77932 659934 77988
rect 659990 77932 660058 77988
rect 660114 77932 660182 77988
rect 660238 77932 660306 77988
rect 660362 77932 660430 77988
rect 660486 77932 660554 77988
rect 660610 77932 660678 77988
rect 660734 77932 660802 77988
rect 660858 77932 660926 77988
rect 660982 77932 661050 77988
rect 661106 77932 661174 77988
rect 661230 77932 661298 77988
rect 661354 77932 661422 77988
rect 661478 77932 661546 77988
rect 661602 77932 661670 77988
rect 661726 77932 662180 77988
rect 662236 77932 662304 77988
rect 662360 77932 662428 77988
rect 662484 77932 662552 77988
rect 662608 77932 662676 77988
rect 662732 77932 662800 77988
rect 662856 77932 662924 77988
rect 662980 77932 663048 77988
rect 663104 77932 663172 77988
rect 663228 77932 663296 77988
rect 663352 77932 663420 77988
rect 663476 77932 663544 77988
rect 663600 77932 663668 77988
rect 663724 77932 663792 77988
rect 663848 77932 663916 77988
rect 663972 77932 664040 77988
rect 664096 77932 664886 77988
rect 664942 77932 665010 77988
rect 665066 77932 665134 77988
rect 665190 77932 665258 77988
rect 665314 77932 665382 77988
rect 665438 77932 665506 77988
rect 665562 77932 665630 77988
rect 665686 77932 665754 77988
rect 665810 77932 665878 77988
rect 665934 77932 666002 77988
rect 666058 77932 666126 77988
rect 666182 77932 666250 77988
rect 666306 77932 666374 77988
rect 666430 77932 666498 77988
rect 666554 77932 666622 77988
rect 666678 77932 666746 77988
rect 666802 77932 667256 77988
rect 667312 77932 667380 77988
rect 667436 77932 667504 77988
rect 667560 77932 667628 77988
rect 667684 77932 667752 77988
rect 667808 77932 667876 77988
rect 667932 77932 668000 77988
rect 668056 77932 668124 77988
rect 668180 77932 668248 77988
rect 668304 77932 668372 77988
rect 668428 77932 668496 77988
rect 668552 77932 668620 77988
rect 668676 77932 668744 77988
rect 668800 77932 668868 77988
rect 668924 77932 668992 77988
rect 669048 77932 669116 77988
rect 669172 77932 669860 77988
rect 669916 77932 669984 77988
rect 670040 77932 670108 77988
rect 670164 77932 670232 77988
rect 670288 77932 670356 77988
rect 670412 77932 670480 77988
rect 670536 77932 670604 77988
rect 670660 77932 670728 77988
rect 670784 77932 670852 77988
rect 670908 77932 670976 77988
rect 671032 77932 671100 77988
rect 671156 77932 671224 77988
rect 671280 77932 671348 77988
rect 671404 77932 671472 77988
rect 671528 77932 671596 77988
rect 671652 77932 699452 77988
rect 699508 77932 699576 77988
rect 699632 77932 699700 77988
rect 699756 77932 699824 77988
rect 699880 77932 699948 77988
rect 700004 77932 700072 77988
rect 700128 77932 700196 77988
rect 700252 77932 700322 77988
rect 77678 77864 700322 77932
rect 77678 77808 77808 77864
rect 77864 77808 77932 77864
rect 77988 77808 78056 77864
rect 78112 77808 78180 77864
rect 78236 77808 78304 77864
rect 78360 77808 78428 77864
rect 78484 77808 78552 77864
rect 78608 77808 94294 77864
rect 94350 77808 94418 77864
rect 94474 77808 104294 77864
rect 104350 77808 104418 77864
rect 104474 77808 124294 77864
rect 124350 77808 124418 77864
rect 124474 77808 134294 77864
rect 134350 77808 134418 77864
rect 134474 77808 144294 77864
rect 144350 77808 144418 77864
rect 144474 77808 154294 77864
rect 154350 77808 154418 77864
rect 154474 77808 164294 77864
rect 164350 77808 164418 77864
rect 164474 77808 174294 77864
rect 174350 77808 174418 77864
rect 174474 77808 184294 77864
rect 184350 77808 184418 77864
rect 184474 77808 194294 77864
rect 194350 77808 194418 77864
rect 194474 77808 204294 77864
rect 204350 77808 204418 77864
rect 204474 77808 214294 77864
rect 214350 77808 214418 77864
rect 214474 77808 224294 77864
rect 224350 77808 224418 77864
rect 224474 77808 234294 77864
rect 234350 77808 234418 77864
rect 234474 77808 244294 77864
rect 244350 77808 244418 77864
rect 244474 77808 254294 77864
rect 254350 77808 254418 77864
rect 254474 77808 264294 77864
rect 264350 77808 264418 77864
rect 264474 77808 294294 77864
rect 294350 77808 294418 77864
rect 294474 77808 304294 77864
rect 304350 77808 304418 77864
rect 304474 77808 314294 77864
rect 314350 77808 314418 77864
rect 314474 77808 324294 77864
rect 324350 77808 324418 77864
rect 324474 77808 334294 77864
rect 334350 77808 334418 77864
rect 334474 77808 344294 77864
rect 344350 77808 344418 77864
rect 344474 77808 354294 77864
rect 354350 77808 354418 77864
rect 354474 77808 364294 77864
rect 364350 77808 364418 77864
rect 364474 77808 374294 77864
rect 374350 77808 374418 77864
rect 374474 77808 384294 77864
rect 384350 77808 384418 77864
rect 384474 77808 394294 77864
rect 394350 77808 394418 77864
rect 394474 77808 404294 77864
rect 404350 77808 404418 77864
rect 404474 77808 414294 77864
rect 414350 77808 414418 77864
rect 414474 77808 424294 77864
rect 424350 77808 424418 77864
rect 424474 77808 434294 77864
rect 434350 77808 434418 77864
rect 434474 77808 444294 77864
rect 444350 77808 444418 77864
rect 444474 77808 454294 77864
rect 454350 77808 454418 77864
rect 454474 77808 464294 77864
rect 464350 77808 464418 77864
rect 464474 77808 474294 77864
rect 474350 77808 474418 77864
rect 474474 77808 484294 77864
rect 484350 77808 484418 77864
rect 484474 77808 494294 77864
rect 494350 77808 494418 77864
rect 494474 77808 504294 77864
rect 504350 77808 504418 77864
rect 504474 77808 514294 77864
rect 514350 77808 514418 77864
rect 514474 77808 524294 77864
rect 524350 77808 524418 77864
rect 524474 77808 534294 77864
rect 534350 77808 534418 77864
rect 534474 77808 544294 77864
rect 544350 77808 544418 77864
rect 544474 77808 554294 77864
rect 554350 77808 554418 77864
rect 554474 77808 592370 77864
rect 592426 77808 592494 77864
rect 592550 77808 592618 77864
rect 592674 77808 592742 77864
rect 592798 77808 592866 77864
rect 592922 77808 592990 77864
rect 593046 77808 593114 77864
rect 593170 77808 624727 77864
rect 624783 77808 624851 77864
rect 624907 77808 632667 77864
rect 632723 77808 632791 77864
rect 632847 77808 640607 77864
rect 640663 77808 640731 77864
rect 640787 77808 648547 77864
rect 648603 77808 648671 77864
rect 648727 77808 657330 77864
rect 657386 77808 657454 77864
rect 657510 77808 657578 77864
rect 657634 77808 657702 77864
rect 657758 77808 657826 77864
rect 657882 77808 657950 77864
rect 658006 77808 658074 77864
rect 658130 77808 658198 77864
rect 658254 77808 658322 77864
rect 658378 77808 658446 77864
rect 658502 77808 658570 77864
rect 658626 77808 658694 77864
rect 658750 77808 658818 77864
rect 658874 77808 658942 77864
rect 658998 77808 659066 77864
rect 659122 77808 659810 77864
rect 659866 77808 659934 77864
rect 659990 77808 660058 77864
rect 660114 77808 660182 77864
rect 660238 77808 660306 77864
rect 660362 77808 660430 77864
rect 660486 77808 660554 77864
rect 660610 77808 660678 77864
rect 660734 77808 660802 77864
rect 660858 77808 660926 77864
rect 660982 77808 661050 77864
rect 661106 77808 661174 77864
rect 661230 77808 661298 77864
rect 661354 77808 661422 77864
rect 661478 77808 661546 77864
rect 661602 77808 661670 77864
rect 661726 77808 662180 77864
rect 662236 77808 662304 77864
rect 662360 77808 662428 77864
rect 662484 77808 662552 77864
rect 662608 77808 662676 77864
rect 662732 77808 662800 77864
rect 662856 77808 662924 77864
rect 662980 77808 663048 77864
rect 663104 77808 663172 77864
rect 663228 77808 663296 77864
rect 663352 77808 663420 77864
rect 663476 77808 663544 77864
rect 663600 77808 663668 77864
rect 663724 77808 663792 77864
rect 663848 77808 663916 77864
rect 663972 77808 664040 77864
rect 664096 77808 664886 77864
rect 664942 77808 665010 77864
rect 665066 77808 665134 77864
rect 665190 77808 665258 77864
rect 665314 77808 665382 77864
rect 665438 77808 665506 77864
rect 665562 77808 665630 77864
rect 665686 77808 665754 77864
rect 665810 77808 665878 77864
rect 665934 77808 666002 77864
rect 666058 77808 666126 77864
rect 666182 77808 666250 77864
rect 666306 77808 666374 77864
rect 666430 77808 666498 77864
rect 666554 77808 666622 77864
rect 666678 77808 666746 77864
rect 666802 77808 667256 77864
rect 667312 77808 667380 77864
rect 667436 77808 667504 77864
rect 667560 77808 667628 77864
rect 667684 77808 667752 77864
rect 667808 77808 667876 77864
rect 667932 77808 668000 77864
rect 668056 77808 668124 77864
rect 668180 77808 668248 77864
rect 668304 77808 668372 77864
rect 668428 77808 668496 77864
rect 668552 77808 668620 77864
rect 668676 77808 668744 77864
rect 668800 77808 668868 77864
rect 668924 77808 668992 77864
rect 669048 77808 669116 77864
rect 669172 77808 669860 77864
rect 669916 77808 669984 77864
rect 670040 77808 670108 77864
rect 670164 77808 670232 77864
rect 670288 77808 670356 77864
rect 670412 77808 670480 77864
rect 670536 77808 670604 77864
rect 670660 77808 670728 77864
rect 670784 77808 670852 77864
rect 670908 77808 670976 77864
rect 671032 77808 671100 77864
rect 671156 77808 671224 77864
rect 671280 77808 671348 77864
rect 671404 77808 671472 77864
rect 671528 77808 671596 77864
rect 671652 77808 699452 77864
rect 699508 77808 699576 77864
rect 699632 77808 699700 77864
rect 699756 77808 699824 77864
rect 699880 77808 699948 77864
rect 700004 77808 700072 77864
rect 700128 77808 700196 77864
rect 700252 77808 700322 77864
rect 77678 77678 700322 77808
rect 699322 75423 701085 75490
rect 699322 75367 699497 75423
rect 699553 75367 699797 75423
rect 699853 75367 700097 75423
rect 700153 75367 701085 75423
rect 699322 75290 701085 75367
rect 701565 75090 701885 75490
rect 697922 75008 701885 75090
rect 697922 74952 698060 75008
rect 698116 74952 698360 75008
rect 698416 74952 698660 75008
rect 698716 74952 701885 75008
rect 697922 74890 701885 74952
<< end >>
