magic
tech gf180mcuC
magscale 1 10
timestamp 1670739833
use caravel_logo  caravel_logo
timestamp 0
transform 1 0 243800 0 1 800
box -746 93 9893 10266
use caravel_motto  caravel_motto
timestamp 0
transform 1 0 294800 0 1 3400
box 1867530 75278 1885498 77962
use caravel_power_routing  caravel_power_routing
timestamp 0
transform 1 0 0 0 1 0
box 70000 70000 706000 944000
use caravel_core  chip_core
timestamp 0
transform 1 0 71000 0 1 71000
box -800 -900 634800 872800
use copyright_block  copyright_block
timestamp 0
transform 1 0 130000 0 1 1600
box -158 -6016 17950 2312
use open_source  open_source
timestamp 0
transform 1 0 187800 0 1 2400
box 540 2880 14316 8010
use chip_io  padframe
timestamp 0
transform 1 0 0 0 1 0
box 0 0 776000 1014000
use user_id_textblock  user_id_textblock
timestamp 0
transform 1 0 52000 0 1 800
box 960 890 40783 9962
<< properties >>
string FIXED_BBOX 0 0 778000 1020000
<< end >>
