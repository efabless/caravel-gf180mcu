magic
tech gf180mcuD
magscale 1 10
timestamp 1655304105
<< pwell >>
rect -1066 -432 1066 432
<< mvnmos >>
rect -802 -224 -662 176
rect -558 -224 -418 176
rect -314 -224 -174 176
rect -70 -224 70 176
rect 174 -224 314 176
rect 418 -224 558 176
rect 662 -224 802 176
<< mvndiff >>
rect -890 163 -802 176
rect -890 -211 -877 163
rect -831 -211 -802 163
rect -890 -224 -802 -211
rect -662 163 -558 176
rect -662 -211 -633 163
rect -587 -211 -558 163
rect -662 -224 -558 -211
rect -418 163 -314 176
rect -418 -211 -389 163
rect -343 -211 -314 163
rect -418 -224 -314 -211
rect -174 163 -70 176
rect -174 -211 -145 163
rect -99 -211 -70 163
rect -174 -224 -70 -211
rect 70 163 174 176
rect 70 -211 99 163
rect 145 -211 174 163
rect 70 -224 174 -211
rect 314 163 418 176
rect 314 -211 343 163
rect 389 -211 418 163
rect 314 -224 418 -211
rect 558 163 662 176
rect 558 -211 587 163
rect 633 -211 662 163
rect 558 -224 662 -211
rect 802 163 890 176
rect 802 -211 831 163
rect 877 -211 890 163
rect 802 -224 890 -211
<< mvndiffc >>
rect -877 -211 -831 163
rect -633 -211 -587 163
rect -389 -211 -343 163
rect -145 -211 -99 163
rect 99 -211 145 163
rect 343 -211 389 163
rect 587 -211 633 163
rect 831 -211 877 163
<< mvpsubdiff >>
rect -1034 328 1034 400
rect -1034 284 -962 328
rect -1034 -284 -1021 284
rect -975 -284 -962 284
rect 962 284 1034 328
rect -1034 -328 -962 -284
rect 962 -284 975 284
rect 1021 -284 1034 284
rect 962 -328 1034 -284
rect -1034 -341 1034 -328
rect -1034 -387 -918 -341
rect 918 -387 1034 -341
rect -1034 -400 1034 -387
<< mvpsubdiffcont >>
rect -1021 -284 -975 284
rect 975 -284 1021 284
rect -918 -387 918 -341
<< polysilicon >>
rect -802 255 -662 268
rect -802 209 -789 255
rect -675 209 -662 255
rect -802 176 -662 209
rect -558 255 -418 268
rect -558 209 -545 255
rect -431 209 -418 255
rect -558 176 -418 209
rect -314 255 -174 268
rect -314 209 -301 255
rect -187 209 -174 255
rect -314 176 -174 209
rect -70 255 70 268
rect -70 209 -57 255
rect 57 209 70 255
rect -70 176 70 209
rect 174 255 314 268
rect 174 209 187 255
rect 301 209 314 255
rect 174 176 314 209
rect 418 255 558 268
rect 418 209 431 255
rect 545 209 558 255
rect 418 176 558 209
rect 662 255 802 268
rect 662 209 675 255
rect 789 209 802 255
rect 662 176 802 209
rect -802 -268 -662 -224
rect -558 -268 -418 -224
rect -314 -268 -174 -224
rect -70 -268 70 -224
rect 174 -268 314 -224
rect 418 -268 558 -224
rect 662 -268 802 -224
<< polycontact >>
rect -789 209 -675 255
rect -545 209 -431 255
rect -301 209 -187 255
rect -57 209 57 255
rect 187 209 301 255
rect 431 209 545 255
rect 675 209 789 255
<< metal1 >>
rect -1021 341 1021 387
rect -1021 284 -975 341
rect 975 284 1021 341
rect -800 209 -789 255
rect -675 209 -664 255
rect -556 209 -545 255
rect -431 209 -420 255
rect -312 209 -301 255
rect -187 209 -176 255
rect -68 209 -57 255
rect 57 209 68 255
rect 176 209 187 255
rect 301 209 312 255
rect 420 209 431 255
rect 545 209 556 255
rect 664 209 675 255
rect 789 209 800 255
rect -877 163 -831 174
rect -877 -222 -831 -211
rect -633 163 -587 174
rect -633 -222 -587 -211
rect -389 163 -343 174
rect -389 -222 -343 -211
rect -145 163 -99 174
rect -145 -222 -99 -211
rect 99 163 145 174
rect 99 -222 145 -211
rect 343 163 389 174
rect 343 -222 389 -211
rect 587 163 633 174
rect 587 -222 633 -211
rect 831 163 877 174
rect 831 -222 877 -211
rect -1021 -341 -975 -284
rect 975 -341 1021 -284
rect -1021 -387 -918 -341
rect 918 -387 1021 -341
<< properties >>
string FIXED_BBOX -998 -364 998 364
string gencell nmos_6p0
string library gf180mcu
string parameters w 2 l 0.7 m 1 nf 7 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.6 wmin 0.3 full_metal 1 compatible {nmos_3p3 nmos_6p0 nmos_6p0_nat}
<< end >>
