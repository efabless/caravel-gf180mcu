magic
tech gf180mcuC
magscale 1 10
timestamp 1671334272
<< mimcap >>
rect -1100 920 900 1000
rect -1100 -920 -1020 920
rect 820 -920 900 920
rect -1100 -1000 900 -920
<< mimcapcontact >>
rect -1020 -920 820 920
<< metal4 >>
rect -1220 1031 1220 1120
rect -1220 1000 1070 1031
rect -1220 -1000 -1100 1000
rect 900 -1000 1070 1000
rect -1220 -1031 1070 -1000
rect 1158 -1031 1220 1031
rect -1220 -1120 1220 -1031
<< via4 >>
rect 1070 -1031 1158 1031
<< metal5 >>
rect 1008 1031 1220 1094
rect -1100 920 900 1000
rect -1100 -920 -1020 920
rect 820 -920 900 920
rect -1100 -1000 900 -920
rect 1008 -1031 1070 1031
rect 1158 -1031 1220 1031
rect 1008 -1094 1220 -1031
<< properties >>
string FIXED_BBOX -1180 -1080 980 1080
string MASKHINTS_CAP_LENGTH -1100 -1000 900 -900
string gencell mim_2p0fF
string library gf180mcu
string parameters w 10.00 l 10.00 val 3.3k carea 25.00 cperi 20.00 nx 1 ny 1 dummy 0 square 0 lmin 5.00 wmin 5.00 lmax 100.0 wmax 100.0 dc 0 bconnect 1 tconnect 1
<< end >>
