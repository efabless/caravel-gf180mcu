magic
tech gf180mcuC
magscale 1 10
timestamp 1670255469
use caravel_power_routing  caravel_power_routing
timestamp 0
transform 1 0 0 0 1 0
box 0 0 1 1
use caravel_core  chip_core
timestamp 0
transform 1 0 71000 0 1 71000
box -800 -844 634800 872800
use chip_io  padframe
timestamp 0
transform 1 0 0 0 1 0
box 0 0 776000 1014000
<< properties >>
string FIXED_BBOX 0 0 778000 1020000
<< end >>
