VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO spare_logic_block
  CLASS BLOCK ;
  FOREIGN spare_logic_block ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 70.000 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 12.775 7.540 14.375 59.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 28.725 7.540 30.325 59.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 44.675 7.540 46.275 59.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 60.625 7.540 62.225 59.100 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 5.300 13.830 69.180 15.430 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 5.300 27.410 69.180 29.010 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 5.300 40.990 69.180 42.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 5.300 54.570 69.180 56.170 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 20.750 7.540 22.350 59.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 36.700 7.540 38.300 59.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 52.650 7.540 54.250 59.100 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 5.300 20.620 69.180 22.220 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 5.300 34.200 69.180 35.800 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 5.300 47.780 69.180 49.380 ;
    END
  END VSS
  PIN spare_xfq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 23.800 4.000 24.360 ;
    END
  END spare_xfq[0]
  PIN spare_xfq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 66.920 0.000 67.480 4.000 ;
    END
  END spare_xfq[1]
  PIN spare_xi[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 33.320 66.000 33.880 70.000 ;
    END
  END spare_xi[0]
  PIN spare_xi[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 26.600 0.000 27.160 4.000 ;
    END
  END spare_xi[1]
  PIN spare_xi[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 71.000 10.360 75.000 10.920 ;
    END
  END spare_xi[2]
  PIN spare_xi[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 50.680 4.000 51.240 ;
    END
  END spare_xi[3]
  PIN spare_xib
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 71.000 3.640 75.000 4.200 ;
    END
  END spare_xib
  PIN spare_xmx[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 73.640 0.000 74.200 4.000 ;
    END
  END spare_xmx[0]
  PIN spare_xmx[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 71.000 50.680 75.000 51.240 ;
    END
  END spare_xmx[1]
  PIN spare_xna[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -0.280 66.000 0.280 70.000 ;
    END
  END spare_xna[0]
  PIN spare_xna[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 40.040 0.000 40.600 4.000 ;
    END
  END spare_xna[1]
  PIN spare_xno[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 17.080 4.000 17.640 ;
    END
  END spare_xno[0]
  PIN spare_xno[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 53.480 0.000 54.040 4.000 ;
    END
  END spare_xno[1]
  PIN spare_xz[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 71.000 57.400 75.000 57.960 ;
    END
  END spare_xz[0]
  PIN spare_xz[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 37.240 4.000 37.800 ;
    END
  END spare_xz[10]
  PIN spare_xz[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 13.160 0.000 13.720 4.000 ;
    END
  END spare_xz[11]
  PIN spare_xz[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 66.920 66.000 67.480 70.000 ;
    END
  END spare_xz[12]
  PIN spare_xz[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 46.760 66.000 47.320 70.000 ;
    END
  END spare_xz[13]
  PIN spare_xz[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 71.000 37.240 75.000 37.800 ;
    END
  END spare_xz[14]
  PIN spare_xz[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 60.200 66.000 60.760 70.000 ;
    END
  END spare_xz[15]
  PIN spare_xz[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 10.360 4.000 10.920 ;
    END
  END spare_xz[16]
  PIN spare_xz[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 71.000 64.120 75.000 64.680 ;
    END
  END spare_xz[17]
  PIN spare_xz[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 13.160 66.000 13.720 70.000 ;
    END
  END spare_xz[18]
  PIN spare_xz[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 -0.280 4.000 0.280 ;
    END
  END spare_xz[19]
  PIN spare_xz[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 40.040 66.000 40.600 70.000 ;
    END
  END spare_xz[1]
  PIN spare_xz[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 71.000 43.960 75.000 44.520 ;
    END
  END spare_xz[20]
  PIN spare_xz[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 6.440 66.000 7.000 70.000 ;
    END
  END spare_xz[21]
  PIN spare_xz[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3.640 4.000 4.200 ;
    END
  END spare_xz[22]
  PIN spare_xz[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 60.200 0.000 60.760 4.000 ;
    END
  END spare_xz[23]
  PIN spare_xz[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 53.480 66.000 54.040 70.000 ;
    END
  END spare_xz[24]
  PIN spare_xz[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 71.000 17.080 75.000 17.640 ;
    END
  END spare_xz[25]
  PIN spare_xz[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 6.440 0.000 7.000 4.000 ;
    END
  END spare_xz[26]
  PIN spare_xz[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 19.880 0.000 20.440 4.000 ;
    END
  END spare_xz[27]
  PIN spare_xz[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 57.400 4.000 57.960 ;
    END
  END spare_xz[28]
  PIN spare_xz[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 71.000 23.800 75.000 24.360 ;
    END
  END spare_xz[29]
  PIN spare_xz[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 33.320 0.000 33.880 4.000 ;
    END
  END spare_xz[2]
  PIN spare_xz[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 43.960 4.000 44.520 ;
    END
  END spare_xz[30]
  PIN spare_xz[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 73.640 66.000 74.200 70.000 ;
    END
  END spare_xz[3]
  PIN spare_xz[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 19.880 66.000 20.440 70.000 ;
    END
  END spare_xz[4]
  PIN spare_xz[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 26.600 66.000 27.160 70.000 ;
    END
  END spare_xz[5]
  PIN spare_xz[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 46.760 0.000 47.320 4.000 ;
    END
  END spare_xz[6]
  PIN spare_xz[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 30.520 4.000 31.080 ;
    END
  END spare_xz[7]
  PIN spare_xz[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 64.120 4.000 64.680 ;
    END
  END spare_xz[8]
  PIN spare_xz[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 71.000 30.520 75.000 31.080 ;
    END
  END spare_xz[9]
  OBS
      LAYER Metal1 ;
        RECT 5.600 6.590 74.110 64.530 ;
      LAYER Metal2 ;
        RECT -0.140 65.700 0.140 66.000 ;
        RECT 0.580 65.700 6.140 66.780 ;
        RECT 7.300 65.700 12.860 66.780 ;
        RECT 14.020 65.700 19.580 66.780 ;
        RECT 20.740 65.700 26.300 66.780 ;
        RECT 27.460 65.700 33.020 66.780 ;
        RECT 34.180 65.700 39.740 66.780 ;
        RECT 40.900 65.700 46.460 66.780 ;
        RECT 47.620 65.700 53.180 66.780 ;
        RECT 54.340 65.700 59.900 66.780 ;
        RECT 61.060 65.700 66.620 66.780 ;
        RECT 67.780 65.700 73.340 66.780 ;
        RECT -0.140 63.700 74.060 65.700 ;
        RECT 0.000 4.300 74.060 63.700 ;
        RECT 0.000 0.580 6.140 4.300 ;
        RECT 4.300 0.140 6.140 0.580 ;
        RECT 4.000 0.000 6.140 0.140 ;
        RECT 7.300 0.000 12.860 4.300 ;
        RECT 14.020 0.000 19.580 4.300 ;
        RECT 20.740 0.000 26.300 4.300 ;
        RECT 27.460 0.000 33.020 4.300 ;
        RECT 34.180 0.000 39.740 4.300 ;
        RECT 40.900 0.000 46.460 4.300 ;
        RECT 47.620 0.000 53.180 4.300 ;
        RECT 54.340 0.000 59.900 4.300 ;
        RECT 61.060 0.000 66.620 4.300 ;
        RECT 67.780 0.000 73.340 4.300 ;
        RECT 4.000 -0.140 5.740 0.000 ;
      LAYER Metal3 ;
        RECT 4.300 63.820 70.700 64.540 ;
        RECT 0.370 58.260 71.820 63.820 ;
        RECT 4.300 57.100 70.700 58.260 ;
        RECT 0.370 51.540 71.820 57.100 ;
        RECT 4.300 50.380 70.700 51.540 ;
        RECT 0.370 44.820 71.820 50.380 ;
        RECT 4.300 43.660 70.700 44.820 ;
        RECT 0.370 38.100 71.820 43.660 ;
        RECT 4.300 36.940 70.700 38.100 ;
        RECT 0.370 31.380 71.820 36.940 ;
        RECT 4.300 30.220 70.700 31.380 ;
        RECT 0.370 24.660 71.820 30.220 ;
        RECT 4.300 23.500 70.700 24.660 ;
        RECT 0.370 17.940 71.820 23.500 ;
        RECT 4.300 16.780 70.700 17.940 ;
        RECT 0.370 11.220 71.820 16.780 ;
        RECT 4.300 10.060 70.700 11.220 ;
        RECT 0.370 4.500 71.820 10.060 ;
        RECT 4.300 3.780 70.700 4.500 ;
      LAYER Metal1 ;
        RECT 0 0 75 70 ;
      LAYER Metal2 ;
        RECT 2 2 73 68 ;
      LAYER Metal3 ;
        RECT 2 2 73 68 ;
      LAYER Metal3 ;
        RECT 2 2 73 68 ;
      LAYER Metal4 ;
        RECT 15 0 55 75 ;
      LAYER Metal5 ;
        RECT 0 0 70 75 ;
  END
END spare_logic_block
END LIBRARY

