* NGSPICE file created from housekeeping.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_4 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 D RN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_4 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_4 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 D SETN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_3 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_3 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_4 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlya_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlya_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1 D RN CLKN Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_20 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_20 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_4 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffsnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffsnq_2 D SETN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_20 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_20 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_2 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_4 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffnsnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffnsnq_1 D SETN CLKN Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tieh abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tieh Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 D RN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_20 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_20 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlya_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlya_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_4 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_4 A1 A2 B1 B2 ZN VDD VSS
.ends

.subckt housekeeping VDD VSS debug_in debug_mode debug_oeb debug_out irq[0] irq[1]
+ irq[2] mask_rev_in[0] mask_rev_in[10] mask_rev_in[11] mask_rev_in[12] mask_rev_in[13]
+ mask_rev_in[14] mask_rev_in[15] mask_rev_in[16] mask_rev_in[17] mask_rev_in[18]
+ mask_rev_in[19] mask_rev_in[1] mask_rev_in[20] mask_rev_in[21] mask_rev_in[22] mask_rev_in[23]
+ mask_rev_in[24] mask_rev_in[25] mask_rev_in[26] mask_rev_in[27] mask_rev_in[28]
+ mask_rev_in[29] mask_rev_in[2] mask_rev_in[30] mask_rev_in[31] mask_rev_in[3] mask_rev_in[4]
+ mask_rev_in[5] mask_rev_in[6] mask_rev_in[7] mask_rev_in[8] mask_rev_in[9] mgmt_gpio_in[0]
+ mgmt_gpio_in[10] mgmt_gpio_in[11] mgmt_gpio_in[12] mgmt_gpio_in[13] mgmt_gpio_in[14]
+ mgmt_gpio_in[15] mgmt_gpio_in[16] mgmt_gpio_in[17] mgmt_gpio_in[18] mgmt_gpio_in[19]
+ mgmt_gpio_in[1] mgmt_gpio_in[20] mgmt_gpio_in[21] mgmt_gpio_in[22] mgmt_gpio_in[23]
+ mgmt_gpio_in[24] mgmt_gpio_in[25] mgmt_gpio_in[26] mgmt_gpio_in[27] mgmt_gpio_in[28]
+ mgmt_gpio_in[29] mgmt_gpio_in[2] mgmt_gpio_in[30] mgmt_gpio_in[31] mgmt_gpio_in[32]
+ mgmt_gpio_in[33] mgmt_gpio_in[34] mgmt_gpio_in[35] mgmt_gpio_in[36] mgmt_gpio_in[37]
+ mgmt_gpio_in[3] mgmt_gpio_in[4] mgmt_gpio_in[5] mgmt_gpio_in[6] mgmt_gpio_in[7]
+ mgmt_gpio_in[8] mgmt_gpio_in[9] mgmt_gpio_oeb[0] mgmt_gpio_oeb[10] mgmt_gpio_oeb[11]
+ mgmt_gpio_oeb[12] mgmt_gpio_oeb[13] mgmt_gpio_oeb[14] mgmt_gpio_oeb[15] mgmt_gpio_oeb[16]
+ mgmt_gpio_oeb[17] mgmt_gpio_oeb[18] mgmt_gpio_oeb[19] mgmt_gpio_oeb[1] mgmt_gpio_oeb[20]
+ mgmt_gpio_oeb[21] mgmt_gpio_oeb[22] mgmt_gpio_oeb[23] mgmt_gpio_oeb[24] mgmt_gpio_oeb[25]
+ mgmt_gpio_oeb[26] mgmt_gpio_oeb[27] mgmt_gpio_oeb[28] mgmt_gpio_oeb[29] mgmt_gpio_oeb[2]
+ mgmt_gpio_oeb[30] mgmt_gpio_oeb[31] mgmt_gpio_oeb[32] mgmt_gpio_oeb[33] mgmt_gpio_oeb[34]
+ mgmt_gpio_oeb[35] mgmt_gpio_oeb[36] mgmt_gpio_oeb[37] mgmt_gpio_oeb[3] mgmt_gpio_oeb[4]
+ mgmt_gpio_oeb[5] mgmt_gpio_oeb[6] mgmt_gpio_oeb[7] mgmt_gpio_oeb[8] mgmt_gpio_oeb[9]
+ mgmt_gpio_out[0] mgmt_gpio_out[10] mgmt_gpio_out[11] mgmt_gpio_out[12] mgmt_gpio_out[13]
+ mgmt_gpio_out[14] mgmt_gpio_out[15] mgmt_gpio_out[16] mgmt_gpio_out[17] mgmt_gpio_out[18]
+ mgmt_gpio_out[19] mgmt_gpio_out[1] mgmt_gpio_out[20] mgmt_gpio_out[21] mgmt_gpio_out[22]
+ mgmt_gpio_out[23] mgmt_gpio_out[24] mgmt_gpio_out[25] mgmt_gpio_out[26] mgmt_gpio_out[27]
+ mgmt_gpio_out[28] mgmt_gpio_out[29] mgmt_gpio_out[2] mgmt_gpio_out[30] mgmt_gpio_out[31]
+ mgmt_gpio_out[32] mgmt_gpio_out[33] mgmt_gpio_out[34] mgmt_gpio_out[35] mgmt_gpio_out[36]
+ mgmt_gpio_out[37] mgmt_gpio_out[3] mgmt_gpio_out[4] mgmt_gpio_out[5] mgmt_gpio_out[6]
+ mgmt_gpio_out[7] mgmt_gpio_out[8] mgmt_gpio_out[9] pad_flash_clk pad_flash_clk_oe
+ pad_flash_csb pad_flash_csb_oe pad_flash_io0_di pad_flash_io0_do pad_flash_io0_ie
+ pad_flash_io0_oe pad_flash_io1_di pad_flash_io1_do pad_flash_io1_ie pad_flash_io1_oe
+ pll90_sel[0] pll90_sel[1] pll90_sel[2] pll_bypass pll_dco_ena pll_div[0] pll_div[1]
+ pll_div[2] pll_div[3] pll_div[4] pll_ena pll_sel[0] pll_sel[1] pll_sel[2] pll_trim[0]
+ pll_trim[10] pll_trim[11] pll_trim[12] pll_trim[13] pll_trim[14] pll_trim[15] pll_trim[16]
+ pll_trim[17] pll_trim[18] pll_trim[19] pll_trim[1] pll_trim[20] pll_trim[21] pll_trim[22]
+ pll_trim[23] pll_trim[24] pll_trim[25] pll_trim[2] pll_trim[3] pll_trim[4] pll_trim[5]
+ pll_trim[6] pll_trim[7] pll_trim[8] pll_trim[9] porb pwr_ctrl_out qspi_enabled reset
+ ser_rx ser_tx serial_clock serial_data_1 serial_data_2 serial_load serial_resetn
+ spi_csb spi_enabled spi_sck spi_sdi spi_sdo spi_sdoenb spimemio_flash_clk spimemio_flash_csb
+ spimemio_flash_io0_di spimemio_flash_io0_do spimemio_flash_io0_oeb spimemio_flash_io1_di
+ spimemio_flash_io1_do spimemio_flash_io1_oeb spimemio_flash_io2_di spimemio_flash_io2_do
+ spimemio_flash_io2_oeb spimemio_flash_io3_di spimemio_flash_io3_do spimemio_flash_io3_oeb
+ trap uart_enabled user_clock wb_ack_o wb_adr_i[0] wb_adr_i[10] wb_adr_i[11] wb_adr_i[12]
+ wb_adr_i[13] wb_adr_i[14] wb_adr_i[15] wb_adr_i[16] wb_adr_i[17] wb_adr_i[18] wb_adr_i[19]
+ wb_adr_i[1] wb_adr_i[20] wb_adr_i[21] wb_adr_i[22] wb_adr_i[23] wb_adr_i[24] wb_adr_i[25]
+ wb_adr_i[26] wb_adr_i[27] wb_adr_i[28] wb_adr_i[29] wb_adr_i[2] wb_adr_i[30] wb_adr_i[31]
+ wb_adr_i[3] wb_adr_i[4] wb_adr_i[5] wb_adr_i[6] wb_adr_i[7] wb_adr_i[8] wb_adr_i[9]
+ wb_clk_i wb_cyc_i wb_dat_i[0] wb_dat_i[10] wb_dat_i[11] wb_dat_i[12] wb_dat_i[13]
+ wb_dat_i[14] wb_dat_i[15] wb_dat_i[16] wb_dat_i[17] wb_dat_i[18] wb_dat_i[19] wb_dat_i[1]
+ wb_dat_i[20] wb_dat_i[21] wb_dat_i[22] wb_dat_i[23] wb_dat_i[24] wb_dat_i[25] wb_dat_i[26]
+ wb_dat_i[27] wb_dat_i[28] wb_dat_i[29] wb_dat_i[2] wb_dat_i[30] wb_dat_i[31] wb_dat_i[3]
+ wb_dat_i[4] wb_dat_i[5] wb_dat_i[6] wb_dat_i[7] wb_dat_i[8] wb_dat_i[9] wb_dat_o[0]
+ wb_dat_o[10] wb_dat_o[11] wb_dat_o[12] wb_dat_o[13] wb_dat_o[14] wb_dat_o[15] wb_dat_o[16]
+ wb_dat_o[17] wb_dat_o[18] wb_dat_o[19] wb_dat_o[1] wb_dat_o[20] wb_dat_o[21] wb_dat_o[22]
+ wb_dat_o[23] wb_dat_o[24] wb_dat_o[25] wb_dat_o[26] wb_dat_o[27] wb_dat_o[28] wb_dat_o[29]
+ wb_dat_o[2] wb_dat_o[30] wb_dat_o[31] wb_dat_o[3] wb_dat_o[4] wb_dat_o[5] wb_dat_o[6]
+ wb_dat_o[7] wb_dat_o[8] wb_dat_o[9] wb_rstn_i wb_sel_i[0] wb_sel_i[1] wb_sel_i[2]
+ wb_sel_i[3] wb_stb_i wb_we_i
X_05903_ _09624_/A1 _11560_/Q _05906_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10669__A1 _10883_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06883_ _06902_/A2 _11094_/Q _06884_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09671_ _09672_/A2 _11570_/Q _09672_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08622_ _08622_/A1 _08622_/A2 _08624_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05834_ _05647_/I _05668_/I _11033_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_39_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11570__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08553_ _08553_/A1 _08553_/A2 _08647_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05765_ _07006_/A2 _08839_/A2 _05766_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07504_ _07938_/A2 _07513_/I _07505_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08484_ _08484_/A1 _08484_/A2 _08485_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input108_I wb_adr_i[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06727__I _11358_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07435_ input101/Z input100/Z _07437_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05696_ _09549_/A1 _11538_/Q _05697_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05848__A1 _08940_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10841__A1 _10883_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09039__A1 _06867_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11322__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_3_3__f_wb_clk_i_I clkbuf_0_wb_clk_i/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07366_ _07366_/I _11234_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_182_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06317_ _08846_/A1 input61/Z _06318_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07297_ _07297_/I _07844_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__08262__A2 _07609_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09105_ _06855_/Z _09114_/A2 _09105_/B _09106_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06248_ _09449_/A1 _11500_/Q _06252_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input73_I mgmt_gpio_in[9] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09036_ _06863_/Z _09039_/A2 _09036_/B _09037_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06273__A1 _08839_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06179_ _06324_/A1 _11588_/Q _07391_/A1 _11243_/Q _06181_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09211__A1 _09158_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11491__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06025__A1 input68/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06025__B2 input39/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07773__A1 _08592_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09938_ _09938_/A1 _09938_/A2 _09938_/B _09940_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09869_ _09927_/A2 _09946_/A1 _09902_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__11561__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05839__A1 _06266_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11313__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11693_ _11693_/D _11693_/RN input68/Z _11693_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__10832__A1 _10924_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10713_ _11416_/Q _10888_/A1 _11408_/Q _10889_/A1 _10713_/C _10717_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_10644_ _10644_/A1 _10644_/A2 _10644_/A3 _10644_/A4 _10645_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_9_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10575_ _10897_/B1 _11461_/Q _10578_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11444__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09450__A1 _09472_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11342__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10060__A2 _11412_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09202__A1 _09121_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11459__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10899__A1 _10899_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06016__A1 _09144_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11492__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07764__A1 _07722_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11127_ _11127_/D _11683_/CLK _11127_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11058_ _11058_/D _11058_/RN input68/Z _11058_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10009_ _10042_/A2 _10265_/A3 _10135_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__11552__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05550_ _05550_/I _11696_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10823__A1 _10914_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08492__A2 _07564_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11304__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07220_ _07240_/A1 _07220_/A2 _07220_/B _07221_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07151_ _11196_/Q _05927_/Z _07151_/B _07151_/C _07152_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__09441__A1 _09187_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06255__A1 _08825_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06102_ _06102_/A1 _06619_/B _06102_/B _06103_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07082_ _07083_/A2 _11152_/Q _07083_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06033_ _09750_/A1 _11599_/Q _06034_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11000__A1 _11000_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07984_ _07984_/I _08649_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
X_09723_ _09723_/I _11586_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06935_ _06837_/Z _06938_/A2 _06935_/B _06936_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09654_ _09121_/I _09672_/A2 _09654_/B _09655_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06866_ _06866_/I _11085_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11543__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08605_ _08603_/Z _07844_/B _08605_/B _08606_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05817_ _06217_/I _08839_/A2 _05818_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11215__CLK _11672_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09585_ _09154_/Z _09597_/A2 _09585_/B _09586_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_06797_ _06797_/I _09121_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_08536_ _08536_/I _08629_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05748_ _06394_/A1 input10/Z _05749_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10814__A1 _10906_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08467_ split8/Z _07722_/I _08467_/B _08468_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05679_ _05732_/I _05669_/I _05803_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_23_464 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08398_ _08398_/A1 _08397_/Z _11255_/Q _07297_/I _08399_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_07418_ _07418_/I _11249_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06494__A1 _06491_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11365__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07349_ _07349_/A1 _06904_/Z _07354_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09432__A1 _09125_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06192__I _06192_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output277_I _11076_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10042__A2 _10042_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10360_ _10360_/A1 _11142_/Q _10362_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_151_336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10291_ _11514_/Q _10369_/A2 _10369_/B1 _11506_/Q _10294_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_128_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09019_ _09019_/I _11363_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09735__A2 _11590_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09499__A1 _09499_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11534__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08171__A1 _08490_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09671__A1 _09672_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10805__B2 _11466_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10281__A2 _10359_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11676_ _11676_/D input162/Z _06687_/A2 _11676_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10627_ _10627_/A1 _10627_/A2 _10627_/A3 _10627_/A4 _10645_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__09974__A2 _10030_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10558_ _10558_/A1 _10924_/A1 _10558_/B _10560_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10033__A2 _10351_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07985__A1 _08355_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06788__A2 _05633_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10489_ _11611_/Q _10915_/A1 _11571_/Q _10911_/A1 _10489_/C _10492_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__07737__A1 _07885_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11238__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06720_ _06786_/A1 _06753_/A1 _06720_/B _06721_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08162__A1 _08162_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06651_ input80/Z input82/Z _06652_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05602_ input58/Z _05515_/I _05603_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06712__A2 input68/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06582_ input99/Z input98/Z _06583_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09370_ _09370_/I _11473_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11388__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08321_ _08321_/I _08593_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09662__A1 _09672_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05533_ _05539_/A1 _05533_/A2 _05537_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08252_ _08281_/A1 _07885_/I _08528_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07203_ _11315_/Q _05924_/Z _07203_/B _07205_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_158_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08183_ _08183_/A1 _08183_/A2 _08189_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06228__A1 _07412_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07134_ _11168_/Q _07137_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_9_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_07065_ _07065_/I _11147_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xoutput231 _11097_/Q mgmt_gpio_out[28] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput220 _11166_/Q mgmt_gpio_out[18] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput253 _06721_/Z pad_flash_io0_do VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput242 _11184_/Q mgmt_gpio_out[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_06016_ _09144_/A1 _11407_/Q _06018_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07728__A1 _07593_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput275 _11074_/Q pll_trim[11] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput286 _11289_/Q pll_trim[21] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput264 _11273_/Q pll_div[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput297 _11071_/Q pll_trim[8] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_59_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07967_ _08449_/B _08609_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input36_I mgmt_gpio_in[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06400__A1 _08839_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09706_ _09722_/A2 _11581_/Q _09707_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06918_ _06918_/I _11104_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07898_ _07685_/I _07680_/I _07899_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__08153__A1 _08161_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09637_ _09647_/A2 _11559_/Q _09638_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06164__B1 _11445_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07900__A1 split21/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06849_ _06847_/Z _06869_/A2 _06849_/B _06850_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09568_ _09572_/A2 _11537_/Q _09569_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08519_ _08519_/A1 _08519_/A2 _08519_/B _08520_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_11530_ _11530_/D _11686_/RN _06705_/Z _11530_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__08616__B _08616_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09499_ _09499_/A1 _09015_/Z _09522_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__09653__A1 _09672_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11461_ _11461_/D _11686_/RN _06705_/Z _11461_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__05690__A2 _05805_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10412_ _10412_/A1 _10412_/A2 _10422_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11392_ _11392_/D _11686_/RN _06705_/Z _11392_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__10015__A2 _11419_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10343_ _10343_/A1 _10382_/A2 _10343_/B _10343_/C _10345_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_10274_ _10353_/A1 _11370_/Q _10276_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07195__A2 _05925_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09961__I _09961_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11530__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08144__A1 split7/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05902__B1 _11544_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09644__A1 _09241_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11680__CLK _06687_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11659_ _11659_/D input76/Z _11663_/CLK _11659_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__11060__CLK input68/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08870_ _07431_/Z _08888_/A2 _08870_/B _08871_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07821_ _07821_/I _08600_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__06933__A2 _06904_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08135__A1 _08434_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07752_ _07752_/I _08242_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__11275__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07683_ _08285_/B _08285_/A2 _07684_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06703_ _11683_/Q _11023_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08686__A2 _08686_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09883__A1 _09876_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06634_ input77/Z input93/Z _06635_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09422_ _09270_/Z _09422_/A2 _09422_/B _09423_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09353_ _09372_/A2 _11468_/Q _09354_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09635__A1 _09154_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08304_ _08580_/A2 _08345_/A2 _08304_/B _08498_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06565_ _11640_/Q _10425_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__08438__A2 split8/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06735__I _11518_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06496_ _06496_/A1 _06496_/A2 _11062_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05516_ _06466_/B _06610_/A3 _05517_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09284_ _09297_/A2 _11446_/Q _09285_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_176_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08235_ _08235_/A1 _08235_/A2 _08236_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08166_ _08202_/A1 _07535_/I _08467_/B _08174_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_07117_ _07117_/A1 _07151_/B _07117_/B _07118_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11403__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08097_ _08106_/A1 _08169_/A2 _08098_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07566__I _07566_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07048_ _08786_/A1 _06217_/Z _06871_/Z _07053_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__11553__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10705__B1 _11616_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08999_ _08999_/I _11357_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08677__A2 _08677_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10961_ _11221_/Q _11025_/A2 _11028_/A1 _08493_/B _10965_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06137__B1 _05925_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06688__A1 _11304_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10484__A2 _10427_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10892_ _10892_/A1 _11237_/Q _10893_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08429__A2 _08562_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09626__A1 _09116_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11513_ _11513_/D _11686_/RN _06705_/Z _11513_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_11444_ _11444_/D _11686_/RN _06705_/Z _11444_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__06860__A1 _06869_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11083__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11375_ _11375_/D _11686_/RN _06705_/Z _11375_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10326_ _11228_/Q _10365_/A2 _10365_/B1 _11232_/Q _10329_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_10257_ _10378_/A1 _11553_/Q _10259_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08365__A1 split8/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10188_ _10188_/A1 _10188_/A2 _10189_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10172__A1 _11447_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10475__A2 _10406_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06679__A1 input1/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06350_ _06350_/A1 _06350_/A2 _06350_/A3 _06350_/A4 _06392_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__10227__A2 _11328_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09093__A2 _09114_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11426__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06281_ _06281_/A1 _06281_/A2 _06281_/A3 _06303_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_08020_ _08020_/I _08021_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11576__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09971_ _10007_/A1 _09899_/I _09972_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_6_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08922_ _08938_/A2 _11333_/Q _08923_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07159__A2 _09116_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08853_ _08863_/A2 _11311_/Q _08854_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06906__A2 _11101_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07804_ _08592_/A2 _08329_/B _08596_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input138_I wb_dat_i[17] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08784_ _06867_/Z _08784_/A2 _08784_/B _08785_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05996_ _06396_/A1 input30/Z _05998_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07735_ _07989_/A1 _07994_/A1 _07828_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08659__A2 _08696_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07666_ _08300_/A2 _08045_/A3 _07674_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09405_ _09405_/I _11484_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06617_ _06617_/I _11221_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07597_ _08262_/B _07609_/I _07600_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10218__A2 _10377_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09336_ _09336_/I _11462_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06548_ _11089_/Q _09946_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09267_ _09272_/A2 _11441_/Q _09268_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08218_ _08126_/I _07722_/I _08218_/B _08696_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06479_ _11064_/Q _05515_/I _06479_/B _06479_/C _06480_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_09198_ _09220_/A2 _11419_/Q _09199_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08149_ split8/Z _08481_/B _08567_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08595__A1 _07609_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07398__A2 _06238_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11160_ _11160_/D _11160_/RN input68/Z _11160_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10111_ _10111_/A1 _10111_/A2 _10111_/A3 _10124_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_11091_ _11091_/D input76/Z _11656_/CLK _11091_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10042_ _10042_/A1 _10042_/A2 _10043_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xsplit8 split8/I split8/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08898__A2 _08913_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_74 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_3_7__f_wb_clk_i clkbuf_0_wb_clk_i/Z _06687_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10944_ _10934_/I _11670_/Q _10945_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11449__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10875_ _10919_/A1 _11109_/Q _10877_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05884__A2 _09449_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11599__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06833__A1 _05616_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08822__A2 _11302_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11427_ _11427_/D _11686_/RN _06705_/Z _11427_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_11358_ _11358_/D _11686_/RN _06705_/Z _11358_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__06061__A2 input55/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05939__A3 _05939_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10309_ _11654_/Q _10383_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_11289_ _11289_/D input76/Z _06705_/Z _11289_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__10145__A1 _11478_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10145__B2 _10366_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05850_ _11361_/Q _08990_/A1 _11353_/Q _05723_/Z _05850_/C _05860_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
Xrebuffer17 _07540_/A1 _07495_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06364__A3 _06217_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07520_ split5/I _07522_/I _08095_/A2 _07521_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05781_ _05781_/I _09374_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XANTENNA__05572__A1 input58/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07451_ _07506_/I _07451_/A2 _07996_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__05875__A2 _05924_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07382_ _07081_/Z _07382_/A2 _07382_/B _07383_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06402_ _11101_/Q _06905_/A1 _11323_/Q _08890_/A1 _06402_/C _06406_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_06333_ _06333_/A1 _06333_/A2 _06334_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09121_ _09121_/I _09121_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__07077__A1 _05703_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09066__A2 _09015_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10620__A2 _11478_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09052_ _06851_/Z _09064_/A2 _09052_/B _09053_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06264_ _06398_/A2 input21/Z _06265_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06824__A1 _06835_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08003_ _08002_/Z _08003_/A2 _08039_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06195_ _09624_/A1 _11556_/Q _06200_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10384__A1 _10384_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08329__A1 _08332_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09954_ _09954_/A1 _11631_/Q _09973_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_871 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_09885_ _09898_/A1 _09892_/A2 _11634_/Q _09891_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08905_ _08905_/I _11327_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10136__B2 _10359_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10687__A2 _11543_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07001__A1 _06837_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08836_ _08837_/A2 _11306_/Q _08837_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08767_ _08767_/I _11285_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05979_ _05833_/I _05700_/I _10190_/A1 _06518_/A1 _05836_/I _05980_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_08698_ _08698_/A1 _08698_/A2 _08698_/A3 _08699_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_07718_ _07718_/A1 _07716_/Z _07718_/A3 _07719_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_07649_ _07694_/A1 _07649_/A2 _08537_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10660_ _10910_/A1 _11567_/Q _10663_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09319_ _09241_/Z _09322_/A2 _09319_/B _09320_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_15_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10072__B1 _10369_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10591_ _10914_/B1 _11605_/Q _10593_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06815__A1 _11000_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11212_ _11212_/D _11656_/CLK _11212_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10375__A1 _10375_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11121__CLK _11672_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11143_ _11143_/D _11686_/RN _06705_/Z _11143_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__07240__A1 _07240_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput120 wb_adr_i[30] input120/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06594__A3 input167/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10127__A1 _10092_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11074_ _11074_/D _11686_/RN _06705_/Z _11074_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
Xinput153 wb_dat_i[30] input153/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput131 wb_dat_i[10] input131/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput142 wb_dat_i[20] input142/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10678__A2 _10897_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10025_ _10025_/A1 _09887_/I _10359_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xinput164 wb_sel_i[1] input164/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07543__A2 _07485_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08740__A1 _06855_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11271__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09296__A2 _11450_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10927_ _10927_/A1 _10880_/C _10927_/B _10928_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07846__A3 split16/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10858_ _10904_/A1 _11155_/Q _10863_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_10789_ _10881_/A1 _11662_/Q _10790_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10602__A2 _11541_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06806__A1 _06835_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11095__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10366__A1 _10366_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09220__A2 _09220_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10118__A1 _10374_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06951_ _06941_/I _11114_/Q _06952_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11614__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09670_ _09670_/I _11569_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05902_ _11552_/Q _09599_/A1 _11544_/Q _09574_/A1 _05902_/C _05906_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_140_297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06882_ _06882_/I _11093_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08621_ _08621_/A1 _08621_/A2 _08621_/A3 _08622_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08731__A1 _07431_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05833_ _05833_/I _08839_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_3
X_08552_ _08380_/B _08692_/A2 _08552_/B _08552_/C _08553_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__09287__A2 _11447_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05764_ _05764_/I _09091_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
X_07503_ split16/I _07938_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08483_ _08483_/A1 _08483_/A2 _08484_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07298__A1 _07844_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05695_ _05687_/I _05726_/I _09549_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_07434_ _07434_/I _11253_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09039__A2 _09039_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10841__A2 _11119_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07365_ _07076_/Z _07368_/A2 _07365_/B _07366_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06316_ _07201_/A1 input52/Z _06318_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07296_ _11016_/A1 _07296_/A2 _07297_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_09104_ _09114_/A2 _11391_/Q _09105_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06247_ _09424_/A1 _11492_/Q _06252_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09035_ _09039_/A2 _11369_/Q _09036_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06273__A2 _08839_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11144__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input66_I mgmt_gpio_in[37] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06178_ _05941_/I _05636_/I _07391_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09211__A2 _09220_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10357__A1 _10357_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06025__A2 _05924_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07222__A1 _05924_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10109__A1 _10366_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07773__A2 _08315_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09937_ _09937_/I _11641_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08970__A1 _07431_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11294__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09868_ _09868_/A1 _11630_/Q _09868_/A3 _09868_/B _11630_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XTAP_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_09799_ _09799_/I _11610_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08819_ _08820_/A2 _06266_/I _08820_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output222_I _06671_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09278__A2 _11444_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07289__A1 _07290_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10712_ _10712_/A1 _10712_/A2 _10713_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11692_ _11692_/D _11692_/RN input68/Z _11692_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__10832__A2 _11330_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10643_ _10643_/I _10644_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_42_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10574_ _10897_/A2 _11453_/Q _10578_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10596__A1 _10902_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09450__A2 _11499_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09202__A2 _09220_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10899__A2 _11253_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11637__CLK _11658_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07764__A2 _07761_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11126_ _11126_/D _11683_/CLK _11126_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07516__A2 _07614_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11057_ _11057_/D _11057_/RN input68/Z _11057_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__10520__A1 _10913_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05527__A1 _06610_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10008_ _10014_/A1 _09878_/I _10363_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_07150_ _05927_/Z _09270_/I _07151_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06563__I _06563_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11167__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09441__A2 _09447_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07081_ _09121_/I _07081_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__10587__A1 _10913_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06255__A2 _06238_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06101_ _11265_/Q _05969_/I _06101_/B _06619_/B _06102_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06032_ _06324_/A1 _11591_/Q _06034_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10339__A1 _10378_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11000__A2 _10966_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07204__A1 _07240_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07755__A2 _08490_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09722_ _09270_/Z _09722_/A2 _09722_/B _09723_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07983_ _07983_/A1 _07983_/A2 _07987_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11240__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08704__A1 _05703_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06934_ _06938_/A2 _11109_/Q _06935_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09653_ _09672_/A2 _11564_/Q _09654_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06865_ _06863_/Z _06869_/A2 _06865_/B _06866_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10511__A1 _10514_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09584_ _09597_/A2 _11542_/Q _09585_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06738__I _11590_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08604_ _07844_/B _11257_/Q _08605_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05816_ _05816_/I _09299_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_82_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input120_I wb_adr_i[30] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_06796_ _11691_/Q _05633_/B _06796_/B _06797_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06191__A1 _07092_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08535_ _08535_/A1 _08535_/A2 _08535_/A3 _08536_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05747_ _05747_/I _06394_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_23_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10814__A2 _11546_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05678_ _09775_/A1 _11610_/Q _05678_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08466_ _08466_/A1 _08466_/A2 _08570_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08397_ _08397_/A1 _08460_/B _08397_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_07417_ _07081_/Z _07417_/A2 _07417_/B _07418_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09968__B1 _11515_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07348_ _07348_/I _11229_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11689__CLKN input68/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09432__A2 _09447_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07279_ _07279_/I _11200_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10290_ _10290_/A1 _10290_/A2 _10290_/A3 _10303_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_output172_I _06748_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09018_ _07426_/Z _09039_/A2 _09018_/B _09019_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11231__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05757__A1 _06839_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09499__A2 _09015_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06182__A1 _06192_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_split21_I split21/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10805__A2 _10897_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11675_ _11675_/D input162/Z _06687_/A2 _11675_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__11298__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10626_ _11454_/Q _10897_/A2 _10897_/B1 _11462_/Q _10627_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_127_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10569__A1 _10887_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10557_ _10548_/Z _10924_/A1 _10557_/A3 _10558_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_10488_ _10916_/A1 _11619_/Q _10489_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__05996__A1 _06396_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11470__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07737__A2 _08339_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08934__A1 _08938_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11222__RN input162/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10741__A1 _10919_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11109_ _11109_/D _11686_/RN _06705_/Z _11109_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__08162__A2 _08167_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06650_ _06650_/A1 _11312_/Q _06652_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06173__A1 _05927_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05601_ _11060_/Q _06500_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06581_ input101/Z input100/Z _06583_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09111__A1 _06863_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08320_ _08686_/A2 _07725_/I _08320_/B _08321_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05532_ _05539_/A1 _05532_/A2 _05541_/A2 _05532_/B2 _11700_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_177_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08251_ _08281_/A1 _08251_/A2 _08528_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07202_ _05924_/Z _09116_/I _07203_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08182_ _08182_/I _08183_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_118_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07133_ _07133_/I _11167_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07064_ _06837_/Z _07067_/A2 _07064_/B _07065_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput210 _10613_/A2 mgmt_gpio_oeb[9] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput232 _11098_/Q mgmt_gpio_out[29] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput221 _11167_/Q mgmt_gpio_out[19] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_06015_ _11519_/Q _09499_/A1 _11511_/Q _09474_/A1 _06015_/C _06024_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__09178__A1 _09195_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput243 _11185_/Q mgmt_gpio_out[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA_input168_I wb_we_i VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07728__A2 _08358_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput276 _11075_/Q pll_trim[12] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput254 _06718_/ZN pad_flash_io0_ie VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput265 _11274_/Q pll_div[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__08925__A1 _08938_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10732__A1 _10905_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05739__A1 _08799_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput287 _11290_/Q pll_trim[22] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput298 _11072_/Q pll_trim[9] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_59_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_07966_ _07966_/A1 _07966_/A2 _07971_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06400__A2 _08839_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09705_ _09705_/I _11580_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input29_I mask_rev_in[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06917_ _06843_/Z _06917_/A2 _06917_/B _06918_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07897_ split15/I _08549_/A1 _07903_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09350__A1 _09372_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09636_ _09636_/I _11558_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11443__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10496__B1 _10886_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06848_ _06869_/A2 _11081_/Q _06849_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11332__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09567_ _09567_/I _11536_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05911__A1 _09449_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06779_ _07110_/I _11070_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09498_ _09498_/I _11514_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08518_ _08518_/I _08601_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09102__A1 _06851_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11482__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10799__A1 _10891_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08449_ _08449_/A1 _08010_/I _08449_/B _08450_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_23_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11460_ _11460_/D _11686_/RN _06705_/Z _11460_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_10411_ _10884_/A1 _10903_/A1 _10493_/A1 _10412_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_99_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11391_ _11391_/D _11686_/RN _06705_/Z _11391_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10342_ _10342_/A1 _10342_/A2 _10342_/A3 _10342_/A4 _10343_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__10971__A1 _10966_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10453__I _10453_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09169__A1 _06867_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07719__A2 _08431_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10273_ _11354_/Q _10351_/A2 _11346_/Q _10351_/B2 _10273_/C _10286_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__08916__A1 _08938_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11204__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10723__A1 _10896_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09341__A1 _09187_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05902__B2 _09574_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09644__A2 _09647_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_71 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11658_ _11658_/D input76/Z _11658_/CLK _11658_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_11589_ _11589_/D _11686_/RN _06705_/Z _11589_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__07407__A1 _07076_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10609_ _10609_/A1 _10092_/Z _10610_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11205__CLK _11683_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08907__A1 _06859_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10714__A1 _10883_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07820_ _06587_/I _07999_/A2 _07470_/I _07821_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_07751_ _07751_/A1 _07989_/A2 _07752_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10190__A2 _10382_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11355__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09332__A1 _09125_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06702_ _05616_/C input68/Z _06704_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07682_ _07682_/I _08285_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06633_ _06633_/I _06633_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09421_ _09422_/A2 _11490_/Q _09422_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09352_ _09352_/I _11467_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06564_ _10426_/A2 _10501_/A1 _10433_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__09635__A2 _09647_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08303_ _08676_/I _08303_/A2 _08494_/B _08307_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_05515_ _05515_/I _06466_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_06495_ _06500_/A1 _11061_/Q _06495_/A3 _06496_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_100_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09283_ _09283_/I _11445_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08234_ _08483_/A1 _08614_/A2 _08205_/C _08235_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__09399__A1 _09399_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08165_ _08165_/A1 _08165_/A2 _08484_/A1 _08235_/A2 _08174_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__11682__RN input162/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07116_ _11189_/Q _05927_/Z _07151_/B _07116_/C _07117_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__10548__A4 _10548_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10953__A1 _10934_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08096_ _08096_/I _08169_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11434__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07047_ _07047_/I _11142_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10705__A1 _11624_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09571__A1 _09572_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10705__B2 _10915_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08998_ _06847_/Z _09013_/A2 _08998_/B _08999_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07949_ split6/I _08444_/B _08692_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10960_ input166/Z input168/Z _11028_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06137__A1 input58/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_3_6__f_wb_clk_i clkbuf_0_wb_clk_i/Z _11683_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09619_ _09241_/Z _09622_/A2 _09619_/B _09620_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10891_ _10891_/A1 _11241_/Q _10893_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output302_I _06577_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11397__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09626__A2 _09647_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11512_ _11512_/D _11686_/RN _06705_/Z _11512_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_11443_ _11443_/D _11686_/RN _06705_/Z _11443_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__11228__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10944__A1 _10934_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06073__B1 _09674_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11374_ _11374_/D _11686_/RN _06705_/Z _11374_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__11425__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09972__I _09972_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06612__A2 _06619_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11378__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10325_ _10325_/A1 _10325_/A2 _10325_/A3 _10325_/A4 _10343_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_10256_ _11577_/Q _10377_/A1 _10379_/A1 _11561_/Q _10259_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09562__A1 _09572_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07492__I _07492_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10187_ _10377_/A1 _11575_/Q _10377_/B1 _11567_/Q _10188_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_120_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06128__A1 _06128_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10227__A3 _10265_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06280_ _06280_/A1 _06280_/A2 _06280_/A3 _06280_/A4 _06281_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__06300__A1 _05723_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11664__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06064__B1 input38/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10935__A1 _10935_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11416__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09970_ _09970_/I _10007_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08921_ _08921_/I _11332_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09553__A1 _09572_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08356__A2 _08686_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08852_ _08852_/I _11310_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07803_ _08332_/A1 _08329_/B _08226_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08783_ _08784_/A2 _11291_/Q _08784_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05995_ _08799_/A1 _05995_/A2 _06265_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07734_ _07734_/I _07989_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06119__A1 _11325_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07665_ _07669_/I _07938_/A2 _07890_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09404_ _09121_/Z _09422_/A2 _09404_/B _09405_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06616_ _06616_/A1 _10930_/C _07296_/A2 _06749_/I _06617_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_92_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07596_ _07596_/I _08262_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_13_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05893__A3 _05893_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09335_ _09154_/Z _09347_/A2 _09335_/B _09336_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06547_ _11092_/Q _09945_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__10623__B1 _11486_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input96_I user_clock VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06478_ _06480_/A1 _06478_/A2 _06478_/B _06479_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09266_ _09266_/I _11440_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08217_ split7/Z _08232_/A2 _08217_/B _08475_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11655__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09197_ _09197_/A1 _09015_/Z _09220_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__11520__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08044__A1 _08162_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08148_ _08169_/A1 _08148_/A2 _08481_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10926__A1 _10092_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11407__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09792__A1 _09187_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08079_ _08079_/I split7/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XANTENNA__07398__A3 _06838_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10110_ _10367_/A1 _11477_/Q _10111_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11090_ _11090_/D input76/Z _11665_/CLK _11090_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__09544__A1 _09241_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11670__CLK _11683_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10041_ _10041_/I _10355_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_152_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06358__A1 _07419_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10154__A2 _06556_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09847__A2 _11626_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10943_ _10943_/I _11669_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10874_ _10920_/A1 _11103_/Q _10920_/B1 _11105_/Q _10877_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_43_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_101_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08283__A1 split14/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11646__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08822__A3 _06904_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10127__B _10127_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11426_ _11426_/D input76/Z _06705_/Z _11426_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__09783__A1 _09125_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11357_ _11357_/D _11686_/RN _06705_/Z _11357_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_10308_ _10308_/I _11653_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09535__A1 _09154_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11288_ _11288_/D _11686_/RN _06705_/Z _11288_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__11289__SETN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10145__A2 _10367_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10239_ _10356_/A1 _11409_/Q _10241_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xrebuffer18 _07921_/A1 _08649_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05780_ _06238_/I _05805_/A2 _05781_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09838__A2 _11623_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07450_ _07513_/I split16/I _07451_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_06401_ _10343_/A1 _05614_/I _05833_/I _06401_/B _06402_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_07381_ _07382_/A2 _11239_/Q _07382_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11543__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06332_ _05703_/Z _11685_/Q _11033_/A2 _06333_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__07077__A2 _07412_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10605__B1 _10920_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09120_ _09120_/I _11395_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10081__A1 _10379_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09051_ _09064_/A2 _11374_/Q _09052_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08002_ _08002_/A1 _07470_/I _08002_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_06263_ input35/Z _06394_/A1 input12/Z _06393_/A1 _06263_/C _06265_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__06824__A2 _09187_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06194_ _06194_/A1 _06194_/A2 _06194_/A3 _06194_/A4 _06212_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__11693__CLK input68/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10384__A2 _06556_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08329__A2 _08417_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input150_I wb_dat_i[28] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09526__A1 _09116_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09953_ _10265_/A1 _10265_/A3 _10382_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_861 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_09884_ _09884_/A1 _09884_/A2 _09927_/A2 _09892_/A2 _09902_/I _11633_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_08904_ _06855_/Z _08913_/A2 _08904_/B _08905_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10136__A2 _10359_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_894 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_872 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_08835_ _08835_/I _11305_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08766_ _07431_/Z _08784_/A2 _08766_/B _08767_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09829__A2 _11620_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07717_ _08294_/B _08294_/C _08395_/A2 _07718_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_input11_I mask_rev_in[16] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05978_ _11296_/Q _06518_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11073__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08697_ _08697_/A1 _08697_/A2 _08697_/A3 _08697_/A4 _08698_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_53_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08501__A2 _07727_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07648_ _08400_/B _07694_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07579_ _07579_/A1 _07994_/A1 _08204_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_09318_ _09322_/A2 _11457_/Q _09319_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08265__A1 _08400_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10072__A1 _11508_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10590_ _10914_/A1 _11597_/Q _10593_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11628__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06815__A2 _05633_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09249_ _09272_/A2 _11435_/Q _09250_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11211_ _11211_/D _11656_/CLK _11211_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11142_ _11142_/D _11686_/RN _06705_/Z _11142_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xinput110 wb_adr_i[21] _07457_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11073_ _11073_/D _11686_/RN _06705_/Z _11073_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__10461__I _10461_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput154 wb_dat_i[31] input154/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput143 wb_dat_i[21] input143/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput121 wb_adr_i[31] input121/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput132 wb_dat_i[11] input132/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10024_ _10024_/I _10359_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
Xinput165 wb_sel_i[2] input165/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11416__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11566__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10926_ _10092_/Z _11664_/Q _10926_/B _10926_/C _10927_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_10857_ _10903_/A1 _11151_/Q _10863_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_182 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_10788_ _10092_/Z _11661_/Q _10788_/B _10880_/C _10790_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__06806__A2 _09125_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11409_ _11409_/D input76/Z _06705_/Z _11409_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_98_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_435 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06950_ _06950_/I _11113_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06881_ _06837_/Z _06902_/A2 _06881_/B _06882_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05901_ _05901_/A1 _05901_/A2 _05902_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06990__A1 _10950_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11096__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input3_I debug_out VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10304__C _10304_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08620_ _08620_/A1 _08658_/A1 _08624_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05832_ _05832_/I _11270_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05545__A2 _05519_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08551_ _08608_/A1 _08694_/A2 _08559_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05763_ _08791_/A1 _07006_/A2 _05764_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07502_ _07515_/A1 split16/Z _07510_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08495__A1 _08686_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05694_ _05693_/Z _11530_/Q _05697_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08482_ _08482_/A1 _08482_/A2 _08657_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07433_ _07431_/Z _07433_/A2 _07433_/B _07434_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_167_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07364_ _07368_/A2 _11234_/Q _07365_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08247__A1 split21/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09103_ _09103_/I _11390_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06315_ _05660_/Z _11619_/Q _06318_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07295_ _11025_/B _11016_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_3
XANTENNA__10054__B2 _10351_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06246_ _06246_/A1 _06246_/A2 _06246_/A3 _06246_/A4 _06258_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_09034_ _09034_/I _11368_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09747__A1 _09725_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08460__B _08460_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06177_ _08825_/A2 _11033_/A2 _06181_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07222__A2 _09158_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input59_I mgmt_gpio_in[30] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11439__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09936_ _10428_/B1 _09936_/A2 _09936_/B _09937_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08970__A2 _08988_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05784__A2 _11466_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06981__A1 _06974_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09867_ _09867_/A1 _11630_/Q _09868_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11589__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09798_ _09270_/I _09798_/A2 _09798_/B _09799_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08818_ _08818_/I _11300_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_output215_I _06693_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08749_ _08759_/A2 _11280_/Q _08750_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_26_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10293__A1 _10370_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10711_ _10887_/B1 _11432_/Q _10712_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11691_ _11691_/D _11691_/RN input68/Z _11691_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_9_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08238__A1 _08490_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10642_ _10642_/A1 _10642_/A2 _10427_/B _10642_/B1 _10401_/I _10643_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_9_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10573_ _10573_/A1 _10573_/A2 _10584_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08789__A2 _08827_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10596__A2 _11517_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer9 _08076_/I _08478_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlya_2
XFILLER_5_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09738__A1 _09725_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08410__A1 split15/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07213__A2 _05924_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11125_ _11125_/D _11672_/CLK _11125_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05775__A2 _05775_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11056_ _11056_/D _11056_/RN input68/Z _11056_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__09910__A1 _10387_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10007_ _10007_/A1 _10265_/A3 _10014_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__05527__A2 _05515_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06724__A1 _06724_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10909_ _10909_/A1 _10909_/A2 _10909_/A3 _10909_/A4 _10918_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_32_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09977__A1 _09972_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10036__A1 _10352_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07080_ _07080_/I _11151_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06100_ _10945_/A1 _05969_/I _06101_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06031_ _09775_/A1 _11607_/Q _06034_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09729__A1 _09725_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07982_ split6/Z _07984_/I _07983_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09721_ _09722_/A2 _11586_/Q _09722_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06963__A1 _06941_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06933_ _06933_/A1 _06904_/Z _06938_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09652_ _09652_/I _11563_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08704__A2 _08786_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09901__A1 _09986_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06864_ _06869_/A2 _11085_/Q _06865_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10511__A2 _11323_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09583_ _09583_/I _11541_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06795_ _10979_/A1 _05633_/B _06796_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08603_ _08603_/A1 _08603_/A2 _08603_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05815_ _08791_/A1 _06217_/I _05816_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_08534_ _08355_/I _08417_/B _08534_/B _08534_/C _08535_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA_input113_I wb_adr_i[24] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05746_ _08799_/A1 _05803_/A2 _05747_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10275__A1 _10352_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07140__A1 _05927_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08465_ _08478_/A1 _08462_/I _08465_/B _08466_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05677_ _05677_/I _09775_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
X_08396_ _08396_/A1 _08563_/A2 _08459_/B _08396_/A4 _08397_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_07416_ _07417_/A2 _11249_/Q _07417_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11111__CLK _11672_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09968__B2 _10373_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09968__A1 _11523_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07347_ _07081_/Z _07347_/A2 _07347_/B _07348_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07278_ _06851_/Z _07290_/A2 _07278_/B _07279_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11261__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09017_ _09039_/A2 _11363_/Q _09018_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08190__B _08493_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06229_ _06229_/A1 _06229_/A2 _06229_/A3 _06229_/A4 _06235_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__06954__A1 _10947_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05757__A2 _11086_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09919_ _11639_/Q _11638_/Q _09920_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__11611__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05833__I _05833_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08459__A1 _07720_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_split14_I split21/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11674_ _11674_/D _11683_/CLK _11674_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06485__A3 _06491_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11604__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10625_ _10896_/A1 _11438_/Q _10627_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10556_ _10556_/A1 _10556_/A2 _10556_/A3 _10556_/A4 _10557_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_10487_ _10487_/A1 _10487_/A2 _10487_/A3 _10487_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_5_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11108_ _11108_/D _11686_/RN _06705_/Z _11108_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__06945__A1 _10938_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11039_ _11039_/I _11686_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07370__A1 _07370_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05600_ _05600_/I _05753_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06580_ input103/Z input102/Z _06583_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10257__A1 _10378_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05920__A2 _11432_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11134__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05531_ _06610_/A3 _11698_/Q _11699_/Q _05532_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09111__A2 _09114_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08250_ _08250_/I _08253_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07673__A2 _08095_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08870__A1 _07431_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08181_ _08490_/A1 _08614_/A2 _08181_/A3 _08182_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_07201_ _07201_/A1 _05924_/Z _07201_/B _09015_/I _07240_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XANTENNA__11284__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10009__A1 _10042_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07132_ _07132_/A1 _07151_/B _07132_/B _07133_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06228__A3 _06217_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput200 _10638_/A1 mgmt_gpio_oeb[34] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_07063_ _07067_/A2 _11147_/Q _07064_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06014_ _06014_/A1 _06014_/A2 _06015_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput211 _06675_/Z mgmt_gpio_out[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput222 _06671_/ZN mgmt_gpio_out[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__09178__A2 _11413_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput233 _11183_/Q mgmt_gpio_out[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput244 _11186_/Q mgmt_gpio_out[5] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_160_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07189__A1 _05925_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput266 _11275_/Q pll_div[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput255 _06718_/I pad_flash_io0_oe VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput277 _11076_/Q pll_trim[13] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__05739__A2 _05805_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput299 _11293_/Q pwr_ctrl_out VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput288 _11291_/Q pll_trim[23] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_07965_ split6/I _08449_/B _07966_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08689__A1 _07566_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09704_ _09121_/I _09722_/A2 _09704_/B _09705_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10699__C _10880_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06916_ _06917_/A2 _11104_/Q _06917_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07896_ _08436_/B _08549_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09635_ _09154_/Z _09647_/A2 _09635_/B _09636_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_3_5__f_wb_clk_i clkbuf_0_wb_clk_i/Z _11672_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09125__I _09125_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10496__A1 _10886_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06847_ _09125_/I _06847_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__07361__A1 _07081_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05911__A2 _11504_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09566_ _09187_/Z _09572_/A2 _09566_/B _09567_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06778_ _07110_/I _11069_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09497_ _09270_/Z _09497_/A2 _09497_/B _09498_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08517_ _08517_/A1 _07564_/I _08518_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10248__B2 _11465_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11627__CLK _11665_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05729_ _08940_/A1 _11346_/Q _05730_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09102__A2 _09114_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10799__A2 _11482_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08448_ _08693_/A2 _08448_/A2 _08555_/A2 _08610_/A1 _08448_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_08379_ _08379_/A1 _08450_/A1 _08552_/B _08382_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_10410_ _10410_/I _10493_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_23_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11390_ _11390_/D _11686_/RN _06705_/Z _11390_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10341_ _10341_/A1 _10341_/A2 _10341_/A3 _10342_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08204__I _08204_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09169__A2 _09169_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10272_ _10350_/A1 _10272_/A2 _10273_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10723__A2 _11440_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11157__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09341__A2 _09347_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10487__A1 _10487_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05902__A2 _09599_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11565__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07104__A1 _07081_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10239__A1 _10356_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07655__A2 _08509_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11657_ _11657_/D input76/Z _11658_/CLK _11657_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__11140__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11588_ _11588_/D _11686_/RN _06705_/Z _11588_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__08604__A1 _07844_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10608_ _11325_/Q _10924_/A1 _10608_/B _10608_/C _10609_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_10539_ _10902_/A2 _11524_/Q _10542_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10411__A1 _10884_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06091__A1 _08915_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05738__I _05738_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07158__C _09015_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08907__A2 _08913_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07750_ _08304_/B _08614_/A2 _08678_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09332__A2 _09347_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06701_ _06701_/I _07242_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_07681_ _08386_/A1 _08395_/A2 _07682_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06632_ input77/Z _06632_/A2 _06632_/B _06633_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09420_ _09420_/I _11489_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09351_ _09116_/Z _09372_/A2 _09351_/B _09352_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06563_ _06563_/I _10501_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09096__A1 _07431_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08302_ _08403_/A2 _08302_/A2 _08494_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09282_ _09125_/Z _09297_/A2 _09282_/B _09283_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05514_ _11162_/Q _05515_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__05657__A1 _07201_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08233_ _08233_/A1 _08657_/A2 _08486_/A2 _08241_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06494_ _06491_/B _11062_/Q _06495_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07646__A2 _08509_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11131__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09399__A2 _09015_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08164_ _08483_/A1 _08205_/C _08242_/A1 _08235_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_07115_ _05927_/Z _09116_/I _07116_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08095_ _08095_/A1 _08095_/A2 _08096_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10402__A1 _10915_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06082__A1 _06082_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06082__B2 _06082_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07046_ _06843_/Z _07046_/A2 _07046_/B _07047_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09020__A1 _09039_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input41_I mgmt_gpio_in[14] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10705__A2 _10916_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11198__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08997_ _09013_/A2 _11357_/Q _08998_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07948_ _07964_/A1 _07981_/A2 _08444_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10469__A1 _10406_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07879_ _07873_/Z _08013_/A2 _08562_/A2 _07883_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__06137__A2 _05924_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09618_ _09622_/A2 _11553_/Q _09619_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10890_ _10890_/A1 _10890_/A2 _10890_/A3 _10890_/A4 _10918_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_09549_ _09549_/A1 _09015_/I _09572_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__11370__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07637__A2 _08417_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08834__A1 _07431_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11511_ _11511_/D _11686_/RN _06705_/Z _11511_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__10641__A1 _10913_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11442_ _11442_/D _11686_/RN _06705_/Z _11442_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_171_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11373_ _11373_/D _11686_/RN _06705_/Z _11373_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__08062__A2 _08332_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06073__A1 _11582_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10324_ _11226_/Q _10363_/A2 _11143_/Q _10363_/B2 _10324_/C _10325_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_10255_ _10255_/A1 _10255_/A2 _10255_/A3 _10264_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11189__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09562__A2 _11535_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10186_ _10379_/A1 _11559_/Q _10378_/A1 _11551_/Q _10188_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_38_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06128__A2 _06128_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10880__A1 _10092_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11361__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08109__I _08616_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07628__A2 _07609_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08825__A1 _08825_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10632__A1 _10903_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06064__A1 input67/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08053__A2 split13/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11322__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09250__A1 _09116_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06064__B2 _05925_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08920_ _07431_/Z _08938_/A2 _08920_/B _08921_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10699__A1 _10092_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08851_ _07431_/Z _08863_/A2 _08851_/B _08852_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11472__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07802_ _07802_/I _08329_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
X_05994_ input16/Z _06393_/A1 _06394_/A1 input7/Z _05998_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08782_ _08782_/I _11290_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07733_ _07733_/A1 _07496_/I _07734_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06119__A2 _08890_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07664_ _07664_/I _08285_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05878__A1 _09374_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09403_ _09422_/A2 _11484_/Q _09404_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06615_ _11221_/Q _07296_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11352__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07595_ _07595_/A1 _08531_/B _07600_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05893__A4 _05893_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09334_ _09347_/A2 _11462_/Q _09335_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06546_ _09938_/B _09859_/A1 _06567_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08816__A1 _08820_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10623__B2 _10894_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06477_ _06475_/Z _06477_/A2 _11066_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11104__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09265_ _09187_/Z _09272_/A2 _09265_/B _09266_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08216_ _08216_/A1 _08576_/A2 _08216_/A3 _08617_/A3 _08221_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA_input89_I spimemio_flash_io1_oeb VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09196_ _09196_/I _11418_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08044__A2 _08167_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08147_ _08147_/A1 _08147_/A2 _08147_/A3 _08226_/A1 _08150_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_20_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09792__A2 _09798_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08078_ split12/I _08545_/A2 _08079_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_07029_ _06837_/Z _07032_/A2 _07029_/B _07030_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09544__A2 _09547_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07593__I _07593_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10040_ _10042_/A1 _10040_/A2 _10041_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output245_I _06666_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11591__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07307__A1 _07081_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10942_ _10942_/A1 _10934_/I _10942_/B _10943_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05869__A1 _06324_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11343__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10873_ _10921_/A1 _11101_/Q _10877_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08807__A1 _08820_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10209__A4 _10209_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_364 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08283__A2 _07609_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10614__A1 _11382_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10614__B2 _10883_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11345__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06294__A1 _07006_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08035__A2 _08395_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11425_ _11425_/D input76/Z _06705_/Z _11425_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__09232__A1 _09246_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08586__A3 _08586_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09783__A2 _09798_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11356_ _11356_/D _11686_/RN _06705_/Z _11356_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__11495__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10307_ _10344_/A1 _10880_/C _10307_/B _10308_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09535__A2 _09547_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11287_ _11287_/D input76/Z _06705_/Z _11287_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_10238_ _11385_/Q _10355_/A2 _11377_/Q _10355_/B2 _10238_/C _10247_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_10169_ _10360_/A1 _11431_/Q _10171_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11582__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xrebuffer19 _07857_/A1 _07500_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06847__I _09125_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10853__A1 _10899_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06400_ _08839_/A1 _08839_/A2 _11307_/Q _06401_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_07380_ _07380_/I _11238_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06331_ _09549_/A1 _11531_/Q _06333_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10605__B2 _11349_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10605__A1 _10920_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09471__A1 _09472_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07077__A3 _06871_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06262_ _06262_/A1 _06262_/A2 _06263_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11381__SETN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09050_ _09050_/I _11373_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06285__A1 _09066_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08001_ _08001_/A1 _08005_/A1 _08167_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__10369__B1 _10369_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06193_ _05703_/Z _07412_/A1 _11152_/Q _06194_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__09223__A1 _09246_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11396__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09952_ _09952_/I _10265_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09526__A2 _09547_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08903_ _08913_/A2 _11327_/Q _08904_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_09883_ _09876_/I _09892_/A2 _09884_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_873 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input143_I wb_dat_i[21] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08834_ _07431_/Z _08837_/A2 _08834_/B _08835_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11218__CLK _11666_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08765_ _08784_/A2 _11285_/Q _08766_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07716_ _08430_/A1 _07716_/A2 _07716_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__06760__A2 _08672_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05977_ _11327_/Q _10190_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_167_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08696_ _08217_/B _08696_/A2 _08696_/B _08696_/C _08697_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_07647_ _07647_/A1 _07647_/A2 _08419_/C _08275_/B _07651_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__11325__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11334__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07578_ _08405_/B _08669_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__11368__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06529_ _11224_/Q _08431_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
X_09317_ _09317_/I _11456_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09462__A1 _09472_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08265__A2 _07616_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06276__A1 _06839_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11349__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10072__A2 _10369_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09248_ _09248_/A1 _09015_/Z _09272_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA_output195_I _06082_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09179_ _09125_/Z _09195_/A2 _09179_/B _09180_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09214__A1 _09187_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06028__A1 _05660_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11021__A1 _11019_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11210_ _11210_/D _11656_/CLK _11210_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07776__A1 _07722_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11141_ _11141_/D _11686_/RN _06705_/Z _11141_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xinput111 wb_adr_i[22] input111/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput100 wb_adr_i[12] input100/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11072_ _11072_/D _11686_/RN _06705_/Z _11072_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
Xinput144 wb_dat_i[22] input144/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput133 wb_dat_i[12] input133/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput122 wb_adr_i[3] _07487_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_130_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10023_ _10023_/A1 _10265_/A3 _10024_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput166 wb_sel_i[3] input166/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput155 wb_dat_i[3] input155/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06503__A2 _11059_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11316__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10925_ _10925_/A1 _10092_/I _10923_/Z _10925_/A4 _10926_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_10856_ _11153_/Q _10902_/A2 _11149_/Q _10902_/B2 _10856_/C _10863_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XPHY_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09453__A1 _09472_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_10787_ _10787_/A1 _10092_/Z _10785_/Z _10787_/A4 _10788_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__06267__B2 _11274_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09205__A1 _09125_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11408_ _11408_/D input76/Z _06705_/Z _11408_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__06019__B2 _09171_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06019__A1 _11423_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11339_ _11339_/D _11686_/RN _06705_/Z _11339_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_140_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06880_ _06902_/A2 _11093_/Q _06881_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05900_ _09549_/A1 _11536_/Q _05901_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05831_ _06667_/A2 _06619_/B _05831_/B _05832_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08550_ _08550_/A1 _08550_/A2 _08694_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11510__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05762_ _11330_/Q _08890_/A1 _11291_/Q _08761_/A1 _05762_/C _05775_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_07501_ _07870_/A3 input97/Z _07515_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08481_ _08481_/A1 _08462_/I _08481_/B _08482_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05693_ _05693_/I _05693_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__10826__A1 _10826_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11307__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07432_ _07433_/A2 _11253_/Q _07433_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09444__A1 _09241_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_322 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07363_ _07398_/A1 _08825_/A2 _06871_/Z _07368_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__08247__A2 _07609_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11660__CLK _11663_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09102_ _06851_/Z _09114_/A2 _09102_/B _09103_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06314_ _05927_/I input43/Z _06318_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07294_ _08672_/B _08036_/B _11028_/A2 _11025_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__10054__A2 _10351_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06245_ _07412_/A1 _06238_/Z _11249_/Q _06246_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09033_ _06859_/Z _09039_/A2 _09033_/B _09034_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11003__A1 _08493_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06176_ _11239_/Q _06181_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_2_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10762__B1 _10886_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09935_ _10911_/A1 _10415_/A2 _09935_/B _09936_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06430__A1 _07398_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09866_ _09866_/A1 _09866_/A2 _09867_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08817_ _06863_/Z _08820_/A2 _08817_/B _08818_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11546__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09797_ _09798_/A2 _11610_/Q _09798_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11190__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08748_ _08748_/I _11279_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08679_ _08679_/A1 _08679_/A2 _08691_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_26_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10710_ _10887_/A2 _11424_/Q _10712_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11288__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11690_ _11690_/D _11690_/RN input68/Z _11690_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__09435__A1 _09154_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06249__A1 _08795_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08238__A2 _08656_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10641_ _10913_/A2 _11590_/Q _10644_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10572_ _10572_/A1 _10572_/A2 _10572_/A3 _10572_/A4 _10573_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_122_222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11124_ _11124_/D _11672_/CLK _11124_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06421__A1 _07419_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11055_ _11055_/I _11702_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05775__A3 _05775_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07781__I _08689_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11533__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10006_ _10006_/A1 _10006_/A2 _10006_/A3 _10006_/A4 _10046_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__11537__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09910__A2 _09912_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06724__A2 _11056_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10808__A1 _10900_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09674__A1 _09674_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10908_ _10908_/I _10909_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11683__CLK _11683_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09426__A1 _09116_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10839_ _10839_/A1 _10839_/A2 _10840_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09977__A2 _09876_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06030_ _09800_/A1 _11615_/Q _06034_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06660__A1 _11059_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11063__CLK input68/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07981_ _08015_/A1 _07981_/A2 _07984_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06412__A1 _08799_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09720_ _09720_/I _11585_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06932_ _06932_/I _11108_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07691__I _07691_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06863_ _09241_/I _06863_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__11528__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09651_ _09116_/I _09672_/A2 _09651_/B _09652_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_3_4__f_wb_clk_i clkbuf_0_wb_clk_i/Z _11666_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08704__A3 _06838_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09582_ _09125_/Z _09597_/A2 _09582_/B _09583_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06794_ _11676_/Q _10979_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08602_ _08602_/A1 _11016_/A1 _08603_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05814_ _11426_/Q _09197_/A1 _11418_/Q _09171_/A1 _05814_/C _05827_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_08533_ _08671_/A1 _08687_/A1 _08626_/A1 _08539_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_05745_ _06393_/A1 input19/Z _05749_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09665__A1 _09672_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input106_I wb_adr_i[18] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07140__A2 _09187_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08464_ _08464_/A1 _08464_/A2 _08464_/A3 _08464_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_05676_ _08825_/A2 _05805_/A2 _05677_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08395_ _08395_/A1 _08395_/A2 _08395_/B _08396_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07415_ _07415_/I _11248_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09968__A2 _10373_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07346_ _07347_/A2 _11229_/Q _07347_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07979__A1 split15/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11406__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07277_ _07290_/A2 _11200_/Q _07278_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10983__B1 _08460_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06651__A1 input80/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input71_I mgmt_gpio_in[7] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09016_ _09016_/A1 _09015_/Z _09039_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__06770__I _07110_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06228_ _07412_/A1 _11142_/Q _06217_/Z _06229_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06159_ _06159_/A1 _06159_/A2 _06160_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11556__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06403__A1 _08742_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09918_ _09918_/I _11638_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09849_ _09849_/I _11626_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11519__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07106__I _07110_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09656__A1 _09672_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07131__A2 _05927_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10266__A2 _10092_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11673_ _11673_/D _11683_/CLK _11673_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_10624_ _10895_/A1 _11446_/Q _10627_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06890__A1 _06851_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10018__A2 _10265_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11086__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10555_ _10887_/B1 _11428_/Q _10556_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10486_ _10486_/A1 _10486_/A2 _10486_/A3 _10486_/A4 _10487_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__06642__A1 input83/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08395__A1 _08395_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_11107_ _11107_/D _11686_/RN _06705_/Z _11107_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_11038_ _09121_/I _11038_/A2 _11038_/B _11039_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05905__B1 _09674_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07370__A2 _06238_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09647__A1 _09270_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06855__I _09158_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05530_ _05541_/A2 _11159_/Q _05539_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07122__A2 _07151_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11429__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08180_ _08180_/A1 _08180_/A2 _08180_/A3 _08183_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_07200_ _08865_/A1 _07114_/B _07201_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06881__A1 _06837_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08870__A2 _08888_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10009__A2 _10265_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07131_ _11192_/Q _05927_/Z _07151_/B _07131_/C _07132_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__11579__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput201 _06643_/Z mgmt_gpio_oeb[35] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_07062_ _08795_/A1 _06238_/Z _06871_/Z _07067_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
Xoutput234 _11099_/Q mgmt_gpio_out[30] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput223 _11168_/Q mgmt_gpio_out[20] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_173_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06013_ _09424_/A1 _11495_/Q _06014_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput212 _06655_/Z mgmt_gpio_out[10] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__07189__A2 _09241_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput267 _11276_/Q pll_div[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput256 _11704_/Z pad_flash_io1_do VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput245 _06666_/ZN mgmt_gpio_out[6] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput289 _11087_/Q pll_trim[24] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput278 _11077_/Q pll_trim[14] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_59_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07964_ _07964_/A1 _07964_/A2 _08449_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_07895_ _07930_/A1 _07973_/A2 _08436_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09703_ _09722_/A2 _11580_/Q _09704_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06915_ _06915_/I _11103_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09634_ _09647_/A2 _11558_/Q _09635_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06846_ _06846_/I _11080_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09638__A1 _09158_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09565_ _09572_/A2 _11536_/Q _09566_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06777_ _07110_/I _11068_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09496_ _09497_/A2 _11514_/Q _09497_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08310__A1 _07605_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08516_ _08516_/A1 _08675_/A3 _08642_/A1 _08598_/I _08520_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__07113__A2 _07242_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05728_ _05728_/I _08940_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XANTENNA__06765__I _07110_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08447_ _08447_/I _08610_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05659_ _08825_/A2 _08719_/A2 _05660_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__06872__A1 _08839_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_426 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_08378_ split8/Z _07976_/I _08378_/B _08552_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09810__A1 _09823_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07329_ _07310_/I _11214_/Q _07330_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10340_ _10379_/A1 _11151_/Q _10341_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output275_I _11074_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10271_ _11330_/Q _10304_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10708__B1 _10913_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10184__A1 _10374_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08129__A1 split7/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09629__A1 _09121_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06675__I _06675_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10239__A2 _11409_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09986__I _09986_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_11656_ _11656_/D input76/Z _11656_/CLK _11656_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__09801__A1 _09823_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11587_ _11587_/D _11686_/RN _06705_/Z _11587_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_10607_ _10607_/A1 _10461_/I _10607_/B _10607_/C _10608_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_10538_ _11508_/Q _10900_/A1 _10538_/B _10542_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10411__A2 _10903_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09935__B _09935_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10469_ _10406_/I _10417_/I _09920_/I _10887_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__10175__A1 _10367_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11101__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10478__A2 _10427_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06700_ _06700_/I _06700_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07680_ _07680_/I _08395_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_64_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_06631_ input77/Z input90/Z _06632_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11251__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09350_ _09372_/A2 _11467_/Q _09351_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06562_ _09908_/A2 _11637_/Q _06563_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09096__A2 _09114_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08301_ _08301_/A1 _08590_/A3 _08303_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09281_ _09297_/A2 _11445_/Q _09282_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05513_ _06611_/B2 _06521_/A2 _06460_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05657__A2 input60/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08232_ split7/Z _08232_/A2 _08656_/B _08486_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09896__I _09896_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06493_ _06493_/A1 _11062_/Q _06491_/B _06496_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_08163_ _08163_/I _08483_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08094_ _08094_/A1 _08094_/A2 _08094_/A3 _08094_/A4 _08101_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_07114_ _05656_/I _07114_/A2 _07114_/B _07114_/C _07151_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__10402__A2 _10914_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06606__A1 _10433_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07045_ _07046_/A2 _11142_/Q _07046_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08359__A1 _08043_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10166__A1 _10357_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08996_ _08996_/I _11356_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07947_ _07947_/A1 _08529_/A2 _07947_/A3 _08370_/B _07950_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA_input34_I mask_rev_in[8] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07878_ _07878_/I _08562_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08531__A1 _08355_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10469__A2 _10417_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_09617_ _09617_/I _11552_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06829_ _06835_/A1 _11077_/Q _06830_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09548_ _09548_/I _11530_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_43_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05896__A2 _05969_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11510_ _11510_/D _11686_/RN _06705_/Z _11510_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_09479_ _09121_/Z _09497_/A2 _09479_/B _09480_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10641__A2 _11590_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06845__A1 _06843_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11441_ _11441_/D input76/Z _06705_/Z _11441_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_11372_ _11372_/D _11686_/RN _06705_/Z _11372_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_152_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06073__A2 _09699_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10323_ _10323_/A1 _10323_/A2 _10324_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11124__CLK _11672_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10254_ _10370_/A1 _11497_/Q _10255_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10185_ _10185_/A1 _10185_/A2 _10185_/A3 _10189_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__07022__A1 _06837_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07573__A2 _08509_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11274__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08825__A2 _08825_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11639_ _11639_/D _11686_/RN _11666_/CLK _11639_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__08589__A1 _08589_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07261__A1 _07265_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06064__A2 _05924_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09250__A2 _09272_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10148__A1 _10148_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10148__B2 _10148_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11617__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08850_ _08863_/A2 _11310_/Q _08851_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07801_ _08045_/A3 _07808_/A2 _07802_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08761__A1 _08761_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08781_ _06863_/Z _08784_/A2 _08781_/B _08782_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05993_ _05993_/A1 _05993_/A2 _05993_/A3 _05993_/A4 _05999_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_07732_ _08600_/A2 _08513_/A2 _08298_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07663_ _07663_/A1 _07690_/A2 _07664_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09402_ _09402_/I _11483_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06614_ _11216_/Q _10930_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10320__B2 _10359_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09333_ _09333_/I _11461_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07594_ _07596_/I _08686_/A2 _08531_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_40_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06545_ _06545_/I _09859_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10623__A2 _10894_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06827__A1 _11014_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06476_ _06476_/A1 _06476_/A2 _06477_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09264_ _09272_/A2 _11440_/Q _09265_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08215_ _08616_/B _07722_/I _08215_/B _08617_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09195_ _06867_/Z _09195_/A2 _09195_/B _09196_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08146_ _08434_/A1 _08227_/B _08226_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11147__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08077_ _08161_/A1 _08200_/B _08464_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07252__A1 _07265_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11564__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11297__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07028_ _07032_/A2 _11137_/Q _07029_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07004__A1 _06843_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06358__A3 _06217_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08752__A1 _08759_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08979_ _06855_/Z _08988_/A2 _08979_/B _08980_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11579__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08504__A1 _07508_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10941_ _10934_/I _11669_/Q _10942_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10311__A1 _10350_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_10872_ _10872_/A1 _10872_/A2 _10872_/A3 _10872_/A4 _10879_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XPHY_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10614__A2 _10884_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06818__A1 _06835_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11517__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11687__CLKN input68/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11424_ _11424_/D input76/Z _06705_/Z _11424_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_61_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10378__A1 _10378_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09232__A2 _11430_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07243__A1 _07265_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11355_ _11355_/D _11686_/RN _06705_/Z _11355_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_10306_ _10306_/A1 _06556_/I _10926_/C _10306_/C _10307_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_11286_ _11286_/D input76/Z _06705_/Z _11286_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__08991__A1 _09013_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10237_ _10237_/A1 _10237_/A2 _10238_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08743__A1 _08759_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10168_ _11399_/Q _10359_/A2 _11391_/Q _10359_/B2 _10168_/C _10173_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_66_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10550__A1 _10886_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09299__A2 _09015_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10099_ _10356_/A1 _11405_/Q _10101_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_179_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10853__A2 _11252_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06863__I _09241_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1090 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06809__A1 _10993_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06330_ _05687_/I _05941_/I _07099_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09471__A2 _11506_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11098__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06261_ _08799_/A1 _11272_/Q _08719_/A2 _06262_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_08000_ _08000_/A1 _08006_/A2 _08005_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10369__B2 _11253_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06192_ _06192_/I _07412_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XANTENNA__07234__A1 _07240_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09951_ _10926_/C _10880_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__08982__A1 _06859_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05796__A1 _09424_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08902_ _08902_/I _11326_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_852 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_830 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_09882_ _11633_/Q _09892_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__08734__A1 _06847_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10541__A1 _10905_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05548__A1 _05519_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_874 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_863 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_08833_ _08837_/A2 _11305_/Q _08834_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_896 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input136_I wb_dat_i[15] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08764_ _08764_/I _11284_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05976_ _05976_/I _08726_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
X_07715_ _08294_/B _08294_/C _08490_/A3 _07716_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_08695_ _08695_/I _08697_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07646_ _08276_/B _08509_/A1 _08275_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07577_ _07607_/A1 _07657_/A2 _08405_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05720__A1 _07006_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06528_ _11687_/Q _11172_/Q _06701_/I _06749_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_09316_ _09187_/Z _09322_/A2 _09316_/B _09317_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06773__I _07110_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06276__A2 _11080_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09247_ _09247_/I _11434_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06459_ _06459_/I _11068_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_output188_I _10148_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09178_ _09195_/A2 _11413_/Q _09179_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09214__A2 _09220_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06028__A2 _11623_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08129_ split7/Z _08217_/B _08130_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07225__A1 _07240_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07776__A2 _07508_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08973__A1 _06847_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11140_ _11140_/D _11686_/RN _06705_/Z _11140_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__10780__A1 _10780_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11261__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput101 wb_adr_i[13] input101/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11071_ _11071_/D _11686_/RN _06705_/Z _11071_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__07109__I _07110_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput123 wb_adr_i[4] _07522_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput145 wb_dat_i[23] input145/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput112 wb_adr_i[23] input112/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput134 wb_dat_i[13] input134/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10022_ _10356_/A1 _11403_/Q _10027_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput156 wb_dat_i[4] input156/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput167 wb_stb_i input167/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_3_0__f_wb_clk_i_I clkbuf_0_wb_clk_i/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11312__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10924_ _10924_/A1 _11207_/Q _10925_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05711__A1 _09624_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10855_ _10855_/A1 _10855_/A2 _10856_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10599__A1 _10905_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06267__A2 _08742_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10786_ _10924_/A1 _11329_/Q _10787_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11462__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10138__C _10138_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09205__A2 _09220_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11407_ _11407_/D input76/Z _06705_/Z _11407_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__06019__A2 _09197_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11338_ _11338_/D _11686_/RN _06705_/Z _11338_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__05778__A1 _06238_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10771__A1 _10771_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11252__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11269_ _11269_/D _11269_/RN input68/Z _11269_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_140_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10523__A1 _10899_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_3_3__f_wb_clk_i clkbuf_0_wb_clk_i/Z _11658_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_05830_ _11269_/Q _05969_/I _05830_/B _06619_/B _05831_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_07500_ _07858_/A2 _07500_/A2 _07870_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_05761_ _05761_/A1 _05761_/A2 _05762_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05950__A1 _06839_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09141__A1 _09142_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08480_ _08480_/A1 _08475_/Z _08619_/A2 _08568_/A2 _08480_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_05692_ _05703_/I _06872_/A2 _05693_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_07431_ _09121_/I _07431_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_35_498 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07362_ _07362_/I _11233_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09444__A2 _09447_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06313_ _06313_/A1 _06313_/A2 _06313_/A3 _06313_/A4 _06329_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_09101_ _09114_/A2 _11390_/Q _09102_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07293_ _07293_/I _07300_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_30_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06244_ _07398_/A1 _06238_/Z _11245_/Q _06246_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09032_ _09039_/A2 _11368_/Q _09033_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06175_ _06175_/A1 _06175_/A2 _06175_/A3 _06175_/A4 _06187_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__07207__A1 _05924_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07758__A2 _08242_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11243__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05769__A1 _09041_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10762__A1 _10886_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09934_ _09934_/I _10415_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06430__A2 _07006_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09865_ _09865_/A1 _09865_/A2 _09866_/A2 _09866_/A1 _11629_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_08816_ _08820_/A2 _11300_/Q _08817_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06768__I _07110_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09796_ _09796_/I _11609_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11335__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08747_ _07431_/Z _08759_/A2 _08747_/B _08748_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05959_ _06396_/A1 input31/Z _05962_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09132__A1 _09142_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08678_ _08678_/A1 _08678_/A2 _08678_/A3 _08678_/A4 _08679_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_53_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07629_ _08415_/B _08417_/A2 _07631_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11485__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10640_ _10913_/B2 _11582_/Q _10644_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09435__A2 _09447_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08238__A3 _08242_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06249__A2 _06238_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10571_ _10888_/A1 _11413_/Q _10572_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_166_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11482__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09199__A1 _09116_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10753__A1 _10911_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11234__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11123_ _11123_/D _11672_/CLK _11123_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06421__A2 _07006_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11054_ _11055_/I _11701_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09371__A1 _09372_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10505__A1 _10905_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10005_ _11491_/Q _10370_/A1 _10371_/A1 _11483_/Q _10006_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_76_332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06185__A1 _09775_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06678__I _06678_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11380__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05932__A1 _08846_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09123__A1 _09121_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09674__A2 _09015_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10907_ _10907_/A1 _10907_/A2 _10908_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_498 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11395__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09426__A2 _09447_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10838_ _10887_/B1 _11141_/Q _10839_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10769_ _10895_/A1 _11449_/Q _10771_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10992__A1 _10966_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11473__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11208__CLK _11656_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06660__A2 input67/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08937__A1 _08938_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11225__RN input162/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10744__A1 _10744_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07980_ _07980_/A1 _07980_/A2 _08648_/A2 _08650_/A3 _07983_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__11358__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06412__A2 _11295_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06931_ _06843_/Z _06931_/A2 _06931_/B _06932_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09362__A1 _09372_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09650_ _09672_/A2 _11563_/Q _09651_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08601_ _08601_/A1 _08601_/A2 _08601_/A3 _08601_/A4 _08602_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_06862_ _06862_/I _11084_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11348__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09581_ _09597_/A2 _11541_/Q _09582_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06793_ _06793_/I _11071_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05813_ _05813_/A1 _05813_/A2 _05814_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08532_ _08532_/A1 _08532_/A2 _08532_/A3 _08626_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05744_ _05744_/I _06393_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__09114__A1 _06867_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08463_ _08474_/A1 _08200_/B _08464_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06479__A2 _05515_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07414_ _07076_/Z _07417_/A2 _07414_/B _07415_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05675_ _05732_/I _09724_/A1 _05805_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_08394_ _08394_/A1 _08545_/A2 _08395_/B _08459_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07345_ _07345_/I _11228_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07979__A2 _08380_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07276_ _07276_/I _11199_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06100__A1 _10945_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11464__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09015_ _09015_/I _09015_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_20
XANTENNA__10983__A1 _08431_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06227_ _07398_/A1 _11140_/Q _06217_/Z _06229_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_input64_I mgmt_gpio_in[35] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08928__A1 _08938_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06651__A2 input82/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08043__I _08043_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06158_ _09117_/A1 _11397_/Q _06159_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06089_ _08726_/A1 _11276_/Q _06092_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06403__A2 _11278_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09917_ _09917_/A1 _09927_/A2 _10407_/A1 _09902_/I _09918_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__09353__A1 _09372_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09848_ _09270_/I _09848_/A2 _09848_/B _09849_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06167__A1 _10942_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05914__A1 _11520_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09779_ _09798_/A2 _11604_/Q _09780_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05914__B2 _09474_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09105__A1 _06855_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10266__A3 _10266_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11672_ _11672_/D _11672_/CLK _11672_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10623_ _11494_/Q _10894_/A2 _11486_/Q _10894_/B2 _10623_/C _10627_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__07419__A1 _05703_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06890__A2 _06902_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08092__A1 _08161_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10554_ _10887_/A2 _11420_/Q _10556_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11455__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10974__A1 _11016_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10485_ _10891_/A1 _11475_/Q _10486_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08919__A1 _08938_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10726__A1 _10899_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11500__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11207__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08395__A2 _08395_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11106_ _11106_/D _11686_/RN _06705_/Z _11106_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__09344__A1 _09241_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11650__CLK _11665_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11037_ _11038_/A2 _11686_/Q _11038_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07370__A3 _06871_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09647__A2 _09647_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10662__B1 _10913_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06881__A2 _06902_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07130_ _05927_/Z _09154_/I _07131_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06871__I _09015_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11446__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11180__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07061_ _07061_/I _11146_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11272__SETN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput235 _11100_/Q mgmt_gpio_out[31] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput224 _11169_/Q mgmt_gpio_out[21] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput202 _06639_/Z mgmt_gpio_oeb[36] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_06012_ _09449_/A1 _11503_/Q _06014_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput213 _11176_/Q mgmt_gpio_out[11] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_160_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08386__A2 _08632_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput246 _11188_/Q mgmt_gpio_out[7] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput268 _11277_/Q pll_div[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput257 _06755_/ZN pad_flash_io1_ie VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_141_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput279 _11078_/Q pll_trim[15] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_07963_ _07963_/A1 _07963_/A2 _08446_/C _08610_/A3 _07966_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__09335__A1 _09154_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11287__SETN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07894_ _07894_/I _07973_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09702_ _09702_/I _11579_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06914_ _06837_/Z _06917_/A2 _06914_/B _06915_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09633_ _09633_/I _11557_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07897__A1 split15/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06845_ _06843_/Z _06869_/A2 _06845_/B _06846_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09564_ _09564_/I _11535_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09638__A2 _09647_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08515_ _08204_/I _07827_/I _08515_/B _08598_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06776_ _07110_/I _11067_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09495_ _09495_/I _11513_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05727_ _07006_/A2 _05995_/A2 _05728_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08446_ _08010_/I _07959_/I _08446_/B _08446_/C _08447_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05658_ _05645_/I _09724_/A1 _08719_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_08377_ _08351_/I _08686_/A1 _08449_/B _08450_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__11685__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06872__A2 _06872_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05589_ _05616_/C _11257_/Q _05589_/B _05590_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07328_ _07328_/A1 _07328_/A2 _11213_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09810__A2 _11614_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08074__A1 _08434_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11523__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10956__A1 _10934_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07259_ _06859_/Z _07265_/A2 _07259_/B _07260_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_output170_I _11295_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10270_ _11653_/Q _10344_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08377__A2 _08686_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09574__A1 _09574_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10708__B2 _11592_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11673__CLK _11683_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output268_I _11277_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10184__A2 _11535_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06388__A1 _07419_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09326__A1 _09116_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07888__A1 _07685_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10487__A3 _10487_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09629__A2 _09647_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06312__A1 _08791_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11676__RN input162/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11655_ _11655_/D input76/Z _11665_/CLK _11655_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_11586_ _11586_/D _11686_/RN _06705_/Z _11586_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__10427__B _10427_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10947__A1 _10947_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10606_ _10922_/A1 _11357_/Q _10919_/A1 _11365_/Q _10607_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07812__A1 _07722_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10537_ _10537_/A1 _10537_/A2 _10537_/A3 _10537_/A4 _10538_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_6_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10468_ _10468_/A1 _10468_/A2 _10468_/A3 _10467_/Z _10487_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__09565__A1 _09572_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10175__A2 _11479_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06379__A1 _07370_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10399_ _10427_/B _10503_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_69_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11600__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06630_ _11313_/Q _06632_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_25_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06561_ _11636_/Q _09908_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11546__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08300_ _08339_/A1 _08300_/A2 _08358_/A2 _08590_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06492_ _06500_/A1 _11061_/Q _06493_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05512_ _05532_/A2 _05533_/A2 _11698_/Q _06521_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09280_ _09280_/I _11444_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06303__A1 _06259_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08231_ _08434_/A1 _08380_/B _08332_/A1 _08656_/B _08657_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08162_ _08162_/A1 _08167_/A1 _08163_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10938__A1 _10938_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07803__A1 _08332_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08093_ split7/I _08659_/A1 _08094_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11696__CLK input68/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07113_ _05656_/I _07242_/A2 _07114_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_109_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10402__A3 _10883_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06606__A2 _09934_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05814__B1 _11418_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07044_ _07044_/I _11141_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09556__A1 _09572_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08359__A2 _08512_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input166_I wb_sel_i[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08995_ _07431_/Z _09013_/A2 _08995_/B _08996_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07946_ split15/I _08352_/B _08370_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05593__A2 _06466_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input27_I mask_rev_in[30] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11076__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07877_ _08519_/A1 _08358_/A2 _07878_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10469__A3 _09920_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09616_ _09187_/Z _09622_/A2 _09616_/B _09617_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06828_ _11696_/Q _05633_/B _06828_/B _09241_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA__06776__I _07110_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10874__B1 _10920_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09547_ _09270_/Z _09547_/A2 _09547_/B _09548_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06759_ _06759_/I _11219_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10626__B1 _10897_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09478_ _09497_/A2 _11508_/Q _09479_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11658__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08429_ _08294_/B _08562_/A2 _08430_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06845__A2 _06869_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11440_ _11440_/D input76/Z _06705_/Z _11440_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__09795__A1 _09241_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11371_ _11371_/D _11686_/RN _06705_/Z _11371_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_50_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10322_ _10361_/A1 _11139_/Q _10323_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09547__A1 _09270_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10253_ _10371_/A1 _11489_/Q _10255_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06460__B _06466_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10184_ _10374_/A1 _11535_/Q _10185_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11419__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11569__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08522__A2 _08522_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11649__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10093__A1 _10350_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08038__A1 split12/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11638_ _11638_/D _11686_/RN _11666_/CLK _11638_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__07310__I _07310_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08589__A2 _08677_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06049__B1 _11510_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09786__A1 _09154_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09946__B _11645_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11569_ _11569_/D _11686_/RN _06705_/Z _11569_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__09538__A1 _09158_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08210__A1 _08434_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08210__B2 _08332_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11099__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07013__A2 _06904_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07800_ _07800_/A1 _07800_/A2 _08509_/C _07800_/A4 _07805_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__08761__A2 _06838_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08780_ _08784_/A2 _11290_/Q _08781_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07731_ _08005_/A2 _07999_/A2 _07470_/I _08513_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_05992_ _11335_/Q _08915_/A1 _08940_/A1 _11343_/Q _05993_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09710__A1 _09154_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08513__A2 _08513_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07662_ _08280_/B _08417_/A2 _08540_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09401_ _09116_/Z _09422_/A2 _09401_/B _09402_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07593_ _07593_/I _08686_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_3
X_06613_ _06613_/I _11161_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10320__A2 _10359_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09332_ _09125_/Z _09347_/A2 _09332_/B _09333_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06544_ _09938_/A1 _11628_/Q _06545_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_500 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06827__A2 _05633_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06475_ _06476_/A1 _06476_/A2 _06475_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_09263_ _09263_/I _11439_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08214_ _08214_/I _08216_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09194_ _09195_/A2 _11418_/Q _09195_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08145_ _08161_/A1 _08227_/B _08147_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09777__A1 _09116_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09529__A1 _09121_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08076_ _08076_/I _08161_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
X_07027_ _06217_/Z _11033_/A2 _06871_/Z _07032_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__10139__A2 _11430_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08978_ _08988_/A2 _11351_/Q _08979_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07929_ _08438_/B _07964_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_152_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09701__A1 _09116_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10940_ _10940_/A1 _10940_/A2 _11668_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output300_I _06408_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_10871_ _10871_/A1 _10871_/A2 _10871_/A3 _10871_/A4 _10872_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XPHY_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_322 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08268__A1 _08400_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_355 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_101_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06818__A2 _09158_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06294__A3 _11033_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11423_ _11423_/D input76/Z _06705_/Z _11423_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__11241__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11354_ _11354_/D _11686_/RN _06705_/Z _11354_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_11285_ _11285_/D input76/Z _06705_/Z _11285_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_10305_ _10305_/A1 _06556_/I _10306_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10236_ _10352_/A1 _11361_/Q _10237_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_3_2__f_wb_clk_i clkbuf_0_wb_clk_i/Z _11665_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08743__A2 _11278_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05557__A2 _05519_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09940__B2 _09922_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06754__A1 _06514_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11391__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10167_ _10167_/A1 _10167_/A2 _10168_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10098_ _11381_/Q _10355_/A2 _11373_/Q _10355_/B2 _10098_/C _10107_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_74_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1091 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06809__A2 _05633_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10066__A1 _11444_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06260_ _06396_/A1 input15/Z _06262_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_163_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10369__A2 _10369_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06191_ _07092_/A1 _11156_/Q _06194_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07234__A2 _11187_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09950_ _09950_/A1 _10047_/B _10926_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__08982__A2 _08988_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06993__A1 _06974_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08901_ _06851_/Z _08913_/A2 _08901_/B _08902_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_853 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_842 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_831 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_820 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_09881_ _09898_/A1 _11633_/Q _09884_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_875 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_864 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_08832_ _08832_/I _11304_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_08763_ _07426_/Z _08784_/A2 _08763_/B _08764_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05975_ _08839_/A1 _05995_/A2 _05976_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input129_I wb_cyc_i VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07714_ _07714_/I _08490_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XANTENNA__08498__A1 _07570_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08694_ _08694_/A1 _08694_/A2 _08694_/A3 _08699_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_07645_ _08276_/B _08417_/A2 _08419_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07576_ _07576_/I _07657_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11114__CLK _11672_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05720__A2 _05803_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09315_ _09322_/A2 _11456_/Q _09316_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06527_ _06527_/I _06701_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_166_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input94_I trap VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09246_ _06867_/Z _09246_/A2 _09246_/B _09247_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06458_ _06458_/A1 _06458_/A2 _06459_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06389_ _08825_/A1 _06238_/Z _11153_/Q _06390_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__07885__I _07885_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09177_ _09177_/I _11412_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08128_ _08161_/A1 _08217_/B _08475_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08059_ _08084_/A1 _08095_/A1 _08142_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08973__A2 _08988_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06984__A1 _06974_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10780__A2 _10780_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11070_ _11070_/D _11070_/RN input68/Z _11070_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xinput102 wb_adr_i[14] input102/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10021_ _10135_/A1 _09887_/I _10356_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xinput135 wb_dat_i[14] input135/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput113 wb_adr_i[24] input113/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput124 wb_adr_i[5] _07447_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_102_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09922__A1 _10642_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput168 wb_we_i input168/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput146 wb_dat_i[24] input146/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput157 wb_dat_i[5] input157/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10296__A1 _10375_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07161__A1 _07197_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10923_ _10923_/A1 _10923_/A2 _10923_/A3 _10923_/A4 _10923_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__05711__A2 _11562_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10854_ _10900_/A1 _11147_/Q _10855_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_169_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11607__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09989__A1 _09896_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10048__A1 _11323_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_10785_ _10785_/A1 _10785_/A2 _10785_/A3 _10785_/A4 _10785_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XPHY_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08413__A1 _07616_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11406_ _11406_/D input76/Z _06705_/Z _11406_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__10220__A1 _10377_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11337_ _11337_/D _11686_/RN _06705_/Z _11337_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__05778__A2 _05803_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10771__A2 _10771_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06975__A1 _10935_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06204__I _06204_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11268_ _11268_/D _11268_/RN input68/Z _11268_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
X_10219_ _10378_/A1 _11552_/Q _10221_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11199_ _11199_/D _11686_/RN _06705_/Z _11199_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_97_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05760_ _06785_/A1 _11078_/Q _05761_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11137__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08575__B _08575_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05691_ _05691_/I _09574_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XANTENNA__10287__B2 _11466_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10826__A3 _10826_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07430_ _07430_/I _11252_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11563__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07361_ _07081_/Z _07361_/A2 _07361_/B _07362_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11287__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06312_ _08791_/A1 _08825_/A2 _11293_/Q _06313_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09100_ _09100_/I _11389_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07292_ _11218_/Q _11222_/D _11220_/Q _11219_/Q _07293_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
XANTENNA__08652__A1 _08692_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09031_ _09031_/I _11367_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06243_ _09374_/A1 _11476_/Q _06246_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06174_ _07201_/A1 input53/Z _06175_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07207__A2 _09121_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10211__A1 _10367_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11501__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09933_ _10642_/A1 _10427_/B _10911_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__09904__A1 _09927_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09864_ _09864_/A1 _09868_/A3 _09866_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_08815_ _08815_/I _11299_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11516__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09795_ _09241_/I _09798_/A2 _09795_/B _09796_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07391__A1 _07391_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08746_ _08759_/A2 _11279_/Q _08747_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05958_ input17/Z _06393_/A1 _06394_/A1 input8/Z _05962_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10278__A1 _10356_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08677_ _08304_/B _08677_/A2 _08678_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05889_ _09248_/A1 _11441_/Q _05891_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07628_ _08415_/B _07609_/Z _07631_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06784__I _07114_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08891__A1 _08913_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07559_ _07575_/A1 _07590_/A1 _07560_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output298_I _11072_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10570_ _10887_/A2 _11421_/Q _10572_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10450__A1 _11411_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10450__B2 _10883_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09229_ _09246_/A2 _11429_/Q _09230_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09199__A2 _09220_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10202__A1 _10357_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06957__A1 _10950_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11122_ _11122_/D _11672_/CLK _11122_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11053_ _11055_/I _11700_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06709__A1 _11057_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10004_ _09996_/I _09876_/I _10371_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__07382__A1 _07081_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05932__A2 input66/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09123__A2 _09142_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10906_ _10906_/A1 _11686_/Q _10907_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08882__A1 _06859_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11170__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05696__A1 _09549_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10837_ _10887_/A2 _11139_/Q _10839_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08634__A1 _08460_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08634__B2 _08493_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10768_ _10896_/A1 _11441_/Q _10771_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10441__A1 _10900_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10699_ _10092_/Z _11659_/Q _10699_/B _10880_/C _10701_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__06948__A1 _06941_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10744__A2 _10092_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06412__A3 _08799_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06930_ _06931_/A2 _11108_/Q _06931_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input1_I debug_mode VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08600_ _08600_/A1 _08600_/A2 _08623_/A2 _08519_/B _08600_/C _08601_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_06861_ _06859_/Z _06869_/A2 _06861_/B _06862_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09580_ _09580_/I _11540_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06792_ _06835_/A1 _09116_/I _06792_/B _06793_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05812_ _09117_/A1 _11402_/Q _05813_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08531_ _08355_/I _08262_/B _08531_/B _08532_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07125__A1 _05927_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05743_ _07398_/A1 _08799_/A1 _05744_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09114__A2 _09114_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08462_ _08462_/I _08474_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05674_ _05590_/I _05674_/A2 _05732_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10680__A1 _10899_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07413_ _07417_/A2 _11248_/Q _07414_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08873__A1 _06847_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_285 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08393_ _08395_/A1 _08545_/A2 _08393_/B _08563_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08625__A1 _08686_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07344_ _07076_/Z _07347_/A2 _07344_/B _07345_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07428__A2 _11252_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07275_ _06847_/Z _07290_/A2 _07275_/B _07276_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_163_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09014_ _09014_/I _11362_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06100__A2 _05969_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06226_ _09171_/A1 _11412_/Q _06229_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06157_ _09144_/A1 _11405_/Q _06159_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input57_I mgmt_gpio_in[29] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06088_ _08803_/A1 _11297_/Q _06092_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11302__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09916_ _09916_/A1 _09916_/A2 _09917_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06779__I _07110_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09847_ _09848_/A2 _11626_/Q _09848_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11452__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05616__C _05616_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06167__A2 _05969_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05914__A2 _09499_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09778_ _09778_/I _11603_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_output213_I _11176_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08729_ _08729_/I _11273_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09105__A2 _09114_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05678__A1 _09775_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10120__B1 _10377_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11671_ _11671_/D _11683_/CLK _11671_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11152__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08616__A1 split8/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10622_ _10622_/A1 _10622_/A2 _10623_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07419__A2 _07419_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10553_ _10888_/A1 _11412_/Q _10556_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10484_ _10484_/A1 _10427_/B _10891_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__10187__B1 _10377_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05850__B2 _05723_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09041__A1 _09041_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10726__A2 _11504_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06689__I _06689_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05602__A1 input58/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11105_ _11105_/D _11686_/RN _06705_/Z _11105_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_78_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09344__A2 _09347_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11036_ _11036_/I _11685_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05905__A2 _09699_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11391__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07658__A2 _08686_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11143__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_462 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07060_ _06843_/Z _07060_/A2 _07060_/B _07061_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11325__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07830__A2 _08677_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06011_ _11487_/Q _09399_/A1 _11479_/Q _09374_/A1 _06011_/C _06024_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
Xoutput225 _11170_/Q mgmt_gpio_out[22] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput203 _06636_/Z mgmt_gpio_oeb[37] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__10178__B1 _10369_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput214 _11177_/Q mgmt_gpio_out[12] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__09032__A1 _09039_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput236 _06646_/ZN mgmt_gpio_out[32] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput247 _06662_/Z mgmt_gpio_out[8] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput258 _06755_/I pad_flash_io1_oe VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__11475__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput269 _11271_/Q pll_ena VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_07962_ split15/Z _08375_/B _08610_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09701_ _09116_/I _09722_/A2 _09701_/B _09702_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07893_ _07917_/A1 split13/Z _07894_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06149__A2 _11461_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09335__A2 _09347_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06913_ _06917_/A2 _11103_/Q _06914_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09632_ _09125_/I _09647_/A2 _09632_/B _09633_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06844_ _06869_/A2 _11080_/Q _06845_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09563_ _09158_/Z _09572_/A2 _09563_/B _09564_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11382__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09099__A1 _06847_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08514_ _08333_/I _08514_/A2 _08514_/A3 _08642_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_130_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06775_ _07110_/I _11066_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input111_I wb_adr_i[22] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09494_ _09241_/Z _09497_/A2 _09494_/B _09495_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08846__A1 _08846_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05726_ _05726_/I _05995_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
X_05657_ _07201_/A1 input60/Z _05662_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08445_ _08445_/A1 _08445_/A2 _08555_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10653__A1 _10092_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11134__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08376_ _08376_/A1 _08140_/I _08610_/A3 _08446_/B _08379_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_05588_ _06490_/B1 _05515_/I _05588_/B _05616_/C _05589_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__10405__A1 _10417_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06872__A3 _06871_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07327_ _07310_/I _11213_/Q _07328_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10956__A2 _11674_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09271__A1 _09272_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06085__A1 _06839_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07258_ _07265_/A2 _11194_/Q _07259_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07189_ _05925_/Z _09241_/I _07190_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06209_ _05703_/Z _11686_/Q _11033_/A2 _06211_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__09023__A1 _09039_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10708__A2 _10913_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09574__A2 _09015_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07585__A1 _08339_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06388__A2 _06238_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output330_I _11668_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09326__A2 _09347_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07337__A1 _07076_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05899__A1 _05693_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10892__A1 _10892_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08837__A1 _07426_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_split12_I split12/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06312__A2 _08825_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11654_ _11654_/D input76/Z _11665_/CLK _11654_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__11348__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10605_ _10920_/A1 _11341_/Q _10920_/B1 _11349_/Q _10607_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10494__I _10494_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11585_ _11585_/D _11686_/RN _06705_/Z _11585_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__08065__A2 _08043_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11347__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09262__A1 _09158_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10536_ _10903_/A1 _11556_/Q _10537_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11498__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10467_ _10467_/A1 _10467_/A2 _10467_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__06379__A2 _06238_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10398_ _06563_/I _09920_/I _10400_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_11019_ _10966_/Z _11019_/A2 _11019_/A3 _11019_/A4 _11019_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__06000__A1 _05693_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10883__A1 _10883_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06560_ _06560_/I _10426_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_06491_ _06479_/C _06500_/B1 _06491_/B _06500_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_05511_ _11699_/Q _05533_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08230_ _08225_/Z _08567_/B _08479_/A1 _08482_/A1 _08233_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__06303__A2 _06265_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08161_ _08161_/A1 _08656_/B _08484_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09253__A1 _09121_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08092_ _08161_/A1 _08659_/A1 _08094_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07112_ _05927_/Z _06701_/I _07114_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10402__A4 _10910_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05814__A1 _11426_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05814__B2 _09171_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07043_ _06837_/Z _07046_/A2 _07043_/B _07044_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input159_I wb_dat_i[7] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08994_ _09013_/A2 _11356_/Q _08995_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07945_ split21/I _08352_/B _07947_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07876_ _07876_/A1 _07876_/A2 _08013_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_09615_ _09622_/A2 _11552_/Q _09616_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06827_ _11014_/A1 _05633_/B _06828_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10874__A1 _10920_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09546_ _09547_/A2 _11530_/Q _09547_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06758_ _06760_/A1 _07296_/A2 _06759_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08819__A1 _08820_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09477_ _09477_/I _11507_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05709_ _05703_/I _08719_/A2 _05710_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11107__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06689_ _06689_/I _06689_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08493__B _08493_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08428_ _08428_/A1 _08544_/A3 _08428_/A3 _08431_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_08359_ _08043_/I _08512_/I _08359_/B _08549_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__11640__CLK _11666_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09795__A2 _09798_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11370_ _11370_/D _11686_/RN _06705_/Z _11370_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA_output280_I _11284_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05805__A1 _06217_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10321_ _10360_/A1 _11141_/Q _10323_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09547__A2 _09547_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08512__I _08512_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10252_ _11513_/Q _10369_/A2 _10369_/B1 _11505_/Q _10255_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_10183_ _10375_/A1 _11543_/Q _10185_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_3_1__f_wb_clk_i clkbuf_0_wb_clk_i/Z _11656_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__11594__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06230__A1 _09144_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06781__A2 _05633_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07730__A1 _07570_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10865__A1 _10911_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11346__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11170__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10617__A1 _10887_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11706_ input66/Z _11706_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08286__A2 _08395_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06297__A1 _06192_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11637_ _11637_/D _11686_/RN _11658_/CLK _11637_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__11286__SETN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09235__A1 _09246_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11568_ _11568_/D _11686_/RN _06705_/Z _11568_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__06049__A1 _11518_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06049__B2 _09474_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09786__A2 _09798_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07797__A1 _07722_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10519_ _10914_/A1 _11596_/Q _10522_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11499_ _11499_/D _11686_/RN _06705_/Z _11499_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__09538__A2 _09547_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11585__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07730_ _07570_/I _07822_/I _08600_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05991_ _05991_/I _08915_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__11513__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05980__B1 _11282_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09710__A2 _09722_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10399__I _10427_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10856__B2 _10902_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07661_ _08280_/B _07609_/Z _07684_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11337__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09400_ _09422_/A2 _11483_/Q _09401_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07592_ _07607_/A1 _07694_/A2 _07596_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06612_ _06612_/A1 _06619_/A1 _06466_/B _05509_/I _06613_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_09331_ _09347_/A2 _11461_/Q _09332_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06543_ _11627_/Q _09938_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10608__A1 _11325_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09474__A1 _09474_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11663__CLK _11663_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06288__A1 _09016_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06474_ _05515_/I _06610_/A3 _06474_/B _06476_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09262_ _09158_/Z _09272_/A2 _09262_/B _09263_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08029__A2 _07885_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08213_ split7/I _08232_/A2 _08213_/B _08214_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09193_ _09193_/I _11417_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09226__A1 _09246_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08144_ split7/Z _08227_/B _08147_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09777__A2 _09798_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11033__A1 _05703_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07788__A1 _08592_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08075_ split12/I _08395_/A1 _08076_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__09529__A2 _09547_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07026_ _07026_/I _11136_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08201__A2 _08242_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10544__B1 _10920_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11576__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07960__A1 _08355_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08977_ _08977_/I _11350_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11193__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07928_ _07928_/A1 _08365_/B _08442_/C _07928_/A4 _07932_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_07859_ input105/Z _06591_/I input106/Z _07470_/I _07859_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__09701__A2 _09722_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11328__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_10870_ _10915_/A1 _11234_/Q _10916_/A1 _11230_/Q _10871_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_09529_ _09121_/Z _09547_/A2 _09529_/B _09530_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08268__A2 _08686_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09465__A1 _09472_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06279__A1 _08761_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_356 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09217__A1 _06863_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11422_ _11422_/D input76/Z _06705_/Z _11422_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__07779__A1 _08328_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11353_ _11353_/D _11686_/RN _06705_/Z _11353_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_11284_ _11284_/D _11686_/RN _06705_/Z _11284_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_10304_ _10304_/A1 _10382_/A2 _10304_/B _10304_/C _10306_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_152_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10235_ _10353_/A1 _11369_/Q _10237_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11536__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06203__A1 _05703_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11567__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10166_ _10357_/A1 _11415_/Q _10167_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10097_ _10097_/A1 _10097_/A2 _10098_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11686__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11319__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10838__A1 _10887_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10999_ _10966_/Z _10999_/A2 _11000_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09456__A1 _09472_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1092 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1081 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1070 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09208__A1 _09154_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06190_ _05687_/I _05742_/I _07092_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11066__CLK input68/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_09880_ _09880_/I _11632_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08900_ _08913_/A2 _11326_/Q _08901_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_843 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_832 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_821 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_08831_ _06847_/Z _08837_/A2 _08831_/B _08832_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11558__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_876 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_865 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06745__A2 input71/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_898 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_887 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_08762_ _08784_/A2 _11284_/Q _08763_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05974_ _05974_/A1 _05974_/A2 _11268_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08693_ _08693_/A1 _08693_/A2 _08693_/A3 _08693_/A4 _08694_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__08498__A2 _07748_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07713_ _07839_/A2 _07751_/A1 _07714_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10829__A1 _10921_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07644_ _08276_/B _07609_/Z _07647_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_497 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07170__A2 _05925_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09447__A1 _09270_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07575_ _07575_/A1 _07525_/I _07576_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09314_ _09314_/I _11455_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06526_ _06526_/A1 _11349_/Q _06527_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__11409__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09245_ _09246_/A2 _11434_/Q _09246_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06457_ _06457_/I _06458_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11006__A1 _10966_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input87_I spimemio_flash_io0_oeb VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06388_ _07419_/A2 _06238_/Z _11149_/Q _06390_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09176_ _09121_/Z _09195_/A2 _09176_/B _09177_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08127_ _08434_/A1 _08217_/B _08224_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09158__I _09158_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11559__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08058_ _08058_/I _08095_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06433__A1 _09016_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07009_ _07009_/I _11131_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10020_ _10357_/A1 _11411_/Q _10027_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput136 wb_dat_i[15] input136/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput114 wb_adr_i[25] input114/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput103 wb_adr_i[15] input103/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput125 wb_adr_i[6] _07513_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__09922__A2 _09935_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput147 wb_dat_i[25] input147/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput158 wb_dat_i[6] input158/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10296__A2 _11546_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10922_ _10922_/A1 _11108_/Q _10923_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09438__A1 _09158_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10853_ _10899_/A1 _11252_/Q _10855_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06466__B _06466_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09989__A2 _09878_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10048__A2 _10382_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10784_ _10921_/A1 _11337_/Q _10785_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08110__A1 _08434_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11089__CLK _11663_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09610__A1 _09154_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11405_ _11405_/D input76/Z _06705_/Z _11405_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_11336_ _11336_/D _11686_/RN _06705_/Z _11336_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__06424__A1 _08915_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08177__A1 _08490_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11267_ _11267_/D _11267_/RN input68/Z _11267_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
X_10218_ _11576_/Q _10377_/A1 _10379_/A1 _11560_/Q _10221_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_11198_ _11198_/D _11686_/RN _06705_/Z _11198_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__07924__A1 split15/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_364 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10149_ _11494_/Q _10370_/A1 _11486_/Q _10371_/A1 _10149_/C _10152_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_121_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07152__A2 _07151_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05690_ _05703_/I _05805_/A2 _05691_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10826__A4 _10826_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09429__A1 _09121_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_07360_ _07361_/A2 _11233_/Q _07361_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06311_ _08825_/A1 _08825_/A2 _11303_/Q _06313_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_07291_ _07291_/I _11204_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09030_ _06855_/Z _09039_/A2 _09030_/B _09031_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06242_ _09399_/A1 _11484_/Q _06246_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11701__CLK input68/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06173_ _05927_/I input44/Z _06175_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09601__A1 _09116_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10211__A2 _11480_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06415__A1 _06785_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09932_ _09932_/I _10427_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__06966__A2 _06904_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06179__B1 _07391_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09863_ _11627_/Q _11628_/Q _11629_/Q _09868_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_640 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_09794_ _09798_/A2 _11609_/Q _09795_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05926__B1 _05925_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input141_I wb_dat_i[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08814_ _06859_/Z _08820_/A2 _08814_/B _08815_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07391__A2 _06904_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08745_ _08745_/I _11278_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09668__A1 _09672_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05957_ _05957_/A1 _05957_/A2 _05957_/A3 _05967_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08340__A1 _08632_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08676_ _08676_/I _08678_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10278__A2 _11410_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05888_ _11409_/Q _09144_/A1 _11401_/Q _09117_/A1 _05888_/C _05893_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__11231__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07627_ _08686_/B _08415_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_13_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07558_ _07558_/I _07607_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08891__A2 _11323_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06509_ _06510_/A2 _11057_/Q _06510_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07489_ _07489_/I _07836_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__08643__A2 split5/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06654__A1 _06786_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output193_I _10146_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10450__A2 _10888_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11381__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09228_ _09228_/I _11428_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09159_ _09169_/A2 _11407_/Q _09160_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06406__A1 _06406_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11121_ _11121_/D _11672_/CLK _11121_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11052_ _11055_/I _11699_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10003_ _09996_/I _09973_/I _10370_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__06709__A2 input67/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09659__A1 _09672_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08331__A1 _08686_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10905_ _10905_/A1 _11158_/Q _10907_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06893__A1 _06855_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10836_ _10836_/A1 _10836_/A2 _11663_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08882__A2 _08888_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10767_ _11497_/Q _10894_/A2 _11489_/Q _10894_/B2 _10767_/C _10771_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__08634__A2 _08634_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10698_ _10698_/A1 _10092_/Z _10696_/Z _10698_/A4 _10699_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__06645__A1 input80/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05999__A3 _05999_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10729__B1 _11520_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08398__B2 _07297_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11319_ _11319_/D input76/Z _06705_/Z _11319_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__11104__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05620__A2 _05515_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09898__A1 _09898_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06860_ _06869_/A2 _11084_/Q _06861_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05811_ _05811_/I _09117_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XANTENNA__05923__A3 _05923_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11254__CLK _06687_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06791_ _06835_/A1 _11071_/Q _06792_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08530_ _08530_/I _08532_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05742_ _05742_/I _07398_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_3
X_05673_ _05673_/A1 _05673_/A2 _05683_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08461_ split12/Z _08614_/A2 _08462_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__07125__A2 _09125_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07412_ _07412_/A1 _06238_/Z _06838_/Z _07417_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__06884__A1 _06843_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08873__A2 _08888_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08392_ _08392_/A1 _08392_/A2 _08613_/A3 _08456_/B _08396_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__09822__A1 _09823_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08625__A2 _08686_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07343_ _07347_/A2 _11228_/Q _07344_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07274_ _07290_/A2 _11199_/Q _07275_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09013_ _06867_/Z _09013_/A2 _09013_/B _09014_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06225_ _09197_/A1 _11420_/Q _06229_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06156_ _11517_/Q _09499_/A1 _11509_/Q _09474_/A1 _06156_/C _06165_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__10196__B2 _10351_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06087_ _06087_/A1 _06087_/A2 _06087_/A3 _06087_/A4 _06093_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_09915_ _09912_/I _10407_/A1 _09916_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_09846_ _09846_/I _11625_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10499__A2 _10387_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_470 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_09777_ _09116_/I _09798_/A2 _09777_/B _09778_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06989_ _06989_/A1 _06989_/A2 _11125_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08728_ _07426_/Z _08740_/A2 _08728_/B _08729_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07116__A2 _05927_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08313__A1 _07508_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08659_ _08659_/A1 _08696_/A2 _08660_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output206_I _06082_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10120__A1 _10377_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11670_ _11670_/D _11683_/CLK _11670_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09813__A1 _09823_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08616__A2 _07727_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10621_ _10892_/A1 _11470_/Q _10622_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07419__A3 _06838_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06627__A1 input92/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10552_ _11436_/Q _10896_/A1 _11380_/Q _10884_/A1 _10552_/C _10556_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_182_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11127__CLK _11683_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10483_ _10892_/A1 _11467_/Q _10486_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10187__A1 _10377_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05850__A2 _08990_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09041__A2 _09015_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_180 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05602__A2 _05515_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11104_ _11104_/D _11686_/RN _06705_/Z _11104_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_150_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11035_ _09116_/I _11038_/A2 _11035_/B _11036_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11277__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08552__A1 _08380_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10111__A1 _10111_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11500__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10662__A2 _10913_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10819_ _10911_/A1 _11578_/Q _10820_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09804__A1 _09823_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11515__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10965__A3 _07297_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06010_ _06010_/A1 _06010_/A2 _06011_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput226 _11171_/Q mgmt_gpio_out[23] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput215 _06693_/Z mgmt_gpio_out[13] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_126_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput204 _06726_/ZN mgmt_gpio_oeb[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput237 _06649_/ZN mgmt_gpio_out[33] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_160_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput248 _06658_/ZN mgmt_gpio_out[9] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput259 _11281_/Q pll90_sel[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__07043__A1 _06837_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07961_ split14/Z _08375_/B _08446_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07594__A2 _08686_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08791__A1 _08791_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09700_ _09722_/A2 _11579_/Q _09701_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06912_ _06912_/A1 _06904_/Z _06917_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07892_ _07892_/I _07917_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09631_ _09647_/A2 _11557_/Q _09632_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06843_ _09121_/I _06843_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_28_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10350__A1 _10350_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09562_ _09572_/A2 _11535_/Q _09563_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06774_ _07110_/I _11065_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08513_ _08572_/A2 _08513_/A2 _08514_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09099__A2 _09114_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05725_ _07006_/A2 _06872_/A2 _05991_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_09493_ _09497_/A2 _11513_/Q _09494_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08846__A2 _06904_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10102__B2 _10359_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08444_ _08449_/A1 _08010_/I _08444_/B _08445_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05656_ _05656_/I _07201_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XANTENNA_input104_I wb_adr_i[16] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06857__A1 _06855_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08375_ _08383_/A1 _08355_/I _08375_/B _08446_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05587_ _11062_/Q _05515_/I _05588_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10405__A2 _10427_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07326_ _10950_/A1 _07326_/A2 _07328_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07257_ _07257_/I _11193_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_151_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07188_ _07188_/I _11178_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06208_ _09549_/A1 _11532_/Q _06211_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08231__B1 _08332_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06139_ _08846_/A1 input63/Z _06141_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_3_0__f_wb_clk_i clkbuf_0_wb_clk_i/Z _11663_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07034__A1 _07398_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08534__A1 _08355_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09829_ _09848_/A2 _11620_/Q _09830_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05899__A2 _11528_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06848__A1 _06869_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06312__A3 _11293_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11653_ _11653_/D input76/Z _11665_/CLK _11653_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10604_ _10604_/A1 _10604_/A2 _10604_/A3 _10604_/A4 _10608_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_80_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11584_ _11584_/D _11686_/RN _06705_/Z _11584_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__09262__A2 _09272_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10535_ _10910_/A1 _11564_/Q _10537_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10466_ _10894_/B2 _11483_/Q _10467_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07025__A1 _06843_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10397_ _10433_/A1 _10406_/I _10883_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_69_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10580__A1 _10894_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_0_wb_clk_i_I wb_clk_i VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11018_ _08431_/B input136/Z _08460_/B input145/Z _11019_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10332__A1 _10370_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07879__A3 _08562_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08540__A4 _08540_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06490_ _06490_/A1 _05588_/B _06490_/B1 _06479_/C _11063_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05510_ _11700_/Q _05532_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06839__A1 _06839_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06303__A3 _06303_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08160_ split7/Z _08656_/B _08165_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07111_ _11164_/Q _07117_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09253__A2 _09272_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07264__A1 _07265_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08091_ _08434_/A1 _08659_/A1 _08094_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11442__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05814__A2 _09197_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07042_ _07046_/A2 _11141_/Q _07043_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11469__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11592__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10571__A1 _10888_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08993_ _08993_/I _11355_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07944_ _08355_/I _08352_/B _08529_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07875_ _07875_/A1 _08006_/A2 _07875_/A3 _07876_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06826_ _11681_/Q _11014_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09614_ _09614_/I _11551_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09545_ _09545_/I _11529_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06757_ _06757_/I _11220_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08819__A2 _06266_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_05708_ _09649_/A1 _11570_/Q _05712_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06688_ _11304_/Q _06688_/A2 _06688_/B _06689_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10626__A2 _10897_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09476_ _09116_/Z _09497_/A2 _09476_/B _09477_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08427_ _08541_/A3 _08541_/A2 _08428_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05639_ _05605_/I _05639_/A2 _09724_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_08358_ _08623_/A2 _08358_/A2 _08512_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07255__A1 _07265_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08289_ _08289_/I _08541_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07309_ _11219_/Q input162/Z _07310_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_166_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output273_I _11079_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05805__A2 _05805_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10320_ _11133_/Q _10359_/A2 _11131_/Q _10359_/B2 _10320_/C _10325_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_10251_ _10251_/A1 _10251_/A2 _10251_/A3 _10264_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08755__A1 _08759_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10182_ _10373_/A1 _11519_/Q _10373_/B1 _11527_/Q _10185_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10314__A1 _10352_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07144__I _11170_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11315__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10617__A2 _11422_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11705_ input65/Z _11705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11465__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11636_ _11636_/D _11686_/RN _11658_/CLK _11636_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XANTENNA__09235__A2 _11431_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06049__A2 _09499_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11567_ _11567_/D _11686_/RN _06705_/Z _11567_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__07246__A1 _07265_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07797__A2 _08639_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10518_ _11612_/Q _10915_/A1 _11572_/Q _10911_/A1 _10518_/C _10522_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_10_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08994__A1 _09013_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11498_ _11498_/D _11686_/RN _06705_/Z _11498_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10449_ _10449_/A1 _10449_/A2 _10449_/A3 _10450_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08746__A1 _08759_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10553__A1 _10888_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06221__A2 _11444_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05990_ _08990_/A1 _11359_/Q _05993_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05980__A1 _11277_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05980__B2 _08742_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09171__A1 _09171_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10856__A2 _10902_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07660_ _07660_/I _08280_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__07721__A2 _08339_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07591_ _07591_/I _07694_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06611_ _06611_/A1 _11690_/Q _11688_/Q _06466_/B _06611_/B2 _11162_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_09330_ _09330_/I _11460_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06542_ _06542_/I _09938_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10608__A2 _10924_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09474__A2 _09015_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09261_ _09272_/A2 _11439_/Q _09262_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08212_ _08575_/B _07722_/I _08212_/B _08576_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06473_ _06497_/A1 _11065_/Q _06473_/A3 _06476_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09192_ _06863_/Z _09195_/A2 _09192_/B _09193_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08143_ _08478_/B _08227_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11033__A2 _11033_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07237__A1 _05924_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08074_ _08434_/A1 _08200_/B _08081_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08985__A1 _06863_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05799__A1 _09449_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11273__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07025_ _06843_/Z _07025_/A2 _07025_/B _07026_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10792__A1 _10887_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06460__A2 _06619_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08737__A1 _06851_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11331__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10544__A1 _10922_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input32_I mask_rev_in[6] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08976_ _06851_/Z _08988_/A2 _08976_/B _08977_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11338__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07927_ _08355_/I _08367_/B _07928_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09162__A1 _09169_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07858_ _07858_/A1 _07858_/A2 _07857_/Z _07860_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__11488__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07789_ _07789_/A1 _07789_/A2 _08320_/B _07789_/A4 _07790_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_06809_ _10993_/A1 _05633_/B _06810_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09528_ _09547_/A2 _11524_/Q _09529_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_324 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09465__A2 _11504_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_09459_ _09472_/A2 _11502_/Q _09460_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08673__B1 _08493_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09217__A2 _09220_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11421_ _11421_/D input76/Z _06705_/Z _11421_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__07779__A2 _08315_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08976__A1 _06851_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11352_ _11352_/D _11686_/RN _06705_/Z _11352_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10303_ _10303_/A1 _10303_/A2 _10303_/A3 _10303_/A4 _10304_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__10783__A1 _10922_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11283_ _11283_/D input76/Z _06705_/Z _11283_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__10535__A1 _10910_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08728__A1 _07426_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10234_ _11353_/Q _10351_/A2 _11345_/Q _10351_/B2 _10234_/C _10247_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__07400__A1 _07076_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06203__A2 _07419_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10165_ _10356_/A1 _11407_/Q _10167_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10096_ _10352_/A1 _11357_/Q _10097_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10299__B1 _10377_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08900__A1 _08913_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10998_ _10998_/A1 _10998_/A2 _10998_/A3 _10999_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__09456__A2 _11501_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1082 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1071 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1060 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1093 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09208__A2 _09220_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11619_ _11619_/D _11686_/RN _06705_/Z _11619_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__07219__A1 _07240_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08967__A1 _07426_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11255__RN input162/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10526__A1 _10894_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08719__A1 _08799_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_844 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_833 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_08830_ _08837_/A2 _11304_/Q _08831_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_877 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_855 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_888 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_08761_ _08761_/A1 _06838_/Z _08784_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__09144__A1 _09144_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05973_ _05584_/I _11268_/Q _05974_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08692_ _08692_/A1 _08692_/A2 _08692_/B _08692_/C _08693_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_07712_ _08426_/A1 _08294_/C _08430_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11630__CLK _11665_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xrepeater345 input76/Z _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
X_07643_ _07643_/I _08276_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__09447__A2 _09447_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07574_ _07574_/A1 _08403_/A2 _07574_/A3 _08258_/B _07583_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_09313_ _09158_/Z _09322_/A2 _09313_/B _09314_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06525_ input67/Z _11303_/Q _06526_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06130__A1 _09624_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09244_ _09244_/I _11433_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06456_ _06456_/A1 _06456_/A2 _06457_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11494__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09175_ _09195_/A2 _11412_/Q _09176_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10214__B1 _10369_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08126_ _08126_/I _08217_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
X_06387_ _09474_/A1 _11507_/Q _06390_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10765__A1 _10892_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11246__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08057_ _08057_/A1 _08057_/A2 _08058_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10780__A4 _10780_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07008_ _06837_/Z _07011_/A2 _07008_/B _07009_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11160__CLK input68/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08186__A2 _08394_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_214 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput115 wb_adr_i[26] input115/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput104 wb_adr_i[16] _07863_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput126 wb_adr_i[7] _07449_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput148 wb_dat_i[26] input148/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput159 wb_dat_i[7] input159/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput137 wb_dat_i[16] input137/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_output236_I _06646_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11285__SETN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08959_ _08963_/A2 _11345_/Q _08960_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09135__A1 _09142_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09902__I _09902_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10921_ _10921_/A1 _11102_/Q _10923_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09438__A2 _09447_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10852_ _10852_/A1 _10852_/A2 _10852_/A3 _10852_/A4 _10872_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_10783_ _10922_/A1 _11361_/Q _10785_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06121__A1 _08940_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_358 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11503__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05880__B1 _11465_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09610__A2 _09622_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11237__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11404_ _11404_/D _11686_/RN _06705_/Z _11404_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__10756__A1 _10887_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11335_ _11335_/D _11686_/RN _06705_/Z _11335_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_137_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11266_ _11266_/D _11266_/RN input68/Z _11266_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XANTENNA__09374__A1 _09374_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10217_ _10217_/A1 _10217_/A2 _10217_/A3 _10226_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11653__CLK _11665_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10508__A1 _10889_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06188__A1 _09599_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11197_ _11197_/D _11686_/RN _06705_/Z _11197_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__05935__A1 _09775_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10148_ _10148_/A1 _10001_/I _09998_/I _10148_/B2 _10149_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_10079_ _10079_/A1 _10079_/A2 _10079_/A3 _10084_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__09126__A1 _09142_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09429__A2 _09447_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_07290_ _06867_/Z _07290_/A2 _07290_/B _07291_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06310_ _05925_/Z input72/Z _06313_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06241_ _06241_/A1 _06241_/A2 _06241_/A3 _06241_/A4 _06258_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__10995__A1 _11016_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11183__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06172_ _05660_/Z _11620_/Q _08846_/A1 input62/Z _06175_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09601__A2 _09622_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11228__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06415__A2 _11071_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09931_ _10428_/B1 _11640_/Q _09932_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09365__A1 _09372_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06179__A1 _06324_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09862_ _09866_/A2 _11627_/Q _11628_/Q _09865_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_652 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_09793_ _09793_/I _11608_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05926__A1 input69/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08813_ _08820_/A2 _11299_/Q _08814_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_674 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05926__B2 input40/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input134_I wb_dat_i[13] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11400__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08744_ _07426_/Z _08759_/A2 _08744_/B _08745_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05956_ _09041_/A1 _11376_/Q _05957_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08675_ _08675_/A1 _08675_/A2 _08675_/A3 _08675_/A4 _08680_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_05887_ _05887_/A1 _05887_/A2 _05888_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10683__B1 _11519_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08340__A2 _08614_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07626_ _07626_/A1 _07626_/A2 _07631_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_26_468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07557_ _07511_/I _07614_/A1 _07558_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11526__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06508_ _06446_/I _06604_/B _11163_/Q _06668_/C _11058_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_07488_ _07552_/A1 input119/Z _07489_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_158_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06654__A2 _11059_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06439_ _06392_/Z _06439_/A2 _06439_/A3 _06439_/A4 _10935_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_09227_ _09121_/Z _09246_/A2 _09227_/B _09228_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09158_ _09158_/I _09158_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__11219__RN input162/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output186_I _06048_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10738__A1 _10921_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11676__CLK _06687_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08109_ _08616_/B _08213_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_107_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09089_ _06867_/Z _09089_/A2 _09089_/B _09090_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_174_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11120_ _11120_/D _11686_/RN _06705_/Z _11120_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__09356__A1 _09372_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11051_ _11055_/I _11698_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10002_ _10369_/A2 _11507_/Q _10006_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10910__A1 _10910_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09108__A1 _06859_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11056__CLK input68/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06342__A1 _09674_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10904_ _10904_/A1 _11156_/Q _10909_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06893__A2 _06902_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10835_ _10881_/A1 _11663_/Q _10836_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10766_ _10766_/A1 _10766_/A2 _10767_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11458__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10697_ _10924_/A1 _11327_/Q _10698_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06645__A2 input81/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10729__A1 _11528_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10729__B2 _10902_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09347__A1 _09270_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11630__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11318_ _11318_/D input76/Z _06705_/Z _11318_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__08711__I _11050_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11249_ _11249_/D _11686_/RN _06705_/Z _11249_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__11270__CLKN input68/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05810_ _06217_/I _06872_/A2 _05811_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06790_ _06790_/I _09116_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__05923__A4 _05923_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05741_ _05940_/A1 _05741_/A2 _05742_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11549__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08460_ _08460_/A1 _08460_/A2 _08460_/B _08522_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05672_ _09750_/A1 _11602_/Q _05673_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08391_ _07492_/I _08204_/I _08391_/B _08456_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07411_ _07411_/I _11247_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07342_ _07419_/A2 _06217_/Z _06871_/Z _07347_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__06884__A2 _06902_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10968__A1 _08493_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11449__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07273_ _07273_/I _11198_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11699__CLK input68/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06224_ _06224_/A1 _06224_/A2 _06224_/A3 _06224_/A4 _06235_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_09012_ _09013_/A2 _11362_/Q _09013_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08389__A2 _08395_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06155_ _06155_/A1 _06155_/A2 _06156_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10196__A2 _10351_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11621__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06086_ _08761_/A1 _11287_/Q _06087_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09338__A1 _09158_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09914_ _11638_/Q _10407_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09845_ _09241_/I _09848_/A2 _09845_/B _09846_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11079__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_09776_ _09798_/A2 _11603_/Q _09777_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06988_ _06974_/I _11125_/Q _06989_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05939_ _05939_/A1 _05939_/A2 _05939_/A3 _05939_/A4 _05968_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_08727_ _08740_/A2 _11273_/Q _08728_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08313__A2 _08686_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06324__A1 _06324_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08658_ _08658_/A1 _08658_/A2 _08662_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09510__A1 _09154_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07609_ _07609_/I _07609_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_169_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08589_ _08589_/A1 _08677_/A2 _08590_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08077__A1 _08161_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10620_ _10891_/A1 _11478_/Q _10622_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06627__A2 input77/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10551_ _10551_/A1 _10551_/A2 _10552_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10482_ _10414_/I _10427_/B _10892_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_154_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09329__A1 _09121_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11612__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11103_ _11103_/D _11686_/RN _06705_/Z _11103_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_11034_ _11038_/A2 _11685_/Q _11035_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08552__A2 _08692_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06315__A1 _05660_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09501__A1 _09116_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10647__B1 _10920_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11679__RN input162/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10818_ _10910_/A1 _11570_/Q _10820_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10749_ _10914_/B1 _11609_/Q _10750_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05826__B1 _11450_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09568__A1 _09572_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10178__A2 _10369_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput216 _06689_/Z mgmt_gpio_out[14] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput205 _06727_/ZN mgmt_gpio_oeb[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput227 _11093_/Q mgmt_gpio_out[24] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput238 _11311_/Q mgmt_gpio_out[34] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__08240__A1 _07837_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10192__B _10880_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput249 _06713_/ZN pad_flash_clk VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_07960_ _08355_/I _08375_/B _07963_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11221__CLK _11683_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08791__A2 _08825_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06911_ _06911_/I _11102_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07891_ _07891_/I _07930_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06003__B1 _11543_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09630_ _09630_/I _11556_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11371__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06842_ _06842_/I _11079_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09561_ _09561_/I _11534_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06773_ _07110_/I _11064_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08512_ _08512_/I _08572_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_82_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05724_ _11338_/Q _10272_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_70_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09492_ _09492_/I _11512_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10102__A2 _10359_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06306__A1 _05584_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08443_ _08443_/A1 _08558_/A1 _08608_/A3 _08448_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_05655_ _08825_/A2 _08799_/A2 _05656_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__06857__A2 _06869_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08374_ _08371_/Z _08445_/A1 _08554_/B _08376_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_05586_ _11063_/Q _06490_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07806__A1 _08696_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10405__A3 _09920_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07325_ _07325_/A1 _07325_/A2 _11212_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07256_ _06855_/Z _07265_/A2 _07256_/B _07257_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11622__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10810__B1 _11522_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11042__I _11050_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09559__A1 _09572_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06207_ _05693_/Z _11524_/Q _06211_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_155_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07187_ _07197_/A1 _07187_/A2 _07187_/B _07188_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10169__A2 _11431_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06138_ input45/Z _05927_/I _07201_/A1 input54/Z _06141_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08231__B2 _08656_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08231__A1 _08434_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11637__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input62_I mgmt_gpio_in[33] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07034__A2 _06217_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06069_ _11542_/Q _10634_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05596__A2 _05633_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09828_ _09828_/I _11619_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09759_ _09759_/I _11597_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08298__A1 _07586_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05520__A2 _06610_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11652_ _11652_/D input76/Z _11665_/CLK _11652_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__09798__A1 _09270_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10603_ _10603_/A1 _10603_/A2 _10603_/A3 _10603_/A4 _10604_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_80_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11583_ _11583_/D _11686_/RN _06705_/Z _11583_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__11244__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10534_ _10904_/A1 _11548_/Q _10537_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10465_ _10389_/I _10427_/B _10894_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_6_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08222__A1 split7/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10396_ _10425_/A2 _10428_/B1 _10406_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_145_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05587__A2 _05515_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11394__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09722__A1 _09270_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11017_ _08493_/B input154/Z _11019_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07605__I _07605_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10096__A1 _10352_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06839__A2 _06838_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09789__A1 _09158_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07110_ _07110_/I _11163_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08461__A1 split12/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08090_ _08090_/A1 _08090_/A2 _08094_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07041_ _07412_/A1 _06217_/Z _06871_/Z _07046_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_133_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10020__A1 _10357_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05578__A2 _06786_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10571__A2 _11413_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08992_ _07426_/Z _09013_/A2 _08992_/B _08993_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07943_ _08557_/B _08352_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_68_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07874_ _07874_/A1 _06587_/I _07876_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09713__A1 _09158_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09613_ _09158_/Z _09622_/A2 _09613_/B _09614_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06825_ _06825_/I _11076_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_43_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09544_ _09241_/Z _09547_/A2 _09544_/B _09545_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06756_ _06760_/A1 _08036_/B _06757_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11117__CLK _11672_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05750__A2 _06396_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06687_ _11304_/Q _06687_/A2 _06688_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09475_ _09497_/A2 _11507_/Q _09476_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05707_ _05707_/I _09649_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XANTENNA__10087__A1 _10087_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08426_ _08426_/A1 _08280_/B _08544_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05638_ _05638_/I _05924_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
X_08357_ _08359_/B _08357_/A2 _08357_/B _08439_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05569_ _05569_/I _11691_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06058__A3 _06058_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08288_ _08614_/A2 _08623_/A2 _08294_/B _08290_/C _08289_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_07308_ _07308_/I _11207_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07239_ _07240_/A1 _11188_/Q _07240_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10250_ _10367_/A1 _11481_/Q _10251_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10011__A1 _10030_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output266_I _11275_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08755__A2 _11282_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10181_ _10181_/A1 _10181_/A2 _10181_/A3 _10189_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__10560__B _10880_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09704__A1 _09121_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06518__A1 _06518_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07191__A1 _07197_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10078__A1 _10374_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11704_ input88/Z _11704_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08256__I split21/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11635_ _11635_/D _11686_/RN _11658_/CLK _11635_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_11566_ _11566_/D _11686_/RN _06705_/Z _11566_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_128_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10250__A1 _10367_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10517_ _10517_/A1 _10517_/A2 _10518_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08205__B split12/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11497_ _11497_/D _11686_/RN _06705_/Z _11497_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_143_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10002__A1 _10369_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10448_ _10903_/A1 _11555_/Q _10449_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10379_ _10379_/A1 _11152_/Q _10380_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10553__A2 _11412_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10305__A2 _06556_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09171__A2 _09015_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07182__A1 _07197_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07590_ _07590_/A1 _08095_/A2 _07591_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06610_ _05509_/I _06610_/A2 _06610_/A3 _06610_/B _11163_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__10069__A1 _10366_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06541_ _09865_/A2 _06541_/A2 _06542_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06472_ _06478_/A2 _06466_/B _06473_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09260_ _09260_/I _11438_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08211_ _08211_/A1 _08471_/B _08570_/A2 _08216_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__05496__A1 _05969_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11018__B1 _08460_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09191_ _09195_/A2 _11417_/Q _09192_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08142_ _08142_/A1 _08142_/A2 _08478_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11033__A3 _06838_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08434__A1 _08434_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07237__A2 _09270_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08073_ _08073_/I _08200_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__08985__A2 _08988_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05799__A2 _11506_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06996__A1 _06974_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07024_ _07025_/A2 _11136_/Q _07025_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10792__A2 _11434_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input164_I wb_sel_i[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08975_ _08988_/A2 _11350_/Q _08976_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07926_ _07926_/I _08355_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA_input25_I mask_rev_in[29] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09162__A2 _11408_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07857_ _07857_/A1 _07857_/A2 _07857_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_06808_ _11678_/Q _10993_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07788_ _08592_/A2 _08592_/B _07789_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09527_ _09527_/I _11523_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06739_ input69/Z input95/Z _06740_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XPHY_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_358 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_09458_ _09458_/I _11501_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_169_335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08673__A1 _08673_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09389_ _09389_/I _11479_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08409_ _08409_/A1 _08626_/A2 _08412_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_8_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07228__A2 _05924_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11420_ _11420_/D input76/Z _06705_/Z _11420_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_177_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08976__A2 _08988_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11351_ _11351_/D _11686_/RN _06705_/Z _11351_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10302_ _10302_/A1 _10302_/A2 _10302_/A3 _10303_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_125_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06987__A1 _10947_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11282_ _11282_/D _11686_/RN _06705_/Z _11282_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_10_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06739__A1 input69/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10233_ _10350_/A1 _10233_/A2 _10234_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_126_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10164_ _11383_/Q _10355_/A2 _11375_/Q _10355_/B2 _10164_/C _10173_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__10299__A1 _10377_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11453__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07155__I _11050_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10095_ _10353_/A1 _11365_/Q _10097_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07164__A1 _05925_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11432__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08900__A2 _11326_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10997_ _08431_/B input133/Z _08460_/B input142/Z _10998_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11468__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11582__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1083 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1061 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1050 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_182 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1094 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_11618_ _11618_/D _11686_/RN _06705_/Z _11618_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__08714__I _11050_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10223__A1 _10374_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08967__A2 _08988_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11549_ _11549_/D _11686_/RN _06705_/Z _11549_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__06978__A1 _10938_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05650__A1 _08795_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_801 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08719__A2 _08719_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_823 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_867 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_856 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_845 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_878 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_08760_ _08760_/I _11283_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05972_ _10950_/A1 _06304_/A2 _06619_/B _05972_/C _05974_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08691_ _08691_/A1 _08691_/A2 _08691_/A3 _08700_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_07711_ _07711_/A1 _07711_/A2 _07718_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09144__A2 _09015_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07642_ _07642_/A1 _08628_/C _07647_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06902__A1 _06867_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11191__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07573_ _08248_/B _08509_/A1 _08258_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09312_ _09322_/A2 _11455_/Q _09313_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06524_ _06524_/I _11159_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06130__A2 _11557_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06455_ _06455_/I _11069_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09243_ _09241_/Z _09246_/A2 _09243_/B _09244_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10462__A1 _10921_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06386_ _09499_/A1 _11515_/Q _06390_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09174_ _09174_/I _11411_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10214__B2 _11504_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08125_ _08125_/A1 _08696_/C _08130_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11050__I _11050_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09080__A1 _06855_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11305__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08056_ _07995_/I _07675_/B _08057_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07630__A2 _08509_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05641__A1 _08825_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07007_ _07011_/A2 _11131_/Q _07008_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput105 wb_adr_i[17] input105/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput116 wb_adr_i[27] _06595_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput127 wb_adr_i[8] input127/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11455__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput149 wb_dat_i[27] input149/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput138 wb_dat_i[17] input138/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08958_ _08958_/I _11344_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07909_ _07909_/I _08361_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_08889_ _08889_/I _11322_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09135__A2 _11400_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10920_ _10920_/A1 _11104_/Q _10920_/B1 _11106_/Q _10923_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10150__B1 _09965_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08894__A1 _08913_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10851_ _11228_/Q _10897_/A2 _10897_/B1 _11232_/Q _10852_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11182__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10782_ _10920_/A1 _11345_/Q _10920_/B1 _11353_/Q _10785_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_52_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_11403_ _11403_/D _11686_/RN _06705_/Z _11403_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_125_213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10756__A2 _11425_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09071__A1 _07431_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07621__A2 _08417_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06054__I _11438_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11334_ _11334_/D _11686_/RN _06705_/Z _11334_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_11265_ _11265_/D _11265_/RN input68/Z _11265_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XANTENNA__09374__A2 _09015_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10216_ _10370_/A1 _11496_/Q _10217_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10508__A2 _11403_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11196_ _11196_/D _11686_/RN _06705_/Z _11196_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10147_ _11574_/Q _10377_/A1 _11566_/Q _10377_/B1 _10147_/C _10152_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_153_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10078_ _10374_/A1 _11532_/Q _10079_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08885__A1 _06863_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11173__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10692__A1 _10921_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08637__A1 _07566_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10444__A1 _10444_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06240_ _07370_/A1 _06238_/Z _11237_/Q _06241_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11328__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06112__A2 _11304_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_06171_ input47/Z _05924_/I _05925_/I input73/Z _06175_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_171_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07612__A2 _08509_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09930_ _11641_/Q _10428_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__11478__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09861_ _09861_/I _11628_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_642 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_09792_ _09187_/I _09798_/A2 _09792_/B _09793_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05926__A2 _05924_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08812_ _08812_/I _11298_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_675 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_08743_ _08759_/A2 _11278_/Q _08744_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05955_ _09016_/A1 _11368_/Q _05957_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09117__A2 _09015_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input127_I wb_adr_i[8] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08674_ _07566_/I _07537_/I _08674_/B _08675_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08876__A1 _06851_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05886_ _09171_/A1 _11417_/Q _05887_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10683__B2 _10902_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11045__I _11050_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11164__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07625_ _08686_/B _08686_/A2 _07626_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07556_ _08589_/A1 _08345_/A2 _08403_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08628__A1 _08355_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06507_ _11058_/Q _06668_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_34_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07487_ _07487_/I _07552_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10986__A2 _10966_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07300__A1 _05616_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input92_I spimemio_flash_io3_do VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09226_ _09246_/A2 _11428_/Q _09227_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06438_ _06438_/A1 _06438_/A2 _06438_/A3 _06438_/A4 _06439_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XANTENNA__05862__A1 _09549_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09157_ _09157_/I _11406_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06369_ _06217_/Z _11033_/A2 _11137_/Q _06370_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_08108_ _08108_/A1 _08108_/A2 _08113_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09088_ _09089_/A2 _11386_/Q _09089_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output179_I _06731_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08039_ _08039_/I _08167_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_11050_ _11050_/I _11697_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10001_ _10001_/I _10369_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__10910__A2 _11262_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09108__A2 _09114_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08867__A1 _07426_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10903_ _10903_/A1 _11152_/Q _10909_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11155__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10834_ _10092_/Z _11662_/Q _10834_/B _10880_/C _10836_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08095__A2 _08095_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10765_ _10892_/A1 _11473_/Q _10766_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10696_ _10696_/A1 _10696_/A2 _10696_/A3 _10696_/A4 _10696_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__11620__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05853__A1 _06396_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10729__A2 _10902_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11317_ _11317_/D input76/Z _06705_/Z _11317_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_4_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09347__A2 _09347_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11248_ _11248_/D _11686_/RN _06705_/Z _11248_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__07358__A1 _07076_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11179_ _11179_/D _11686_/RN _06705_/Z _11179_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__06030__A1 _09800_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11394__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05740_ _05740_/I _06398_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__11146__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05671_ _05636_/I _05726_/I _09750_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__10665__A1 _10887_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08390_ _08560_/I _08390_/A2 _08390_/A3 _08613_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11150__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07410_ _07081_/Z _07410_/A2 _07410_/B _07411_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07341_ _07341_/I _11227_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07272_ _07081_/Z _07290_/A2 _07272_/B _07273_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_12_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06223_ _08825_/A1 _11233_/Q _06217_/Z _06224_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11284__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05844__A1 _08761_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09011_ _09011_/I _11361_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09035__A1 _09039_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08389__A3 _08656_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06154_ _09449_/A1 _11501_/Q _06155_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10653__B _10653_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06085_ _06839_/A1 _11082_/Q _06087_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09338__A2 _09347_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09913_ _10394_/A2 _11638_/Q _09916_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09844_ _09848_/A2 _11625_/Q _09845_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11385__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09775_ _09775_/A1 _09015_/I _09798_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__06572__A2 _08036_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06987_ _10947_/A1 _06990_/A2 _06989_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_160_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05938_ _05938_/A1 _05938_/A2 _05938_/A3 _05938_/A4 _05939_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_08726_ _08726_/A1 _06904_/Z _08740_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_73_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05869_ _06324_/A1 _11593_/Q _05871_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10656__A1 _10914_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08657_ _08657_/A1 _08657_/A2 _08657_/A3 _08658_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__09510__A2 _09522_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11137__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07608_ _08625_/B _08247_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_26_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08588_ _08588_/A1 _08588_/A2 _08588_/A3 _08638_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_169_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07539_ _08249_/B _07539_/A2 _07539_/A3 _07544_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__06088__A1 _08803_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11643__CLK _11665_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output296_I _11086_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10550_ _10886_/B2 _11388_/Q _10551_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10481_ _10897_/A2 _11451_/Q _10486_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09026__A1 _09039_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05835__A1 _08839_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09209_ _09209_/I _11422_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10592__B1 _10916_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09329__A2 _09347_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06260__A1 _06396_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11102_ _11102_/D _11686_/RN _06705_/Z _11102_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_11033_ _05703_/Z _11033_/A2 _06838_/Z _11038_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_78_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06012__A1 _09449_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10895__A1 _10895_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11376__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11173__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09501__A2 _09522_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10647__A1 _10920_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10647__B2 _11350_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06315__A2 _11619_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10817_ _10817_/A1 _10817_/A2 _10817_/A3 _10817_/A4 _10826_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__09265__A1 _09187_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07815__A2 _08495_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10748_ _10914_/A1 _11601_/Q _10750_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11300__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09017__A1 _09039_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10679_ _10679_/A1 _10679_/A2 _10679_/A3 _10679_/A4 _10691_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xoutput217 _06685_/Z mgmt_gpio_out[15] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput206 _06082_/A1 mgmt_gpio_oeb[5] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput228 _11094_/Q mgmt_gpio_out[25] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput239 _06652_/ZN mgmt_gpio_out[35] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__08240__A2 _07492_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06251__A1 _07427_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08791__A3 _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06910_ _06843_/Z _06910_/A2 _06910_/B _06911_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07890_ _07890_/A1 _07890_/A2 _07890_/B _07891_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06003__B2 _09574_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11516__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11367__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06841_ _06837_/Z _06869_/A2 _06841_/B _06842_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10886__B2 _10886_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09560_ _09154_/Z _09572_/A2 _09560_/B _09561_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06772_ _07110_/I _11063_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09491_ _09187_/Z _09497_/A2 _09491_/B _09492_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08511_ _07572_/I _07802_/I _08511_/B _08511_/C _08675_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__10638__A1 _10638_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11119__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05723_ _05723_/I _05723_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08442_ _08442_/A1 _07920_/I _08442_/B _08442_/C _08608_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08700__B1 _11016_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11666__CLK _11666_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05654_ _05645_/I _05669_/I _08799_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_90_180 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08373_ split8/Z _07959_/I _08373_/B _08554_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05585_ _11205_/Q _05616_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XANTENNA__09256__A1 _09125_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07324_ _07310_/I _11212_/Q _07325_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07255_ _07265_/A2 _11193_/Q _07256_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10810__A1 _11530_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05817__A1 _06217_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10810__B2 _10902_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06206_ _06206_/A1 _06206_/A2 _06206_/A3 _06206_/A4 _06212_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__09559__A2 _11534_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07186_ _07197_/A1 _11178_/Q _07187_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_172_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08231__A2 _08380_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06137_ input58/Z _05924_/I _05925_/I input37/Z _06141_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07034__A3 _06871_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06242__A1 _09399_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06068_ _11550_/Q _10146_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input55_I mgmt_gpio_in[27] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08788__B _11292_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11196__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09827_ _09116_/I _09848_/A2 _09827_/B _09828_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07742__A1 _08589_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11358__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09758_ _09125_/I _09773_/A2 _09758_/B _09759_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_285 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10629__A1 _10900_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08709_ _07431_/Z _08709_/A2 _08709_/B _08710_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08298__A2 _08495_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09689_ _09689_/I _11575_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_output309_I _06725_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11530__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11651_ _11651_/D input76/Z _11665_/CLK _11651_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_11582_ _11582_/D _11686_/RN _06705_/Z _11582_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__09798__A2 _09798_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10602_ _10906_/A1 _11541_/Q _10603_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10533_ _10906_/A1 _11540_/Q _10537_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_167_285 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_435 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10464_ _10894_/A2 _11491_/Q _10467_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10395_ _10484_/A1 _09934_/I _10914_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_6_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11539__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06233__A1 _06217_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05992__B1 _08940_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09722__A2 _09722_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11016_ _11016_/A1 input159/Z _11019_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10868__A1 _10914_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08717__I _11050_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11521__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09238__A1 _09246_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09789__A2 _09798_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11069__CLK input68/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08461__A2 _08614_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07040_ _07040_/I _11140_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09410__A1 _09154_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10020__A2 _11411_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08991_ _09013_/A2 _11355_/Q _08992_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07942_ _07942_/A1 _07942_/A2 _07947_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07873_ _07880_/A1 _08012_/A1 _07873_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__09713__A2 _09722_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10859__A1 _10905_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09612_ _09622_/A2 _11551_/Q _09613_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06824_ _06835_/A1 _09187_/I _06824_/B _06825_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09543_ _09547_/A2 _11529_/Q _09544_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06755_ _06755_/I _06755_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09474_ _09474_/A1 _09015_/Z _09497_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_06686_ _11179_/Q _06688_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05706_ _05703_/I _08799_/A2 _05707_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10087__A2 _06556_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11512__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05637_ _07419_/A2 _08825_/A2 _05638_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08425_ _08425_/A1 _08425_/A2 _08428_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06160__B1 _11413_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09229__A1 _09246_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08356_ _08351_/I _08686_/A1 _08436_/B _08437_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05568_ _06786_/A1 _05519_/I _05568_/B _05569_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07307_ _07081_/Z _07307_/A2 _07307_/B _07308_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08287_ _08540_/A3 _08630_/B _08630_/C _08292_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05499_ _05499_/I _11702_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07238_ _11322_/Q _05924_/Z _07238_/B _07240_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09401__A1 _09116_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07169_ _05925_/Z _09125_/I _07170_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10011__A2 _10265_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10180_ _10370_/A1 _11495_/Q _10181_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09704__A2 _09722_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06518__A2 _06266_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09468__A1 _09472_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11503__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11211__CLK _11656_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11027__A1 _11027_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11634_ _11634_/D _11686_/RN _11658_/CLK _11634_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__09640__A1 _09647_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11565_ _11565_/D _11686_/RN _06705_/Z _11565_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_11496_ _11496_/D _11686_/RN _06705_/Z _11496_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10516_ _10916_/A1 _11620_/Q _10517_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11361__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10447_ _10884_/A1 _11379_/Q _10449_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07954__A1 split15/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10378_ _10378_/A1 _11156_/Q _10380_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_151_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07616__I _07616_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06509__A2 _11057_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09459__A1 _09472_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06540_ _11630_/Q _06541_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_33_320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11636__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06471_ _06469_/Z _06471_/A2 _11067_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08210_ _08434_/A1 _08659_/A1 _08209_/B _08332_/A1 _08570_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11018__A1 _08431_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10926__B _10926_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09190_ _09190_/I _11416_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09631__A1 _09647_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08141_ _08141_/A1 _08618_/C _08147_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08072_ _08106_/A1 _08148_/A2 _08073_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07023_ _07023_/I _11135_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08198__A1 split12/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07945__A1 split21/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input157_I wb_dat_i[5] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08974_ _08974_/I _11349_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07925_ split21/I _08367_/B _08442_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11048__I _11050_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07856_ input127/Z split16/I _07857_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08370__A1 split8/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07787_ _08328_/B1 _08505_/B _08320_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11234__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input18_I mask_rev_in[22] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06807_ _06807_/I _11073_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06738_ _11590_/Q _06738_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09526_ _09116_/Z _09547_/A2 _09526_/B _09527_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09457_ _09125_/Z _09472_/A2 _09457_/B _09458_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06684__A1 _11305_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08673__A2 _08460_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08408_ _08419_/A1 _07596_/I _08408_/B _08408_/C _08626_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__11009__A1 _11016_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_06669_ _11058_/Q input38/Z _11056_/Q _06671_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09388_ _09158_/Z _09397_/A2 _09388_/B _09389_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10480__A2 _10427_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11384__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09622__A1 _09270_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08339_ _08339_/A1 _08347_/A1 _08339_/B _08641_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_11350_ _11350_/D _11686_/RN _06705_/Z _11350_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10301_ _10379_/A1 _11562_/Q _10302_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11281_ _11281_/D _11686_/RN _06705_/Z _11281_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_105_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07936__A1 _08355_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10232_ _11652_/Q _10305_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10163_ _10163_/A1 _10163_/A2 _10164_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10094_ _11349_/Q _10351_/A2 _11341_/Q _10351_/B2 _10094_/C _10107_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__07164__A2 _09121_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06372__B1 _07427_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_253 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10996_ _08493_/B input150/Z _10998_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1040 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1073 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1062 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1051 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1095 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1084 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10471__A2 _10406_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09613__A1 _09158_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11617_ _11617_/D _11686_/RN _06705_/Z _11617_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_30_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11548_ _11548_/D _11686_/RN _06705_/Z _11548_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__10759__B1 _11409_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11479_ _11479_/D _11686_/RN _06705_/Z _11479_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_143_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11107__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05650__A2 _08825_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08719__A3 _06838_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_835 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07927__A1 _08355_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_868 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_857 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_07710_ _07710_/A1 _08430_/A2 _07711_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11257__CLK _11683_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_879 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05971_ _06304_/A2 _06040_/A1 _05972_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08690_ _08690_/A1 _08690_/A2 _08690_/A3 _08690_/A4 _08691_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_07641_ _07643_/I _08686_/A2 _08628_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_25_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07572_ _07572_/I _08509_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XANTENNA__06902__A2 _06902_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07081__I _09121_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09311_ _09311_/I _11454_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06523_ _06610_/A3 _06611_/B2 _06523_/B _06524_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_15_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09852__A1 _10092_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09242_ _09246_/A2 _11433_/Q _09243_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06454_ _06454_/A1 _06454_/A2 _06455_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09604__A1 _09121_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06385_ _06385_/A1 _06385_/A2 _06385_/A3 _06385_/A4 _06391_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_09173_ _09116_/Z _09195_/A2 _09173_/B _09174_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10214__A2 _10369_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08124_ split8/I _08126_/I _08696_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09080__A2 _09089_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08055_ _08055_/A1 _08055_/A2 _08084_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05641__A2 _08839_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07006_ _07419_/A2 _07006_/A2 _06871_/Z _07011_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
Xinput117 wb_adr_i[28] _06597_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput106 wb_adr_i[18] input106/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_142_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput139 wb_dat_i[18] input139/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput128 wb_adr_i[9] input128/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08957_ _06859_/Z _08963_/A2 _08957_/B _08958_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07908_ _07930_/A1 _07981_/A2 _07909_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08888_ _06867_/Z _08888_/A2 _08888_/B _08889_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07146__A2 _05927_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07839_ _07989_/A1 _07839_/A2 _07840_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10150__A1 _10634_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10150__B2 _10634_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10410__I _10410_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10850_ _10896_/A1 _11143_/Q _10852_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08894__A2 _11324_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09509_ _09522_/A2 _11518_/Q _09510_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_169_111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10781_ _10919_/A1 _11369_/Q _10785_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_145 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08036__B _08036_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11402_ _11402_/D _11686_/RN _06705_/Z _11402_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__06409__A1 _08795_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10205__A2 _11432_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09071__A2 _09089_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11333_ _11333_/D _11686_/RN _06705_/Z _11333_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__05632__A2 _05515_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11264_ _11264_/D _11264_/RN input68/Z _11264_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
X_10215_ _10371_/A1 _11488_/Q _10217_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11195_ _11195_/D _11686_/RN _06705_/Z _11195_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_133_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10146_ _09972_/I _10146_/A2 _09876_/I _10146_/B1 _09975_/I _10147_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_10077_ _10375_/A1 _11540_/Q _10079_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07137__A2 _07151_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06896__A1 _06859_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08885__A2 _08888_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10979_ _10979_/A1 _10966_/Z _10979_/B _10980_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10444__A2 _10506_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06648__A1 input80/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06170_ _06170_/A1 _06170_/A2 _11265_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09860_ _09868_/A1 _09860_/A2 _09938_/A2 _09866_/A2 _09861_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__07076__I _09116_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_09791_ _09798_/A2 _11608_/Q _09792_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08811_ _06847_/Z _08820_/A2 _08811_/B _08812_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_654 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_08742_ _08742_/A1 _06904_/Z _08759_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_05954_ _11392_/Q _09091_/A1 _09066_/A1 _11384_/Q _05957_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_687 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08325__A1 _08686_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08673_ _08673_/A1 _08460_/B _08493_/B _08673_/B2 _08673_/C _08682_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_07624_ _07640_/A1 _07657_/A2 _08686_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06887__A1 _06847_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08876__A2 _08888_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05885_ _09197_/A1 _11425_/Q _05887_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10683__A2 _10902_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09825__A1 _05660_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07555_ _07555_/I _08345_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_13_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07486_ _07663_/A1 _07690_/A2 _07486_/A3 _08249_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__10435__A2 _09934_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06506_ _11160_/Q _06604_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09225_ _09225_/I _11427_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06437_ _06437_/A1 _06437_/A2 _06437_/A3 _06437_/A4 _06438_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA_input85_I spimemio_flash_csb VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11452__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09156_ _09154_/Z _09169_/A2 _09156_/B _09157_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06368_ _07370_/A1 _11135_/Q _06217_/Z _06370_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__07064__A1 _06837_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08107_ split8/I _08616_/B _08108_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09087_ _09087_/I _11385_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11422__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08800__A2 _11295_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06299_ _07398_/A1 _07006_/A2 _11108_/Q _06301_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_08038_ split12/I _08423_/A2 _08573_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__06811__A1 _06835_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11467__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11572__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10000_ _10000_/A1 _10040_/A2 _10001_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10371__A1 _10371_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09989_ _09896_/I _09878_/I _10367_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_88_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08867__A2 _08888_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10902_ _11154_/Q _10902_/A2 _11150_/Q _10902_/B2 _10902_/C _10909_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__09816__A1 _09823_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11405__SETN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10833_ _10833_/A1 _10092_/Z _10831_/Z _10833_/A4 _10834_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_10764_ _10891_/A1 _11481_/Q _10766_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_10695_ _10919_/A1 _11367_/Q _10696_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_172_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07055__A1 _05703_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11316_ _11316_/D _11686_/RN _06705_/Z _11316_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__11091__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11247_ _11247_/D _11686_/RN _06705_/Z _11247_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_11178_ _11178_/D _11686_/RN _06705_/Z _11178_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10129_ _10129_/I _11648_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10114__A1 _10371_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05670_ _05940_/A2 _05699_/A2 _05726_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__06869__A1 _06867_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10665__A2 _11431_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09807__A1 _09823_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07340_ _07081_/Z _07340_/A2 _07340_/B _07341_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07294__A1 _08672_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07271_ _07290_/A2 _11198_/Q _07272_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11445__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06097__A2 _06396_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09010_ _06863_/Z _09013_/A2 _09010_/B _09011_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_163_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06222_ _07419_/A2 _11229_/Q _06217_/Z _06224_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06153_ _09424_/A1 _11493_/Q _06155_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07046__A1 _06843_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11595__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10653__C _10880_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06084_ _06785_/A1 _11074_/Q _06087_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07349__A2 _06904_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09912_ _09912_/I _10394_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_09843_ _09843_/I _11624_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10353__A1 _10353_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06021__A2 _11431_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_462 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_09774_ _09774_/I _11602_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06986_ _06986_/I _11124_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05780__A1 _06238_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05937_ _09750_/A1 _11600_/Q _05938_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08725_ _08725_/I _11272_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05868_ _05868_/A1 _05868_/A2 _05868_/A3 _05868_/A4 _05894_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_08656_ _08656_/A1 _08696_/A2 _08656_/B _08657_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08587_ _07609_/Z _08592_/A2 _08587_/B _08588_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07607_ _07607_/A1 _07527_/I _08625_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05799_ _09449_/A1 _11506_/Q _05800_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07538_ _08294_/C _08592_/A2 _07539_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09274__A2 _09015_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07469_ _07689_/A2 _07689_/A1 _07540_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10480_ _10480_/A1 _10427_/B _10897_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA_output191_I _10634_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09026__A2 _11366_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05835__A2 _11033_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09208_ _09154_/Z _09220_/A2 _09208_/B _09209_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output289_I _11087_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09139_ _06863_/Z _09142_/A2 _09139_/B _09140_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09982__B1 _10377_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07588__A2 _08509_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10592__B2 _11621_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10592__A1 _10915_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11101_ _11101_/D _11686_/RN _06705_/Z _11101_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_118_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11032_ _11032_/A1 _11032_/A2 _11032_/B1 _07300_/C _11684_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08537__A1 _08686_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10895__A2 _11227_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11318__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11468__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10816_ _10816_/I _10817_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_13_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09265__A2 _09272_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10747_ _10747_/A1 _10747_/A2 _11661_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10678_ _11455_/Q _10897_/A2 _10897_/B1 _11463_/Q _10679_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xoutput207 _10137_/B2 mgmt_gpio_oeb[6] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput229 _11095_/Q mgmt_gpio_out[26] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput218 _11164_/Q mgmt_gpio_out[16] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__06251__A2 _11253_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08791__A4 _06904_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06003__A2 _09599_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10335__A1 _10374_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07200__A1 _08865_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06840_ _06869_/A2 _11079_/Q _06841_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10886__A2 _10886_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06771_ _07110_/I _11062_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05762__A1 _11330_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05762__B2 _08761_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09490_ _09497_/A2 _11512_/Q _09491_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08510_ _08510_/A1 _08596_/A1 _08516_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10638__A2 _10416_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05722_ _07006_/A2 _05805_/A2 _05723_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08441_ _08442_/A1 _08607_/B _08441_/B _08441_/C _08558_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08700__A1 _08431_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08700__B2 _08700_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05653_ _05605_/I _05610_/I _05669_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08372_ _08351_/I _08686_/A1 _08444_/B _08445_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05584_ _05584_/I _06619_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XANTENNA__09256__A2 _09272_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07323_ _10947_/A1 _07326_/A2 _07325_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07254_ _07254_/I _11192_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10810__A2 _10902_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05817__A2 _08839_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06205_ _05703_/Z _08825_/A1 _11247_/Q _06206_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_07185_ _11202_/Q _05925_/Z _07185_/B _07187_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06136_ _11549_/Q _09599_/A1 _11541_/Q _09574_/A1 _06136_/C _06148_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__10574__A1 _10897_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06067_ _06067_/A1 _06067_/A2 _06067_/A3 _06099_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_input48_I mgmt_gpio_in[20] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09192__A1 _06863_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09826_ _09848_/A2 _11619_/Q _09827_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_3_5__f_wb_clk_i_I clkbuf_0_wb_clk_i/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07742__A2 _08490_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09757_ _09773_/A2 _11597_/Q _09758_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06969_ _06969_/I _11119_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11610__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10629__A2 _11510_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08708_ _08709_/A2 _11262_/Q _08709_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09688_ _09158_/I _09697_/A2 _09688_/B _09689_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output204_I _06726_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08639_ _07566_/I _07537_/I _08639_/B _08640_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_11650_ _11650_/D input76/Z _11665_/CLK _11650_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_11581_ _11581_/D _11686_/RN _06705_/Z _11581_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__07258__A1 _07265_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10601_ _10904_/A1 _11549_/Q _10603_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10532_ _10532_/A1 _10532_/A2 _10532_/A3 _10532_/A4 _10548_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_80_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08470__A3 _08586_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11294__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10463_ _10463_/A1 _10427_/B _10894_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__08758__A1 _08759_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10394_ _10460_/A1 _10394_/A2 _10484_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__10565__A1 _10884_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06233__A2 _11033_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11140__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11015_ _11015_/I _11681_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10317__A1 _10356_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10868__A2 _11238_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11290__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09238__A2 _11432_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07249__A1 _07265_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08997__A1 _09013_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06472__A2 _06466_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08749__A1 _08759_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10005__B1 _10371_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09410__A2 _09422_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07421__A1 _07076_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08990_ _08990_/A1 _06838_/Z _09013_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_07941_ split6/I _08557_/B _07942_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11633__CLK _11658_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05983__A1 _08761_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07872_ _07872_/I _08012_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09611_ _09611_/I _11550_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_18_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06823_ _06835_/A1 _11076_/Q _06824_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_09542_ _09542_/I _11528_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06754_ _06514_/B _06754_/A2 _06754_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05705_ _05705_/I _09674_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_83_468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09473_ _09473_/I _11506_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06685_ _06685_/I _06685_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08424_ _08540_/A1 _08540_/A2 _08540_/A4 _08425_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05636_ _05636_/I _08825_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_4
XANTENNA_input102_I wb_adr_i[14] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06160__A1 _11421_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05567_ _05519_/I _11691_/Q _05568_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08355_ _08355_/I _08686_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__06160__B2 _09171_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08988__A1 _06867_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07306_ _07307_/A2 _11207_/Q _07307_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08286_ _08294_/B _08395_/A2 _08280_/B _08630_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_109_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05498_ _06786_/A1 _05498_/A2 _05498_/B _05499_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11276__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10795__A1 _10883_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07237_ _05924_/Z _09270_/I _07238_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11163__CLK input68/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07168_ _07168_/I _11174_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09401__A2 _09422_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07412__A1 _07412_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06119_ _11325_/Q _08890_/A1 _06119_/B _06119_/C _06128_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_182_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07099_ _07099_/A1 _06904_/Z _07104_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09165__A1 _09169_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09809_ _09809_/I _11613_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08912__A1 _08913_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11200__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07722__I _07722_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09468__A2 _11505_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11702_ _11702_/D _11702_/RN input68/Z _11702_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__11027__A2 _08036_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11633_ _11633_/D _11686_/RN _11658_/CLK _11633_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_24_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08979__A1 _06855_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09640__A2 _11560_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11506__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11564_ _11564_/D _11686_/RN _06705_/Z _11564_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__10786__A1 _10924_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11495_ _11495_/D _11686_/RN _06705_/Z _11495_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10515_ _10914_/B1 _11604_/Q _10517_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10446_ _10904_/A1 _11547_/Q _10449_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07403__A1 _07081_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10538__A1 _11508_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11656__CLK _11656_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08600__B1 _08623_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10377_ _10377_/A1 _11146_/Q _10377_/B1 _11262_/Q _10380_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_2_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05965__A1 _08940_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09156__A1 _09154_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08903__A1 _08913_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10710__A1 _10887_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06142__A1 _09775_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06470_ _06470_/A1 _06468_/Z _06471_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08140_ _08140_/I _08618_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_119_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11186__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09631__A2 _11557_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10777__A1 _10900_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11258__RN input162/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08071_ _08071_/I _08148_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_119_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07022_ _06837_/Z _07025_/A2 _07022_/B _07023_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08198__A2 _08242_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10529__A1 _10897_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05956__A1 _09041_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08973_ _06847_/Z _08988_/A2 _08973_/B _08974_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07924_ split15/I _08367_/B _08365_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11430__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07855_ _07855_/A1 _07855_/A2 _07858_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05708__A1 _09649_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07786_ _08696_/A2 _08505_/B _07789_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06381__A1 _09374_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06806_ _06835_/A1 _09125_/I _06806_/B _06807_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_45_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09525_ _09547_/A2 _11523_/Q _09526_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06737_ _11574_/Q _10642_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_36_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09456_ _09472_/A2 _11501_/Q _09457_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11529__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06133__A1 _05693_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06668_ _11182_/Q _06701_/I _06668_/B _06668_/C _06671_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XPHY_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11497__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_08407_ _08528_/A1 _08403_/Z _08532_/A1 _08409_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05619_ _11064_/Q _05515_/I _05620_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06599_ _06599_/A1 _06599_/A2 _06599_/A3 _06599_/A4 _06600_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_09387_ _09397_/A2 _11479_/Q _09388_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09622__A2 _09622_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08338_ _08517_/A1 _07555_/I _08339_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05892__B1 _11449_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11249__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10768__A1 _10896_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11679__CLK _06687_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10408__I _10408_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08269_ _08269_/A1 _08687_/A2 _08274_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07633__A1 _07635_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06436__A2 _11119_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10300_ _10378_/A1 _11554_/Q _10302_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11280_ _11280_/D input76/Z _06705_/Z _11280_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10231_ _10231_/A1 _10231_/A2 _11651_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10162_ _10352_/A1 _11359_/Q _10163_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_145 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09138__A1 _09142_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10093_ _10350_/A1 _10607_/A1 _10094_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11059__CLK input68/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06372__A1 _09424_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06372__B2 _11252_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08361__A2 _08355_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10995_ _11016_/A1 input156/Z _10998_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1030 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09310__A1 _09154_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11488__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1052 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1041 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06124__A1 _09041_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1096 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1085 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09613__A2 _09622_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11616_ _11616_/D _11686_/RN _06705_/Z _11616_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__10759__A1 _11417_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10208__B1 _11440_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05700__I _05700_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07624__A1 _07640_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11547_ _11547_/D _11686_/RN _06705_/Z _11547_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__10759__B2 _10889_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11478_ _11478_/D _11686_/RN _06705_/Z _11478_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__11660__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08232__B _08656_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10429_ _10429_/A1 _10429_/A2 _10514_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06531__I _11219_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_825 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07627__I _08686_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_847 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_836 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09129__A1 _09142_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05970_ _11267_/Q _06040_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_07640_ _07640_/A1 _07527_/I _07643_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08352__A2 _08355_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06363__A1 _07398_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07571_ _08339_/A1 _08494_/A2 _07572_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_09310_ _09154_/Z _09322_/A2 _09310_/B _09311_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06522_ _06612_/A1 _11161_/Q _06523_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09301__A1 _09116_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11479__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06115__A1 _06839_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09852__A2 _09935_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09241_ _09241_/I _09241_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_06453_ _06458_/A2 _11069_/Q _06454_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_33_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05874__B1 _07201_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06384_ _07398_/A1 _06238_/Z _11244_/Q _06385_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__06706__I _11486_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09172_ _09195_/A2 _11411_/Q _09173_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08123_ _08156_/A2 _08142_/A2 _08126_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07615__A1 _07640_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09604__A2 _09622_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08054_ _08054_/A1 _08054_/A2 _08055_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09368__A1 _09372_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07005_ _07005_/I _11130_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11651__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05929__A1 _05660_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput118 wb_adr_i[29] input118/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput107 wb_adr_i[19] _06591_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__11201__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10922__A1 _10922_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput129 wb_cyc_i input129/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input30_I mask_rev_in[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08956_ _08963_/A2 _11344_/Q _08957_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07907_ _07907_/A1 _07917_/A1 _07981_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08887_ _08888_/A2 _11322_/Q _08888_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09540__A1 _09547_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08343__A2 _08677_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07838_ _08519_/B _08519_/A1 _07843_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11351__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06354__A1 _08786_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10150__A2 _09961_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09508_ _09508_/I _11517_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07769_ _08592_/A2 _07774_/A2 _07771_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10780_ _10780_/A1 _10780_/A2 _10780_/A3 _10780_/A4 _10787_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__10989__A1 _08493_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06106__A1 _06396_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_09439_ _09439_/I _11495_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06657__A2 input68/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_11401_ _11401_/D input76/Z _06705_/Z _11401_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__06409__A2 _08799_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11642__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11332_ _11332_/D _11686_/RN _06705_/Z _11332_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__09359__A1 _09372_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11263_ _11263_/D _11263_/RN input68/Z _11263_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
X_11194_ _11194_/D _11686_/RN _06705_/Z _11194_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10214_ _11512_/Q _10369_/A2 _10369_/B1 _11504_/Q _10217_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11635__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10145_ _11478_/Q _10367_/A1 _11470_/Q _10366_/A1 _10145_/C _10152_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__10913__B2 _10913_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10076_ _10373_/A1 _11516_/Q _10373_/B1 _11524_/Q _10079_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09531__A1 _09547_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08334__A2 _08513_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06345__A1 _09624_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06896__A2 _06902_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10978_ _10966_/Z _10978_/A2 _10979_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06648__A2 input79/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07131__B _07151_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08270__A1 split14/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11224__CLK _11683_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11633__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09770__A1 _09241_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10904__A1 _10904_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08810_ _08820_/A2 _11298_/Q _08811_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_09790_ _09790_/I _11607_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11374__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_644 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_677 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_08741_ _08741_/I _11277_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05953_ _05953_/A1 _05953_/A2 _05953_/A3 _05953_/A4 _05967_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08325__A2 _08639_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05884_ _11505_/Q _09449_/A1 _11497_/Q _09424_/A1 _05884_/C _05893_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__06336__A1 _05703_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08672_ _08672_/A1 _08688_/A3 _08672_/B _08673_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09522__A1 _09270_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10668__B1 _10886_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07623_ _07623_/A1 _07623_/A2 _08413_/C _08268_/B _07626_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__06887__A2 _06902_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09825__A2 _09015_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07554_ _07579_/A1 _07839_/A2 _07555_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07485_ _07485_/I _07486_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06505_ _06505_/A1 _06604_/A1 _11059_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09224_ _09116_/Z _09246_/A2 _09224_/B _09225_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10840__B1 _11135_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06436_ _06966_/A1 _11119_/Q _06437_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09155_ _09169_/A2 _11406_/Q _09156_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06367_ _09117_/A1 _11395_/Q _06370_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08106_ _08106_/A1 _08142_/A1 _08616_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09086_ _06863_/Z _09089_/A2 _09086_/B _09087_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input78_I ser_tx VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06298_ _08990_/A1 _11356_/Q _06933_/A1 _11110_/Q _06301_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11624__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08037_ _08037_/A1 _08037_/A2 _08194_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06811__A2 _11074_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08800__A3 _06904_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09761__A1 _09154_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09988_ _10366_/A1 _11467_/Q _09991_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08939_ _08939_/I _11338_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09513__A1 _09158_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10901_ _10901_/A1 _10901_/A2 _10902_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06327__A1 _09750_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05515__I _05515_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09816__A2 _11616_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10832_ _10924_/A1 _11330_/Q _10833_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10763_ _10763_/A1 _10763_/A2 _10763_/A3 _10763_/A4 _10780_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_12_143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11247__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10694_ _10922_/A1 _11359_/Q _10696_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07055__A2 _08795_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06802__A2 _05633_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11615__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11315_ _11315_/D _11686_/RN _06705_/Z _11315_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__11397__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11246_ _11246_/D _11686_/RN _06705_/Z _11246_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_11177_ _11177_/D _11686_/RN _06705_/Z _11177_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__09752__A1 _09116_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11589__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10128_ _10154_/A1 _10880_/C _10128_/B _10129_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09504__A1 _09121_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07126__B _07151_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10059_ _10356_/A1 _11404_/Q _10061_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10114__A2 _11485_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06869__A2 _06869_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10822__B1 _10916_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07270_ _07270_/I _11197_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07294__A2 _08036_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06221_ _09274_/A1 _11444_/Q _06224_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08243__A1 _08545_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06152_ _11485_/Q _09399_/A1 _11477_/Q _09374_/A1 _06152_/C _06165_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__11606__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06083_ _08742_/A1 _11281_/Q _06087_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09911_ _09911_/A1 _09935_/B _09922_/B _10404_/A1 _11637_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06006__B1 _09674_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09842_ _09187_/I _09848_/A2 _09842_/B _09843_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_09773_ _09270_/I _09773_/A2 _09773_/B _09774_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_284 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_474 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_06985_ _10945_/A1 _06974_/I _06985_/B _06986_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input132_I wb_dat_i[11] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08724_ _07431_/Z _08724_/A2 _08724_/B _08725_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_05936_ _06324_/A1 _11592_/Q _05938_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05780__A2 _05805_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06309__A1 _05924_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08655_ _08655_/A1 _08655_/A2 _08673_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05867_ _11569_/Q _09649_/A1 _09624_/A1 _11561_/Q _05868_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08586_ _08586_/A1 _08586_/A2 _08586_/A3 _08586_/A4 _08690_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_07606_ _07606_/A1 _07606_/A2 _07613_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_81_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07537_ _07537_/I _08592_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_05798_ _05798_/I _09449_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
X_07468_ _07478_/A1 _08006_/A2 _07689_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07399_ _07403_/A2 _11244_/Q _07400_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06419_ _06419_/A1 _06419_/A2 _06419_/A3 _06439_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_09207_ _09220_/A2 _11422_/Q _09208_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09138_ _09142_/A2 _11401_/Q _09139_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10416__I _10416_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09982__A1 _10377_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11100_ _11100_/D _11686_/RN _06705_/Z _11100_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_118_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09069_ _09069_/I _11379_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11031_ _11684_/Q _11032_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08537__A2 _08686_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10344__A2 _06556_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10815_ _10815_/A1 _10815_/A2 _10816_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05523__A2 _06619_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06720__A1 _06786_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10746_ _10881_/A1 _11661_/Q _10747_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10677_ _10896_/A1 _11439_/Q _10679_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10032__A1 _10350_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput208 _10137_/A1 mgmt_gpio_oeb[7] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput219 _11165_/Q mgmt_gpio_out[17] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_99_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11229_ _11229_/D _11686_/RN _06705_/Z _11229_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__07635__I _07635_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11451__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06770_ _07110_/I _11061_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05762__A2 _08890_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11412__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05721_ _05721_/I _08990_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XANTENNA__10099__A1 _10356_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05652_ _05927_/I input51/Z _05662_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08440_ _08435_/Z _08653_/A1 _08550_/A2 _08443_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_90_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06711__A1 _06514_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08371_ _08433_/A1 _08371_/A2 _08558_/A2 _08692_/B _08371_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
X_05583_ _11701_/Q _11161_/Q _05584_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__11562__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07267__A2 _06838_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07322_ _07322_/I _11211_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07253_ _06851_/Z _07265_/A2 _07253_/B _07254_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07184_ _05925_/Z _09187_/I _07185_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06204_ _06204_/I _08825_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_06135_ _06135_/A1 _06135_/A2 _06136_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10023__A1 _10023_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06066_ _06324_/A1 _11590_/Q _09750_/A1 _11598_/Q _06067_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11404__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09716__A1 _09187_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08519__A2 _08519_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09825_ _05660_/Z _09015_/I _09848_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__09192__A2 _09195_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09756_ _09756_/I _11596_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06968_ _06837_/Z _06971_/A2 _06968_/B _06969_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11419__SETN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_09687_ _09697_/A2 _11575_/Q _09688_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08707_ _08707_/I _11261_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05919_ _09248_/A1 _11440_/Q _05921_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11092__CLK _11663_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06899_ _06863_/Z _06902_/A2 _06899_/B _06900_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08638_ _08638_/A1 _08638_/A2 _08638_/A3 _08638_/A4 _08691_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__06702__A1 _05616_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08569_ _08620_/A1 _08569_/A2 _08662_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10600_ _10903_/A1 _11557_/Q _10603_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11580_ _11580_/D _11686_/RN _06705_/Z _11580_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__10262__A1 _10375_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10531_ _10892_/A1 _11468_/Q _10532_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06624__I _11534_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10462_ _10921_/A1 _11331_/Q _10468_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10393_ _10393_/I _10460_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__09955__A1 _09973_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08758__A2 _11283_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10565__A2 _11381_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09707__A1 _09125_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11014_ _11014_/A1 _10966_/Z _11014_/B _11015_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_77_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05992__A2 _08915_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10317__A2 _11135_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07194__A1 _05925_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11435__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11705__I input65/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11585__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05703__I _05703_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10253__A1 _10371_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10729_ _11528_/Q _10902_/A2 _11520_/Q _10902_/B2 _10729_/C _10736_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__10005__A1 _11491_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05680__A1 _08825_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_324 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07940_ _07964_/A1 _07973_/A2 _08557_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05983__A2 _11288_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07871_ _07871_/A1 _07871_/A2 _07872_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09610_ _09154_/Z _09622_/A2 _09610_/B _09611_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06822_ _11695_/Q _05633_/B _06822_/B _09187_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_09541_ _09187_/Z _09547_/A2 _09541_/B _09542_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_95_285 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06753_ _06753_/A1 _06754_/A2 _06753_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05704_ _05703_/Z _08839_/A2 _05705_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09472_ _09270_/Z _09472_/A2 _09472_/B _09473_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06684_ _11305_/Q _06684_/A2 _06684_/B _06685_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_36_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08423_ _08285_/B _08423_/A2 _08540_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05635_ _05718_/A1 _05776_/A2 _05636_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__06160__A2 _09197_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08354_ _08656_/A1 _08367_/B split15/I _08361_/B _08548_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05566_ _05566_/I _11692_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08988__A2 _08988_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07305_ _07305_/I _11206_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08285_ _07455_/Z _08285_/A2 _08285_/B _08540_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06999__A1 _08795_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05497_ _05498_/A2 _11702_/Q _05498_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11308__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07236_ _07236_/I _11187_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07167_ _07197_/A1 _07167_/A2 _07167_/B _07168_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_172_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07412__A2 _06238_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06118_ _06118_/A1 _06118_/A2 _06118_/A3 _06119_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_input60_I mgmt_gpio_in[31] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11458__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07098_ _07098_/I _11156_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_78_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06049_ _11518_/Q _09499_/A1 _11510_/Q _09474_/A1 _06049_/C _06058_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__07176__A1 _07197_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09165__A2 _11409_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09808_ _09125_/I _09823_/A2 _09808_/B _09809_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07715__A3 _08490_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08912__A2 _11330_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09739_ _09158_/I _09725_/Z _09739_/B _09740_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10483__A1 _10892_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11701_ _11701_/D _11701_/RN input68/Z _11701_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_11632_ _11632_/D _11686_/RN _11666_/CLK _11632_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XANTENNA__08979__A2 _08988_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10235__A1 _10353_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11563_ _11563_/D _11686_/RN _06705_/Z _11563_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__10786__A2 _11329_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11494_ _11494_/D _11686_/RN _06705_/Z _11494_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_6_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10514_ _10514_/I _10924_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__05662__A1 _05662_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10445_ _10445_/I _10888_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_10_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10538__A2 _10900_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10376_ _10376_/A1 _10376_/A2 _10376_/A3 _10381_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__06611__B1 _06466_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07167__A1 _07197_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09156__A2 _09169_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10710__A2 _11424_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06914__A1 _06837_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_285 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10474__A1 _10896_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09092__A1 _09114_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08070_ _08095_/A1 split13/Z _08071_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11600__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07021_ _07025_/A2 _11135_/Q _07022_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10514__I _10514_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08972_ _08988_/A2 _11349_/Q _08973_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07923_ _07923_/A1 _07923_/A2 _07928_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07158__A1 _07201_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07854_ _07854_/A1 _07854_/A2 _07855_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06805_ _06835_/A1 _11073_/Q _06806_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11194__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07785_ _07785_/A1 _07785_/A2 _07789_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09524_ _05693_/Z _09015_/I _09547_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_06736_ _11558_/Q _10146_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_09455_ _09455_/I _11500_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06667_ _06701_/I _06667_/A2 _06668_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06133__A2 _11525_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08406_ _08406_/A1 _08406_/A2 _08532_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_101_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05618_ _11065_/Q _06480_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__11130__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07330__A1 _10954_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06598_ _06598_/A1 input118/Z _06599_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09386_ _09386_/I _11478_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08337_ _08600_/A1 _08332_/B _08517_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05549_ _05549_/A1 _05519_/I _05549_/B _05550_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09083__A1 _06859_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08268_ _08400_/A1 _08686_/B _08268_/B _08687_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07633__A2 _08686_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11280__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11282__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07219_ _07240_/A1 _11184_/Q _07220_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08199_ _08199_/I _08232_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_10230_ _10881_/A1 _11651_/Q _10231_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output264_I _11273_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10161_ _10353_/A1 _11367_/Q _10163_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10092_ _10092_/I _10092_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__08897__A1 _08913_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06372__A2 _11491_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11185__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10994_ _10994_/I _11678_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1020 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1053 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1042 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07321__A1 _10945_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1097 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1086 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10208__A1 _11448_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11623__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11615_ _11615_/D _11686_/RN _06705_/Z _11615_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__09074__A1 _06847_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11546_ _11546_/D _11686_/RN _06705_/Z _11546_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_168_393 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10759__A2 _10888_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11477_ _11477_/D _11686_/RN _06705_/Z _11477_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_143_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10428_ _10428_/A1 _10428_/A2 _10428_/B1 _10428_/B2 _10429_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_10359_ _11134_/Q _10359_/A2 _11132_/Q _10359_/B2 _10359_/C _10364_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__06060__A1 _05927_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_848 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_837 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10144__B1 _09986_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08888__A1 _06867_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11176__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10695__A1 _10919_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07570_ _07570_/I _08494_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11153__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06521_ _05509_/I _06521_/A2 _06612_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10447__A1 _10884_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07312__A1 _07310_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09240_ _09240_/I _11432_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06452_ _06452_/I _11070_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05874__B2 input59/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06383_ _07412_/A1 _06238_/Z _11248_/Q _06385_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09171_ _09171_/A1 _09015_/Z _09195_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_08122_ _08122_/A1 _08218_/B _08472_/C _08122_/A4 _08125_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_08053_ _08057_/A1 split13/Z _08055_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_147_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11100__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07004_ _06843_/Z _07004_/A2 _07004_/B _07005_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07379__A1 _07076_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input162_I wb_rstn_i VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05929__A2 _11624_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput108 wb_adr_i[1] _07496_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08955_ _08955_/I _11343_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput119 wb_adr_i[2] input119/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__08328__B1 _08328_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07906_ split6/I _07921_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XANTENNA_input23_I mask_rev_in[27] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08879__A1 _06855_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08886_ _08886_/I _11321_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10135__B1 _10615_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09540__A2 _11528_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07837_ _07837_/I _08519_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__10686__A1 _10905_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11167__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07768_ _08328_/B1 _08587_/B _08310_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09507_ _09125_/Z _09522_/A2 _09507_/B _09508_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06719_ _06753_/A1 input86/Z _06720_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07699_ _07839_/A2 _07699_/A2 _07700_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11646__CLK _11663_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_09438_ _09158_/Z _09447_/A2 _09438_/B _09439_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05865__A1 _09699_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09369_ _09241_/Z _09372_/A2 _09369_/B _09370_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08803__A1 _08803_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11400_ _11400_/D input76/Z _06705_/Z _11400_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__06409__A3 _06408_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05617__A1 _05616_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10610__A1 _10092_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11331_ _11331_/D _11686_/RN _06705_/Z _11331_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_125_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11262_ _11262_/D _11686_/RN _06705_/Z _11262_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_21_74 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06290__A1 _08795_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11193_ _11193_/D _11686_/RN _06705_/Z _11193_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10213_ _10213_/A1 _10213_/A2 _10213_/A3 _10226_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_10144_ _10144_/A1 _09985_/I _09986_/I _10144_/B2 _10145_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__10913__A2 _10913_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07790__A1 _08332_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11176__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10075_ _10075_/A1 _10075_/A2 _10075_/A3 _10084_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__09531__A2 _11525_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11158__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10677__A1 _10896_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06079__I _11366_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10977_ _10977_/A1 _10977_/A2 _10977_/A3 _10978_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_15_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_5 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11330__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05856__A1 _09016_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10601__A1 _10904_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11529_ _11529_/D _11686_/RN _06705_/Z _11529_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__08270__A2 _07609_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08022__A2 _08204_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11519__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06033__A1 _09750_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_612 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09770__A2 _09773_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_08740_ _06855_/Z _08740_/A2 _08740_/B _08741_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05952_ _06785_/A1 _11076_/Q _05953_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_678 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_05883_ _05883_/A1 _05883_/A2 _05884_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08671_ _08671_/A1 _08671_/A2 _08688_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11149__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11669__CLK _11683_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09522__A2 _09522_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10668__A1 _10886_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06336__A2 _07412_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07622_ _08264_/B _08509_/A1 _08268_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07553_ _07553_/I _07839_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07484_ _08358_/A2 split5/Z _07485_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06504_ _06502_/I _11688_/Q _06604_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_166_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09223_ _09246_/A2 _11427_/Q _09224_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09038__A1 _09039_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11321__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10840__B2 _10889_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06435_ _08795_/A1 _07006_/A2 _11129_/Q _06437_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09154_ _09154_/I _09154_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_08105_ _08105_/A1 _08215_/B _08471_/C _08105_/A4 _08108_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_06366_ _09144_/A1 _11403_/Q _06370_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06297_ _06192_/I _05719_/I _06933_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09085_ _09089_/A2 _11385_/Q _09086_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput90 spimemio_flash_io2_do input90/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08036_ _08036_/A1 _08036_/A2 _08036_/B _08037_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09210__A1 _09220_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11199__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09761__A2 _09773_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09987_ _09896_/I _09959_/I _10366_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_08938_ _06867_/Z _08938_/A2 _08938_/B _08939_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09513__A2 _09522_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10659__B2 _10915_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10659__A1 _11623_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08869_ _08888_/A2 _11316_/Q _08870_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10900_ _10900_/A1 _11148_/Q _10901_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11560__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10831_ _10831_/A1 _10831_/A2 _10831_/A3 _10831_/A4 _10831_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_10762_ _10886_/B2 _11393_/Q _10886_/A2 _11401_/Q _10763_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09029__A1 _09039_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11312__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10693_ _10920_/A1 _11343_/Q _10920_/B1 _11351_/Q _10696_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_8_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08252__A2 _07885_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07055__A3 _06871_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11314_ _11314_/D _11686_/RN _06705_/Z _11314_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_141_506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11245_ _11245_/D _11686_/RN _06705_/Z _11245_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_106_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06015__A1 _11519_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09201__A1 _09220_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06015__B2 _09474_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11176_ _11176_/D _11686_/RN _06705_/Z _11176_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__09752__A2 _09773_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10127_ _10092_/Z _11647_/Q _10127_/B _10926_/C _10128_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__09504__A2 _09522_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10058_ _11380_/Q _10355_/A2 _11372_/Q _10355_/B2 _10058_/C _10067_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__11551__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09268__A1 _09241_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07818__A2 _08339_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10822__A1 _10915_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05829__A1 _10957_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11303__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10822__B2 _11626_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06220_ _09299_/A1 _11452_/Q _06224_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09440__A1 _09447_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08243__A2 _08490_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06151_ _06151_/A1 _06151_/A2 _06152_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06254__A1 _09474_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06082_ _06082_/A1 _05771_/I _05728_/I _06082_/B2 _06082_/C _06093_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__11341__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09910_ _10387_/I _09912_/I _09911_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10338__B1 _10377_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09841_ _09848_/A2 _11624_/Q _09842_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11491__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_431 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06557__A2 _10092_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10889__A1 _10889_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09772_ _09773_/A2 _11602_/Q _09773_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06984_ _06974_/I _11124_/Q _06985_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_464 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_05935_ _09775_/A1 _11608_/Q _05938_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08723_ _08724_/A2 _11272_/Q _08724_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_497 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06309__A2 input36/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08654_ _08694_/A3 _08694_/A2 _08655_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05866_ _09674_/A1 _11577_/Q _05868_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input125_I wb_adr_i[6] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11542__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08585_ _07609_/Z _08315_/B _08586_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05797_ _06238_/I _08799_/A2 _05798_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07605_ _07605_/I _07606_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09259__A1 _09154_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07536_ _08339_/A1 _08614_/A2 _07537_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_41_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10813__A1 _10905_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07467_ _07471_/A1 _07471_/A2 _07478_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA_input90_I spimemio_flash_io2_do VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09206_ _09206_/I _11421_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07398_ _07398_/A1 _06238_/Z _06838_/Z _07403_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_06418_ _06418_/A1 _06418_/A2 _06418_/A3 _06418_/A4 _06419_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__09431__A1 _09447_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08234__A2 _08614_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06349_ _06349_/A1 _06349_/A2 _06349_/A3 _06349_/A4 _06350_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_09137_ _09137_/I _11400_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06245__A1 _07412_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09068_ _07426_/Z _09089_/A2 _09068_/B _09069_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08019_ _07837_/I _08391_/B _08612_/I _08020_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_output177_I _06056_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06796__A2 _05633_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11030_ _11030_/A1 _11030_/A2 _11030_/A3 _11032_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_76_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11214__CLK _11672_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10814_ _10906_/A1 _11546_/Q _10815_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06720__A2 _06753_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10804__A1 _10896_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10745_ _10092_/Z _11660_/Q _10745_/B _10880_/C _10747_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_43_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10676_ _10895_/A1 _11447_/Q _10679_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11364__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09422__A1 _09270_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput209 _10613_/B1 mgmt_gpio_oeb[8] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_11228_ _11228_/D _11686_/RN _06705_/Z _11228_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_4_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11159_ _11159_/D _07106_/ZN input68/Z _11159_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_82_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05720_ _07006_/A2 _05803_/A2 _05721_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10099__A2 _11405_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06172__B1 _08846_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05651_ _05651_/I _05927_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__08161__A1 _08161_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08370_ split8/I _08444_/B _08370_/B _08692_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06711__A2 input84/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07321_ _10945_/A1 _07310_/I _07321_/B _07322_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05582_ _11270_/Q _06667_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07252_ _07265_/A2 _11192_/Q _07253_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09413__A1 _09158_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07183_ _07183_/I _11177_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06203_ _05703_/Z _07419_/A2 _11251_/Q _06206_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06134_ _09549_/A1 _11533_/Q _06135_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06227__A1 _07398_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10023__A2 _10265_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06065_ _11614_/Q _09800_/A1 _09775_/A1 _11606_/Q _06067_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08431__B _08431_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09716__A2 _09722_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06730__I _11422_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09824_ _09824_/I _11618_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09755_ _09121_/I _09773_/A2 _09755_/B _09756_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11237__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06967_ _06971_/A2 _11119_/Q _06968_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06898_ _06902_/A2 _11099_/Q _06899_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09686_ _09686_/I _11574_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08706_ _07426_/Z _08709_/A2 _08706_/B _08707_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05918_ _11424_/Q _09197_/A1 _11416_/Q _09171_/A1 _05918_/C _05923_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__08152__A1 split7/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08637_ _07566_/I _07537_/I _08637_/B _08638_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05849_ _10233_/A2 _05991_/I _05849_/B _05850_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_64_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11573__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06702__A2 input68/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11387__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05910__B1 _11480_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08568_ _08568_/A1 _08568_/A2 _08569_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07519_ split13/I _08095_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08499_ _08499_/I _08588_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10262__A2 _11545_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10530_ _10897_/A2 _11452_/Q _10532_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_182_214 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11588__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10461_ _10461_/I _10921_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__09404__A1 _09121_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10014__A2 _09876_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06218__A1 _08786_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10392_ _10392_/A1 _10407_/A1 _10393_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09707__A2 _09722_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06640__I input80/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11013_ _10966_/Z _11013_/A2 _11014_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08391__A1 _07492_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07194__A2 _09270_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11506__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09891__B2 _09902_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09643__A1 _09647_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10253__A2 _11489_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10728_ _10728_/A1 _10728_/A2 _10729_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10659_ _11623_/Q _10916_/A1 _11615_/Q _10915_/A1 _10659_/C _10663_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__06209__A1 _05703_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10005__A2 _10370_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05680__A2 _05803_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10961__B1 _11028_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07870_ _07870_/A1 _07471_/B _07870_/A3 _07871_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__07185__A2 _05925_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10713__B1 _11408_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06821_ _11007_/A1 _05633_/B _06822_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09540_ _09547_/A2 _11528_/Q _09541_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06752_ input76/Z _06754_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09471_ _09472_/A2 _11506_/Q _09472_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05703_ _05703_/I _05703_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_06683_ _11305_/Q input96/Z _06684_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08422_ _08422_/A1 _08666_/A2 _08666_/A1 _08664_/A3 _08425_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_05634_ _05716_/A1 _05715_/I _05776_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_08353_ _08353_/I _08433_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09634__A1 _09647_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05565_ _05565_/A1 _05519_/I _05565_/B _05566_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08284_ _08284_/A1 _08540_/A1 _08282_/Z _08666_/A1 _08292_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__10244__A2 _11425_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07304_ _07076_/Z _07307_/A2 _07304_/B _07305_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06999__A2 _07006_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05496_ _05969_/I _11159_/Q _05498_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07235_ _07240_/A1 _07235_/A2 _07235_/B _07236_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07166_ _07197_/A1 _11174_/Q _07167_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07097_ _07081_/Z _07097_/A2 _07097_/B _07098_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06117_ _08761_/A1 _11286_/Q _06118_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06048_ _10148_/B2 _05798_/I _05795_/I _06048_/B2 _06049_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__07412__A3 _06838_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input53_I mgmt_gpio_in[25] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08373__A1 split8/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07176__A2 _11176_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07999_ _08003_/A2 _07999_/A2 _08001_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10180__A1 _10370_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09807_ _09823_/A2 _11613_/Q _09808_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09738_ _09725_/Z _11591_/Q _09739_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09669_ _09241_/Z _09672_/A2 _09669_/B _09670_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06136__B1 _11541_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06687__A1 _11304_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11700_ _11700_/D _11700_/RN input68/Z _11700_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_91_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09625__A1 _09647_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11631_ _11631_/D _11686_/RN _11666_/CLK _11631_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_11562_ _11562_/D _11686_/RN _06705_/Z _11562_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_24_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06439__A1 _06392_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10513_ _10513_/A1 _10047_/B _10513_/A3 _10559_/A1 _10880_/C _11656_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_155_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11493_ _11493_/D _11686_/RN _06705_/Z _11493_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_10444_ _10444_/A1 _10506_/A2 _10445_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_170_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10375_ _10375_/A1 _11686_/Q _10376_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11402__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11552__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08116__A1 split8/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06127__B1 _11381_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09616__A1 _09187_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11403__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07020_ _07370_/A1 _06217_/Z _06871_/Z _07025_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__11082__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08971_ _08971_/I _11348_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07922_ _07922_/I _07923_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07853_ input103/Z _07863_/I _07854_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07158__A2 _05925_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10162__A1 _10352_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06804_ _06804_/I _09125_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__06905__A2 _06904_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07784_ _07722_/I _08689_/B _07785_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08107__A1 split8/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06735_ _11518_/Q _06735_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09523_ _09523_/I _11522_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_43_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_09454_ _09121_/Z _09472_/A2 _09454_/B _09455_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10465__A2 _10427_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06666_ _06666_/A1 _06666_/A2 _06666_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09385_ _09154_/Z _09397_/A2 _09385_/B _09386_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_08405_ _08419_/A1 _07586_/I _08405_/B _08406_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05617_ _05616_/C _11258_/Q _05617_/B _05802_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__07330__A2 _07310_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06597_ _06597_/I _06598_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09607__A1 _09125_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08336_ _08336_/A1 _08675_/A2 _08336_/A3 _08642_/A3 _08342_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__07881__A3 _07885_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05548_ _05519_/I _11696_/Q _05549_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09083__A2 _09089_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07094__A1 _07076_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08267_ _08263_/Z _08413_/B _08529_/A4 _08269_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11425__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08830__A2 _11304_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08198_ split12/Z _08242_/A1 _08199_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06841__A1 _06837_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07218_ _11318_/Q _05924_/Z _07218_/B _07220_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07149_ _11171_/Q _07152_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_145_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11575__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_464 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10160_ _11351_/Q _10351_/A2 _11343_/Q _10351_/B2 _10160_/C _10173_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_10091_ _11648_/Q _10154_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_19_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08897__A2 _11325_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10993_ _10993_/A1 _10966_/Z _10993_/B _10994_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08649__A2 _08692_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06109__B1 _08742_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1021 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1010 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10456__A2 _10506_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1065 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1054 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1032 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07321__A2 _07310_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1098 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1087 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_11614_ _11614_/D _11686_/RN _06705_/Z _11614_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__09074__A2 _09089_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11545_ _11545_/D _11686_/RN _06705_/Z _11545_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__07085__A1 _08825_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11476_ _11476_/D _11686_/RN _06705_/Z _11476_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_10427_ _10427_/A1 _09912_/I _10427_/B _10428_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08585__A1 _07609_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_816 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_10358_ _10358_/A1 _10358_/A2 _10359_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06060__A2 input46/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10289_ _10367_/A1 _11482_/Q _10290_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_827 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10144__B2 _10144_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10144__A1 _10144_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08888__A2 _08888_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06899__A1 _06863_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06363__A3 _06217_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06520_ _06520_/I _06577_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10447__A2 _11379_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11448__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06451_ _06451_/A1 _06458_/A2 _06451_/B _06452_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05874__A2 _05927_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06382_ _09399_/A1 _11483_/Q _06385_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09170_ _09170_/I _11410_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08121_ split7/I _08220_/B _08122_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11357__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08052_ _08054_/A1 _07522_/I _08057_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10080__B1 _10377_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11598__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06823__A1 _06835_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07003_ _07004_/A2 _11130_/Q _07004_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput109 wb_adr_i[20] _07470_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_input155_I wb_dat_i[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08954_ _06855_/Z _08963_/A2 _08954_/B _08955_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08328__A1 _07593_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07905_ _08545_/A1 _08519_/A2 split6/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__08879__A2 _08888_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08885_ _06863_/Z _08888_/A2 _08885_/B _08886_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10686__A2 _11535_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07836_ _07836_/A1 _07989_/A1 _07837_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07767_ _07530_/I _07752_/I _08328_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA_input16_I mask_rev_in[20] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06354__A3 _06217_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09506_ _09522_/A2 _11517_/Q _09507_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10438__A2 _09934_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06718_ _06718_/I _06718_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08500__A1 _08509_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07698_ _08294_/B _08614_/A2 _08290_/C _07704_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09437_ _09447_/A2 _11495_/Q _09438_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06649_ _06649_/A1 _06649_/A2 _06649_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05865__A2 _11585_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09368_ _09372_/A2 _11473_/Q _09369_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_177_180 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08319_ _08332_/A1 _08417_/A2 _08505_/B _08593_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07067__A1 _06843_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09299_ _09299_/A1 _09015_/Z _09322_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__05617__A2 _11258_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08803__A2 _06904_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11330_ _11330_/D input76/Z _06705_/Z _11330_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_108_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11261_ _11261_/D _11686_/RN _06705_/Z _11261_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__06290__A2 _07006_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11192_ _11192_/D _11686_/RN _06705_/Z _11192_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10212_ _10366_/A1 _11472_/Q _10213_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10374__A1 _10374_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10143_ _10143_/A1 _10143_/A2 _10143_/A3 _10143_/A4 _10153_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__08319__A1 _08332_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10074_ _10370_/A1 _11492_/Q _10075_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10677__A2 _11439_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09819__A1 _09823_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10976_ _08431_/B input161/Z _08460_/B input138/Z _10977_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06805__A1 _06835_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11528_ _11528_/D _11686_/RN _06705_/Z _11528_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__11094__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11459_ _11459_/D _11686_/RN _06705_/Z _11459_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__06281__A2 _06281_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07230__A1 _07240_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11120__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input8_I mask_rev_in[13] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10117__A1 _10375_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05792__A1 _06238_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05951_ _08761_/A1 _11289_/Q _05953_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_679 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_05882_ _09474_/A1 _11513_/Q _05883_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08670_ _08403_/Z _07582_/I _08670_/A3 _08670_/A4 _08671_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__05544__A1 _05519_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07621_ _08264_/B _08417_/A2 _08413_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07552_ _07552_/A1 input119/Z _07553_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06503_ _06611_/A1 _11059_/Q _06505_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07483_ _08495_/B _08358_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_34_462 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09222_ _09222_/A1 _09015_/Z _09246_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__09038__A2 _11370_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10840__A2 _10888_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06434_ _09041_/A1 _11371_/Q _06437_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_147_320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09153_ _09153_/I _11405_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06365_ _06365_/A1 _06365_/A2 _06365_/A3 _06365_/A4 _06371_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_181_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08104_ split7/I _08209_/B _08105_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06733__I _11478_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09084_ _09084_/I _11384_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06296_ _06296_/A1 _06296_/A2 _06296_/A3 _06302_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xinput91 spimemio_flash_io2_oeb input91/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08035_ _08395_/B _08395_/A1 _08036_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput80 spi_enabled input80/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09210__A2 _11423_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10356__A1 _10356_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07564__I _07564_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07772__A2 _08696_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09986_ _09986_/I _10365_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__10108__B2 _11461_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08937_ _08938_/A2 _11338_/Q _08938_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11613__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10659__A2 _10916_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08868_ _08868_/I _11315_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07819_ _07819_/A1 _08514_/A2 _08335_/A1 _07819_/A4 _07826_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__08721__A1 _07426_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08799_ _08799_/A1 _08799_/A2 _08801_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10830_ _10919_/A1 _11370_/Q _10831_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10761_ _10883_/A1 _11377_/Q _10763_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_157_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10692_ _10921_/A1 _11335_/Q _10696_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10044__B1 _10355_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10595__A1 _10902_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06643__I _06643_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11313_ _11313_/D _11686_/RN _06705_/Z _11313_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_11244_ _11244_/D _11686_/RN _06705_/Z _11244_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__11143__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06015__A2 _09499_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07212__A1 _05924_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11175_ _11175_/D _11686_/RN _06705_/Z _11175_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__11293__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05774__B2 _09066_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08960__A1 _06863_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10126_ _10107_/Z _10092_/Z _10126_/A3 _10126_/A4 _10127_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_10057_ _10057_/A1 _10057_/A2 _10058_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_180_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09268__A2 _09272_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10959_ input168/Z input163/Z _11025_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05829__A2 _05969_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_498 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10586__A1 _10913_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06150_ _09349_/A1 _11469_/Q _06151_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06254__A2 _11508_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06081_ _05723_/Z _11350_/Q _06082_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06006__A2 _09699_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10338__A1 _10377_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10338__B2 _11261_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11636__CLK _11658_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09840_ _09840_/I _11623_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10889__A2 _11136_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09771_ _09771_/I _11601_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06983_ _06983_/I _11123_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06557__A3 _06577_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08951__A1 _06851_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05765__A1 _07006_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05934_ _09800_/A1 _11616_/Q _05938_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08722_ _08722_/I _11271_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_498 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_08653_ _08653_/A1 _08653_/A2 _07911_/I _08653_/A4 _08694_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_05865_ _09699_/A1 _11585_/Q _05868_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05796_ _09424_/A1 _11498_/Q _05800_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07604_ _07593_/I _07774_/A2 _07605_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08584_ _08584_/A1 _08431_/B _08460_/B _08584_/B2 _08584_/C _08603_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA_input118_I wb_adr_i[29] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06728__I _11382_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09259__A2 _09272_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07535_ _07535_/I _08614_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_07466_ _07865_/A1 _07463_/Z _07466_/A3 _07471_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_139_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06417_ _08761_/A1 _11284_/Q _06418_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09205_ _09125_/Z _09220_/A2 _09205_/B _09206_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_167_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07397_ _07397_/I _11243_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11166__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10577__A1 _10895_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06348_ _05703_/Z _08786_/A1 _11261_/Q _06349_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_input83_I spi_sdoenb VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09136_ _06859_/Z _09142_/A2 _09136_/B _09137_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10026__B1 _10359_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06245__A2 _06238_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06279_ _08761_/A1 _11285_/Q _06280_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09067_ _09089_/A2 _11379_/Q _09068_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08018_ _08562_/A1 _08632_/A2 _08649_/B _08612_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_78_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09195__A1 _06867_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output337_I _11674_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07745__A2 split13/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09969_ _11634_/Q _11633_/Q _09970_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__08942__A1 _07426_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11230__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10813_ _10905_/A1 _11538_/Q _10815_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11509__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11297__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10744_ _10744_/A1 _10092_/Z _10742_/Z _10744_/A4 _10745_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_10675_ _11495_/Q _10894_/A2 _11487_/Q _10894_/B2 _10675_/C _10679_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__10568__A1 _10889_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09422__A2 _09422_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07433__A1 _07431_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11659__CLK _11663_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05995__A1 _08799_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11227_ _11227_/D _11686_/RN _06705_/Z _11227_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__07736__A2 _08495_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11158_ _11158_/D _11686_/RN _06705_/Z _11158_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10109_ _10366_/A1 _11469_/Q _10111_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11221__RN input162/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_435 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10740__A1 _10922_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11089_ _11089_/D input76/Z _11663_/CLK _11089_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__06172__A1 _05660_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08161__A2 _08656_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05650_ _08795_/A1 _08825_/A2 _05651_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06172__B2 input62/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05581_ _05581_/I _11687_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11189__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10256__B1 _10379_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09110__A1 _09114_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07320_ _07310_/I _11211_/Q _07321_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07251_ _07251_/I _11191_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07182_ _07197_/A1 _07182_/A2 _07182_/B _07183_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06202_ _09699_/A1 _11580_/Q _06206_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09413__A2 _09422_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06133_ _05693_/Z _11525_/Q _06135_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07424__A1 _07081_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06064_ input67/Z _05924_/I input38/Z _05925_/I _06064_/C _06067_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__05986__A1 _09016_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09823_ _09270_/I _09823_/A2 _09823_/B _09824_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10731__A1 _10903_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09754_ _09773_/A2 _11596_/Q _09755_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06966_ _06966_/A1 _06904_/Z _06971_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06897_ _06897_/I _11098_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09685_ _09154_/I _09697_/A2 _09685_/B _09686_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08705_ _08709_/A2 _11261_/Q _08706_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05917_ _05917_/A1 _05917_/A2 _05918_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08636_ _08636_/I _08638_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05848_ _08940_/A1 _11345_/Q _05849_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05910__A1 _11488_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05910__B2 _09374_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08567_ _08567_/A1 _08696_/A2 _08567_/B _08567_/C _08568_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_05779_ _05779_/I _09399_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XANTENNA__09101__A1 _09114_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07518_ _07524_/A2 split13/Z _07521_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08498_ _07570_/I _07748_/I _08498_/B _08498_/C _08499_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_07449_ _07449_/I split16/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_10460_ _10460_/A1 _10506_/A2 _10460_/A3 _10461_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__09404__A2 _09422_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_09119_ _09116_/Z _09142_/A2 _09119_/B _09120_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10391_ _10391_/I _10915_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XANTENNA__09955__A3 _10265_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09168__A1 _09169_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11012_ _11012_/A1 _11012_/A2 _11012_/A3 _11013_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08915__A1 _08915_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08391__A2 _08204_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11203__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10722__A1 _10895_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05729__A1 _08940_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09340__A1 _09347_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06154__A1 _09449_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11331__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09891__A2 _10023_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09643__A2 _11561_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11481__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10727_ _10900_/A1 _11512_/Q _10728_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10658_ _10658_/A1 _10658_/A2 _10659_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10589_ _10589_/A1 _10589_/A2 _10589_/A3 _10589_/A4 _10589_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__05968__A1 _05968_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10961__B2 _08493_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11442__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09159__A1 _09169_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08906__A1 _08913_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10713__B2 _10889_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06820_ _11680_/Q _11007_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06751_ _06751_/I _11217_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09470_ _09470_/I _11505_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09331__A1 _09347_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06682_ _11180_/Q _06684_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05702_ _05702_/I _09699_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XANTENNA__06145__A1 _09750_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08421_ split15/Z _08283_/B _08664_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05633_ _05633_/A1 _05633_/A2 _05633_/B _05715_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08352_ _08383_/A1 _08355_/I _08352_/B _08353_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05564_ _05519_/I _11692_/Q _05565_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08283_ split14/Z _07609_/Z _08283_/B _08666_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05495_ _05526_/A1 _11070_/Q _05969_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_07303_ _07307_/A2 _11206_/Q _07304_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06999__A3 _06871_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07234_ _07240_/A1 _11187_/Q _07235_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11681__RN input162/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07165_ _11198_/Q _05925_/Z _07165_/B _07167_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07837__I _07837_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07096_ _07097_/A2 _11156_/Q _07097_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05959__A1 _06396_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06116_ _06785_/A1 _11073_/Q _06118_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11204__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06047_ _11494_/Q _06048_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11433__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input46_I mgmt_gpio_in[19] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07998_ _07998_/A1 _07470_/I _08003_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06384__A1 _07398_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09806_ _09806_/I _11612_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11354__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09737_ _09737_/I _11590_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06949_ _10942_/A1 _06941_/I _06949_/B _06950_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09322__A1 _09270_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09668_ _09672_/A2 _11569_/Q _09669_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06136__B2 _09574_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06687__A2 _06687_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08619_ _08619_/A1 _08619_/A2 _08658_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09599_ _09599_/A1 _09015_/I _09622_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_11630_ _11630_/D input76/Z _11665_/CLK _11630_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_24_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11561_ _11561_/D _11686_/RN _06705_/Z _11561_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__06439__A2 _06439_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10512_ _11656_/Q _10559_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_11492_ _11492_/D _11686_/RN _06705_/Z _11492_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_10443_ _11539_/Q _10906_/A1 _11499_/Q _10899_/A1 _10443_/C _10451_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_40_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10374_ _10374_/A1 _11158_/Q _10376_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06072__B1 _09624_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11424__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08364__A2 _08355_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08116__A2 _08575_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09313__A1 _09158_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10459__B1 _10919_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06127__B2 _09066_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09616__A2 _09622_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10631__B1 _11518_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11227__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11663__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11415__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11572__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11377__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08970_ _07431_/Z _08988_/A2 _08970_/B _08971_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07921_ _07921_/A1 _08367_/B _07922_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07852_ input101/Z input102/Z _07854_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06366__A1 _09144_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06803_ _11692_/Q _05633_/B _06803_/B _06804_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11587__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput1 debug_mode input1/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09522_ _09270_/Z _09522_/A2 _09522_/B _09523_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07783_ _07783_/A1 _08504_/C _08317_/B _07783_/A4 _07785_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__08107__A2 _08616_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09304__A1 _09121_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06734_ _11510_/Q _10148_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_36_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09453_ _09472_/A2 _11500_/Q _09454_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06665_ input78/Z input95/Z _06666_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06669__A2 input38/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09384_ _09397_/A2 _11478_/Q _09385_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_319 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10870__B1 _10916_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05616_ _06490_/B1 _06466_/B _05616_/B _05616_/C _05617_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08404_ split15/I _08419_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input100_I wb_adr_i[12] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06596_ _06596_/A1 input115/Z _06599_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09607__A2 _09622_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08335_ _08335_/A1 _08335_/A2 _08642_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05547_ _11695_/Q _05549_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11525__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08266_ _08266_/I _08529_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08197_ _08434_/A1 _08200_/B _08659_/A1 _08332_/A1 _08660_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11654__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06841__A2 _06869_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07217_ _05924_/Z _09154_/I _07218_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07148_ _07148_/I _11170_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09791__A1 _09798_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11406__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10925__A1 _10925_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07079_ _07076_/Z _07083_/A2 _07079_/B _07080_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_120_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10090_ _10090_/A1 _10090_/A2 _11647_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09543__A1 _09547_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10153__A2 _10382_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10992_ _10966_/Z _10992_/A2 _10993_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05580__A2 _06619_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06109__A1 _11275_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1022 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1011 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08347__B _11025_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1055 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1033 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_74 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1099 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1088 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1077 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1066 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_11613_ _11613_/D _11686_/RN _06705_/Z _11613_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_11544_ _11544_/D _11686_/RN _06705_/Z _11544_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_168_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07085__A2 _06238_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10613__B1 _10613_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06832__A2 _05633_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11475_ _11475_/D _11686_/RN _06705_/Z _11475_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__11645__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10426_ _11637_/Q _10426_/A2 _10428_/B2 _10426_/B2 _10426_/C _10428_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__08585__A2 _08315_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09782__A1 _09798_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06045__B1 _11478_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10916__A1 _10916_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_817 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_10357_ _10357_/A1 _11138_/Q _10358_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10288_ _10366_/A1 _11474_/Q _10290_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_839 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_828 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09534__A1 _09547_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06348__A1 _05703_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06899__A2 _06902_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06556__I _06556_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06450_ _06454_/A1 _11070_/Q _06451_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_21_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06381_ _09374_/A1 _11475_/Q _06385_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08120_ _08161_/A1 _08220_/B _08472_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08273__A1 split14/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08051_ _08051_/I _08169_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10080__A1 _10377_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06823__A2 _11076_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07002_ _07002_/I _11129_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09773__A1 _09270_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10383__A2 _06556_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08953_ _08963_/A2 _11343_/Q _08954_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07904_ _08359_/B _08545_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XANTENNA__09525__A1 _09547_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input148_I wb_dat_i[26] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06339__A1 _09699_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08884_ _08888_/A2 _11321_/Q _08885_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10135__A2 _10615_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07835_ _07835_/I _08519_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
X_07766_ _07766_/A1 _08500_/C _07766_/A3 _07766_/A4 _07771_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_09505_ _09505_/I _11516_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06717_ _06717_/I _06718_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09436_ _09436_/I _11494_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07697_ _07697_/I _08290_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10843__B1 _10886_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06648_ input80/Z input79/Z _06649_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_06579_ input105/Z _07863_/I _06583_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09367_ _09367_/I _11472_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11542__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08318_ _08318_/A1 _08690_/A3 _08322_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08264__A1 split14/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09298_ _09298_/I _11450_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08249_ _07682_/I _07685_/I _08249_/B _08250_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11627__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07297__I _07297_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11260_ _11260_/D input162/Z _11666_/CLK _11260_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_11191_ _11191_/D _11686_/RN _06705_/Z _11191_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__08567__A2 _08696_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11692__CLK input68/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10211_ _10367_/A1 _11480_/Q _10213_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09764__A1 _09158_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10142_ _11446_/Q _10363_/A2 _11438_/Q _10363_/B2 _10142_/C _10143_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
Xoutput190 _06625_/ZN mgmt_gpio_oeb[25] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__09516__A1 _09187_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08319__A2 _08417_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10073_ _10371_/A1 _11484_/Q _10075_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10126__A2 _10092_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05553__A2 _05519_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11072__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10975_ _08493_/B input147/Z _10977_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_43_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08255__A1 _08400_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11618__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11527_ _11527_/D _11686_/RN _06705_/Z _11527_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_7_320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06805__A2 _11073_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10062__B2 _10359_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11458_ _11458_/D _11686_/RN _06705_/Z _11458_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__09755__A1 _09121_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10409_ _10506_/A2 _10501_/A2 _10410_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11011__B1 _08460_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11389_ _11389_/D _11686_/RN _06705_/Z _11389_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XTAP_603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09507__A1 _09125_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10117__A2 _11541_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05792__A2 _08839_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05950_ _06839_/A1 _11084_/Q _05953_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_05881_ _09499_/A1 _11521_/Q _05883_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11415__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07620_ _08264_/B _07609_/Z _07623_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08730__A2 _11274_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07551_ _07551_/I _07579_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__06741__A1 input63/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06502_ _06502_/I _06611_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07482_ _07808_/A2 _07793_/A2 _08495_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__11565__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08494__A1 _08589_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09221_ _09221_/I _11426_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06433_ _09016_/A1 _11363_/Q _06437_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09152_ _09125_/Z _09169_/A2 _09152_/B _09153_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06364_ _07412_/A1 _11141_/Q _06217_/Z _06365_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11609__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08103_ _08161_/A1 _08209_/B _08471_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10053__A1 _10350_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08797__A2 _08827_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09083_ _06859_/Z _09089_/A2 _09083_/B _09084_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06295_ _08940_/A1 _11340_/Q _06296_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08034_ _08034_/A1 _08034_/A2 _08036_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xinput81 spi_sck input81/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput70 mgmt_gpio_in[6] input70/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput92 spimemio_flash_io3_do input92/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_150_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08549__A2 _08692_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06024__A3 _06024_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10356__A2 _11136_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09985_ _09985_/I _10365_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__10271__I _11330_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08936_ _08936_/I _11337_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_76_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11095__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08867_ _07426_/Z _08888_/A2 _08867_/B _08868_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07818_ _08347_/A1 _08339_/A1 _07819_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08798_ _08798_/I _11294_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07749_ _08304_/B _08580_/A2 _07754_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10760_ _10884_/A1 _11385_/Q _10763_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09419_ _09241_/Z _09422_/A2 _09419_/B _09420_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10292__A1 _10371_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10691_ _10691_/A1 _10691_/A2 _10691_/A3 _10691_/A4 _10698_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_12_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08237__A1 split12/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10044__A1 _11379_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08788__A2 _07114_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10595__A2 _11525_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06799__A1 _06835_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11312_ _11312_/D _11686_/RN _06705_/Z _11312_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_11243_ _11243_/D _11686_/RN _06705_/Z _11243_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__11341__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11174_ _11174_/D _11686_/RN _06705_/Z _11174_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__07212__A2 _09125_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11438__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06971__A1 _06843_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05774__A2 _09091_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08960__A2 _08963_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10125_ _10265_/A1 _11325_/Q _10265_/A3 _10126_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11356__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10056_ _10352_/A1 _11356_/Q _10057_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11588__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10958_ _10958_/I _11674_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_466 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10889_ _10889_/A1 _11136_/Q _10890_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10586__A2 _11581_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09976__A1 _10379_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06080_ _11342_/Q _06082_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08400__A1 _08400_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07203__A2 _05924_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09770_ _09241_/I _09773_/A2 _09770_/B _09771_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06982_ _10942_/A1 _06974_/I _06982_/B _06983_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_466 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_500 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08951__A2 _08963_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05765__A2 _08839_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05933_ _05933_/A1 _05933_/A2 _05933_/A3 _05933_/A4 _05939_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_08721_ _07426_/Z _08724_/A2 _08721_/B _08722_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_08652_ _08692_/A2 _08361_/B _08653_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09900__A1 _09952_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05864_ _11553_/Q _09599_/A1 _11545_/Q _09574_/A1 _05864_/C _05868_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_07603_ _08637_/B _07774_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__06714__A1 _11056_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05795_ _05795_/I _09424_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
X_08583_ _08583_/A1 _08493_/B _08584_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_07534_ _07751_/A1 _07994_/A1 _07535_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08467__A1 split8/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07465_ _07465_/I _07466_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10274__A1 _10353_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06416_ _08839_/A1 _11087_/Q _06872_/A2 _06418_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09204_ _09220_/A2 _11421_/Q _09205_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06493__A3 _06491_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07396_ _07081_/Z _07396_/A2 _07396_/B _07397_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10026__A1 _10359_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06347_ _05703_/Z _08795_/A1 _11145_/Q _06349_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_5_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_09135_ _09142_/A2 _11400_/Q _09136_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10577__A2 _11445_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input76_I porb VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06278_ _08839_/A1 _11088_/Q _06872_/A2 _06280_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09066_ _09066_/A1 _09015_/Z _09089_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__09719__A1 _09241_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08017_ _08562_/A1 _08017_/A2 _08391_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09195__A2 _09195_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09968_ _11523_/Q _10373_/B1 _11515_/Q _10373_/A1 _09968_/C _09983_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__06402__B1 _11323_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08942__A2 _08963_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08919_ _08938_/A2 _11332_/Q _08920_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09899_ _09899_/I _10265_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_4
XFILLER_168_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10812_ _10903_/A1 _11562_/Q _10817_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10743_ _10924_/A1 _11328_/Q _10744_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11110__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07130__A1 _05927_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07681__A2 _08395_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10674_ _10674_/A1 _10674_/A2 _10675_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05692__A1 _05703_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09965__I _09965_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_3_2__f_wb_clk_i_I clkbuf_0_wb_clk_i/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10568__A2 _11405_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11260__CLK _11666_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07485__I _07485_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05995__A2 _05995_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07197__A1 _07197_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11226_ _11226_/D _11686_/RN _06705_/Z _11226_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_4_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11157_ _11157_/D _11686_/RN _06705_/Z _11157_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_67_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_10108_ _11453_/Q _10365_/A2 _10365_/B1 _11461_/Q _10111_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_11088_ _11088_/D _11686_/RN _06705_/Z _11088_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_63_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10039_ _10039_/I _10042_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06172__A2 _11620_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08449__A1 _08449_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05580_ _05509_/I _06619_/A1 _05580_/A3 _05581_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_51_506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10256__B2 _11561_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07250_ _06847_/Z _07265_/A2 _07250_/B _07251_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05683__A1 _05683_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07181_ _07197_/A1 _11177_/Q _07182_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11603__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06201_ _09674_/A1 _11572_/Q _06206_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06132_ _11581_/Q _09699_/A1 _11573_/Q _09674_/A1 _06132_/C _06148_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_8_470 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10559__A2 _06556_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06227__A3 _06217_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06063_ _06063_/A1 _06063_/A2 _06063_/A3 _06063_/A4 _06064_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_09822_ _09823_/A2 _11618_/Q _09823_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10731__A2 _11560_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09753_ _09753_/I _11595_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06935__A1 _06837_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08704_ _05703_/Z _08786_/A1 _06838_/Z _08709_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_06965_ _06965_/I _11118_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input130_I wb_dat_i[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06896_ _06859_/Z _06902_/A2 _06896_/B _06897_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09684_ _09697_/A2 _11574_/Q _09685_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05916_ _09117_/A1 _11400_/Q _05917_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08635_ _07844_/B _11258_/Q _08646_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10495__A1 _10410_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05847_ _11337_/Q _10233_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08566_ _08566_/A1 _08475_/Z _08620_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11133__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07517_ split5/I _07522_/I _07524_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05910__A2 _09399_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05778_ _06238_/I _05803_/A2 _05779_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08497_ _08678_/A1 _08590_/A2 _08497_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__07112__A1 _05927_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07448_ _07522_/I split13/I _07506_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__08860__A1 _06855_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07379_ _07076_/Z _07382_/A2 _07379_/B _07380_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_13_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11283__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09118_ _09142_/A2 _11395_/Q _09119_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10390_ _10456_/A1 _10415_/A2 _10391_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output182_I _06044_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06218__A3 _06217_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09049_ _06847_/Z _09064_/A2 _09049_/B _09050_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_150_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07179__A1 _05925_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09168__A2 _11410_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11011_ _08431_/B input135/Z _08460_/B input144/Z _11012_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08915__A2 _06838_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10722__A2 _11448_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_285 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06926__A1 _07398_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09340__A2 _11464_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06154__A2 _11501_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07351__A1 _07076_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09891__A3 _09927_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11626__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10238__B2 _10355_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10726_ _10899_/A1 _11504_/Q _10728_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07654__A2 _08417_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08851__A1 _07431_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10657_ _10914_/B1 _11607_/Q _10658_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05665__A1 _08825_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10588_ _10911_/A1 _11573_/Q _10589_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06209__A3 _11033_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05968__A2 _05968_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10961__A2 _11025_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06090__A1 _08890_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08906__A2 _11328_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11209_ _11209_/D _11656_/CLK _11209_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10713__A2 _10888_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06917__A1 _06843_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11156__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06750_ _06760_/A1 _11028_/A2 _06751_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_95_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09331__A2 _11461_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05701_ _05703_/I _08791_/A1 _05702_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06681_ _06681_/I _06681_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_182 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08420_ _08414_/Z _08420_/A2 _08627_/I _08538_/A1 _08422_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_05632_ _11066_/Q _05515_/I _05633_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07342__A1 _07419_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07893__A2 split13/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10229__A1 _10092_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08351_ _08351_/I _08383_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_05563_ _11691_/Q _05565_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09095__A1 _09114_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08282_ _08666_/A3 _08664_/A2 _08282_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__07645__A2 _08417_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07302_ _08839_/A1 _07419_/A2 _06871_/Z _07307_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_05494_ _05576_/C _06456_/A2 _05526_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11130__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07233_ _11321_/Q _05924_/Z _07233_/B _07235_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07164_ _05925_/Z _09121_/I _07165_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08070__A2 split13/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07095_ _07095_/I _11155_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06115_ _06839_/A1 _11081_/Q _06118_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_172_293 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06046_ _11502_/Q _10148_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06081__A1 _05723_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07997_ _07997_/A1 _07997_/A2 _07997_/A3 _07998_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA_input39_I mgmt_gpio_in[12] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06384__A2 _06238_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09805_ _09121_/I _09823_/A2 _09805_/B _09806_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11197__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09736_ _09154_/I _09725_/Z _09736_/B _09737_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06948_ _06941_/I _11113_/Q _06949_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09667_ _09667_/I _11568_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06879_ _07201_/A1 _06838_/Z _06902_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__06136__A2 _09599_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08618_ _08227_/B _08696_/A2 _08618_/B _08618_/C _08619_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_131_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11649__CLK _11665_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07333__A1 _10957_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09598_ _09598_/I _11546_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08549_ _08549_/A1 _08692_/A2 _08549_/B _08549_/C _08550_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_24_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09086__A1 _06863_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05895__A1 _10954_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11560_ _11560_/D _11686_/RN _06705_/Z _11560_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__07636__A2 _07609_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06439__A3 _06439_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10640__A1 _10913_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_repeater345_I input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10511_ _10514_/I _11323_/Q _10513_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_155_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11491_ _11491_/D _11686_/RN _06705_/Z _11491_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__08633__B _08672_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10442_ _10442_/A1 _10442_/A2 _10442_/A3 _10443_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_10373_ _10373_/A1 _11150_/Q _10373_/B1 _11154_/Q _10376_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11179__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09010__A1 _06863_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11188__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10459__A1 _10922_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06127__A2 _09091_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07324__A1 _07310_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09077__A1 _06851_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05886__A1 _09171_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11360__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10631__A1 _11526_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10709_ _10709_/A1 _10709_/A2 _10709_/A3 _10709_/A4 _10737_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__10631__B2 _10902_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11689_ _11689_/D _11042_/ZN input68/Z _11689_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnsnq_1
XANTENNA__08052__A2 _07522_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07920_ _07920_/I _08367_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_46_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05810__A1 _06217_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09001__A1 _06851_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07851_ _07851_/A1 _07851_/A2 _07855_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11179__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10698__A1 _10698_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07782_ _08592_/A2 _08505_/B _07783_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06802_ _10986_/A1 _05633_/B _06803_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput2 debug_oeb input2/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06366__A2 _11403_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09521_ _09522_/A2 _11522_/Q _09522_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06733_ _11478_/Q _06733_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07315__A1 _07310_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09452_ _09452_/I _11499_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06664_ _06664_/A1 _11187_/Q _06666_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06595_ _06595_/I _06596_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09383_ _09383_/I _11477_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05877__A1 _09399_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_08403_ _08403_/A1 _08403_/A2 _08403_/A3 _08403_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__10870__A1 _10915_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05615_ _06466_/B _11064_/Q _05616_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_358 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11351__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09068__A1 _07426_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08334_ _08347_/A1 _08513_/A2 _08335_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05546_ _05546_/I _11697_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11103__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08265_ _08400_/A1 _07616_/I _08265_/B _08266_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08196_ _08478_/B _07722_/I _08196_/B _08618_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06752__I input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07216_ _07216_/I _11183_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07147_ _07147_/A1 _07151_/B _07147_/B _07148_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_133_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11321__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10925__A2 _10092_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05801__A1 _11522_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07078_ _07083_/A2 _11151_/Q _07079_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06029_ _06029_/A1 _06029_/A2 _06029_/A3 _06029_/A4 _06035_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__05801__B2 _09474_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10138__B1 _11358_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11471__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_214 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10991_ _10991_/A1 _10991_/A2 _10991_/A3 _10992_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11590__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09719_ _09241_/Z _09722_/A2 _09719_/B _09720_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11079__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output312_I _11666_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1001 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1056 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1045 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1034 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1023 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11342__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1089 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_11612_ _11612_/D _11686_/RN _06705_/Z _11612_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__11632__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10613__A1 _10410_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11543_ _11543_/D _11686_/RN _06705_/Z _11543_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__07085__A3 _06871_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10613__B2 _10494_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11474_ _11474_/D _11686_/RN _06705_/Z _11474_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__06293__A1 _08915_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06662__I _06662_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10425_ _10408_/I _10425_/A2 _10426_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06045__B2 _09374_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06045__A1 _11486_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10377__B1 _10377_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09973__I _09973_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_10356_ _10356_/A1 _11136_/Q _10358_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_829 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_10287_ _11458_/Q _10365_/A2 _10365_/B1 _11466_/Q _10290_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09534__A2 _11526_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06348__A2 _08786_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09922__B _09922_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06837__I _09116_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10852__A1 _10852_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05859__B2 _09066_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11333__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06380_ _06380_/A1 _06380_/A2 _06380_/A3 _06380_/A4 _06391_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__08273__A2 _07609_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08050_ _08114_/A1 _08067_/A1 _08067_/A2 _08051_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_119_249 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11344__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06284__A1 _07419_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07001_ _06837_/Z _07004_/A2 _07001_/B _07002_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08025__A2 _08545_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06036__A1 _06036_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07784__A1 _07722_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09773__A2 _09773_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11494__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08952_ _08952_/I _11342_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07903_ _07903_/A1 _07903_/A2 _07903_/A3 _07903_/A4 _07912_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__09525__A2 _11523_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08883_ _08883_/I _11320_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07536__A1 _08339_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07834_ _08600_/A1 _08358_/A2 _07835_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07765_ _07537_/I _07761_/I _07766_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09504_ _09121_/Z _09522_/A2 _09504_/B _09505_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07696_ _07696_/A1 _08541_/A2 _07704_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06716_ _06753_/A1 input87/Z _06717_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05651__I _05651_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09435_ _09154_/Z _09447_/A2 _09435_/B _09436_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11324__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_06647_ _06650_/A1 _11310_/Q _06649_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10843__A1 _10886_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_09366_ _09187_/Z _09372_/A2 _09366_/B _09367_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06578_ _09857_/A1 _09927_/A2 _09950_/A1 _11090_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_08317_ _08686_/A2 _08689_/B _08317_/B _08690_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08264__A2 _07609_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05529_ _06460_/A1 _05529_/A2 _05529_/B _05529_/C _05541_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_09297_ _09270_/Z _09297_/A2 _09297_/B _09298_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08248_ split21/Z _07609_/Z _08248_/B _08403_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06027__A1 _08846_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08179_ _08242_/B _08490_/A3 _08180_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10210_ _11456_/Q _10365_/A2 _10365_/B1 _11464_/Q _10213_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09213__A1 _09220_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11190_ _11190_/D _11686_/RN _06705_/Z _11190_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__09764__A2 _09773_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11020__A1 _10966_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06578__A2 _09927_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output262_I _11292_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10141_ _10141_/A1 _10141_/A2 _10142_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput191 _10634_/A2 mgmt_gpio_oeb[26] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__09516__A2 _09522_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput180 _10144_/B2 mgmt_gpio_oeb[16] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_10072_ _11508_/Q _10369_/A2 _10369_/B1 _11500_/Q _10075_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10126__A3 _10126_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11217__CLK _11672_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10974_ _11016_/A1 input141/Z _10977_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10834__A1 _10092_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11315__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11571__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11367__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11526_ _11526_/D _11686_/RN _06705_/Z _11526_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_11_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10062__A2 _10359_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11457_ _11457_/D _11686_/RN _06705_/Z _11457_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__09204__A1 _09220_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09755__A2 _09773_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10408_ _10408_/I _10501_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11011__A1 _08431_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11388_ _11388_/D _11686_/RN _06705_/Z _11388_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_10339_ _10378_/A1 _11155_/Q _10341_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_604 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10770__B1 _10897_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09507__A2 _09522_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11524__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05880_ _11473_/Q _09349_/A1 _11465_/Q _09324_/A1 _05880_/C _05893_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_120_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11554__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07550_ _07675_/A2 _07733_/A1 _07551_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__06741__A2 input80/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06501_ _05572_/B _05576_/C _06502_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11306__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09691__A1 _09187_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07481_ _07522_/I split13/I _07793_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__11539__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09878__I _09878_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09220_ _06867_/Z _09220_/A2 _09220_/B _09221_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06432_ _06432_/A1 _06432_/A2 _06432_/A3 _06432_/A4 _06438_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__09443__A1 _09447_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09151_ _09169_/A2 _11405_/Q _09152_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06363_ _07398_/A1 _11139_/Q _06217_/Z _06365_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_08102_ _08434_/A1 _08209_/B _08215_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09082_ _09089_/A2 _11384_/Q _09083_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08033_ _07840_/I _07555_/I _08033_/B _08034_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06294_ _07006_/A2 _11106_/Q _11033_/A2 _06296_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xinput60 mgmt_gpio_in[31] input60/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput82 spi_sdo input82/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput71 mgmt_gpio_in[7] input71/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput93 spimemio_flash_io3_oeb input93/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11002__A1 _11016_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input160_I wb_dat_i[8] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06024__A4 _06024_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09984_ _09984_/A1 _10030_/A2 _09985_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07509__A1 _08315_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08935_ _06863_/Z _08938_/A2 _08935_/B _08936_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input21_I mask_rev_in[25] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08866_ _08888_/A2 _11315_/Q _08867_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11545__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07817_ _07570_/I _08495_/B _08347_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_17_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08797_ _08797_/A1 _08827_/A2 _08797_/B _08798_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07748_ _07748_/I _08304_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__09682__A1 _09125_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07679_ _07699_/A2 _07989_/A2 _07680_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10292__A2 _11490_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09418_ _09422_/A2 _11489_/Q _09419_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10690_ _10690_/A1 _10690_/A2 _10690_/A3 _10690_/A4 _10691_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_178_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08237__A2 _08614_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09434__A1 _09447_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09349_ _09349_/A1 _09015_/Z _09372_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_12_147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06248__A1 _09449_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10044__A2 _10355_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11311_ _11311_/D _11686_/RN _06705_/Z _11311_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_126_506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06799__A2 _09121_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11242_ _11242_/D _11686_/RN _06705_/Z _11242_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_164_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11173_ _11173_/D _11686_/RN _06705_/Z _11173_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10124_ _10124_/A1 _10124_/A2 _10124_/A3 _10124_/A4 _10126_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__06420__A1 _09091_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10055_ _10353_/A1 _11364_/Q _10057_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11536__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10807__A1 _10899_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10957_ _10957_/A1 _10934_/I _10957_/B _10958_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10283__A2 _11426_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10888_ _10888_/A1 _11138_/Q _10890_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09425__A1 _09447_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06239__A1 _06238_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10035__A2 _09876_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11509_ _11509_/D _11686_/RN _06705_/Z _11509_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__07739__A1 _08589_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08400__A2 _08686_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06411__A1 _08799_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06981_ _06974_/I _11123_/Q _06982_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_05932_ _08846_/A1 input66/Z _05933_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08720_ _08724_/A2 _11271_/Q _08721_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11527__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08651_ _08651_/A1 _08651_/A2 _08651_/A3 _08651_/A4 _08655_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_05863_ _05863_/A1 _05863_/A2 _05864_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11532__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09900__A2 _10265_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07602_ _07760_/A1 _07793_/A2 _08637_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06714__A2 input89/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10510__A3 _10510_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05794_ _06238_/I _08719_/A2 _05795_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08582_ _08582_/A1 _08582_/A2 _08582_/A3 _08581_/Z _08583_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__05922__B1 _11448_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07533_ _07533_/I _07994_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XANTENNA__08467__A2 _07722_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11682__CLK _06687_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07464_ input100/Z input103/Z _07465_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10274__A2 _11370_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06415_ _06785_/A1 _11071_/Q _06418_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09203_ _09203_/I _11420_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09416__A1 _09187_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07395_ _07396_/A2 _11243_/Q _07396_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09134_ _09134_/I _11399_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_175_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07978__A1 split14/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06346_ _09649_/A1 _11563_/Q _06349_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06277_ _06785_/A1 _11072_/Q _06280_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09065_ _09065_/I _11378_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09719__A2 _09722_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08016_ _08016_/I _08017_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input69_I mgmt_gpio_in[5] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11062__CLK input68/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06402__A1 _11101_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09967_ _09967_/A1 _09967_/A2 _09968_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06402__B2 _08890_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08918_ _08918_/I _11331_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_990 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11518__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09898_ _09898_/A1 _10030_/A1 _09952_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output225_I _11170_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08849_ _08849_/I _11309_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10811_ _10904_/A1 _11554_/Q _10817_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10265__A2 _11329_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10742_ _10742_/A1 _10742_/A2 _10742_/A3 _10742_/A4 _10742_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__07130__A2 _09154_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10673_ _10892_/A1 _11471_/Q _10674_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09407__A1 _09125_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10457__I _10457_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05692__A2 _06872_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07969__A1 split14/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11405__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06641__A1 _11606_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06670__I input75/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11225_ _11225_/D input162/Z _06687_/A2 _11225_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__08394__A1 _08394_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11555__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11156_ _11156_/D _11686_/RN _06705_/Z _11156_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_68_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_11087_ _11087_/D _11686_/RN _06705_/Z _11087_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_10107_ _10107_/A1 _10107_/A2 _10107_/A3 _10107_/A4 _10107_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_67_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08146__A1 _08434_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10038_ _10353_/A1 _11363_/Q _10045_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09646__A1 _09647_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10256__A2 _10377_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07121__A2 _05927_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06200_ _06200_/A1 _06200_/A2 _06200_/A3 _06200_/A4 _06212_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__06880__A1 _06902_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07180_ _11201_/Q _05925_/Z _07180_/B _07182_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10008__A2 _09878_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06131_ _06131_/A1 _06131_/A2 _06132_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11085__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06062_ _08846_/A1 input64/Z _06063_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06632__A1 input77/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10964__B1 _11027_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10716__B1 _10886_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09821_ _09821_/I _11617_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10192__A1 _10192_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09752_ _09116_/I _09773_/A2 _09752_/B _09753_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08137__A1 split7/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05924__I _05924_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08703_ _08703_/I _11260_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06964_ _10957_/A1 _06941_/I _06964_/B _06965_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06895_ _06902_/A2 _11098_/Q _06896_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09683_ _09683_/I _11573_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09885__A1 _09898_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05915_ _09144_/A1 _11408_/Q _05917_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08634_ _08460_/B _08634_/A2 _08634_/B1 _08493_/B _08634_/C _08646_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__10495__A2 _10417_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input123_I wb_adr_i[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05846_ _11329_/Q _08890_/A1 _08803_/A1 _05841_/Z _05846_/C _05860_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__06699__A1 _06266_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09637__A1 _09647_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08565_ _08222_/B _08696_/A2 _08565_/B _08565_/C _08566_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_05777_ _05777_/I _06238_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
X_07516_ _07516_/A1 _07614_/A1 _08400_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11340__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08496_ _08299_/I _08496_/A2 _08590_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07112__A2 _06701_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07447_ _07447_/I split13/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__08860__A2 _08863_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11428__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07378_ _07382_/A2 _11238_/Q _07379_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06329_ _06329_/A1 _06329_/A2 _06329_/A3 _06329_/A4 _06392_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_09117_ _09117_/A1 _09015_/Z _09142_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__11355__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11578__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07586__I _07586_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09048_ _09064_/A2 _11373_/Q _09049_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output175_I _10615_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11010_ _08493_/B input153/Z _11012_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10183__A1 _10375_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07179__A2 _09158_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06926__A2 _07006_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08128__A1 _08161_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09628__A1 _09647_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10238__A2 _10355_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08300__A1 _08339_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10725_ _10725_/A1 _10725_/A2 _10725_/A3 _10725_/A4 _10737_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_9_213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08851__A2 _08863_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10656_ _10914_/A1 _11599_/Q _10658_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05665__A2 _06872_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10587_ _10913_/A2 _11589_/Q _10589_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09800__A1 _09800_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06090__A2 _11326_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11208_ _11208_/D _11656_/CLK _11208_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10174__B2 _11463_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07590__A2 _08095_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08119__A1 _08434_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11139_ _11139_/D _11686_/RN _06705_/Z _11139_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_55_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06680_ _11326_/Q input1/Z _06680_/B _06681_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05700_ _05700_/I _08791_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__07342__A2 _06217_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05631_ _06466_/B _11067_/Q _05633_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08350_ _08545_/A1 _08395_/A1 _08351_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09619__A1 _09241_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05562_ _05562_/I _11693_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07301_ _07301_/I _11205_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08281_ _08281_/A1 _08519_/A2 _08280_/B _08666_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05493_ _11068_/Q _06456_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06853__A1 _06851_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07232_ _05924_/Z _09241_/I _07233_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07163_ _07163_/I _11173_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06114_ _06114_/A1 _06114_/A2 _06114_/A3 _06119_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_145_464 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07094_ _07076_/Z _07097_/A2 _07094_/B _07095_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06045_ _11486_/Q _09399_/A1 _11478_/Q _09374_/A1 _06045_/C _06058_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__06081__A2 _11350_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08358__A1 _08623_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09804_ _09823_/A2 _11612_/Q _09805_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10165__A1 _10356_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07996_ _08054_/A1 _07996_/A2 _07997_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11100__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09735_ _09725_/Z _11590_/Q _09736_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07581__A2 _07593_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05592__A1 _06466_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06947_ _06947_/A1 _06947_/A2 _11112_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_09666_ _09187_/Z _09672_/A2 _09666_/B _09667_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08617_ _08617_/A1 _08617_/A2 _08617_/A3 _08617_/A4 _08697_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_06878_ _06878_/I _11088_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07333__A2 _07310_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09597_ _09270_/Z _09597_/A2 _09597_/B _09598_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11250__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05829_ _10957_/A1 _05969_/I _05830_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08548_ _08435_/Z _07922_/I _08548_/A3 _08548_/A4 _08608_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__09086__A2 _09089_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05895__A2 _05969_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08479_ _08479_/A1 _08479_/A2 _08568_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07097__A1 _07081_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11490_ _11490_/D _11686_/RN _06705_/Z _11490_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__10640__A2 _11582_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10510_ _10510_/A1 _10487_/Z _10510_/A3 _10510_/A4 _10513_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__06844__A1 _06869_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08833__A2 _11305_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10441_ _10900_/A1 _11507_/Q _10442_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_156_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10372_ _10372_/A1 _10372_/A2 _10372_/A3 _10381_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__06072__A2 _09649_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09010__A2 _09013_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08521__A1 _08521_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09077__A2 _09089_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05886__A2 _11417_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10631__A2 _10902_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10708_ _11584_/Q _10913_/B2 _10913_/A2 _11592_/Q _10709_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06835__A1 _06835_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11688_ _11688_/D _11688_/RN input68/Z _11688_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_139_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10639_ _11622_/Q _10916_/A1 _11614_/Q _10915_/A1 _10639_/C _10644_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__11123__CLK _11672_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05810__A2 _06872_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10147__B2 _10377_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09001__A2 _09013_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07850_ input99/Z input100/Z _07851_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10698__A2 _10092_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07781_ _08689_/B _08505_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06801_ _11677_/Q _10986_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11273__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09520_ _09520_/I _11521_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06732_ _11454_/Q _10144_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xinput3 debug_out input3/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09451_ _09116_/Z _09472_/A2 _09451_/B _09452_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06663_ input95/Z _06664_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06594_ _06594_/A1 input129/Z input167/Z _06599_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09382_ _09125_/Z _09397_/A2 _09382_/B _09383_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05877__A2 _11489_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08402_ split15/Z _08248_/B _08403_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09068__A2 _09089_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05614_ _05614_/I _07419_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_177_320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08333_ _08333_/I _08336_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05545_ _05545_/A1 _05519_/I _05545_/B _05546_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07079__A1 _07076_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08264_ split14/Z _07609_/Z _08264_/B _08413_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05629__A2 _05515_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08195_ _08195_/I _11254_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07215_ _07240_/A1 _07215_/A2 _07215_/B _07216_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07146_ _11195_/Q _05927_/Z _07151_/B _07146_/C _07147_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_07077_ _05703_/Z _07412_/A1 _06871_/Z _07083_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_06028_ _05660_/Z _11623_/Q _06029_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input51_I mgmt_gpio_in[23] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput340 _11213_/Q wb_dat_o[5] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__11616__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05801__A2 _09499_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10138__A1 _11366_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10138__B2 _10352_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09718_ _09722_/A2 _11585_/Q _09719_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07979_ split15/Z _08380_/B _08650_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10990_ _08431_/B input132/Z _08460_/B input140/Z _10991_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_142_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1013 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1002 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_09649_ _09649_/A1 _09015_/I _09672_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_35_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1046 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1024 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1068 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1057 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_11611_ _11611_/D _11686_/RN _06705_/Z _11611_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_42_178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06817__A1 _06835_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11542_ _11542_/D _11686_/RN _06705_/Z _11542_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_168_364 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10613__A2 _10613_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11473_ _11473_/D _11686_/RN _06705_/Z _11473_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__11146__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10424_ _11636_/Q _11641_/Q _10426_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07242__A1 _05927_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06045__A2 _09399_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10377__B2 _11262_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10377__A1 _10377_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08990__A1 _08990_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10355_ _11130_/Q _10355_/A2 _11120_/Q _10355_/B2 _10355_/C _10364_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_151_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_819 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11296__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10286_ _10286_/A1 _10286_/A2 _10286_/A3 _10286_/A4 _10304_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__05556__A1 _05519_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06348__A3 _11261_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07545__A2 split16/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08742__A1 _08742_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10301__A1 _10379_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05859__A2 _09091_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11097__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07481__A1 _07522_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06284__A2 _07006_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07000_ _07004_/A2 _11129_/Q _07001_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06036__A2 _06036_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11639__CLK _11666_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09222__A2 _09015_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07784__A2 _08689_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08951_ _06851_/Z _08963_/A2 _08951_/B _08952_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08981__A1 _08988_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07902_ _07926_/I _08549_/A1 _07903_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08882_ _06859_/Z _08888_/A2 _08882_/B _08883_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07536__A2 _08614_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07833_ _07833_/A1 _07833_/A2 _07843_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10540__A1 _10902_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07764_ _07722_/I _07761_/I _07766_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09503_ _09522_/A2 _11516_/Q _09504_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07695_ _07691_/I _07697_/I _07492_/I _08541_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_06715_ _06715_/I _06755_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09434_ _09447_/A2 _11494_/Q _09435_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_06646_ _06646_/A1 _06646_/A2 _06646_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11169__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09365_ _09372_/A2 _11472_/Q _09366_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06577_ _06577_/A1 _06556_/I _09950_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08316_ _08316_/A1 _08586_/A2 _08504_/B _08318_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09296_ _09297_/A2 _11450_/Q _09297_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05528_ _06446_/I _05528_/A2 _05501_/Z _06491_/B _05529_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA_input99_I wb_adr_i[11] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08247_ split21/Z _07609_/Z _08247_/B _08411_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06027__A2 input65/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08178_ _08240_/B _08242_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07224__A1 _07240_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09213__A2 _11424_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10359__B2 _10359_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07129_ _11167_/Q _07132_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07775__A2 _08586_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput170 _11295_/Q irq[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__08972__A1 _08988_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10140_ _10361_/A1 _11422_/Q _10141_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput192 _10634_/B2 mgmt_gpio_oeb[27] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput181 _10144_/A1 mgmt_gpio_oeb[17] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_10071_ _10071_/A1 _10071_/A2 _10071_/A3 _10084_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11260__RN input162/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08724__A1 _07431_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08639__B _08639_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10531__A1 _10892_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10973_ _10973_/I _11675_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10295__B1 _10373_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11525_ _11525_/D _11686_/RN _06705_/Z _11525_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_11456_ _11456_/D _11686_/RN _06705_/Z _11456_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__09204__A2 _11421_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07215__A1 _07240_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10407_ _10407_/A1 _11639_/Q _10408_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11387_ _11387_/D _11686_/RN _06705_/Z _11387_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_112_426 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10338_ _10377_/A1 _11145_/Q _10377_/B1 _11261_/Q _10341_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08963__A1 _06867_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_616 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10770__B2 _11465_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11251__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07518__A2 split13/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10269_ _10269_/I _11652_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07480_ _07513_/I split16/I _07808_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06500_ _06500_/A1 _05603_/B _06500_/B1 _06479_/C _11060_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09691__A2 _09697_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11311__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05701__A1 _05703_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06431_ _06933_/A1 _11109_/Q _06432_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09150_ _09150_/I _11404_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06362_ _09171_/A1 _11411_/Q _06365_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11461__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08101_ _08101_/A1 _08101_/A2 _08105_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09081_ _09081_/I _11383_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06293_ _08915_/A1 _11332_/Q _06912_/A1 _11104_/Q _06296_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_174_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08032_ _08032_/A1 _08032_/A2 _08032_/A3 _08034_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xinput50 mgmt_gpio_in[22] input50/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput61 mgmt_gpio_in[32] input61/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11490__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput72 mgmt_gpio_in[8] input72/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput94 trap input94/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput83 spi_sdoenb input83/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11078__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05927__I _05927_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09983_ _09983_/A1 _09983_/A2 _09983_/A3 _09983_/A4 _10046_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__08954__A1 _06855_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input153_I wb_dat_i[30] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11242__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10761__A1 _10883_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08934_ _08938_/A2 _11337_/Q _08935_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07509__A2 split5/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08706__A1 _07426_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09903__B1 _10265_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10513__B2 _10880_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10513__A1 _10513_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08865_ _08865_/A1 _06838_/Z _08888_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_07816_ _07816_/A1 _08513_/A2 _08335_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06193__A1 _05703_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08796_ _08797_/A1 _07114_/C _11294_/Q _08797_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07747_ _07747_/A1 _07808_/A1 _07748_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input14_I mask_rev_in[19] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07678_ _08438_/C _08438_/B _08386_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__09682__A2 _09697_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06629_ _06629_/I _06629_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09417_ _09417_/I _11488_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_498 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_09348_ _09348_/I _11466_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10229__B _10229_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09279_ _09121_/Z _09297_/A2 _09279_/B _09280_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_11310_ _11310_/D _11686_/RN _06705_/Z _11310_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__11481__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09198__A1 _09220_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11241_ _11241_/D _11686_/RN _06705_/Z _11241_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_11172_ _11172_/D _11172_/RN input68/Z _11172_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__08945__A1 _07431_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10752__A1 _10910_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10123_ _10123_/A1 _10123_/A2 _10123_/A3 _10124_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11233__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10054_ _11348_/Q _10351_/A2 _11340_/Q _10351_/B2 _10054_/C _10067_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__06184__A1 _07398_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11334__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09122__A1 _09142_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10807__A2 _11506_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10956_ _10934_/I _11674_/Q _10957_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11484__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10887_ _11140_/Q _10887_/A2 _10887_/B1 _11142_/Q _10890_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09425__A2 _11491_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11472__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11508_ _11508_/D _11686_/RN _06705_/Z _11508_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__09189__A1 _09187_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11439_ _11439_/D input76/Z _06705_/Z _11439_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__11224__RN input162/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10743__A1 _10924_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06980_ _06980_/A1 _06980_/A2 _11122_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_435 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06411__A2 _08839_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05931_ _06197_/I _05636_/I _08846_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA_input6_I mask_rev_in[11] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06175__A1 _06175_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08650_ _08650_/A1 _08650_/A2 _08650_/A3 _08651_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05862_ _09549_/A1 _11537_/Q _05863_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07601_ _07601_/I _07760_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08581_ _08581_/A1 _08182_/I _08491_/I _08581_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_05793_ _05793_/I _09474_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_81_335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09113__A1 _09114_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07532_ _07532_/I _07751_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07463_ input127/Z input99/Z _07463_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06414_ _06839_/A1 _11079_/Q _06418_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09202_ _09121_/Z _09220_/A2 _09202_/B _09203_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09416__A2 _09422_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07394_ _07394_/I _11242_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07427__A1 _07427_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_09133_ _06855_/Z _09142_/A2 _09133_/B _09134_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06345_ _09624_/A1 _11555_/Q _06349_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07978__A2 _08380_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10982__A1 _08493_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06276_ _06839_/A1 _11080_/Q _06280_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09064_ _06867_/Z _09064_/A2 _09064_/B _09065_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05989__A1 _05723_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08015_ _08015_/A1 _08015_/A2 _08016_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11463__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11207__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09966_ _10375_/A1 _11539_/Q _09967_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11357__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_980 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09897_ _09984_/A1 _09898_/A1 _09986_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08917_ _07426_/Z _08938_/A2 _08917_/B _08918_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_991 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_08848_ _07426_/Z _08863_/A2 _08848_/B _08849_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06166__A1 _06166_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08779_ _08779_/I _11289_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09104__A1 _09114_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10810_ _11530_/Q _10902_/A2 _11522_/Q _10902_/B2 _10810_/C _10817_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__10265__A3 _10265_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10741_ _10919_/A1 _11368_/Q _10742_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_159_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10672_ _10891_/A1 _11479_/Q _10674_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09407__A2 _09422_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11523__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08091__A1 _08434_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11454__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06641__A2 input80/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11224_ _11224_/D input162/Z _11683_/CLK _11224_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__10725__A1 _10725_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11206__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09591__A1 _09187_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08394__A2 _08545_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11155_ _11155_/D _11686_/RN _06705_/Z _11155_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_11086_ _11086_/D _11686_/RN _06705_/Z _11086_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_10106_ _11445_/Q _10363_/A2 _11437_/Q _10363_/B2 _10106_/C _10107_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__09343__A1 _09347_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10037_ _10039_/I _09973_/I _10353_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__06157__A1 _09144_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05904__A1 _09649_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09646__A2 _11562_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10939_ _10934_/I _11668_/Q _10940_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08118__I _08575_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_172_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08082__A1 split12/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06130_ _09624_/A1 _11557_/Q _06131_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06061_ _07201_/A1 input55/Z _06063_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10964__B2 _08460_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10964__A1 _08431_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08909__A1 _08913_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10716__B2 _11400_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10716__A1 _10886_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09582__A1 _09125_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09820_ _09241_/I _09823_/A2 _09820_/B _09821_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06396__A1 _06396_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09751_ _09773_/A2 _11595_/Q _09752_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06963_ _06941_/I _11118_/Q _06964_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10192__A2 _06556_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05914_ _11520_/Q _09499_/A1 _11512_/Q _09474_/A1 _05914_/C _05923_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__09334__A1 _09347_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08702_ _08702_/A1 _07844_/B _08702_/B _08703_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06894_ _06894_/I _11097_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09682_ _09125_/I _09697_/A2 _09682_/B _09683_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08633_ _08633_/A1 _08633_/A2 _08672_/B _08634_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05845_ _05845_/A1 _05845_/A2 _05845_/A3 _05846_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_08564_ _08564_/A1 _08564_/A2 _08563_/Z _08584_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05776_ _05776_/A1 _05776_/A2 _05777_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input116_I wb_adr_i[27] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07515_ _07515_/A1 _07515_/A2 _07614_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08495_ _08686_/A2 _07537_/I _08495_/B _08496_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_120_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07446_ _07997_/A2 _07997_/A3 _07846_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__06320__A1 _09775_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11684__RN input162/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07377_ _08825_/A2 _11033_/A2 _06838_/Z _07382_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__06771__I _07110_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06328_ _06328_/A1 _06328_/A2 _06328_/A3 _06328_/A4 _06329_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_09116_ _09116_/I _09116_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA_input81_I spi_sck VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09047_ _09047_/I _11372_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06259_ _06259_/A1 _06259_/A2 _06259_/A3 _06259_/A4 _06259_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__10707__A1 _10911_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06387__A1 _09474_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10183__A2 _11543_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06926__A3 _06871_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09949_ _11646_/Q _10086_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09325__A1 _09347_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06139__A1 _08846_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07107__I _07110_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11675__RN input162/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10724_ _11456_/Q _10897_/A2 _10897_/B1 _11464_/Q _10725_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06311__A1 _08825_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10655_ _10655_/A1 _10655_/A2 _11659_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11522__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06681__I _06681_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10586_ _10913_/B2 _11581_/Q _10589_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09800__A2 _09015_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11477__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06378__A1 _06238_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11672__CLK _11672_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08367__A2 _08355_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11207_ _11207_/D _11686_/RN _06705_/Z _11207_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_11138_ _11138_/D _11686_/RN _06705_/Z _11138_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__09316__A1 _09187_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11069_ _11069_/D _11069_/RN input68/Z _11069_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_48_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05630_ _05630_/A1 _05630_/A2 _05633_/B _11260_/Q _05716_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07342__A3 _06871_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09619__A2 _09622_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05561_ _05561_/A1 _05519_/I _05561_/B _05562_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07300_ _05616_/C _11216_/Q _07300_/B _07300_/C _07301_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08280_ split14/Z _07609_/Z _08280_/B _08540_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05492_ _11069_/Q _05576_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11666__RN input162/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06853__A2 _06869_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07231_ _07231_/I _11186_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07162_ _07197_/A1 _07162_/A2 _07162_/B _07163_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06066__B1 _09750_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11418__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06113_ _08803_/A1 _11298_/Q _06114_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07093_ _07097_/A2 _11155_/Q _07094_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06044_ _06044_/A1 _05786_/I _05783_/I _10144_/A1 _06045_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__08358__A2 _08358_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09803_ _09803_/I _11611_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06369__A1 _06217_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07995_ _07995_/I _08054_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XANTENNA__09307__A1 _09125_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09734_ _09734_/I _11589_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06946_ _06941_/I _11112_/Q _06947_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09665_ _09672_/A2 _11568_/Q _09666_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06877_ _06843_/Z _06877_/A2 _06877_/B _06878_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08616_ split8/Z _07727_/I _08616_/B _08617_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05828_ _05828_/A1 _05828_/A2 _05828_/A3 _10957_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__06766__I _07110_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09596_ _09597_/A2 _11546_/Q _09597_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08547_ _08692_/A2 _08367_/B _08548_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05603__C _05616_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05759_ _05759_/I _06785_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XANTENNA__11545__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08294__A1 _08395_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08478_ _08478_/A1 _08462_/I _08478_/B _08479_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07429_ _07426_/Z _07433_/A2 _07429_/B _07430_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06844__A2 _11080_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11657__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10440_ _10440_/A1 _10427_/B _10900_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_136_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06057__B1 _11446_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11409__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output285_I _11288_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09794__A1 _09798_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11695__CLK input68/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10371_ _10371_/A1 _11245_/Q _10372_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09546__A1 _09547_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08349__A2 _07297_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10156__A2 _10880_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07021__A2 _11135_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06780__A1 _05616_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11075__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08521__A2 _11016_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08285__A1 _07455_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10707_ _10911_/A1 _11576_/Q _10709_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11648__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06835__A2 _09270_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08037__A1 _08037_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11687_ _11687_/D _11687_/RN input68/Z _11687_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
X_10638_ _10638_/A1 _10416_/I _10638_/B _10639_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10919__A1 _10919_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09785__A1 _09798_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10569_ _10887_/B1 _11429_/Q _10572_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10395__A2 _09934_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09537__A1 _09547_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10147__A2 _10377_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11418__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07780_ _07793_/A1 _07808_/A1 _08689_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06800_ _06800_/I _11072_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06731_ _11446_/Q _06731_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xinput4 mask_rev_in[0] input4/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09450_ _09472_/A2 _11499_/Q _09451_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11568__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08401_ _08401_/A1 _08250_/I _08528_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06523__A1 _06610_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06662_ _06662_/I _06662_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07866__A4 split16/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06593_ input121/Z input120/Z _06594_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09381_ _09397_/A2 _11477_/Q _09382_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05613_ _05753_/A1 _05940_/A1 _05614_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08332_ _08332_/A1 _08417_/A2 _08332_/B _08333_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05544_ _05519_/I _11697_/Q _05545_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08276__A1 split14/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08263_ _08411_/A1 _08263_/A2 _08263_/A3 _08408_/B _08263_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__11639__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07214_ _07240_/A1 _11183_/Q _07215_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08194_ _08194_/A1 _08194_/A2 _08194_/B _08195_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07145_ _05927_/Z _09241_/I _07146_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09776__A1 _09798_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07076_ _09116_/I _07076_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_06027_ _08846_/A1 input65/Z _06029_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09528__A1 _09547_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput330 _11668_/Q wb_dat_o[25] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput341 _11214_/Q wb_dat_o[6] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA_input44_I mgmt_gpio_in[17] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10138__A2 _10353_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11098__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07978_ split14/Z _08380_/B _08648_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09717_ _09717_/I _11584_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05565__A2 _05519_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06762__A1 _06701_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06929_ _06929_/I _11107_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09700__A1 _09722_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09648_ _09648_/I _11562_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1003 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06514__A1 _06446_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1025 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1014 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_09579_ _09121_/Z _09597_/A2 _09579_/B _09580_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_output200_I _10638_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1069 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_11610_ _11610_/D _11686_/RN _06705_/Z _11610_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_1058 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_11541_ _11541_/D _11686_/RN _06705_/Z _11541_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__10074__A1 _10370_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10613__A3 _10417_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06817__A2 _11075_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08019__A1 _07837_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11472_ _11472_/D _11686_/RN _06705_/Z _11472_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__09767__A1 _09187_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06164__C _06164_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10423_ _11637_/Q _11638_/Q _10428_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07242__A2 _07242_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10354_ _10354_/A1 _10354_/A2 _10355_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09519__A1 _09241_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08990__A2 _06838_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10285_ _11450_/Q _10363_/A2 _11442_/Q _10363_/B2 _10285_/C _10286_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__08742__A2 _06904_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06753__A1 _06753_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10301__A2 _11562_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08258__A1 _08400_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07481__A2 split13/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09758__A1 _09125_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07233__A2 _05924_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11240__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08950_ _08963_/A2 _11342_/Q _08951_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07901_ _07685_/I _07700_/I _07926_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08881_ _08888_/A2 _11320_/Q _08882_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07832_ _07827_/I _07570_/I _07833_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08733__A2 _11275_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11390__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09502_ _09502_/I _11515_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07763_ _07763_/I _08500_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07694_ _07694_/A1 _07694_/A2 _07697_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10828__B1 _10920_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06714_ _11056_/Q input89/Z _06715_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09433_ _09433_/I _11493_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06645_ input80/Z input81/Z _06646_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08249__A1 _07682_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09364_ _09364_/I _11471_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_08315_ _08332_/A1 _08417_/A2 _08315_/B _08504_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06576_ _09935_/B _09927_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__10056__A1 _10352_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09295_ _09295_/I _11449_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05527_ _06610_/A3 _05515_/I _06491_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_08246_ _08246_/A1 _08246_/A2 _08246_/B _08349_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08177_ _08490_/A1 _08181_/A3 _08240_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07128_ _07128_/I _11166_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_284 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10359__A2 _10359_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08421__A1 split15/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07059_ _07060_/A2 _11146_/Q _07060_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08972__A2 _11349_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput193 _10146_/A2 mgmt_gpio_oeb[28] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput182 _06044_/A1 mgmt_gpio_oeb[18] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_153_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10070_ _10367_/A1 _11476_/Q _10071_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output248_I _06658_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput171 _06746_/Z irq[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_47_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10972_ _10972_/A1 _10966_/Z _10972_/B _10973_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_474 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10295__B2 _11530_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10295__A1 _10373_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11113__CLK _11672_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10047__A1 _10047_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09988__A1 _10366_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11524_ _11524_/D _11686_/RN _06705_/Z _11524_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_144_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11455_ _11455_/D _11686_/RN _06705_/Z _11455_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__06671__B1 _11056_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10406_ _10406_/I _10506_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
X_11386_ _11386_/D _11686_/RN _06705_/Z _11386_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10337_ _10337_/A1 _10337_/A2 _10337_/A3 _10342_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08963__A2 _08963_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_606 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10770__A2 _10897_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10268_ _10305_/A1 _10880_/C _10268_/B _10269_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_639 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10199_ _10199_/A1 _10199_/A2 _10200_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_179_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06430_ _07398_/A1 _07006_/A2 _11107_/Q _06432_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__05701__A2 _08791_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10038__A1 _10353_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11606__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06361_ _09197_/A1 _11419_/Q _06365_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08100_ _08100_/I _08101_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06292_ _05941_/I _05719_/I _06912_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09080_ _06855_/Z _09089_/A2 _09080_/B _09081_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08031_ _08031_/I _08032_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_147_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput40 mgmt_gpio_in[13] input40/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput51 mgmt_gpio_in[23] input51/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput62 mgmt_gpio_in[33] input62/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput73 mgmt_gpio_in[9] input73/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput84 spimemio_flash_clk input84/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput95 uart_enabled input95/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10210__B2 _11464_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09982_ _10377_/A1 _11571_/Q _10377_/B1 _11563_/Q _09983_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08954__A2 _08963_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08933_ _08933_/I _11336_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08864_ _08864_/I _11314_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input146_I wb_dat_i[24] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09903__B2 _09922_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07815_ _07555_/I _08495_/B _07816_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06193__A2 _07412_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08795_ _08795_/A1 _08799_/A1 _08797_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07746_ _07746_/I _07808_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11136__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10277__B2 _10355_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07677_ _07907_/A1 _07892_/I _08438_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09416_ _09187_/Z _09422_/A2 _09416_/B _09417_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06628_ _06628_/A1 input77/Z _06628_/B _06629_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06774__I _07110_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08890__A1 _08890_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09347_ _09270_/Z _09347_/A2 _09347_/B _09348_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06559_ _10392_/A1 _11638_/Q _06560_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11286__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09278_ _09297_/A2 _11444_/Q _09279_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10229__C _10880_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08229_ _08079_/I _08199_/I _08481_/B _08482_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_11240_ _11240_/D _11686_/RN _06705_/Z _11240_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__09198__A2 _11419_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11171_ _11171_/D _11686_/RN _06705_/Z _11171_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__06405__B1 _08803_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10201__A1 _10356_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08945__A2 _08963_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10122_ _10378_/A1 _11549_/Q _10123_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10053_ _10350_/A1 _10053_/A2 _10054_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06708__A1 _06753_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06184__A2 _08825_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10955_ _10955_/I _11673_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11629__CLK _11665_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08881__A1 _08888_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10886_ _11134_/Q _10886_/A2 _11132_/Q _10886_/B2 _10886_/C _10890_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__06239__A3 _11033_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11507_ _11507_/D _11686_/RN _06705_/Z _11507_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_117_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10934__I _10934_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08404__I split15/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11438_ _11438_/D _11686_/RN _06705_/Z _11438_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__09189__A2 _09195_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11369_ _11369_/D _11686_/RN _06705_/Z _11369_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_98_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_403 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10743__A2 _11328_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06411__A3 input94/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06859__I _09187_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05930_ _05930_/A1 _05940_/A1 _06197_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__11159__CLK input68/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_05861_ _05693_/Z _11529_/Q _05863_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08164__A3 _08242_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08580_ _08243_/B _08580_/A2 _08582_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07372__A1 _07076_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07600_ _07600_/A1 _07600_/A2 _08408_/C _08260_/B _07606_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_07531_ _07675_/A2 input97/Z _07532_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05792_ _06238_/I _08839_/A2 _05793_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_293 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07462_ _07462_/A1 _07462_/A2 _07865_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08872__A1 _08888_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07393_ _07076_/Z _07396_/A2 _07393_/B _07394_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09201_ _09220_/A2 _11420_/Q _09202_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06413_ _06413_/A1 _06413_/A2 _06413_/A3 _06413_/A4 _06419_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_06344_ _06344_/A1 _06344_/A2 _06350_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09132_ _09142_/A2 _11399_/Q _09133_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10431__A1 _10444_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07427__A2 _06904_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09063_ _09064_/A2 _11378_/Q _09064_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06275_ _06275_/A1 _06275_/A2 _06275_/A3 _06275_/A4 _06281_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_08014_ _08014_/I _08562_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__06938__A1 _06843_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09965_ _09965_/I _10375_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_970 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06769__I _07110_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09896_ _09896_/I _09984_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08916_ _08938_/A2 _11331_/Q _08917_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_981 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_08847_ _08863_/A2 _11309_/Q _08848_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06166__A2 _06166_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07363__A1 _07398_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08778_ _06859_/Z _08784_/A2 _08778_/B _08779_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07115__A1 _05927_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07729_ _08054_/A2 _07808_/A2 _07822_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08863__A1 _06859_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10740_ _10922_/A1 _11360_/Q _10742_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11151__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10670__A1 _10884_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10671_ _10671_/A1 _10671_/A2 _10671_/A3 _10671_/A4 _10691_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_43_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11223_ _11223_/D input162/Z _11683_/CLK _11223_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__10186__B1 _10378_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11301__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09591__A2 _09597_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11154_ _11154_/D _11686_/RN _06705_/Z _11154_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_68_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11085_ _11085_/D input76/Z _06705_/Z _11085_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_10105_ _10105_/A1 _10105_/A2 _10106_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09343__A2 _11465_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10489__B2 _10911_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10036_ _10352_/A1 _11355_/Q _10045_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11451__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07354__A1 _07081_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06157__A2 _11405_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10929__I _11666_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11077__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11390__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10938_ _10938_/A1 _10950_/A2 _10940_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08854__A1 _06847_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10661__A1 _10911_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11142__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10869_ _10914_/A1 _11242_/Q _10871_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_157_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06060_ _05927_/I input46/Z _06063_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10964__A2 _11029_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06093__A1 _06093_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08909__A2 _11329_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05840__A1 _06266_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09582__A2 _09597_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09750_ _09750_/A1 _09015_/I _09773_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_06962_ _06962_/I _11117_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09681_ _09697_/A2 _11573_/Q _09682_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05913_ _05913_/A1 _05913_/A2 _05914_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08701_ _07844_/B _11260_/Q _08702_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06893_ _06855_/Z _06902_/A2 _06893_/B _06894_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08632_ _08294_/B _08632_/A2 _08290_/C _08633_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_94_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05844_ _08761_/A1 _11290_/Q _05845_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08563_ _08563_/A1 _08563_/A2 _08563_/A3 _08563_/A4 _08563_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_05775_ _05775_/A1 _05775_/A2 _05775_/A3 _05775_/A4 _05828_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__09098__A1 _09114_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07514_ _07888_/A2 _07506_/I _08046_/B _07515_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08494_ _08589_/A1 _08494_/A2 _08494_/B _08494_/C _08678_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA_input109_I wb_adr_i[20] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07445_ _07445_/I _07997_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XANTENNA__05659__A1 _08825_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10652__A1 _10652_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10247__A4 _10247_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11133__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07376_ _07376_/I _11237_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06327_ _09750_/A1 _11595_/Q _06328_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09115_ _09115_/I _11394_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06258_ _06258_/A1 _06258_/A2 _06258_/A3 _06258_/A4 _06259_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__06084__A1 _06785_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input74_I pad_flash_io0_di VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11324__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09046_ _07431_/Z _09064_/A2 _09046_/B _09047_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06189_ _09574_/A1 _11540_/Q _06194_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11474__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09948_ _09948_/I _11645_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_180_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06139__A2 input63/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09879_ _09898_/A1 _10040_/A2 _09927_/A2 _11632_/Q _09902_/I _09880_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_38_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10891__A1 _10891_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09089__A1 _06867_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08300__A3 _08358_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10723_ _10896_/A1 _11440_/Q _10725_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06311__A2 _08825_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10654_ _10881_/A1 _11659_/Q _10655_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10585_ _10910_/A1 _11565_/Q _10589_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09261__A1 _09272_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05822__A1 _06217_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09013__A1 _06867_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11206_ _11206_/D _11686_/RN _06705_/Z _11206_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__07575__A1 _07575_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11137_ _11137_/D _11686_/RN _06705_/Z _11137_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_95_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07327__A1 _07310_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11068_ _11068_/D _11068_/RN input68/Z _11068_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_91_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10019_ _10019_/I _10357_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_36_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_358 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05560_ _05519_/I _11693_/Q _05561_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10634__B2 _10634_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05491_ input58/Z _06786_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_07230_ _07240_/A1 _07230_/A2 _07230_/B _07231_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11347__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07161_ _07197_/A1 _11173_/Q _07162_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10608__B _10608_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09252__A1 _09272_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06066__A1 _06324_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06112_ _08829_/A1 _11304_/Q _06114_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11497__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07092_ _07092_/A1 _06904_/Z _07097_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06043_ _11462_/Q _10144_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09004__A1 _06855_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09802_ _09116_/I _09823_/A2 _09802_/B _09803_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_5_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06369__A2 _11033_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07994_ _07994_/A1 _07551_/I _07995_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_09733_ _09125_/I _09725_/Z _09733_/B _09734_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06945_ _10938_/A1 _06957_/A2 _06947_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07318__A1 _10942_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09664_ _09664_/I _11567_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06876_ _06877_/A2 _11088_/Q _06877_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10468__A4 _10467_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09595_ _09595_/I _11545_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08615_ _08693_/A1 _08615_/A2 _08615_/A3 _08615_/A4 _08634_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_05827_ _05827_/A1 _05827_/A2 _05827_/A3 _05827_/A4 _05828_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__11354__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10873__A1 _10921_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08546_ _08546_/I _08692_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_05758_ _08791_/A1 _08799_/A1 _05759_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09491__A1 _09187_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08477_ _08477_/I _08619_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05689_ _05689_/I _09599_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XANTENNA__10625__A1 _10896_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11106__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07428_ _07433_/A2 _11252_/Q _07429_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07359_ _07359_/I _11232_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09243__A1 _09241_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10370_ _10370_/A1 _11249_/Q _10372_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output180_I _10144_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output278_I _11077_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09029_ _09039_/A2 _11367_/Q _09030_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09546__A2 _11530_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07557__A1 _07511_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11593__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07309__A1 _11219_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06780__A2 _11687_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10864__A1 _10910_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11345__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06532__A2 _08672_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09482__A1 _09125_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10706_ _10910_/A1 _11568_/Q _10709_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11686_ _11686_/D _11686_/RN _06705_/Z _11686_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__06048__A1 _10148_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10637_ _10914_/B1 _11606_/Q _10638_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06048__B2 _06048_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09785__A2 _11606_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10568_ _10889_/A1 _11405_/Q _10572_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10499_ _10499_/A1 _10387_/I _10902_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_150_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11584__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06867__I _09270_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06730_ _11422_/Q _06730_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xinput5 mask_rev_in[10] input5/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06661_ _11059_/Q _06661_/A2 _06661_/B _06662_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10610__C _10880_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11336__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08400_ _08400_/A1 _08686_/A2 _08400_/B _08400_/C _08401_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_05612_ _05612_/I _05940_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
X_06592_ _06592_/A1 _06592_/A2 input114/Z _06599_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09380_ _09380_/I _11476_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08331_ _08686_/A2 _08674_/B _08331_/B _08675_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05543_ _11696_/Q _05545_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08276__A2 _07609_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08262_ split21/Z _07609_/Z _08262_/B _08408_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07213_ _11317_/Q _05924_/Z _07213_/B _07215_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08028__A2 _08677_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08193_ _07297_/I _11254_/Q _08194_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06039__A1 _10947_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07144_ _11170_/Q _07147_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07787__A1 _08328_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07075_ _07075_/I _11150_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06026_ input48/Z _05927_/Z _07201_/A1 input56/Z _06029_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_145_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09528__A2 _11524_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput331 _11669_/Q wb_dat_o[26] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput320 _11121_/Q wb_dat_o[16] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput342 _11215_/Q wb_dat_o[7] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_160_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10543__B1 _10921_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07977_ _08355_/I _08380_/B _07980_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11575__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input37_I mgmt_gpio_in[10] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11461__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09716_ _09187_/I _09722_/A2 _09716_/B _09717_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06762__A2 _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06928_ _06837_/Z _06931_/A2 _06928_/B _06929_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06777__I _07110_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11512__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10846__A1 _10892_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11327__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09647_ _09270_/Z _09647_/A2 _09647_/B _09648_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06859_ _09187_/I _06859_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_1004 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1037 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11476__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1026 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1015 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_09578_ _09597_/A2 _11540_/Q _09579_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1059 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1048 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_08529_ _08411_/Z _08529_/A2 _07618_/I _08529_/A4 _08687_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__11662__CLK _11663_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11540_ _11540_/D _11686_/RN _06705_/Z _11540_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__06278__A1 _08839_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11471_ _11471_/D _11686_/RN _06705_/Z _11471_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_129_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09216__A1 _09220_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09767__A2 _09773_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10422_ _10422_/A1 _10914_/A1 _10916_/A1 _10904_/A1 _10429_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__07778__A1 _08696_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10353_ _10353_/A1 _11110_/Q _10354_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09519__A2 _09522_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07242__A3 _09015_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05789__B1 _11482_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10782__B1 _10920_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10284_ _10284_/A1 _10284_/A2 _10285_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11566__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06202__A1 _09699_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11429__SETN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11192__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10837__A1 _10887_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11318__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06269__A1 _06694_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11669_ _11669_/D _11683_/CLK _11669_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09207__A1 _09220_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11014__A1 _11014_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09758__A2 _09773_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07769__A1 _08592_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06441__A1 _05584_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07900_ split21/I _08549_/A1 _07903_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08880_ _08880_/I _11319_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11535__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07831_ _07831_/A1 _07831_/A2 _07831_/A3 _07833_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_110_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09501_ _09116_/Z _09522_/A2 _09501_/B _09502_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07762_ _08696_/A2 _08587_/B _07763_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09694__A1 _09241_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07693_ _08630_/A2 _07660_/I _07696_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11685__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10828__A1 _10920_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11309__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06713_ _06713_/A1 _06713_/A2 _06713_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09432_ _09125_/Z _09447_/A2 _09432_/B _09433_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_497 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06644_ _06650_/A1 _11309_/Q _06646_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09363_ _09158_/Z _09372_/A2 _09363_/B _09364_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06575_ _11091_/Q _09935_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09446__A1 _09447_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08249__A2 _07685_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08314_ _08314_/I _08586_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05526_ _05526_/A1 _05575_/A1 _05528_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09997__A2 _10042_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09294_ _09241_/Z _09297_/A2 _09294_/B _09295_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08245_ _07990_/I _08185_/I _08245_/B _08246_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08176_ _08490_/A1 _08176_/A2 _08180_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06680__A1 _11326_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07127_ _07127_/A1 _07151_/B _07127_/B _07128_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_137_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11065__CLK input68/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07058_ _07058_/I _11145_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xoutput194 _10146_/B1 mgmt_gpio_oeb[29] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput183 _06733_/ZN mgmt_gpio_oeb[19] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_06009_ _09349_/A1 _11471_/Q _06010_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput172 _06748_/Z irq[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_10971_ _10966_/Z _10971_/A2 _10972_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10819__A1 _10911_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09685__A1 _09154_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10295__A2 _11522_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07160__A2 _05925_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09437__A1 _09447_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10047__A2 _10382_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11523_ _11523_/D _11686_/RN _06705_/Z _11523_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__11408__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11454_ _11454_/D _11686_/RN _06705_/Z _11454_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__06671__B2 _06724_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10405_ _10417_/I _10427_/B _09920_/I _10903_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__11558__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11385_ _11385_/D _11686_/RN _06705_/Z _11385_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10336_ _10375_/A1 _11685_/Q _10337_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_10267_ _10092_/Z _11651_/Q _10267_/B _10926_/C _10268_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08176__A1 _08490_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10198_ _10352_/A1 _11360_/Q _10199_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09676__A1 _09116_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07151__A2 _05927_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09428__A1 _09447_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09979__A2 _10040_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06360_ _06360_/A1 _06360_/A2 _06360_/A3 _06360_/A4 _06371_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__11088__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06291_ _06291_/A1 _06291_/A2 _06291_/A3 _06302_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_08030_ _08459_/C _08563_/A1 _08031_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput30 mask_rev_in[4] input30/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput52 mgmt_gpio_in[24] input52/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput63 mgmt_gpio_in[34] input63/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput41 mgmt_gpio_in[14] input41/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput96 user_clock input96/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput85 spimemio_flash_csb input85/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09600__A1 _09622_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput74 pad_flash_io0_di input74/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09981_ _09972_/I _09959_/I _10377_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__06414__A1 _06839_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08932_ _06859_/Z _08938_/A2 _08932_/B _08933_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08167__A1 _08167_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09903__A2 _09935_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08863_ _06859_/Z _08863_/A2 _08863_/B _08864_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07914__A1 split21/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07814_ _08696_/A2 _08332_/B _08514_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08794_ _08794_/I _11293_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input139_I wb_dat_i[18] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07745_ _07675_/B split13/Z _07746_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10277__A2 _10355_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07142__A2 _07151_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07676_ _07858_/A2 _07676_/A2 _07892_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09415_ _09422_/A2 _11488_/Q _09416_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06627_ input92/Z input77/Z _06628_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09419__A1 _09241_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08890__A2 _06838_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09346_ _09347_/A2 _11466_/Q _09347_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06558_ _11639_/Q _10392_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06489_ _06489_/A1 _06491_/B _06489_/A3 _06490_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09277_ _09277_/I _11443_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05509_ _05509_/I _06611_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_148_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08228_ _08228_/I _08479_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06653__A1 _11059_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11700__CLK input68/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08159_ _08159_/I _08656_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_146_391 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11170_ _11170_/D _11686_/RN _06705_/Z _11170_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_106_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output260_I _11282_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06405__A1 _11306_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06405__B2 _11645_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10201__A2 _11408_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10121_ _10379_/A1 _11557_/Q _10123_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10052_ _11332_/Q _10053_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06708__A2 input85/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07381__A2 _11239_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10268__A2 _10880_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10954_ _10954_/A1 _10934_/I _10954_/B _10955_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11230__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10885_ _10885_/A1 _10885_/A2 _10886_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06892__A1 _06902_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11506_ _11506_/D _11686_/RN _06705_/Z _11506_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__09830__A1 _09121_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10976__B1 _08460_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11380__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11292__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10440__A2 _10427_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11437_ _11437_/D input76/Z _06705_/Z _11437_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_140_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11368_ _11368_/D _11686_/RN _06705_/Z _11368_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_10319_ _10319_/A1 _10319_/A2 _10320_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08149__A1 split8/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_426 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_11299_ _11299_/D input76/Z _06705_/Z _11299_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_85_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05860_ _05860_/A1 _05860_/A2 _05860_/A3 _05860_/A4 _05894_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__09649__A1 _09649_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05791_ _05791_/I _09499_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
X_07530_ _07530_/I _08339_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_4
X_07461_ input128/Z input102/Z _07462_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06883__A1 _06902_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07392_ _07396_/A2 _11242_/Q _07393_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09200_ _09200_/I _11419_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06412_ _08799_/A1 _11295_/Q _08799_/A2 _06413_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06343_ _05703_/Z _07419_/A2 _11250_/Q _06344_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09131_ _09131_/I _11398_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06635__A1 _11622_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09062_ _09062_/I _11377_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06274_ _08839_/A1 _07419_/A2 _11207_/Q _06275_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_08013_ _08013_/A1 _08013_/A2 _08014_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07060__A1 _06843_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10195__A1 _10350_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09964_ _10018_/A1 _09899_/I _09965_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11103__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_971 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_09895_ _10030_/A1 _09899_/I _09896_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__09888__A1 _09898_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08915_ _08915_/A1 _06838_/Z _08938_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_982 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10498__A2 _10417_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08846_ _08846_/A1 _06904_/Z _08863_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__07363__A2 _08825_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11253__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08777_ _08784_/A2 _11289_/Q _08778_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05989_ _05723_/Z _11351_/Q _05993_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07115__A2 _09116_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07728_ _07593_/I _08358_/A2 _07738_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08863__A2 _08863_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07659_ _07659_/A1 _08663_/B _07684_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06874__A1 _06837_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10670_ _10884_/A1 _11383_/Q _10671_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10670__A2 _11383_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09329_ _09121_/Z _09347_/A2 _09329_/B _09330_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_159_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10422__A2 _10914_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11222_ _11222_/D input162/Z _11666_/CLK _11222_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__10186__A1 _10379_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11153_ _11153_/D _11686_/RN _06705_/Z _11153_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_68_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09879__A1 _09898_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11084_ _11084_/D input76/Z _06705_/Z _11084_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_10104_ _10361_/A1 _11421_/Q _10105_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10489__A2 _10915_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09879__B2 _09902_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10035_ _10039_/I _09876_/I _10352_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_48_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10110__A1 _10367_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10937_ _10937_/A1 _10937_/A2 _11667_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08854__A2 _08863_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06865__A1 _06863_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_10868_ _10914_/B1 _11238_/Q _10871_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10799_ _10891_/A1 _11482_/Q _10801_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_470 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07290__A1 _06867_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11126__CLK _11683_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10177__A1 _10177_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_180 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06961_ _10954_/A1 _06941_/I _06961_/B _06962_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11276__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05912_ _09424_/A1 _11496_/Q _05913_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09680_ _09680_/I _11572_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08700_ _08431_/B _08700_/A2 _11016_/A1 _08700_/B2 _08700_/C _08702_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_11642__346 _11642_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__tieh
X_06892_ _06902_/A2 _11097_/Q _06893_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08542__A1 _07691_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08631_ _08631_/A1 _08631_/A2 _08631_/A3 _08633_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_05843_ _06785_/A1 _11077_/Q _05845_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08562_ _08562_/A1 _08562_/A2 _08563_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05774_ _11394_/Q _09091_/A1 _11386_/Q _09066_/A1 _05774_/C _05775_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_07513_ _07513_/I _08046_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08493_ _08493_/A1 _08493_/A2 _08493_/A3 _08493_/B _08522_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_07444_ _07444_/A1 _07444_/A2 _07445_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__05659__A2 _08719_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06856__A1 _06869_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10652__A2 _10092_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07375_ _07081_/Z _07375_/A2 _07375_/B _07376_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06326_ _07391_/A1 _11242_/Q _06328_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09114_ _06867_/Z _09114_/A2 _09114_/B _09115_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07281__A1 _06855_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06257_ _06257_/A1 _06257_/A2 _06257_/A3 _06257_/A4 _06258_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__06084__A2 _11074_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09045_ _09064_/A2 _11372_/Q _09046_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input67_I mgmt_gpio_in[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11619__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06188_ _09599_/A1 _11548_/Q _06194_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10168__B2 _10359_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08781__A1 _06863_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09947_ _09947_/A1 _09947_/A2 _11092_/Q _06608_/B _09948_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_49_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_790 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_09878_ _09878_/I _10040_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10340__A1 _10379_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08829_ _08829_/A1 _06904_/Z _08837_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__05633__B _05633_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09089__A2 _09089_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10722_ _10895_/A1 _11448_/Q _10725_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08836__A2 _11306_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11149__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10653_ _10092_/Z _11658_/Q _10653_/B _10880_/C _10655_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_70_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10584_ _10584_/A1 _10578_/Z _10583_/Z _10604_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_139_464 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07272__A1 _07081_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09261__A2 _11439_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05822__A2 _08799_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11299__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09013__A2 _09013_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10159__A1 _10350_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11205_ _11205_/D input162/Z _11683_/CLK _11205_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XANTENNA__06378__A3 _11033_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07575__A2 _07525_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08772__A1 _06851_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11136_ _11136_/D _11686_/RN _06705_/Z _11136_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_11067_ _11067_/D _11067_/RN input68/Z _11067_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__10331__A1 _10371_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10018_ _10018_/A1 _10265_/A3 _10019_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_145 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08827__A2 _08827_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10634__A2 _10634_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07160_ _11197_/Q _05925_/Z _07160_/B _07162_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10398__A1 _06563_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06066__A2 _11590_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07091_ _07091_/I _11154_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06111_ _06111_/I _08829_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
X_06042_ _11470_/Q _06044_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09004__A2 _09013_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07015__A1 _06837_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09801_ _09823_/A2 _11611_/Q _09802_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08763__A1 _07426_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10343__C _10343_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07993_ _07993_/A1 _08388_/B _08021_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09732_ _09725_/Z _11589_/Q _09733_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10570__A1 _10887_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08515__A1 _08204_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06944_ _06944_/A1 _06944_/A2 _11111_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07318__A2 _07310_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09663_ _09158_/I _09672_/A2 _09663_/B _09664_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06875_ _06875_/I _11087_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09594_ _09241_/Z _09597_/A2 _09594_/B _09595_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08614_ _08393_/B _08614_/A2 _08615_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05826_ _11458_/Q _09299_/A1 _11450_/Q _09274_/A1 _05826_/C _05827_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA_input121_I wb_adr_i[31] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10873__A2 _11101_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08545_ _08545_/A1 _08545_/A2 _08546_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05757_ _06839_/A1 _11086_/Q _05761_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06829__A1 _06835_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09491__A2 _09497_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08476_ _08134_/I _08462_/I _08476_/B _08476_/C _08477_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05688_ _05703_/I _05803_/A2 _05689_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10625__A2 _11438_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07427_ _07427_/A1 _06904_/Z _07433_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05501__A1 _06610_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07358_ _07076_/Z _07361_/A2 _07358_/B _07359_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06309_ _05924_/Z input36/Z _06313_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09243__A2 _09246_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11441__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07289_ _07290_/A2 _11204_/Q _07290_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09028_ _09028_/I _11366_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11076__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07006__A1 _07419_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11591__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07557__A2 _07614_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05568__A1 _06786_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07309__A2 input162/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10313__A1 _10353_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10864__A2 _11261_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09482__A2 _09497_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07493__A1 _08519_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10705_ _11624_/Q _10916_/A1 _11616_/Q _10915_/A1 _10705_/C _10709_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_11685_ _11685_/D _11686_/RN _06705_/Z _11685_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10636_ _10636_/A1 _10636_/A2 _10636_/A3 _10636_/A4 _10645_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_139_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10567_ _10567_/A1 _10567_/A2 _10567_/A3 _10567_/A4 _10573_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_10498_ _10499_/A1 _10417_/I _10902_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__11281__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10552__B2 _10884_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06220__A2 _11452_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11119_ _11119_/D _11686_/RN _06705_/Z _11119_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xinput6 mask_rev_in[11] input6/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06660_ _11059_/Q input67/Z _06661_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11314__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05611_ _05646_/A1 _05639_/A2 _05612_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06591_ _06591_/I _06592_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05731__B2 _05723_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08330_ _08330_/A1 _08596_/A3 _08511_/B _08336_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05542_ _05542_/I _11698_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10607__A2 _10461_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11464__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07484__A1 _08358_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08261_ _08261_/I _08263_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_32_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07212_ _05924_/Z _09125_/I _07213_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08192_ _08192_/A1 _08246_/B _08194_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07143_ _07143_/I _11169_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xoutput310 _11705_/Z spimemio_flash_io2_di VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_07074_ _06843_/Z _07074_/A2 _07074_/B _07075_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08984__A1 _08988_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput332 _11670_/Q wb_dat_o[27] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_06025_ input68/Z _05924_/Z _05925_/Z input39/Z _06029_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xoutput321 _11122_/Q wb_dat_o[17] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput343 _11111_/Q wb_dat_o[8] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__10791__A1 _10887_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10543__A1 _10920_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07976_ _07976_/I _08380_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
X_09715_ _09722_/A2 _11584_/Q _09716_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06927_ _06931_/A2 _11107_/Q _06928_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09646_ _09647_/A2 _11562_/Q _09647_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06858_ _06858_/I _11083_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1038 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1016 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1005 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_09577_ _09577_/I _11539_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06789_ _08787_/A2 _08787_/A3 _06790_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05809_ _09144_/A1 _11410_/Q _05813_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05722__A1 _07006_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1049 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_08528_ _08528_/A1 _08528_/A2 _08528_/A3 _08528_/A4 _08671_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_42_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08459_ _07720_/I _08033_/B _08459_/B _08459_/C _08460_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_11_502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06278__A2 _11088_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_11470_ _11470_/D _11686_/RN _06705_/Z _11470_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA_output290_I _11088_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09216__A2 _11425_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10421_ _10471_/A1 _10427_/B _10904_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__07227__A1 _05924_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07778__A2 _08315_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05789__A1 _11490_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08975__A1 _08988_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10352_ _10352_/A1 _11108_/Q _10354_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05789__B2 _09374_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10782__A1 _10920_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09924__B1 _09927_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10283_ _10361_/A1 _11426_/Q _10284_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10534__A1 _10904_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11337__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05961__A1 _08799_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09152__A1 _09125_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11487__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05713__A1 _11586_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05713__B2 _09674_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_11668_ _11668_/D _11672_/CLK _11668_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09207__A2 _11422_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11014__A2 _10966_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11599_ _11599_/D _11686_/RN _06705_/Z _11599_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10619_ _10619_/A1 _10619_/A2 _10619_/A3 _10619_/A4 _10645_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_182_370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10222__B1 _10373_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08966__A1 _08988_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10773__A1 _10903_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11254__RN input162/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10525__A1 _10891_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07830_ _08341_/B _08677_/A2 _07831_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09391__A1 _09187_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07761_ _07761_/I _08587_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09500_ _09522_/A2 _11515_/Q _09501_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05952__A1 _06785_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06712_ _11056_/Q input68/Z _06713_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09694__A2 _09697_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07692_ _08294_/B split5/Z _08630_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06643_ _06643_/I _06643_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09431_ _09447_/A2 _11493_/Q _09432_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05704__A1 _05703_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09362_ _09372_/A2 _11471_/Q _09363_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06574_ _06574_/A1 _06556_/I _09857_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08313_ _07508_/I _08686_/A2 _08313_/B _08314_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05525_ _05576_/B _05575_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09293_ _09297_/A2 _11449_/Q _09294_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08244_ _08244_/A1 _08581_/A1 _08492_/B _08246_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_08175_ _08170_/I _07492_/I _08176_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06680__A2 input1/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07209__A1 _07240_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07126_ _11191_/Q _05927_/Z _07151_/B _07126_/C _07127_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_137_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08957__A1 _06859_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10764__A1 _10891_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11245__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07057_ _06837_/Z _07060_/A2 _07057_/B _07058_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08709__A1 _07431_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10516__A1 _10916_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06008_ _09324_/A1 _11463_/Q _06010_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput173 _06681_/Z mgmt_gpio_oeb[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput184 _06678_/Z mgmt_gpio_oeb[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput195 _06082_/B2 mgmt_gpio_oeb[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__06196__A1 _09649_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09382__A1 _09125_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07959_ _07959_/I _08375_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_46_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10970_ _10970_/A1 _10970_/A2 _10970_/A3 _10971_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__09685__A2 _09697_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09629_ _09121_/I _09647_/A2 _09629_/B _09630_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_output303_I _05947_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07448__A1 _07522_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11522_ _11522_/D _11686_/RN _06705_/Z _11522_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_7_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11453_ _11453_/D _11686_/RN _06705_/Z _11453_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_10404_ _10404_/A1 _11636_/Q _10417_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__08948__A1 _06847_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11236__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11384_ _11384_/D _11686_/RN _06705_/Z _11384_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10335_ _10374_/A1 _11157_/Q _10337_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10266_ _10247_/Z _10092_/I _10266_/A3 _10266_/A4 _10267_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_608 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06187__A1 _06187_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10197_ _10353_/A1 _11368_/Q _10199_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05934__A1 _09800_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09676__A2 _09697_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05698__B1 _11546_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10443__B1 _11499_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06290_ _08795_/A1 _07006_/A2 _11130_/Q _06291_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11460__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput31 mask_rev_in[5] input31/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput20 mask_rev_in[24] input20/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput53 mgmt_gpio_in[25] input53/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput64 mgmt_gpio_in[35] input64/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11502__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput42 mgmt_gpio_in[15] input42/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05777__I _05777_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput97 wb_adr_i[0] input97/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput86 spimemio_flash_io0_do input86/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11227__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput75 pad_flash_io1_di input75/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07611__A1 _08417_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09980_ _09980_/I _10377_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XANTENNA__06414__A2 _11079_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11475__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08931_ _08938_/A2 _11336_/Q _08932_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08862_ _08863_/A2 _11314_/Q _08863_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11652__CLK _11665_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07813_ _07813_/A1 _07813_/A2 _07819_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_96_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08793_ _07426_/Z _08793_/A2 _08793_/B _08794_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07744_ _07744_/A1 _08494_/C _07754_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_72_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07675_ _07533_/I _07675_/A2 _07675_/B _07676_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06626_ _11314_/Q _06628_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09414_ _09414_/I _11487_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11413__SETN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09419__A2 _09422_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09345_ _09345_/I _11465_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06557_ _06574_/A1 _10092_/I _06577_/A1 _06557_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
X_06488_ _06488_/A1 _06490_/B1 _06489_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09276_ _09116_/Z _09297_/A2 _09276_/B _09277_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input97_I wb_adr_i[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05508_ _06451_/A1 _11068_/Q _05509_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10985__A1 _10966_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11466__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08227_ split7/Z _08232_/A2 _08227_/B _08228_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11428__SETN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11182__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08158_ _08158_/A1 _08158_/A2 _08165_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10737__A1 _10737_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11218__RN input162/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08089_ _08089_/I _08090_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07109_ _07110_/I _11162_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10120_ _10377_/A1 _11573_/Q _10377_/B1 _11565_/Q _10123_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_10051_ _11324_/Q _10558_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07905__A2 _08519_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06169__A1 _05584_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09107__A1 _09114_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10953_ _10934_/I _11673_/Q _10954_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_10884_ _10884_/A1 _11130_/Q _10885_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11525__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11505_ _11505_/D _11686_/RN _06705_/Z _11505_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__07841__A1 _08545_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11457__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10976__A1 _08431_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11436_ _11436_/D input76/Z _06705_/Z _11436_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__09594__A1 _09241_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08397__A2 _08460_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11675__CLK _06687_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11367_ _11367_/D _11686_/RN _06705_/Z _11367_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_10318_ _10357_/A1 _11137_/Q _10319_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09346__A1 _09347_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_11298_ _11298_/D input76/Z _06705_/Z _11298_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10249_ _10366_/A1 _11473_/Q _10251_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09897__A2 _09898_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10900__A1 _10900_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05790_ _08791_/A1 _06238_/I _05791_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09649__A2 _09015_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07460_ input98/Z input101/Z _07462_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06332__A1 _05703_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07391_ _07391_/A1 _06904_/Z _07396_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06411_ _08799_/A1 _08839_/A2 input94/Z _06413_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_147_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06342_ _09674_/A1 _11571_/Q _06344_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09130_ _06851_/Z _09142_/A2 _09130_/B _09131_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11448__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10967__A1 _11016_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09061_ _06863_/Z _09064_/A2 _09061_/B _09062_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08012_ _08012_/A1 _07457_/I _08013_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06635__A2 input77/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06273_ _08839_/A1 _08839_/A2 _11308_/Q _06275_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__10719__A1 _10892_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09585__A1 _09154_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09963_ _09887_/I _09878_/I _10018_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input151_I wb_dat_i[29] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11620__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09337__A1 _09347_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08914_ _08914_/I _11330_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_961 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_950 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_09894_ _11635_/Q _09899_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_994 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_983 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_972 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_08845_ _08845_/I _11308_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07363__A3 _06871_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08776_ _08776_/I _11288_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07727_ _07727_/I _08696_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XANTENNA_input12_I mask_rev_in[17] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05988_ _11391_/Q _09091_/A1 _11383_/Q _09066_/A1 _05988_/C _05993_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__11548__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07658_ _07660_/I _08686_/A2 _08663_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07589_ _07589_/A1 _07589_/A2 _07589_/A3 _08255_/B _07595_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_06609_ _06609_/I _11091_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09328_ _09347_/A2 _11460_/Q _09329_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11698__CLK input68/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11439__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10422__A3 _10916_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09259_ _09154_/Z _09272_/A2 _09259_/B _09260_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09576__A1 _09116_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11221_ _11221_/D input162/Z _11683_/CLK _11221_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_11152_ _11152_/D _11686_/RN _06705_/Z _11152_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__09328__A1 _09347_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10103_ _10360_/A1 _11429_/Q _10105_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09879__A2 _10040_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11083_ _11083_/D _11686_/RN _06705_/Z _11083_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_68_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10034_ _10034_/A1 _10265_/A3 _10039_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_48_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11078__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06011__B1 _11479_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09500__A1 _09522_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06314__A1 _05927_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10110__A2 _11477_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10936_ _10934_/I _11667_/Q _10937_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11678__RN input162/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10867_ _11246_/Q _10913_/A2 _11250_/Q _10913_/B2 _10867_/C _10871_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__06865__A2 _06869_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_293 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_10798_ _10798_/A1 _10798_/A2 _10798_/A3 _10798_/A4 _10826_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__06078__B1 _11358_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07814__A1 _08696_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07290__A2 _07290_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11419_ _11419_/D input76/Z _06705_/Z _11419_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__11602__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09319__A1 _09241_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06960_ _06941_/I _11117_/Q _06961_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06891_ _06891_/I _11096_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05911_ _09449_/A1 _11504_/Q _05913_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input4_I mask_rev_in[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08542__A2 _07492_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08630_ _07660_/I _08630_/A2 _08630_/B _08630_/C _08631_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05842_ _06839_/A1 _11085_/Q _05845_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08561_ _08561_/A1 _08561_/A2 _08613_/A1 _08564_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_05773_ _05773_/A1 _05773_/A2 _05774_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07512_ split5/I _07888_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08492_ _08185_/I _07564_/I _08492_/B _08492_/C _08493_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__06305__A1 _05969_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07443_ _06591_/I input106/Z _07444_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07374_ _07375_/A2 _11237_/Q _07375_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09113_ _09114_/A2 _11394_/Q _09114_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06325_ _08825_/A2 _11238_/Q _11033_/A2 _06328_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_30_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07281__A2 _07290_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06256_ _07419_/A2 _06238_/I _11150_/Q _06257_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09044_ _09044_/I _11371_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06187_ _06187_/A1 _06187_/A2 _06187_/A3 _06259_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__10168__A2 _10359_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11220__CLK _11672_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08781__A2 _08784_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09946_ _09946_/A1 _11092_/Q _11645_/Q _09947_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06792__A1 _06835_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09730__A1 _09121_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09877_ _11632_/Q _11631_/Q _09878_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08828_ _08828_/I _11303_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11370__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11291__SETN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08759_ _06859_/Z _08759_/A2 _08759_/B _08760_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08297__A1 _08204_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10721_ _11496_/Q _10894_/A2 _11488_/Q _10894_/B2 _10721_/C _10725_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__08049__A1 _08315_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10267__B _10267_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10652_ _10652_/A1 _10092_/Z _10650_/Z _10652_/A4 _10653_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__09797__A1 _09798_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10583_ _10583_/A1 _10583_/A2 _10583_/A3 _10583_/A4 _10583_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_166_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07272__A2 _07290_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09549__A1 _09549_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11204_ _11204_/D _11686_/RN _06705_/Z _11204_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_141_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07024__A2 _11136_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08772__A2 _08784_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11135_ _11135_/D _11686_/RN _06705_/Z _11135_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_95_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11066_ _11066_/D _11066_/RN input68/Z _11066_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__09721__A1 _09722_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08524__A2 _07844_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10017_ _11443_/Q _10363_/A2 _11435_/Q _10363_/B2 _10017_/C _10027_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__08288__A1 _08614_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10095__A1 _10353_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10919_ _10919_/A1 _11110_/Q _10923_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09788__A1 _09798_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07090_ _07081_/Z _07090_/A2 _07090_/B _07091_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10398__A2 _09920_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06110_ _08839_/A1 _08795_/A1 _06111_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11243__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06041_ _06041_/I _11267_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08212__A1 _08575_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07992_ _08385_/I _08357_/A2 _08388_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09800_ _09800_/A1 _09015_/I _09823_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__09960__A1 _10042_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08763__A2 _08784_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09731_ _09731_/I _11588_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06943_ _06941_/I _11111_/Q _06944_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11393__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10570__A2 _11421_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09712__A1 _09722_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09662_ _09672_/A2 _11567_/Q _09663_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06874_ _06837_/Z _06877_/A2 _06874_/B _06875_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09593_ _09597_/A2 _11545_/Q _09594_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08613_ _08613_/A1 _08613_/A2 _08613_/A3 _08615_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_05825_ _05825_/A1 _05825_/A2 _05826_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08544_ _08544_/A1 _08291_/I _08544_/A3 _08544_/A4 _08584_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA_input114_I wb_adr_i[25] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05756_ _05756_/I _06839_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_08475_ _08475_/A1 _08475_/A2 _08475_/A3 _08475_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_05687_ _05687_/I _05703_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__06829__A2 _11077_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10087__B _10880_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07426_ _09116_/I _07426_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__09779__A1 _09798_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07357_ _07361_/A2 _11232_/Q _07358_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06308_ _06308_/I _11264_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07288_ _07288_/I _11203_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09027_ _06851_/Z _09039_/A2 _09027_/B _09028_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06239_ _06238_/Z _11241_/Q _11033_/A2 _06241_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__07006__A2 _07006_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05568__A2 _05519_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output333_I _11671_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09703__A1 _09722_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09929_ _09929_/I _11640_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_171_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11116__CLK _11672_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10077__A1 _10375_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_split15_I split15/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07493__A2 _08358_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10704_ _10704_/A1 _10704_/A2 _10705_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11684_ _11684_/D input162/Z _06687_/A2 _11684_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10635_ _10635_/I _10636_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_139_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10566_ _10886_/A2 _11397_/Q _10567_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10497_ _10503_/A2 _10501_/A2 _10499_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_11118_ _11118_/D _11672_/CLK _11118_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10552__A2 _10896_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11049_ _11050_/I _11696_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xinput7 mask_rev_in[12] input7/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10304__A2 _10382_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06508__A1 _06446_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07181__A1 _07197_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05610_ _05610_/I _05639_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06590_ input106/Z input113/Z _06592_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10068__A1 _11452_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05731__A2 _08990_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11609__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05541_ _05541_/A1 _05541_/A2 _05541_/B _05542_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07484__A2 split5/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08681__A1 _08681_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08260_ _08400_/A1 _08625_/B _08260_/B _08261_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08191_ _08191_/I _08246_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07211_ _07211_/I _11182_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07142_ _07142_/A1 _07151_/B _07142_/B _07143_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07073_ _07074_/A2 _11150_/Q _07074_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput300 _06408_/Z reset VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__10240__A1 _10357_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput311 _11706_/Z spimemio_flash_io3_di VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput333 _11671_/Q wb_dat_o[28] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_06024_ _06024_/A1 _06024_/A2 _06024_/A3 _06024_/A4 _06035_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_133_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput322 _11123_/Q wb_dat_o[18] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput344 _11112_/Q wb_dat_o[9] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__10791__A2 _11426_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09933__A1 _10642_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08736__A2 _11276_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07975_ _07975_/A1 _08552_/C _07980_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09714_ _09714_/I _11583_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06926_ _07398_/A1 _07006_/A2 _06871_/Z _06931_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__11139__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09645_ _09645_/I _11561_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06857_ _06855_/Z _06869_/A2 _06857_/B _06858_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07172__A1 _07197_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05808_ _05808_/I _09144_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XTAP_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1017 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1006 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_09576_ _09116_/Z _09597_/A2 _09576_/B _09577_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06788_ _10972_/A1 _05633_/B _08787_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05722__A2 _05805_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10059__A1 _10356_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_08527_ _08527_/I _08528_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05739_ _08799_/A1 _05805_/A2 _05740_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11289__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08458_ _08458_/A1 _08564_/A2 _08563_/A3 _08460_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__06278__A3 _06872_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07409_ _07410_/A2 _11247_/Q _07410_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08389_ _08562_/A1 _08395_/A1 _08656_/B _08390_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_10420_ _10493_/A2 _10427_/A1 _10471_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA_clkbuf_3_7__f_wb_clk_i_I clkbuf_0_wb_clk_i/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07227__A2 _09187_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08975__A2 _11350_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10351_ _11106_/Q _10351_/A2 _11104_/Q _10351_/B2 _10351_/C _10364_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__05789__A2 _09399_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10282_ _10360_/A1 _11434_/Q _10284_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08727__A2 _11273_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05961__A2 _11033_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09152__A2 _09169_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_71 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05713__A2 _09699_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06910__A1 _06843_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08663__A1 _08355_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10470__A1 _10887_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11667_ _11667_/D _11683_/CLK _11667_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11598_ _11598_/D _11686_/RN _06705_/Z _11598_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__08415__A1 split15/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10618_ _10887_/B1 _11430_/Q _10619_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07218__A2 _05924_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10222__A1 _10373_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10222__B2 _11528_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10549_ _10889_/A1 _11404_/Q _10886_/A2 _11396_/Q _10551_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10773__A2 _11561_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09915__A1 _09912_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09391__A2 _09397_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07760_ _07760_/A1 _08054_/A2 _07761_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_2_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10289__A1 _10367_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05952__A2 _11076_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06711_ _06514_/B input84/Z _06713_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09430_ _09430_/I _11492_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07691_ _07691_/I _08294_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XANTENNA__11431__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09270__I _09270_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05704__A2 _08839_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06901__A1 _06902_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06642_ input83/Z _06650_/A1 _06642_/B _06643_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11190__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09361_ _09361_/I _11470_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06573_ _06573_/I _11223_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08312_ _08312_/A1 _08500_/B _08638_/A3 _08502_/A1 _08316_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_09292_ _09292_/I _11448_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05524_ _11070_/Q _11159_/Q _05576_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11581__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08243_ _08545_/A2 _08490_/A3 _08243_/B _08492_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_32_182 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08174_ _08174_/A1 _08174_/A2 _08174_/A3 _08180_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_07125_ _05927_/Z _09125_/I _07126_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10213__A1 _10213_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08957__A2 _08963_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07056_ _07060_/A2 _11145_/Q _07057_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11040__I _11050_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06968__A1 _06837_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06007_ _06007_/A1 _06007_/A2 _06007_/A3 _06007_/A4 _06035_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xoutput185 _06706_/ZN mgmt_gpio_oeb[20] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA_input42_I mgmt_gpio_in[15] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10516__A2 _11620_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput174 _10615_/A2 mgmt_gpio_oeb[10] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput196 _10642_/B1 mgmt_gpio_oeb[30] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__09382__A2 _09397_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07393__A1 _07076_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07958_ _07958_/A1 _08554_/C _07963_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07145__A1 _05927_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07889_ _07889_/I split15/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_28_466 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06909_ _06910_/A2 _11102_/Q _06910_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09628_ _09647_/A2 _11556_/Q _09629_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09559_ _09572_/A2 _11534_/Q _09560_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11181__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08645__A1 _08645_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07448__A2 split13/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11521_ _11521_/D _11686_/RN _06705_/Z _11521_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_11452_ _11452_/D _11686_/RN _06705_/Z _11452_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_10403_ _10440_/A1 _10406_/I _10884_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_11383_ _11383_/D _11686_/RN _06705_/Z _11383_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__10204__B2 _10359_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10204__A1 _11400_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08948__A2 _08963_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09070__A1 _09089_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10334_ _10373_/A1 _11149_/Q _10373_/B1 _11153_/Q _10337_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11304__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07620__A2 _07609_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05631__A1 _06466_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10265_ _10265_/A1 _11329_/Q _10265_/A3 _10266_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_10196_ _11352_/Q _10351_/A2 _11344_/Q _10351_/B2 _10196_/C _10209_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__11454__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07384__A1 _06238_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05934__A2 _11616_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10286__A4 _10286_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08884__A1 _08888_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05698__B2 _09574_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07603__I _08637_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10691__A1 _10691_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10443__B2 _10899_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput10 mask_rev_in[15] input10/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput21 mask_rev_in[25] input21/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput54 mgmt_gpio_in[26] input54/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput43 mgmt_gpio_in[16] input43/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05870__A1 _09750_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput32 mask_rev_in[6] input32/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput98 wb_adr_i[10] input98/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput65 mgmt_gpio_in[36] input65/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput87 spimemio_flash_io0_oeb input87/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput76 porb input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
XANTENNA__09061__A1 _06863_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05622__A1 _08684_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08930_ _08930_/I _11335_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08861_ _08861_/I _11313_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07812_ _07722_/I _08674_/B _07813_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07375__A1 _07081_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08792_ _08793_/A2 _11293_/Q _08793_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07743_ _07743_/I _08494_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07674_ _07674_/A1 _07674_/A2 _07907_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08875__A1 _08888_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06625_ _11526_/Q _06625_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09413_ _09158_/Z _09422_/A2 _09413_/B _09414_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07513__I _07513_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09344_ _09241_/Z _09347_/A2 _09344_/B _09345_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_12_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06556_ _06556_/I _10092_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_33_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06487_ _06487_/I _11064_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09275_ _09297_/A2 _11443_/Q _09276_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05507_ _05507_/I _06451_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08226_ _08226_/A1 _08226_/A2 _08567_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11327__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05861__A1 _05693_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08157_ split8/Z _08159_/I _08158_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10737__A2 _10737_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07108_ _07110_/I _11161_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09052__A1 _06851_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08088_ _08656_/A1 _08659_/A1 _08089_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11477__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07039_ _06843_/Z _07039_/A2 _07039_/B _07040_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10050_ _10050_/I _11646_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output246_I _11188_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11597__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05916__A2 _11400_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10952_ _10952_/A1 _10952_/A2 _11672_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08866__A1 _08888_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10673__A1 _10892_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11154__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10883_ _10883_/A1 _11120_/Q _10885_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10425__A1 _10408_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09291__A1 _09187_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11504_ _11504_/D _11686_/RN _06705_/Z _11504_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__07841__A2 _08677_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11435_ _11435_/D _11686_/RN _06705_/Z _11435_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__09043__A1 _07426_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09594__A2 _09597_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11366_ _11366_/D _11686_/RN _06705_/Z _11366_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__05604__A1 _05616_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11297_ _11297_/D input76/Z _06705_/Z _11297_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_10317_ _10356_/A1 _11135_/Q _10319_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09346__A2 _11466_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10248_ _11457_/Q _10365_/A2 _10365_/B1 _11465_/Q _10251_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05907__A2 _11464_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10179_ _10371_/A1 _11487_/Q _10181_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11393__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08857__A1 _06851_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11145__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10664__A1 _10887_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06410_ _08786_/A1 _08799_/A1 _11292_/Q _06413_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_07390_ _07390_/I _11241_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06341_ _06341_/A1 _06341_/A2 _06350_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09282__A1 _09125_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09060_ _09064_/A2 _11377_/Q _09061_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06272_ _06905_/A1 _11102_/Q _06275_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08011_ _08434_/A1 _08386_/A1 _08390_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07832__A2 _07570_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05843__A1 _06785_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09585__A2 _09597_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09962_ _10374_/A1 _11531_/Q _09967_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09337__A2 _11463_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07508__I _07508_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08913_ _06867_/Z _08913_/A2 _08913_/B _08914_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_962 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_951 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_940 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_09893_ _09893_/I _10030_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_995 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_984 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_973 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input144_I wb_dat_i[22] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08844_ _07431_/Z _08844_/A2 _08844_/B _08845_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08775_ _06855_/Z _08784_/A2 _08775_/B _08776_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11384__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05987_ _05987_/A1 _05987_/A2 _05988_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_150_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07726_ _08339_/A1 _08490_/A3 _07727_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__08848__A1 _07426_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07657_ _07694_/A1 _07657_/A2 _07660_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11136__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07588_ _08669_/A2 _08509_/A1 _08255_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06608_ _06557_/Z _06608_/A2 _06608_/B _06609_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09327_ _09327_/I _11459_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06539_ _11629_/Q _09865_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10422__A4 _10904_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09258_ _09272_/A2 _11438_/Q _09259_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output196_I _10642_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08209_ split7/I _08232_/A2 _08209_/B _08471_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09189_ _09187_/Z _09195_/A2 _09189_/B _09190_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09576__A2 _09597_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11220_ _11220_/D input162/Z _11672_/CLK _11220_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_108_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11151_ _11151_/D _11686_/RN _06705_/Z _11151_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10102_ _11397_/Q _10359_/A2 _11389_/Q _10359_/B2 _10102_/C _10107_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_11082_ _11082_/D input76/Z _06705_/Z _11082_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_68_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09879__A3 _09927_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10033_ _11347_/Q _10351_/A2 _11339_/Q _10351_/B2 _10033_/C _10045_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__06011__B2 _09374_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06011__A1 _11487_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10894__B2 _10894_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11375__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08839__A1 _08839_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06314__A2 input43/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09500__A2 _11515_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10935_ _10935_/A1 _10950_/A2 _10937_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10646__A1 _10919_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10866_ _10866_/A1 _10866_/A2 _10867_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09264__A1 _09272_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11642__CLK _11663_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10797_ _10886_/B2 _11394_/Q _10886_/A2 _11402_/Q _10798_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06078__B2 _08990_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06078__A1 _11382_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09016__A1 _09016_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11418_ _11418_/D input76/Z _06705_/Z _11418_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__08712__I _11050_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11412__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11349_ _11349_/D _11686_/RN _06705_/Z _11349_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_100_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06890_ _06851_/Z _06902_/A2 _06890_/B _06891_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05910_ _11488_/Q _09399_/A1 _11480_/Q _09374_/A1 _05910_/C _05923_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__10334__B1 _10373_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05841_ _05841_/I _05841_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11366__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11427__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08560_ _08560_/I _08561_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11172__CLK input68/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05772_ _09016_/A1 _11370_/Q _05773_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10637__A1 _10914_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07511_ _07511_/I _07516_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08491_ _08491_/I _08493_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07442_ input105/Z _07863_/I _07444_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07373_ _07373_/I _11236_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06324_ _06324_/A1 _11587_/Q _06328_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09112_ _09112_/I _11393_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09255__A1 _09272_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06255_ _08825_/A1 _06238_/Z _11154_/Q _06257_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09043_ _07426_/Z _09064_/A2 _09043_/B _09044_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09007__A1 _06859_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06186_ _06186_/A1 _06186_/A2 _06186_/A3 _06187_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09945_ _06567_/I _09945_/A2 _09947_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09876_ _09876_/I _09898_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06792__A2 _09116_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11515__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09730__A2 _09725_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_781 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_08827_ _08827_/A1 _08827_/A2 _08827_/B _08828_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10876__A1 _10922_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08758_ _08759_/A2 _11283_/Q _08759_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09494__A1 _09241_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10628__A1 _10899_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08297__A2 _07748_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08689_ _07566_/I _07537_/I _08689_/B _08690_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07709_ _08294_/B _08483_/A2 _08430_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11665__CLK _11665_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output209_I _10613_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11109__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10720_ _10720_/A1 _10720_/A2 _10721_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10651_ _10924_/A1 _11326_/Q _10652_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09246__A1 _06867_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10582_ _10891_/A1 _11477_/Q _10583_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10800__A1 _10892_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05807__A1 _05995_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09549__A2 _09015_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11203_ _11203_/D _11686_/RN _06705_/Z _11203_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__06232__A1 _07370_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11134_ _11134_/D _11686_/RN _06705_/Z _11134_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__11195__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11065_ _11065_/D _11065_/RN input68/Z _11065_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__10316__B1 _11119_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09721__A2 _11586_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10016_ _10016_/A1 _10016_/A2 _10017_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10867__B2 _10913_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09485__A1 _09154_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08288__A2 _08623_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10918_ _10918_/A1 _10918_/A2 _10918_/A3 _10918_/A4 _10925_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__06299__A1 _07398_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11520__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10849_ _10895_/A1 _11226_/Q _10852_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06040_ _06040_/A1 _06619_/B _06040_/B _06041_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_172_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11538__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08212__A2 _07722_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07991_ _08386_/A1 _08395_/A1 _08357_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06223__A1 _08825_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09730_ _09121_/I _09725_/Z _09730_/B _09731_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06942_ _10935_/A1 _06957_/A2 _06944_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10858__A1 _10904_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09661_ _09661_/I _11566_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11688__CLK input68/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06873_ _06877_/A2 _11087_/Q _06874_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06526__A2 _11349_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09592_ _09592_/I _11544_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08612_ _08612_/I _08613_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05824_ _09248_/A1 _11442_/Q _05825_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09476__A1 _09116_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08543_ _08294_/C _08543_/A2 _08543_/B _08544_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05755_ _07419_/A2 _08799_/A1 _05756_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input107_I wb_adr_i[19] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10086__A2 _06556_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08474_ _08474_/A1 _08217_/B _08475_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05686_ _05751_/A1 _05776_/A2 _05687_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__11511__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07425_ _07425_/I _11251_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11043__I _11050_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11035__A1 _09116_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07356_ _08825_/A1 _06217_/Z _06871_/Z _07361_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_07287_ _06863_/Z _07290_/A2 _07287_/B _07288_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06307_ _06307_/A1 _06307_/A2 _06307_/B _06308_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11068__CLK input68/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06238_ _06238_/I _06238_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_09026_ _09039_/A2 _11366_/Q _09027_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10794__B1 _11410_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input72_I mgmt_gpio_in[8] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09400__A1 _09422_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06169_ _05584_/I _11265_/Q _06170_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07006__A3 _06871_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11578__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07962__A1 split15/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09928_ _09928_/A1 _09928_/A2 _09929_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10849__A1 _10895_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09859_ _09859_/A1 _09859_/A2 _09860_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06517__A2 _06694_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07190__A2 _05925_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07431__I _09121_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11502__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10703_ _10914_/B1 _11608_/Q _10704_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11683_ _11683_/D input162/Z _11683_/CLK _11683_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__09219__A1 _09220_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10634_ _10504_/I _10634_/A2 _10432_/I _10634_/B2 _10635_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__06491__B _06491_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10565_ _10884_/A1 _11381_/Q _10567_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10496_ _10886_/B2 _11387_/Q _10886_/A2 _11395_/Q _10509_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11569__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06205__A1 _05703_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07953__A1 split21/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06756__A2 _08036_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11117_ _11117_/D _11672_/CLK _11117_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05964__B1 _08990_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11048_ _11050_/I _11695_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xinput8 mask_rev_in[13] input8/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07181__A2 _11177_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05540_ input58/Z _06610_/A3 _05540_/B _05541_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08681__A2 _11016_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11210__CLK _11656_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08190_ _08185_/I _07535_/I _08493_/B _08191_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11017__A1 _08493_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06692__A1 _11306_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07210_ _07240_/A1 _07210_/A2 _07210_/B _07211_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07141_ _11194_/Q _05927_/Z _07151_/B _07141_/C _07142_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_145_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11290__SETN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11360__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07072_ _07072_/I _11149_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xoutput301 _06740_/Z ser_rx VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__10240__A2 _11417_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput334 _11672_/Q wb_dat_o[29] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_126_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput323 _11124_/Q wb_dat_o[19] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_06023_ _11455_/Q _09299_/A1 _11447_/Q _09274_/A1 _06023_/C _06024_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
Xoutput312 _11666_/Q wb_ack_o VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_160_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08197__B2 _08332_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08197__A1 _08434_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09933__A2 _10427_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07944__A1 _08355_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06747__A2 input39/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07974_ split6/Z _07976_/I _08552_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_101_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09697__A1 _09270_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09713_ _09158_/I _09722_/A2 _09713_/B _09714_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06925_ _06925_/I _11106_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09644_ _09241_/Z _09647_/A2 _09644_/B _09645_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06856_ _06869_/A2 _11083_/Q _06857_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05807_ _05995_/A2 _06217_/I _05808_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06787_ _11675_/Q _10972_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09449__A1 _09449_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1029 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1018 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1007 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_09575_ _09597_/A2 _11539_/Q _09576_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08526_ _08686_/A1 _07562_/I _07685_/I _07485_/I _08527_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_23_320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05738_ _05738_/I _08799_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_4
X_08457_ _08562_/A1 _08545_/A2 _08656_/B _08563_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05669_ _05669_/I _05699_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06683__A1 _11305_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07408_ _07408_/I _11246_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08388_ _08453_/A1 _08388_/A2 _08388_/B _08560_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_7_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09621__A1 _09622_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10767__B1 _11489_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07339_ _07340_/A2 _11227_/Q _07340_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output276_I _11075_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06435__A1 _08795_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10350_ _10350_/A1 _10350_/A2 _10351_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09009_ _09013_/A2 _11361_/Q _09010_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10281_ _11402_/Q _10359_/A2 _11394_/Q _10359_/B2 _10281_/C _10286_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__08188__A1 _08490_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07935__A1 split21/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07426__I _09116_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09688__A1 _09158_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11233__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11383__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11666_ _11666_/D input162/Z _11666_/CLK _11666_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_174_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09612__A1 _09622_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11597_ _11597_/D _11686_/RN _06705_/Z _11597_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__08415__A2 _08417_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10617_ _10887_/A2 _11422_/Q _10619_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10222__A2 _11520_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10548_ _10548_/A1 _10548_/A2 _10548_/A3 _10548_/A4 _10548_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
XANTENNA__06426__A1 _08940_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10479_ _10897_/B1 _11459_/Q _10486_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10190__C _10190_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09679__A1 _09121_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10289__A2 _11482_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06710_ _06710_/A1 _06710_/A2 _06710_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07690_ _07690_/A1 _07690_/A2 _07691_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06641_ _11606_/Q input80/Z _06642_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__08103__A1 _08161_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09360_ _09154_/Z _09372_/A2 _09360_/B _09361_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06572_ _06749_/I _08036_/B _06572_/B _06573_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08311_ _08311_/A1 _08411_/A2 _08502_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09291_ _09187_/Z _09297_/A2 _09291_/B _09292_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05523_ _05523_/A1 _06619_/A1 _06446_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_08242_ _08242_/A1 _08490_/A3 _08242_/B _08581_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10997__B1 _08460_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09603__A1 _09622_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08173_ _08487_/I _08621_/A1 _08174_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07124_ _11166_/Q _07127_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06417__A1 _08761_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07090__A1 _07081_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07055_ _05703_/Z _08795_/A1 _06871_/Z _07060_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_06006_ _11583_/Q _09699_/A1 _09674_/A1 _11575_/Q _06007_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11106__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput186 _06048_/B2 mgmt_gpio_oeb[21] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput175 _10615_/B2 mgmt_gpio_oeb[11] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput197 _10642_/A2 mgmt_gpio_oeb[31] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__05928__B1 _07201_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07957_ split6/I _07959_/I _08554_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11256__CLK _11666_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input35_I mask_rev_in[9] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06908_ _06908_/I _11101_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07145__A2 _09241_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07888_ _07685_/I _07888_/A2 _07889_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_55_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09627_ _09627_/I _11555_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05922__C _05922_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06839_ _06839_/A1 _06838_/Z _06869_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_28_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_09558_ _09558_/I _11533_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08509_ _08509_/A1 _08509_/A2 _08509_/B _08509_/C _08596_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_178_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09842__A1 _09187_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11520_ _11520_/D _11686_/RN _06705_/Z _11520_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_09489_ _09489_/I _11511_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10452__A2 _10506_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11451_ _11451_/D _11686_/RN _06705_/Z _11451_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_10402_ _10915_/A1 _10914_/B1 _10883_/A1 _10910_/A1 _10412_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_11382_ _11382_/D input76/Z _06705_/Z _11382_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__10204__A2 _10359_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10333_ _10333_/A1 _10333_/A2 _10333_/A3 _10342_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_10264_ _10264_/A1 _10264_/A2 _10264_/A3 _10264_/A4 _10266_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_120_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10195_ _10350_/A1 _10195_/A2 _10196_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07384__A2 _11033_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_71 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07136__A2 _05927_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05698__A2 _09599_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10691__A2 _10691_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06895__A1 _06902_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10310__I _11101_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09833__A1 _09125_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10443__A2 _10906_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08715__I _11050_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11649_ _11649_/D input76/Z _11665_/CLK _11649_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xinput22 mask_rev_in[26] input22/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput11 mask_rev_in[16] input11/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput55 mgmt_gpio_in[27] input55/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput44 mgmt_gpio_in[17] input44/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11129__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput33 mask_rev_in[7] input33/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput66 mgmt_gpio_in[37] input66/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput88 spimemio_flash_io1_do input88/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09061__A2 _09064_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput77 qspi_enabled input77/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput99 wb_adr_i[11] input99/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11279__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08860_ _06855_/Z _08863_/A2 _08860_/B _08861_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08572__A1 split12/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07811_ _07805_/Z _08511_/C _08331_/B _07811_/A4 _07813_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_08791_ _08791_/A1 _08825_/A2 _11686_/RN _06904_/Z _08793_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_07742_ _08589_/A1 _08490_/A3 _07743_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07127__A2 _07151_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07673_ _07858_/A2 _08095_/A2 _07674_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06624_ _11534_/Q _10634_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09412_ _09422_/A2 _11487_/Q _09413_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06886__A1 _06902_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09343_ _09347_/A2 _11465_/Q _09344_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06555_ _11090_/Q _06556_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__06638__A1 _11614_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06486_ _06479_/C _06486_/A2 _06486_/B _06487_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09274_ _09274_/A1 _09015_/Z _09297_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_05506_ _11070_/Q _11069_/Q _05507_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_33_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08225_ _08618_/B _08225_/A2 _08225_/A3 _08565_/B _08225_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
X_08156_ _08169_/A1 _08156_/A2 _08159_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10198__A1 _10352_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09052__A2 _09064_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07107_ _07110_/I _11160_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_173_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08087_ _08465_/B _08659_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_79_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07038_ _07039_/A2 _11140_/Q _07039_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10370__A1 _10370_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output239_I _06652_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08989_ _08989_/I _11354_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08315__A1 _08332_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10122__A1 _10378_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10951_ _10934_/I _11672_/Q _10952_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06877__A1 _06843_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10882_ _10882_/A1 _10882_/A2 _11664_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08618__A2 _08696_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11503_ _11503_/D _11686_/RN _06705_/Z _11503_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_11_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06055__I _11430_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11434_ _11434_/D input76/Z _06705_/Z _11434_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__09043__A2 _09064_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11421__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11365_ _11365_/D _11686_/RN _06705_/Z _11365_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__05604__A2 _11254_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11296_ _11296_/D input76/Z _06705_/Z _11296_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10316_ _11129_/Q _10355_/A2 _11119_/Q _10355_/B2 _10316_/C _10325_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_429 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11090__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10247_ _10247_/A1 _10247_/A2 _10247_/A3 _10247_/A4 _10247_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__11074__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11571__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10178_ _11511_/Q _10369_/A2 _10369_/B1 _11503_/Q _10181_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10113__A1 _10370_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11089__SETN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06868__A1 _06869_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08857__A2 _08863_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06332__A3 _11033_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10664__A2 _11423_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08609__A2 _08692_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05540__A1 input58/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06674__B _06674_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_06340_ _05703_/Z _08825_/A1 _11246_/Q _06341_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_15_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_06271_ _05833_/I _06204_/I _06905_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08010_ _08010_/I _08434_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XANTENNA__05843__A2 _11077_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09961_ _09961_/I _10374_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__08793__A1 _07426_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08912_ _08913_/A2 _11330_/Q _08913_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_952 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_930 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09892_ _09993_/A1 _09892_/A2 _09893_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_985 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_974 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_963 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10352__A1 _10352_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08843_ _08844_/A2 _11308_/Q _08844_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input137_I wb_dat_i[16] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06020__A2 _11439_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08774_ _08784_/A2 _11288_/Q _08775_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05986_ _09016_/A1 _11367_/Q _05987_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07725_ _07725_/I _08592_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__11046__I _11050_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08848__A2 _08863_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07656_ _07656_/A1 _07656_/A2 _08666_/A2 _08664_/A2 _07659_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__07520__A2 _07522_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07587_ _08669_/A2 _08417_/A2 _07589_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05531__A1 _06610_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06607_ _11089_/Q _11302_/Q _06608_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06538_ _06538_/I _11225_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09326_ _09116_/Z _09347_/A2 _09326_/B _09327_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08355__I _08355_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07284__A1 _06859_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11444__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09257_ _09257_/I _11437_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08208_ _08208_/A1 _08466_/A1 _08211_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06469_ _06470_/A1 _06468_/Z _06469_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_153_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10834__B _10834_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09188_ _09195_/A2 _11416_/Q _09189_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08139_ _08656_/A1 _08609_/B _08140_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07036__A1 _06837_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11594__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07587__A2 _08417_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11150_ _11150_/D _11686_/RN _06705_/Z _11150_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__08784__A1 _06867_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10591__A1 _10914_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10101_ _10101_/A1 _10101_/A2 _10102_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07339__A2 _11227_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11081_ _11081_/D input76/Z _06705_/Z _11081_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_10032_ _10350_/A1 _10032_/A2 _10033_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06011__A2 _09399_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10894__A2 _10894_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05770__A1 _07006_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08839__A2 _08839_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10934_ _10934_/I _10950_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10646__A2 _11366_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10865_ _10911_/A1 _11145_/Q _10866_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_284 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07275__A1 _06847_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06078__A2 _09066_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10796_ _10884_/A1 _11386_/Q _10798_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09264__A2 _11440_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09016__A2 _09015_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11417_ _11417_/D input76/Z _06705_/Z _11417_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_8_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07027__A1 _06217_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08775__A1 _06855_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11348_ _11348_/D _11686_/RN _06705_/Z _11348_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__06513__I _11056_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10582__A1 _10891_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05589__A1 _05616_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06250__A2 _05777_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11279_ _11279_/D _11686_/RN _06705_/Z _11279_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__10334__A1 _10373_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05840_ _06266_/I _10927_/A1 _05840_/B _05841_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11317__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06669__B _11056_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07750__A2 _08614_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07510_ _07510_/A1 _07510_/A2 _07511_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05771_ _05771_/I _09016_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XANTENNA__10637__A2 _11606_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08490_ _08490_/A1 _08656_/B _08490_/A3 _08491_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_62_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07441_ _07441_/A1 _07441_/A2 _07997_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11581__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11467__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07502__A2 split16/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07372_ _07076_/Z _07375_/A2 _07372_/B _07373_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06323_ _06323_/A1 _06323_/A2 _06323_/A3 _06323_/A4 _06329_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_09111_ _06863_/Z _09114_/A2 _09111_/B _09112_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09255__A2 _11437_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11596__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06254_ _09474_/A1 _11508_/Q _06257_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09042_ _09064_/A2 _11371_/Q _09043_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09007__A2 _09013_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06185_ _09775_/A1 _11604_/Q _06186_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07018__A1 _06843_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07519__I split13/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08766__A1 _07431_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09944_ _09945_/A2 _06542_/I _06553_/I _09944_/B1 _09944_/B2 _11644_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_131_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09875_ _09954_/A1 _09958_/A1 _09876_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_793 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_08826_ _08827_/A1 _07114_/C _11303_/Q _08827_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09191__A1 _09195_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08757_ _08757_/I _11282_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05752__A1 _05833_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05969_ _05969_/I _06304_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__09494__A2 _09497_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11549__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07708_ _07720_/I _08495_/B _08483_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08688_ _08688_/A1 _08688_/A2 _08688_/A3 _08700_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_07639_ _07639_/A1 _07639_/A2 _07639_/A3 _08278_/B _07642_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__05504__A1 _06786_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10650_ _10650_/A1 _10650_/A2 _10650_/A3 _10650_/A4 _10650_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_09309_ _09322_/A2 _11454_/Q _09310_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09246__A2 _09246_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10581_ _10894_/B2 _11485_/Q _10583_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05807__A2 _06217_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11202_ _11202_/D _11686_/RN _06705_/Z _11202_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__10564__A1 _10883_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08509__A1 _08509_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06232__A2 _11136_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11133_ _11133_/D _11686_/RN _06705_/Z _11133_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_11064_ _11064_/D _11064_/RN input68/Z _11064_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__09182__A1 _09154_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10316__B2 _10355_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10015_ _10361_/A1 _11419_/Q _10016_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07732__A2 _08513_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10867__A2 _10913_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05743__A1 _07398_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09485__A2 _09497_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10917_ _10917_/A1 _10917_/A2 _10917_/A3 _10917_/A4 _10918_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__06299__A2 _07006_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10848_ _11248_/Q _10894_/A2 _11244_/Q _10894_/B2 _10848_/C _10852_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_10779_ _10779_/A1 _10779_/A2 _10779_/A3 _10779_/A4 _10780_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__10252__B1 _10369_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10555__A1 _10887_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07990_ _07990_/I _08395_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_4_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06941_ _06941_/I _06957_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09660_ _09154_/I _09672_/A2 _09660_/B _09661_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05982__A1 _06839_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09173__A1 _09116_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08611_ _08651_/A3 _08651_/A2 _08615_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_94_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07723__A2 split13/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06872_ _08839_/A1 _06872_/A2 _06871_/Z _06877_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__08920__A1 _07431_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09591_ _09187_/Z _09597_/A2 _09591_/B _09592_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05823_ _05823_/I _09248_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
X_08542_ _07691_/I _07492_/I _08543_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05754_ _06204_/I _05738_/I _08761_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__09476__A2 _09497_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08473_ _08473_/A1 _08576_/A1 _08617_/A2 _08695_/I _08480_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__10491__B1 _10914_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07424_ _07081_/Z _07424_/A2 _07424_/B _07425_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05685_ _05685_/I _05751_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07355_ _07355_/I _11231_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07239__A1 _07240_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07286_ _07290_/A2 _11203_/Q _07287_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08987__A1 _08988_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06306_ _05584_/I _11264_/Q _06307_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06237_ _09349_/A1 _11468_/Q _06241_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10794__A1 _11418_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10794__B2 _10889_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09025_ _09025_/I _11365_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input65_I mgmt_gpio_in[36] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06168_ _11264_/Q _05969_/I _06168_/B _06619_/B _06170_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__10546__A1 _10919_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06099_ _06099_/A1 _06099_/A2 _06099_/A3 _06099_/A4 _10945_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__06214__A2 _11227_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09927_ _10642_/A1 _09927_/A2 _10425_/A2 _09928_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__11632__CLK _11666_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05973__A1 _05584_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09858_ _09866_/A2 _09864_/A1 _09868_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09789_ _09158_/I _09798_/A2 _09789_/B _09790_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08809_ _08809_/I _11297_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05725__A1 _07006_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10702_ _10914_/A1 _11600_/Q _10704_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11682_ _11682_/D input162/Z _06687_/A2 _11682_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__11411__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09219__A2 _11426_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10633_ _10904_/A1 _11550_/Q _10636_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08978__A1 _08988_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10564_ _10883_/A1 _11373_/Q _10567_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10495_ _10410_/I _10417_/I _10886_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__11162__CLK input68/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06205__A2 _08825_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11116_ _11116_/D _11672_/CLK _11116_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09155__A1 _09169_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11047_ _11050_/I _11694_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xinput9 mask_rev_in[14] input9/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08718__I _11050_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06141__A1 _06141_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06238__I _06238_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06692__A2 _06692_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07140_ _05927_/Z _09187_/I _07141_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11505__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08969__A1 _08988_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10776__A1 _10899_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11257__RN input162/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07071_ _06837_/Z _07074_/A2 _07071_/B _07072_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06444__A2 _06446_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10528__A1 _11444_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06022_ _06022_/A1 _06022_/A2 _06023_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput302 _06577_/A1 serial_clock VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput313 _11208_/Q wb_dat_o[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput324 _11209_/Q wb_dat_o[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput335 _11210_/Q wb_dat_o[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__09394__A1 _09241_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11655__CLK _11665_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06701__I _06701_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07973_ _08015_/A1 _07973_/A2 _07976_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09712_ _09722_/A2 _11583_/Q _09713_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09146__A1 _09116_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05955__A1 _09016_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09697__A2 _09697_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06924_ _06843_/Z _06924_/A2 _06924_/B _06925_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06855_ _09158_/I _06855_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_09643_ _09647_/A2 _11561_/Q _09644_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09574_ _09574_/A1 _09015_/I _09597_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_05806_ _05806_/I _09171_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XANTENNA__09449__A2 _09015_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1019 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1008 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_06786_ _06786_/A1 _05616_/C _08787_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08525_ _08525_/I _11256_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05737_ _06192_/I _05738_/I _06396_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__06132__A1 _11581_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08456_ _08519_/A1 _08393_/B _08456_/B _08564_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06132__B2 _09674_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05668_ _05668_/I _05940_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_50_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11496__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08387_ _08387_/I _08388_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06683__A2 input96/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07407_ _07076_/Z _07410_/A2 _07407_/B _07408_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05599_ _05644_/A1 _05674_/A2 _05600_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07338_ _07338_/I _11226_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11185__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10767__B2 _10894_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08424__A3 _08540_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11248__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07632__A1 _07640_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07269_ _07076_/Z _07290_/A2 _07269_/B _07270_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06435__A2 _07006_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05643__B1 _05925_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10519__A1 _10914_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output171_I _06746_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output269_I _11271_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10280_ _10280_/A1 _10280_/A2 _10281_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09008_ _09008_/I _11360_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09385__A1 _09154_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06199__A1 _05703_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05946__A1 _06266_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09688__A2 _09697_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11528__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_71 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06123__B2 _08990_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06123__A1 _11349_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10455__B1 _10920_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11487__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06674__A2 input1/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11665_ _11665_/D input76/Z _11665_/CLK _11665_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_41_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_10616_ _10616_/I _10619_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11365__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11596_ _11596_/D _11686_/RN _06705_/Z _11596_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__11239__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11678__CLK _06687_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10547_ _10547_/A1 _10547_/A2 _10547_/A3 _10547_/A4 _10548_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_10478_ _10478_/A1 _10427_/B _10897_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__08179__A2 _08490_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09376__A1 _09116_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05937__A1 _09750_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09679__A2 _09697_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11058__CLK input68/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06640_ input80/Z _06650_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06362__A1 _09171_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06571_ _11218_/Q _06572_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_17_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08310_ _07605_/I _08310_/A2 _08638_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09290_ _09297_/A2 _11448_/Q _09291_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05522_ _11161_/Q _06619_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
X_08241_ _08241_/A1 _08241_/A2 _08488_/A1 _08244_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__11478__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10997__A1 _08431_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10749__A1 _10914_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08172_ _08490_/A1 _08614_/A2 _08656_/B _08621_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__07614__A1 _07614_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07123_ _07123_/I _11165_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06417__A2 _11284_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_429 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07054_ _07054_/I _11144_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06005_ _09624_/A1 _11559_/Q _06007_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11650__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput176 _06730_/ZN mgmt_gpio_oeb[12] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__07917__A2 _08095_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input167_I wb_stb_i VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput187 _10148_/B2 mgmt_gpio_oeb[22] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput198 _06622_/ZN mgmt_gpio_oeb[32] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__11049__I _11050_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11402__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09119__A1 _09116_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10921__A1 _10921_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07956_ _07964_/A1 _08015_/A2 _07959_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input28_I mask_rev_in[31] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06907_ _06837_/Z _06910_/A2 _06907_/B _06908_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07887_ _07887_/A1 _08549_/C _07903_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06838_ _09015_/I _06838_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09626_ _09116_/I _09647_/A2 _09626_/B _09627_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09557_ _09125_/Z _09572_/A2 _09557_/B _09558_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06769_ _07110_/I _11060_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09488_ _09158_/Z _09497_/A2 _09488_/B _09489_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08508_ _08508_/A1 _08690_/A2 _08508_/A3 _08640_/A2 _08510_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_08439_ _08439_/A1 _08439_/A2 _08550_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08645__A3 _11016_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10988__A1 _11016_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05864__B1 _11545_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06656__A2 _11174_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11450_ _11450_/D _11686_/RN _06705_/Z _11450_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_7_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10401_ _10401_/I _10910_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_109_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11381_ _11381_/D input76/Z _06705_/Z _11381_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_10332_ _10370_/A1 _11248_/Q _10333_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11641__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10263_ _10263_/A1 _10263_/A2 _10263_/A3 _10264_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_2_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11200__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10194_ _10194_/A1 _10194_/A2 _11650_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07384__A3 _06838_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11350__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10140__A2 _11422_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07121__B _07151_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11648_ _11648_/D input76/Z _11658_/CLK _11648_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xinput12 mask_rev_in[17] input12/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05855__B1 _05995_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09597__A1 _09270_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput45 mgmt_gpio_in[18] input45/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11579_ _11579_/D _11686_/RN _06705_/Z _11579_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
Xinput34 mask_rev_in[8] input34/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput23 mask_rev_in[27] input23/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput56 mgmt_gpio_in[28] input56/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput89 spimemio_flash_io1_oeb input89/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput78 ser_tx input78/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput67 mgmt_gpio_in[3] input67/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10903__A1 _10903_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07810_ _08592_/A2 _08332_/B _07811_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08790_ _08790_/I _11292_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07741_ _07738_/Z _08302_/A2 _08590_/A1 _07744_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_96_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09521__A1 _09522_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07672_ _07672_/A1 _07890_/B _08438_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06335__A1 _09599_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09411_ _09411_/I _11486_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06623_ _11566_/Q _10642_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08088__A1 _08656_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09342_ _09342_/I _11464_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06554_ _09859_/A2 _09865_/A2 _11630_/Q _06574_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05505_ _05505_/I _11701_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06638__A2 input77/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06485_ _06489_/A1 _11064_/Q _06491_/B _06486_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09273_ _09273_/I _11442_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08224_ _08134_/I _07722_/I _08224_/B _08565_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05846__B1 _08803_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09588__A1 _09158_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08155_ _08155_/A1 _08155_/A2 _08155_/A3 _08650_/A2 _08158_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__10737__A4 _10737_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07106_ _07110_/I _07106_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11623__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08086_ _08106_/A1 _08156_/A2 _08465_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11223__CLK _11683_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08260__A1 _08400_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06810__A2 _05633_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07037_ _07037_/I _11139_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09760__A1 _09773_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06023__B1 _11447_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08988_ _06867_/Z _08988_/A2 _08988_/B _08989_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11373__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07939_ _07939_/I _07964_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09512__A1 _09522_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08315__A2 _08417_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06326__A1 _07391_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10950_ _10950_/A1 _10950_/A2 _10952_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09609_ _09622_/A2 _11550_/Q _09610_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10881_ _10881_/A1 _11664_/Q _10882_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07720__I _07720_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11502_ _11502_/D _11686_/RN _06705_/Z _11502_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__09579__A1 _09121_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_11433_ _11433_/D input76/Z _06705_/Z _11433_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_11364_ _11364_/D _11686_/RN _06705_/Z _11364_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_11295_ _11295_/D _11686_/RN _06705_/Z _11295_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10315_ _10315_/A1 _10315_/A2 _10316_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_10246_ _11449_/Q _10363_/A2 _11441_/Q _10363_/B2 _10246_/C _10247_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__08554__A2 _08692_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_71 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09751__A1 _09773_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10897__B1 _10897_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10177_ _10177_/A1 _10177_/A2 _10177_/A3 _10189_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_19_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06317__A1 _08846_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07116__B _07151_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09503__A1 _09522_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06868__A2 _11086_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05540__A2 _06610_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1180 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07817__A1 _07570_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10821__B1 _11586_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08490__A1 _08490_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06270_ _08890_/A1 _11324_/Q _06275_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11246__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08242__A1 _08242_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09990__A1 _10367_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09960_ _10042_/A2 _09960_/A2 _09899_/I _09961_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_170_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08911_ _08911_/I _11329_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11396__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09742__A1 _09187_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_953 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_942 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_931 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08545__A2 _08545_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09891_ _09891_/A1 _10023_/A1 _09927_/A2 _09993_/A1 _09902_/I _11634_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XTAP_986 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_975 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_964 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_08842_ _08842_/I _11307_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_997 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_08773_ _08773_/I _11287_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05985_ _09041_/A1 _11375_/Q _05987_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07724_ _07793_/A1 _08054_/A2 _07725_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07655_ _08283_/B _08509_/A1 _08664_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10104__A2 _11421_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07520__A3 _08095_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06606_ _10433_/A1 _09934_/I _06608_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07586_ _07586_/I _08417_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_3
X_09325_ _09347_/A2 _11459_/Q _09326_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06537_ _06749_/I _11028_/A2 _06537_/B _06538_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07284__A2 _07290_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06468_ _06491_/B _11067_/Q _06468_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA_input95_I uart_enabled VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09256_ _09125_/Z _09272_/A2 _09256_/B _09257_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08207_ _08079_/I _08199_/I _08465_/B _08466_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09187_ _09187_/I _09187_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__10834__C _10880_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06399_ _11206_/Q _10343_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08138_ _08138_/A1 _08196_/B _08476_/C _08138_/A4 _08141_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_08069_ _08069_/I _08106_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_134_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09981__A1 _09972_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10406__I _10406_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08784__A2 _08784_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11080_ _11080_/D _11686_/RN _06705_/Z _11080_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA_output251_I _06710_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10100_ _10357_/A1 _11413_/Q _10101_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09733__A1 _09125_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10031_ _11331_/Q _10032_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10343__A2 _10382_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11119__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05770__A2 _08719_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08839__A3 _06838_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10933_ _11222_/D input162/Z _10934_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_10864_ _10910_/A1 _11261_/Q _10866_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_10795_ _10883_/A1 _11378_/Q _10798_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_285 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08472__A1 _08575_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07275__A2 _07290_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_71 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_11416_ _11416_/D input76/Z _06705_/Z _11416_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__07027__A2 _11033_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08775__A2 _08784_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11347_ _11347_/D _11686_/RN _06705_/Z _11347_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__10582__A2 _11477_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06786__A1 _06786_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11278_ _11278_/D _11686_/RN _06705_/Z _11278_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10229_ _10092_/Z _11650_/Q _10229_/B _10880_/C _10231_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05770_ _07006_/A2 _08719_/A2 _05771_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10051__I _11324_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10098__A1 _11381_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_393 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10098__B2 _10355_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07440_ _07440_/A1 _07440_/A2 _07441_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07371_ _07375_/A2 _11236_/Q _07372_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06322_ _07398_/A1 _08825_/A2 _11234_/Q _06323_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09110_ _09114_/A2 _11393_/Q _09111_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09041_ _09041_/A1 _09015_/Z _09064_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_06253_ _09499_/A1 _11516_/Q _06257_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08215__A1 _08616_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06184_ _07398_/A1 _08825_/A2 _11235_/Q _06186_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08766__A2 _08784_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10022__A1 _10356_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09943_ _09943_/I _11643_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09715__A1 _09722_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09874_ _11632_/Q _09954_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_750 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07535__I _07535_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_08825_ _08825_/A1 _08825_/A2 _08827_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09191__A2 _11417_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05968_ _05968_/A1 _05968_/A2 _10950_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input10_I mask_rev_in[15] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08756_ _06855_/Z _08759_/A2 _08756_/B _08757_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05752__A2 _05700_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07707_ _07836_/A1 _07751_/A1 _07720_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05899_ _05693_/Z _11528_/Q _05901_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08687_ _08687_/A1 _08687_/A2 _08687_/A3 _08687_/A4 _08688_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__11411__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07638_ _08417_/B _08509_/A1 _08278_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07569_ _07579_/A1 _07989_/A2 _07570_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09308_ _09308_/I _11453_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11073__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11561__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10580_ _10894_/A2 _11493_/Q _10583_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output299_I _11293_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10261__A1 _10374_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09239_ _09187_/Z _09246_/A2 _09239_/B _09240_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08315__B _08315_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11088__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11201_ _11201_/D _11686_/RN _06705_/Z _11201_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_134_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11132_ _11132_/D _11686_/RN _06705_/Z _11132_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__06232__A3 _06217_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09706__A1 _09722_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11063_ _11063_/D _11063_/RN input68/Z _11063_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__10316__A2 _10355_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10014_ _10014_/A1 _09876_/I _10361_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09182__A2 _09195_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05743__A2 _08799_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11091__CLK _11656_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10916_ _10916_/A1 _11231_/Q _10917_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10847_ _10847_/A1 _10847_/A2 _10848_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10778_ _11529_/Q _10902_/A2 _10902_/B2 _11521_/Q _10779_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07799__A3 _08639_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10252__B2 _11505_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10004__A1 _09996_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06223__A3 _06217_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06940_ _11218_/Q input162/Z _06941_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA_input2_I debug_oeb VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10307__A2 _10880_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09173__A2 _09195_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06871_ _09015_/I _06871_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_08610_ _08610_/A1 _08140_/I _08610_/A3 _08610_/A4 _08651_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__07184__A1 _05925_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05822_ _06217_/I _08799_/A2 _05823_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11434__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08920__A2 _08938_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09590_ _09597_/A2 _11544_/Q _09591_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06931__A1 _06843_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08541_ _08541_/A1 _08541_/A2 _08541_/A3 _08631_/A2 _08544_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_05753_ _05753_/A1 _05753_/A2 _06204_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_82_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11584__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08472_ _08575_/B _08462_/I _08472_/B _08472_/C _08695_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08684__A1 _08684_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05684_ _05802_/A2 _05684_/A2 _05685_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__10491__A1 _10914_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07423_ _07424_/A2 _11251_/Q _07424_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05498__A1 _06786_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07354_ _07081_/Z _07354_/A2 _07354_/B _07355_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08436__A1 _08449_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07239__A2 _11188_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07285_ _07285_/I _11202_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06305_ _05969_/I _11263_/Q _06619_/B _06307_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06236_ _09324_/A1 _11460_/Q _06241_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10794__A2 _10888_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09024_ _06847_/Z _09039_/A2 _09024_/B _09025_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08739__A2 _11277_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06167_ _10942_/A1 _05969_/I _06168_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06098_ _06098_/A1 _06098_/A2 _06098_/A3 _06099_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_input58_I mgmt_gpio_in[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09926_ _09936_/A2 _11640_/Q _09928_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09857_ _09857_/A1 _09945_/A2 _09864_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_09788_ _09798_/A2 _11607_/Q _09789_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08808_ _06851_/Z _08820_/A2 _08808_/B _08809_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05725__A2 _06872_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output214_I _11177_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08739_ _08740_/A2 _11277_/Q _08740_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10701_ _10701_/A1 _10701_/A2 _11660_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11681_ _11681_/D input162/Z _06687_/A2 _11681_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10632_ _10903_/A1 _11558_/Q _10636_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10234__B2 _10351_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10563_ _10886_/B2 _11389_/Q _10567_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11307__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05661__A1 _05660_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07650__A2 _08686_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09927__A1 _10642_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10494_ _10494_/I _10886_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_30_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11580__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11457__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11115_ _11115_/D _11672_/CLK _11115_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11046_ _11050_/I _11693_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05964__A2 _05723_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07166__A1 _07197_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11595__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10473__A1 _10406_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06141__A2 _06141_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11533__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09091__A1 _09091_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10776__A2 _11505_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07070_ _07074_/A2 _11149_/Q _07071_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05652__A1 _05927_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07641__A2 _08686_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06021_ _09222_/A1 _11431_/Q _06022_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10528__A2 _10895_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput325 _11125_/Q wb_dat_o[20] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput314 _11113_/Q wb_dat_o[10] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput303 _05947_/Z serial_data_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__09394__A2 _09397_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput336 _11673_/Q wb_dat_o[30] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__11548__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09711_ _09711_/I _11582_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07972_ _08438_/C _08015_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09146__A2 _09169_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08354__B1 split15/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06923_ _06924_/A2 _11106_/Q _06924_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09642_ _09642_/I _11560_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06854_ _06854_/I _11082_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11193__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09573_ _09573_/I _11538_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06785_ _06785_/A1 _09015_/I _06835_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_05805_ _06217_/I _05805_/A2 _05806_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1009 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_08524_ _08524_/A1 _07844_/B _08524_/B _08525_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05736_ _05776_/A1 _05751_/A2 _05738_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA_input112_I wb_adr_i[23] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08455_ _08455_/A1 _08455_/A2 _08613_/A1 _08458_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__06132__A2 _09699_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05667_ _06324_/A1 _11594_/Q _05673_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10464__A1 _10894_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08386_ _08386_/A1 _08632_/A2 _08387_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07406_ _07410_/A2 _11246_/Q _07407_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05598_ _05598_/I _05674_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10216__A1 _10370_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07337_ _07076_/Z _07340_/A2 _07337_/B _07338_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09082__A1 _09089_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10767__A2 _10894_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05643__A1 input71/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07268_ _07290_/A2 _11197_/Q _07269_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07199_ _05638_/I _06701_/I _08865_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_09007_ _06859_/Z _09013_/A2 _09007_/B _09008_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06219_ _06219_/A1 _06219_/A2 _06219_/A3 _06219_/A4 _06235_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__08188__A3 _08242_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09385__A2 _09397_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06199__A2 _08795_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07396__A1 _07081_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09909_ _11637_/Q _11636_/Q _09912_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__11184__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_split13_I split13/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06123__A2 _05723_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07320__A1 _07310_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10455__A1 _10920_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11664_ _11664_/D input76/Z _11665_/CLK _11664_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XPHY_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05882__A1 _09474_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10615_ _10507_/I _10615_/A2 _10445_/I _10615_/B2 _10616_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_167_360 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11595_ _11595_/D _11686_/RN _06705_/Z _11595_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__09073__A1 _09089_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08820__A1 _07431_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10546_ _10919_/A1 _11364_/Q _10547_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10477_ _10477_/A1 _10477_/A2 _10477_/A3 _10477_/A4 _10487_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__09376__A2 _09397_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08584__B1 _08460_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10930__A2 _11666_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11029_ _11029_/A1 _08672_/B _11030_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08887__A1 _08888_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11175__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10694__A1 _10922_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06362__A2 _11411_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08639__A1 _07566_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06570_ _08460_/B _08036_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_24_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09300__A2 _11451_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10446__A1 _10904_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05521_ _06444_/A1 _11700_/Q _11699_/Q _11698_/Q _05529_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__06114__A2 _06114_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07311__A1 _10935_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08240_ _07837_/I _07492_/I _08240_/B _08488_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05873__A1 _05660_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08171_ _08490_/A1 _08181_/A3 _08580_/A2 _08487_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11622__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07122_ _07122_/A1 _07151_/B _07122_/B _07123_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09064__A1 _06867_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07614__A2 split16/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08811__A1 _06847_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07053_ _06843_/Z _07053_/A2 _07053_/B _07054_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06004_ _09649_/A1 _11567_/Q _06007_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput177 _06056_/B2 mgmt_gpio_oeb[13] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput199 _06738_/ZN mgmt_gpio_oeb[33] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput188 _10148_/A1 mgmt_gpio_oeb[23] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__05928__A2 _05927_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07955_ _07955_/A1 _07955_/A2 _07955_/A3 _08373_/B _07958_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_87_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09119__A2 _09142_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08878__A1 _08888_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06906_ _06910_/A2 _11101_/Q _06907_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07886_ _08359_/B _07886_/A2 _08549_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10685__A1 _10903_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09625_ _09647_/A2 _11555_/Q _09626_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11166__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06837_ _09116_/I _06837_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_09556_ _09572_/A2 _11533_/Q _09557_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11152__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06768_ _07110_/I _11059_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09487_ _09497_/A2 _11511_/Q _09488_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08507_ _07572_/I _07725_/I _08507_/B _08507_/C _08640_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05719_ _05719_/I _07006_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_4
X_06699_ _06266_/I _09944_/B2 _06699_/B _06700_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07302__A1 _08839_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08438_ split6/Z split8/Z _08438_/B _08438_/C _08439_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_23_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08369_ split8/I _08557_/B _08369_/B _08558_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05864__B2 _09574_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09055__A1 _06855_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10400_ _10400_/A1 _10503_/A2 _10401_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11380_ _11380_/D _11686_/RN _06705_/Z _11380_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_10331_ _10371_/A1 _11244_/Q _10333_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06622__I _11582_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10262_ _10375_/A1 _11545_/Q _10263_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10373__B1 _10373_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10193_ _10881_/A1 _11650_/Q _10194_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05919__A2 _11440_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10676__A1 _10895_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11157__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08869__A1 _08888_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10691__A4 _10691_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09294__A1 _09241_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11645__CLK _11658_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10979__A2 _10966_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07844__A2 _11016_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11647_ _11647_/D input76/Z _11663_/CLK _11647_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xinput13 mask_rev_in[18] input13/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05855__B2 _08799_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09046__A1 _07431_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09597__A2 _09597_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput46 mgmt_gpio_in[19] input46/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11578_ _11578_/D _11686_/RN _06705_/Z _11578_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xinput35 mask_rev_in[9] input35/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput24 mask_rev_in[28] input24/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput57 mgmt_gpio_in[29] input57/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10600__A1 _10903_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10529_ _10897_/B1 _11460_/Q _10532_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05607__A1 _06466_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput79 spi_csb input79/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput68 mgmt_gpio_in[4] input68/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__09349__A2 _09015_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06032__A1 _06324_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07740_ _08600_/A2 _08339_/A1 _08590_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10116__B1 _10373_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11175__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07671_ _07938_/A1 _07938_/A3 _07890_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11148__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09521__A2 _11522_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10667__B2 _10889_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09410_ _09154_/Z _09422_/A2 _09410_/B _09411_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06622_ _11582_/Q _06622_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_18_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09341_ _09187_/Z _09347_/A2 _09341_/B _09342_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09285__A1 _09154_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06553_ _06553_/I _09859_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05504_ _06786_/A1 _05504_/A2 _05504_/B _05505_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_52_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06484_ _06497_/A1 _06484_/A2 _06489_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09272_ _09270_/Z _09272_/A2 _09272_/B _09273_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05846__A1 _11329_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06707__I _11057_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08223_ _08476_/B _08225_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_20_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05846__B2 _05841_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11320__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09588__A2 _09597_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08154_ _08434_/A1 _08567_/A1 _08650_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08085_ _08085_/I _08156_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07105_ _07105_/I _11158_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_173_182 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07036_ _06837_/Z _07039_/A2 _07036_/B _07037_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06271__A1 _05833_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input40_I mgmt_gpio_in[13] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11518__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06574__A2 _06556_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08987_ _08988_/A2 _11354_/Q _08988_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07938_ _07938_/A1 _07938_/A2 _07938_/A3 _07939_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_113_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11364__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07869_ _07869_/A1 _07470_/I _07871_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09512__A2 _11519_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11668__CLK _11672_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11139__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09608_ _09608_/I _11549_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_16_439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10880_ _10092_/Z _11663_/Q _10880_/B _10880_/C _10882_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09539_ _09539_/I _11527_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11379__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09276__A1 _09116_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11501_ _11501_/D _11686_/RN _06705_/Z _11501_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_132_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11311__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10830__A1 _10919_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09579__A2 _09597_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11432_ _11432_/D input76/Z _06705_/Z _11432_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_11363_ _11363_/D _11686_/RN _06705_/Z _11363_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_11294_ _11294_/D _11686_/RN _06705_/Z _11294_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10314_ _10352_/A1 _11107_/Q _10315_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11198__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_10245_ _10245_/A1 _10245_/A2 _10246_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10176_ _10366_/A1 _11471_/Q _10177_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11378__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07762__A1 _08696_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_285 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06317__A2 input61/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10649__A1 _10922_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11550__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09267__A1 _09272_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07817__A2 _08495_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10821__B2 _10913_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08490__A2 _08656_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05828__A1 _05828_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11302__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08242__A2 _08490_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06253__A1 _09499_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_910 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_09890_ _11634_/Q _09993_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08910_ _06863_/Z _08913_/A2 _08910_/B _08911_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09742__A2 _09725_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06005__A1 _09624_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_943 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_932 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11369__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10888__A1 _10888_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08841_ _07426_/Z _08844_/A2 _08841_/B _08842_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07753__A1 _08589_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_987 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_965 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_954 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_998 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_05984_ _05984_/A1 _05984_/A2 _05984_/A3 _05984_/A4 _05999_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_08772_ _06851_/Z _08784_/A2 _08772_/B _08773_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07723_ _07675_/B split13/I _08054_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07654_ _08283_/B _08417_/A2 _08666_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06605_ _06605_/I _11160_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07585_ _08339_/A1 _08345_/A2 _07586_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__09258__A1 _09272_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09324_ _09324_/A1 _09015_/Z _09347_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_06536_ _11220_/Q _06537_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_80_397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10812__A1 _10903_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05819__A1 _06217_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06467_ _06497_/A1 _11066_/Q _06478_/B _06470_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09255_ _09272_/A2 _11437_/Q _09256_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08206_ _08660_/A3 _08464_/A1 _08206_/A3 _08206_/A4 _08208_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA_input88_I spimemio_flash_io1_do VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06398_ input20/Z _06398_/A2 _06398_/B _06439_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09186_ _09186_/I _11415_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08137_ split7/Z _08222_/B _08138_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08068_ _08068_/A1 _08114_/A1 _08069_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06244__A1 _07398_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10040__A2 _10040_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11340__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06795__A2 _05633_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07019_ _07019_/I _11134_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10030_ _10030_/A1 _10030_/A2 _10265_/A3 _10350_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XANTENNA__11490__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09733__A2 _09725_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output244_I _11186_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09497__A1 _09270_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10932_ _10932_/I _11666_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10500__B1 _10902_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10863_ _10863_/A1 _10863_/A2 _10863_/A3 _10863_/A4 _10872_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__09249__A1 _09272_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_10794_ _11418_/Q _10888_/A1 _11410_/Q _10889_/A1 _10794_/C _10798_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XPHY_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_253 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10803__A1 _10895_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06483__B2 _05515_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09421__A1 _09422_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08224__A2 _07722_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11415_ _11415_/D input76/Z _06705_/Z _11415_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__07027__A3 _06871_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11599__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11346_ _11346_/D _11686_/RN _06705_/Z _11346_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__06786__A2 _05616_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11277_ _11277_/D _11686_/RN _06705_/Z _11277_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10228_ _10209_/Z _10092_/Z _10228_/A3 _10228_/A4 _10229_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_10159_ _10350_/A1 _10159_/A2 _10160_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_181_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09488__A1 _09158_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10098__A2 _10355_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08160__A1 split7/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06171__B1 _05925_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11213__CLK _11656_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07370_ _07370_/A1 _06238_/Z _06871_/Z _07375_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_06321_ _07349_/A1 _11230_/Q _06323_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09660__A1 _09154_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06252_ _06252_/A1 _06252_/A2 _06252_/A3 _06252_/A4 _06258_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__06474__A1 _05515_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09040_ _09040_/I _11370_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11363__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09412__A1 _09422_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08215__A2 _07722_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06183_ _09800_/A1 _11612_/Q _07349_/A1 _11231_/Q _06186_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_171_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09963__A2 _09878_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06226__A1 _09171_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10022__A2 _11403_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09942_ _09942_/A1 _09944_/B1 _09942_/B _09943_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07726__A1 _08339_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09873_ _09873_/I _11631_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_784 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input142_I wb_dat_i[20] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_762 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_08824_ _08824_/I _11302_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08755_ _08759_/A2 _11282_/Q _08756_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09479__A1 _09121_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07706_ _08543_/B _07710_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05967_ _05967_/A1 _05967_/A2 _05967_/A3 _05967_/A4 _05968_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_08686_ _08686_/A1 _08686_/A2 _08686_/B _08687_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05898_ _05898_/A1 _05898_/A2 _11269_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11514__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07637_ _08417_/B _08417_/A2 _07639_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07568_ _07487_/I input119/Z _07989_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11038__A1 _09121_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09307_ _09125_/Z _09322_/A2 _09307_/B _09308_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06519_ _06519_/A1 _06519_/A2 _06520_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07499_ _07513_/I split13/I _07857_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__09651__A1 _09116_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10797__B1 _10886_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output194_I _10146_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09238_ _09246_/A2 _11432_/Q _09239_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09403__A1 _09422_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10417__I _10417_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09169_ _06867_/Z _09169_/A2 _09169_/B _09170_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10549__B1 _10886_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11200_ _11200_/D _11686_/RN _06705_/Z _11200_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_119_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11131_ _11131_/D _11686_/RN _06705_/Z _11131_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__09706__A2 _11581_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11062_ _11062_/D _11062_/RN input68/Z _11062_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_95_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10013_ _10360_/A1 _11427_/Q _10016_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10721__B1 _11488_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11236__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06940__A2 input162/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11505__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10915_ _10915_/A1 _11235_/Q _10917_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11029__A1 _11029_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10846_ _10892_/A1 _11236_/Q _10847_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11386__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10777_ _10900_/A1 _11513_/Q _10779_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10252__A2 _10369_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10004__A2 _09876_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06208__A1 _09549_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11329_ _11329_/D input76/Z _06705_/Z _11329_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__07708__A1 _07720_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06870_ _06870_/I _11086_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08381__A1 _08656_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07184__A2 _09187_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05821_ _09222_/A1 _11434_/Q _05825_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08540_ _08540_/A1 _08540_/A2 _08540_/A3 _08540_/A4 _08631_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_05752_ _05833_/I _05700_/I _08890_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_05683_ _05683_/A1 _05683_/A2 _05678_/Z _05682_/Z _05714_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_08471_ _08098_/I _08462_/I _08471_/B _08471_/C _08617_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_23_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08684__A2 _07297_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07422_ _07422_/I _11250_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09881__A1 _09898_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06695__A1 _06266_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07353_ _07354_/A2 _11231_/Q _07354_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07284_ _06859_/Z _07290_/A2 _07284_/B _07285_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06715__I _06715_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10243__A2 _11433_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06304_ _10938_/A1 _06304_/A2 _06307_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09023_ _09039_/A2 _11365_/Q _09024_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06235_ _06235_/A1 _06235_/A2 _06235_/A3 _06235_/A4 _06259_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__11109__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06166_ _06166_/A1 _06166_/A2 _06166_/A3 _10942_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_06097_ input29/Z _06396_/A1 input23/Z _06398_/A2 _06097_/C _06098_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__11259__CLK _06687_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09925_ _09925_/I _11639_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09856_ _09856_/I _11627_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07175__A2 _05925_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08807_ _08820_/A2 _11297_/Q _08808_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_09787_ _09787_/I _11606_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06999_ _08795_/A1 _07006_/A2 _06871_/Z _07004_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__08124__A1 split8/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08738_ _08738_/I _11276_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08669_ _08355_/I _08669_/A2 _08670_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output207_I _10137_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09872__A1 _09902_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10700_ _10881_/A1 _11660_/Q _10701_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_11680_ _11680_/D input162/Z _06687_/A2 _11680_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__10482__A2 _10427_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08326__B _08639_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09624__A1 _09624_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10631_ _11526_/Q _10902_/A2 _11518_/Q _10902_/B2 _10631_/C _10636_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_14_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06625__I _11526_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10562_ _10562_/A1 _10562_/A2 _11657_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10234__A2 _10351_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05661__A2 _11626_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10493_ _10493_/A1 _10493_/A2 _10494_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_154_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09927__A2 _09927_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05949__B1 _08803_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11114_ _11114_/D _11672_/CLK _11114_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11045_ _11050_/I _11692_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07166__A2 _11174_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11706__I input66/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_3_4__f_wb_clk_i_I clkbuf_0_wb_clk_i/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06677__A1 _11326_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10473__A2 _06563_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09615__A1 _09622_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_10829_ _10921_/A1 _11338_/Q _10831_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06535__I _08493_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06429__A1 _08990_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09091__A2 _09015_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06020_ _09248_/A1 _11439_/Q _06022_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_160_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput326 _11126_/Q wb_dat_o[21] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput315 _11114_/Q wb_dat_o[11] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput304 _05841_/Z serial_data_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput337 _11674_/Q wb_dat_o[31] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__11401__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07971_ _07971_/A1 _07971_/A2 _07971_/A3 _08378_/B _07975_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__06601__A1 _06616_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09710_ _09154_/I _09722_/A2 _09710_/B _09711_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06922_ _06922_/I _11105_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11072__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11551__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08354__A1 _08656_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09641_ _09187_/Z _09647_/A2 _09641_/B _09642_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06853_ _06851_/Z _06869_/A2 _06853_/B _06854_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_27_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10161__A1 _10353_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09572_ _09270_/Z _09572_/A2 _09572_/B _09573_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06784_ _07114_/C _09015_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_20
XFILLER_55_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05804_ _05804_/I _09197_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_08523_ _07844_/B _08523_/A2 _08524_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05735_ _05735_/I _05776_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11087__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input105_I wb_adr_i[17] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08454_ _08454_/A1 _08454_/A2 _08454_/A3 _08454_/A4 _08613_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__10464__A2 _11491_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05666_ _05666_/I _06324_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__09606__A1 _09622_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08385_ _08385_/I _08453_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07405_ _05703_/Z _08825_/A1 _06838_/Z _07410_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_05597_ _05597_/A1 _05633_/B _05597_/B _05598_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11640__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07336_ _07340_/A2 _11226_/Q _07337_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07267_ _07267_/A1 _06838_/Z _07290_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA_input70_I mgmt_gpio_in[6] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09006_ _09013_/A2 _11360_/Q _09007_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07198_ _07198_/I _11180_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05643__A2 _05924_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06218_ _08786_/A1 _11144_/Q _06217_/Z _06219_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11081__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06840__A1 _06869_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06149_ _09324_/A1 _11461_/Q _06151_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08345__A1 _08490_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09908_ _10404_/A1 _09908_/A2 _10387_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09839_ _09158_/I _09848_/A2 _09839_/B _09840_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_73_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09845__A1 _09241_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06108__B1 _08799_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_11663_ _11663_/D input76/Z _11663_/CLK _11663_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XPHY_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_10614_ _11382_/Q _10884_/A1 _11374_/Q _10883_/A1 _10614_/C _10619_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_11594_ _11594_/D _11686_/RN _06705_/Z _11594_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__09073__A2 _11381_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11424__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08820__A2 _08820_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10545_ _10883_/A1 _11372_/Q _10547_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10476_ _10895_/A1 _11443_/Q _10477_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11574__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08584__B2 _08584_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11028_ _11028_/A1 _11028_/A2 _11030_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06898__A1 _06902_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08887__A2 _11322_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09836__A1 _09154_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05520_ _06611_/B2 _06610_/A3 _06444_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05873__A2 _11625_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08170_ _08170_/I _08181_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_32_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07121_ _11190_/Q _05927_/Z _07151_/B _07121_/C _07122_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__09064__A2 _09064_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08811__A2 _08820_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07052_ _07053_/A2 _11144_/Q _07053_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06003_ _11551_/Q _09599_/A1 _11543_/Q _09574_/A1 _06003_/C _06007_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__08575__A1 split8/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07378__A2 _11238_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput189 _06735_/ZN mgmt_gpio_oeb[24] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput178 _06056_/A1 mgmt_gpio_oeb[14] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_07954_ split15/I _08692_/A1 _08373_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07885_ _07885_/I _07886_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10134__A1 _11350_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06905_ _06905_/A1 _06904_/Z _06910_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09624_ _09624_/A1 _09015_/I _09647_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__06889__A1 _06902_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10134__B2 _10351_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06836_ _06836_/I _11078_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09827__A1 _09116_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09555_ _09555_/I _11532_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06767_ _07110_/I _11058_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09486_ _09486_/I _11510_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08506_ _08593_/A1 _08593_/A4 _08508_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05718_ _05718_/A1 _05751_/A2 _05719_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_06698_ _06266_/I _11297_/Q _06699_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08437_ _08437_/A1 _08437_/A2 _08653_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11447__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05649_ _05649_/I _08795_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_3
XFILLER_62_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07302__A2 _07419_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05864__A2 _09599_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08368_ _08363_/Z _08441_/B _08368_/A3 _08442_/B _08371_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__09055__A2 _09064_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08299_ _08299_/I _08301_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07319_ _07319_/I _11210_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11597__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10330_ _11147_/Q _10369_/A2 _10369_/B1 _11252_/Q _10333_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__05616__A2 _06466_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output274_I _11073_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10261_ _10374_/A1 _11537_/Q _10263_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05519__I _05519_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10373__A1 _10373_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10192_ _10192_/A1 _06556_/I _10880_/C _10192_/C _10194_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__11532__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10676__A2 _11447_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05552__A1 _05519_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11547__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11646_ _11646_/D input76/Z _11663_/CLK _11646_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__09046__A2 _09064_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11577_ _11577_/D _11686_/RN _06705_/Z _11577_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__07057__A1 _06837_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput36 mgmt_gpio_in[0] input36/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput14 mask_rev_in[19] input14/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput25 mask_rev_in[29] input25/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10600__A2 _11557_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10528_ _11444_/Q _10895_/A1 _10528_/B _10532_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xinput47 mgmt_gpio_in[1] input47/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput58 mgmt_gpio_in[2] input58/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput69 mgmt_gpio_in[5] input69/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_182_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11093__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10459_ _10922_/A1 _11355_/Q _10919_/A1 _11363_/Q _10468_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10116__A1 _10373_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10116__B2 _11525_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07670_ _07674_/A2 _08046_/B _07938_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10667__A2 _10888_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06621_ _11598_/Q _10638_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_25_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09340_ _09347_/A2 _11464_/Q _09341_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10419__A2 _09934_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06552_ _09938_/A2 _11627_/Q _06553_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07296__A1 _11016_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09271_ _09272_/A2 _11442_/Q _09272_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05503_ _05504_/A2 _11701_/Q _05504_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08222_ split7/Z _08232_/A2 _08222_/B _08476_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06483_ _06484_/A2 _06483_/A2 _11063_/Q _05515_/I _06486_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__05846__A2 _08890_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08153_ _08161_/A1 _08567_/A1 _08155_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07048__A1 _08786_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08084_ _08084_/A1 _08058_/I _08085_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07104_ _07081_/Z _07104_/A2 _07104_/B _07105_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07599__A2 _08509_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07035_ _07039_/A2 _11139_/Q _07036_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06271__A2 _06204_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10355__B2 _10355_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08986_ _08986_/I _11353_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07220__A1 _07240_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07937_ _07937_/A1 _08369_/B _08441_/C _07937_/A4 _07942_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA_input33_I mask_rev_in[7] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05782__A1 _06238_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07868_ _07870_/A1 _07870_/A3 _07869_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09607_ _09125_/Z _09622_/A2 _09607_/B _09608_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07799_ _07530_/I _07752_/I _08639_/B _07800_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_06819_ _06819_/I _11075_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09538_ _09158_/Z _09547_/A2 _09538_/B _09539_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07287__A1 _06863_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11025__B _11025_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09469_ _09241_/Z _09472_/A2 _09469_/B _09470_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_11500_ _11500_/D _11686_/RN _06705_/Z _11500_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__10291__B1 _10369_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10830__A2 _11370_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11431_ _11431_/D input76/Z _06705_/Z _11431_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__07039__A1 _06843_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08787__A1 _06904_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06633__I _06633_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11362_ _11362_/D _11686_/RN _06705_/Z _11362_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__10594__A1 _10899_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11075__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10313_ _10353_/A1 _11109_/Q _10315_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11293_ _11293_/D _06705_/Z _11293_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_152_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10244_ _10361_/A1 _11425_/Q _10245_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10175_ _10367_/A1 _11479_/Q _10177_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10897__A2 _10897_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11612__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10649__A2 _11358_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07278__A1 _06851_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1182 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_179_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10821__A2 _10913_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05828__A2 _05828_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08490__A3 _08490_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11629_ _11629_/D input76/Z _11665_/CLK _11629_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__08778__A1 _06859_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10585__A1 _10910_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07450__A1 _07513_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11142__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_944 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_911 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07202__A1 _05924_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08840_ _08844_/A2 _11307_/Q _08841_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07753__A2 _08242_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_977 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_966 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08950__A1 _08963_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_999 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05983_ _08761_/A1 _11288_/Q _05984_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08771_ _08784_/A2 _11287_/Q _08772_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11292__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07722_ _07722_/I _08332_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_07653_ _08283_/B _07609_/Z _07656_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05516__A1 _06466_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06604_ _06604_/A1 _11690_/Q _06604_/B _06605_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07584_ _08669_/A2 _07609_/I _07589_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09323_ _09323_/I _11458_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09258__A2 _11438_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06535_ _08493_/B _11028_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__07269__A1 _07076_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10812__A2 _11562_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05819__A2 _08719_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06466_ _06478_/A2 _06480_/A1 _06466_/B _06478_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09254_ _09254_/I _11436_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08205_ _08519_/A2 _08623_/A2 split12/Z _08205_/C _08206_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_21_498 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_09185_ _09158_/Z _09195_/A2 _09185_/B _09186_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08136_ _08161_/A1 _08222_/B _08476_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06397_ _06397_/A1 _06397_/A2 _06397_/A3 _06397_/A4 _06398_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__08769__A1 _06847_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10576__A1 _10896_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08067_ _08067_/A1 _08067_/A2 _08068_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06244__A2 _06238_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10328__A1 _10366_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07018_ _06843_/Z _07018_/A2 _07018_/B _07019_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11635__CLK _11658_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09194__A1 _09195_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08941__A1 _08963_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10879__A2 _10092_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output237_I _06649_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05755__A1 _07419_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08969_ _08988_/A2 _11348_/Q _08970_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09497__A2 _09497_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10931_ _10931_/A1 _10931_/A2 _10931_/B _10932_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10500__B2 _11515_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10500__A1 _11523_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06704__B1 _05616_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06180__A1 _09750_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10862_ _10862_/I _10863_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_10793_ _10793_/A1 _10793_/A2 _10794_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10803__A2 _11450_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_287 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11296__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11165__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11414_ _11414_/D input76/Z _06705_/Z _11414_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__09421__A2 _11490_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11345_ _11345_/D _11686_/RN _06705_/Z _11345_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_11276_ _11276_/D _11686_/RN _06705_/Z _11276_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__09185__A1 _09158_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10227_ _10265_/A1 _11328_/Q _10265_/A3 _10228_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08932__A1 _06859_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11220__RN input162/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05746__A1 _08799_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10158_ _11335_/Q _10159_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10089_ _10881_/A1 _11647_/Q _10090_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09488__A2 _09497_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07499__A1 _07513_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08160__A2 _08656_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06171__A1 input47/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11508__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06320_ _09775_/A1 _11603_/Q _06323_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09660__A2 _09672_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06251_ _07427_/A1 _11253_/Q _06252_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06474__A2 _06610_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11363__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09412__A2 _11487_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06182_ _06192_/I _05636_/I _07349_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_143_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11658__CLK _11658_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06226__A2 _11412_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09941_ _09944_/B1 _09945_/A2 _06520_/I _09922_/B _09942_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__05985__A1 _09041_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09176__A1 _09121_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07726__A2 _08490_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09872_ _09902_/I _09958_/A1 _09872_/B _09873_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08923__A1 _06847_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10730__A1 _10904_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_08823_ _05836_/I _08827_/A2 _08823_/B _08824_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05737__A1 _06192_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_796 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input135_I wb_dat_i[14] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08754_ _08754_/I _11281_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05966_ _10195_/A2 _05991_/I _05966_/B _05966_/C _05967_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__09479__A2 _09497_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07705_ _08630_/A2 _07697_/I _08543_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_38_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08685_ _08685_/I _11259_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05897_ _05584_/I _11269_/Q _05898_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07636_ _08417_/B _07609_/Z _07639_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07567_ _08248_/B _07609_/I _07574_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09306_ _09322_/A2 _11453_/Q _09307_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06518_ _06518_/A1 _06266_/I _06519_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11188__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07498_ _08300_/A2 _07522_/I _07858_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__09651__A2 _09672_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11278__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10797__A1 _10886_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09237_ _09237_/I _11431_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06449_ _06449_/I _06454_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_output187_I _10148_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09168_ _09169_/A2 _11410_/Q _09169_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10549__A1 _10889_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08119_ _08434_/A1 _08220_/B _08218_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07414__A1 _07076_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09099_ _06847_/Z _09114_/A2 _09099_/B _09100_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_11130_ _11130_/D _11686_/RN _06705_/Z _11130_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__11450__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11061_ _11061_/D _11061_/RN input68/Z _11061_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10012_ _10025_/A1 _09970_/I _10360_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__10721__B2 _10894_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11202__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06153__A1 _09424_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10914_ _10914_/A1 _11243_/Q _10914_/B1 _11239_/Q _10917_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__05900__A1 _09549_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11029__A2 _08672_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10845_ _10891_/A1 _11240_/Q _10847_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10776_ _10899_/A1 _11505_/Q _10779_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10788__A1 _10092_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07405__A1 _05703_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11328_ _11328_/D input76/Z _06705_/Z _11328_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_4_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05967__A1 _05967_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11441__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11259_ _11259_/D input162/Z _06687_/A2 _11259_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__07708__A2 _08495_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05820_ _05820_/I _09222_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_67_468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_287 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05751_ _05751_/A1 _05751_/A2 _05833_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__06144__A1 _06324_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05682_ _09800_/A1 _11618_/Q _05682_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08470_ _08214_/I _08470_/A2 _08586_/A3 _08576_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11330__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07421_ _07076_/Z _07424_/A2 _07421_/B _07422_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_90_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07352_ _07352_/I _11230_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06303_ _06259_/Z _06265_/Z _06303_/A3 _06303_/A4 _10938_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__11480__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07283_ _07290_/A2 _11202_/Q _07284_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06234_ _06234_/A1 _06234_/A2 _06234_/A3 _06234_/A4 _06235_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_09022_ _09022_/I _11364_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09397__A1 _09270_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11680__RN input162/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06165_ _06165_/A1 _06165_/A2 _06165_/A3 _06165_/A4 _06166_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__07947__A2 _08529_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06731__I _11446_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10951__A1 _10934_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06096_ _06096_/A1 _06096_/A2 _06097_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09149__A1 _09121_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11432__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09924_ _09936_/A2 _10392_/A1 _09927_/A2 _10440_/A1 _09925_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_09855_ _09866_/A2 _09938_/A1 _09855_/B _09856_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10703__A1 _10914_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08372__A2 _08686_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08806_ _08806_/I _11296_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_571 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_09786_ _09154_/I _09798_/A2 _09786_/B _09787_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06383__A1 _07412_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06998_ _06998_/I _11128_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08737_ _06851_/Z _08740_/A2 _08737_/B _08738_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05949_ _11283_/Q _08742_/A1 _08803_/A1 _05947_/Z _05949_/C _05953_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_121_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08668_ _08668_/I _08670_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07619_ _07619_/A1 _07619_/A2 _07623_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10630_ _10630_/A1 _10630_/A2 _10631_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08599_ _08599_/I _08600_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09624__A2 _09015_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10561_ _10881_/A1 _11657_/Q _10562_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10492_ _10492_/A1 _10492_/A2 _10492_/A3 _10510_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__09388__A1 _09158_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10942__A1 _10942_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11203__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05949__A1 _11283_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05949__B2 _05947_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11423__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06071__B1 _11526_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11113_ _11113_/D _11672_/CLK _11113_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11044_ _11050_/I _11691_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09952__I _09952_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09560__A1 _09154_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06374__A1 _09449_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11353__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10170__A2 _11423_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06677__A2 _06701_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10473__A3 _09920_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10828_ _10920_/A1 _11346_/Q _10920_/B1 _11354_/Q _10831_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_10759_ _11417_/Q _10888_/A1 _11409_/Q _10889_/A1 _10759_/C _10763_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__09379__A1 _09121_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11662__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput316 _11115_/Q wb_dat_o[12] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput305 _06700_/Z serial_load VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_141_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput327 _11127_/Q wb_dat_o[22] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__11414__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput338 _11211_/Q wb_dat_o[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_07970_ split15/Z _08609_/B _08378_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06921_ _06837_/Z _06924_/A2 _06921_/B _06922_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09551__A1 _09116_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09640_ _09647_/A2 _11560_/Q _09641_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06852_ _06869_/A2 _11082_/Q _06853_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09571_ _09572_/A2 _11538_/Q _09572_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06783_ _06783_/I _07114_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_05803_ _06217_/I _05803_/A2 _05804_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08522_ _08522_/A1 _08522_/A2 _08522_/A3 _08522_/A4 _08524_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_05734_ _05802_/A2 _05624_/I _05735_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06117__A1 _08761_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08453_ _08453_/A1 _08562_/A2 _08454_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_07404_ _07404_/I _11245_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05665_ _08825_/A2 _06872_/A2 _05666_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06668__A2 _06701_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08384_ _08454_/A1 _08454_/A2 _08392_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05596_ _08523_/A2 _05633_/B _05597_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06726__I _11350_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07335_ _06213_/Z _06904_/Z _07340_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07266_ _07266_/I _11196_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08290__A1 _08394_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06217_ _06217_/I _06217_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__11653__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09005_ _09005_/I _11359_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11226__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07197_ _07197_/A1 _07197_/A2 _07197_/B _07198_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input63_I mgmt_gpio_in[34] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06840__A2 _11079_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08042__A1 _08614_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06148_ _06148_/A1 _06148_/A2 _06148_/A3 _06166_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__10924__A1 _10924_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06079_ _11366_/Q _06082_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06053__B1 _11414_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09907_ _11637_/Q _10404_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__11376__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09838_ _09848_/A2 _11623_/Q _09839_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_09769_ _09773_/A2 _11601_/Q _09770_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06108__B2 _06108_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_74 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05867__B1 _09624_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06636__I _06636_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11662_ _11662_/D input76/Z _11663_/CLK _11662_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XPHY_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_11593_ _11593_/D _11686_/RN _06705_/Z _11593_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10613_ _10410_/I _10613_/A2 _10417_/I _10613_/B1 _10494_/I _10614_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_10544_ _10922_/A1 _11356_/Q _10920_/B1 _11348_/Q _10547_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11644__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10475_ _10642_/A1 _10406_/I _10895_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_123_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08584__A2 _08431_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10915__A1 _10915_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11027_ _11027_/A1 _08036_/B _11030_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06347__A1 _05703_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07151__B _07151_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10851__B1 _10897_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11249__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07120_ _05927_/Z _09121_/I _07121_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06822__A2 _05633_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07051_ _07051_/I _11143_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11399__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06002_ _06002_/A1 _06002_/A2 _06003_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09772__A1 _09773_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08575__A2 _07727_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10906__A1 _10906_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput179 _06731_/ZN mgmt_gpio_oeb[15] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__10382__A2 _10382_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07953_ split21/Z _08692_/A1 _07955_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_498 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07884_ _07873_/Z _08013_/A2 _08359_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__09524__A1 _05693_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06904_ _09015_/I _06904_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__10134__A2 _10351_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09623_ _09623_/I _11554_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06835_ _06835_/A1 _09270_/I _06835_/B _06836_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05561__A2 _05519_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09554_ _09121_/Z _09572_/A2 _09554_/B _09555_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06766_ _07110_/I _11057_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09485_ _09154_/Z _09497_/A2 _09485_/B _09486_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08505_ _08696_/A2 _08509_/A1 _08505_/B _08593_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05717_ _05717_/I _05751_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
X_06697_ _11644_/Q _09944_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_36_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_08436_ _08449_/A1 _08010_/I _08436_/B _08437_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_168_115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05648_ _05930_/A1 _05753_/A2 _05649_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07302__A3 _06871_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08367_ _08383_/A1 _08355_/I _08367_/B _08442_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05579_ _11702_/Q _11687_/Q _05580_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07318_ _10942_/A1 _07310_/I _07318_/B _07319_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11626__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08298_ _07586_/I _08495_/B _08298_/B _08299_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07249_ _07265_/A2 _11191_/Q _07250_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10070__A1 _10367_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10260_ _10373_/A1 _11521_/Q _10373_/B1 _11529_/Q _10263_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06026__B1 _07201_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09763__A1 _09773_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output267_I _11276_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10191_ _10191_/A1 _06556_/I _10192_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06577__A1 _06577_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09515__A1 _09522_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10125__A2 _11325_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11645_ _11645_/D input76/Z _11658_/CLK _11645_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__11071__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11541__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11576_ _11576_/D _11686_/RN _06705_/Z _11576_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__11617__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput37 mgmt_gpio_in[10] input37/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput26 mask_rev_in[2] input26/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput15 mask_rev_in[1] input15/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput59 mgmt_gpio_in[30] input59/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput48 mgmt_gpio_in[20] input48/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10527_ _10527_/A1 _10527_/A2 _10527_/A3 _10527_/A4 _10528_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_6_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10458_ _10463_/A1 _10406_/I _10919_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__11086__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11691__CLK input68/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09754__A1 _09773_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10389_ _10389_/I _10456_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_123_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07146__B _07151_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09506__A1 _09522_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10116__A2 _11517_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06620_ _06620_/I _11689_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06551_ _11628_/Q _09938_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11071__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09270_ _09270_/I _09270_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_06482_ _11064_/Q _06483_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05502_ _05501_/Z _06456_/A2 _05504_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08221_ _08221_/A1 _08475_/A1 _08221_/A3 _08472_/B _08225_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__08245__A1 _07990_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08152_ split7/Z _08567_/A1 _08155_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07048__A2 _06217_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11608__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08083_ split8/I _08656_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_07103_ _07104_/A2 _11158_/Q _07104_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08796__A2 _07114_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07034_ _07398_/A1 _06217_/Z _06871_/Z _07039_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__09745__A1 _09241_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input165_I wb_sel_i[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10355__A2 _10355_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08985_ _06863_/Z _08988_/A2 _08985_/B _08986_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07936_ _08355_/I _08364_/B _07937_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05782__A2 _06872_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input26_I mask_rev_in[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07867_ _07867_/A1 _07867_/A2 _07870_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11414__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09606_ _09622_/A2 _11549_/Q _09607_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07570__I _07570_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07798_ _07727_/I _08639_/B _08509_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08720__A2 _11271_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06818_ _06835_/A1 _09158_/I _06818_/B _06819_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09537_ _09547_/A2 _11527_/Q _09538_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06749_ _06749_/I _06760_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09468_ _09472_/A2 _11505_/Q _09469_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07287__A2 _07290_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11564__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_474 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06119__C _06119_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10291__B2 _11506_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09399_ _09399_/A1 _09015_/Z _09422_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_08419_ _08419_/A1 _07643_/I _08419_/B _08419_/C _08538_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_11430_ _11430_/D input76/Z _06705_/Z _11430_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_11361_ _11361_/D _11686_/RN _06705_/Z _11361_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_164_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10594__A2 _11501_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06798__A1 _06835_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10312_ _11105_/Q _10351_/A2 _11103_/Q _10351_/B2 _10312_/C _10325_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__09736__A1 _09154_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10880__B _10880_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11292_ _11292_/D _11686_/RN _06705_/Z _11292_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_140_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10346__A2 _10880_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10243_ _10360_/A1 _11433_/Q _10245_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10174_ _11455_/Q _10365_/A2 _10365_/B1 _11463_/Q _10177_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_19_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11094__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06722__A1 _06753_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07278__A2 _07290_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08227__A1 split7/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11628_ _11628_/D input76/Z _11665_/CLK _11628_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_8_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08778__A2 _08784_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_11559_ _11559_/D _11686_/RN _06705_/Z _11559_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__07450__A2 split16/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09727__A1 _09116_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_934 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_923 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_912 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07202__A2 _09116_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_978 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_967 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_956 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_945 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11437__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_989 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_287 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06961__A1 _10954_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05982_ _06839_/A1 _11083_/Q _05984_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08770_ _08770_/I _11286_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07721_ _08580_/A2 _08339_/A1 _07722_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_65_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11587__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07652_ _08537_/B _08283_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__08702__A2 _07844_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05516__A2 _06610_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07583_ _07583_/A1 _07583_/A2 _07589_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06603_ _10931_/A1 _10930_/B _11216_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06534_ _11225_/Q _08493_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
X_09322_ _09270_/Z _09322_/A2 _09322_/B _09323_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_43_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07269__A2 _07290_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06465_ _06484_/A2 _11064_/Q _06478_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10273__B2 _10351_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09253_ _09121_/Z _09272_/A2 _09253_/B _09254_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06734__I _11510_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08204_ _08204_/I _08623_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06396_ _06396_/A1 input4/Z _06397_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09184_ _09195_/A2 _11415_/Q _09185_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08135_ _08434_/A1 _08222_/B _08196_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09966__A1 _10375_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11531__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08769__A2 _08784_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10576__A2 _11437_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08066_ _08066_/A1 _08571_/B _08081_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09718__A1 _09722_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07017_ _07018_/A2 _11134_/Q _07018_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09194__A2 _11418_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06952__A1 _10945_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05755__A2 _08799_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08968_ _08968_/I _11347_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07919_ _07930_/A1 _08015_/A2 _07920_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08899_ _08899_/I _11325_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10930_ _11222_/D _11666_/Q _10930_/B _10930_/C _10931_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__10500__A2 _10902_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06704__A1 _07242_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10861_ _10861_/A1 _10861_/A2 _10862_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_10792_ _10887_/B1 _11434_/Q _10793_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_11413_ _11413_/D input76/Z _06705_/Z _11413_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__07432__A2 _11253_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11344_ _11344_/D _11686_/RN _06705_/Z _11344_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__09709__A1 _09722_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11275_ _11275_/D _11686_/RN _06705_/Z _11275_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_10226_ _10226_/A1 _10226_/A2 _10226_/A3 _10226_/A4 _10228_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__09185__A2 _09195_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07196__A1 _07197_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09724__A4 _07114_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06943__A1 _06941_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10157_ _10157_/I _11649_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05746__A2 _05803_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08932__A2 _08938_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_10088_ _10926_/C _10881_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XANTENNA__07499__A2 split13/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06171__A2 _05924_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07120__A1 _05927_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06250_ _06197_/I _05777_/I _07427_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_30_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05682__A1 _09800_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_285 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06181_ _06181_/A1 _06181_/A2 _06181_/B _06181_/C _06187_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__10558__A2 _10924_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09940_ _09940_/A1 _11092_/Q _09940_/B1 _09922_/B _09944_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_171_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09176__A2 _09195_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07187__A1 _07197_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09871_ _09958_/A1 _09935_/B _09872_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_786 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_08822_ _05836_/I _11302_/Q _06904_/Z _08823_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08923__A2 _08938_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05737__A2 _05738_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_797 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_08753_ _06851_/Z _08759_/A2 _08753_/B _08754_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05965_ _08940_/A1 _11344_/Q _05966_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07704_ _07704_/A1 _07704_/A2 _07704_/A3 _07704_/A4 _07711_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA_input128_I wb_adr_i[9] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06729__I _11414_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08684_ _08684_/A1 _07297_/I _08684_/B _08685_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05896_ _11268_/Q _05969_/I _05896_/B _06619_/B _05898_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_07635_ _07635_/I _08417_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__06162__A2 _11437_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07566_ _07566_/I _07609_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_139_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09305_ _09305_/I _11452_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06517_ _09942_/A1 _06694_/A1 _06519_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10246__A1 _11449_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07497_ _07533_/I _07675_/A2 _08300_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_139_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input93_I spimemio_flash_io3_oeb VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09236_ _09158_/Z _09246_/A2 _09236_/B _09237_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07662__A2 _08417_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06448_ _06458_/A2 _11069_/Q _06449_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11602__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06379_ _07370_/A1 _06238_/Z _11236_/Q _06380_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09167_ _09167_/I _11409_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08118_ _08575_/B _08220_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09098_ _09114_/A2 _11389_/Q _09099_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08049_ _08315_/B _08054_/A1 _08067_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11485__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07295__I _11025_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11060_ _11060_/D _11060_/RN input68/Z _11060_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10011_ _10030_/A2 _10265_/A3 _10025_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__10182__B1 _10373_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07717__A3 _08395_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10721__A2 _10894_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10485__A1 _10891_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09015__I _09015_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06639__I _06639_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10913_ _11247_/Q _10913_/A2 _11251_/Q _10913_/B2 _10913_/C _10917_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__11132__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10844_ _10844_/A1 _10844_/A2 _10844_/A3 _10844_/A4 _10872_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_157_213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10775_ _11545_/Q _10906_/A1 _11537_/Q _10905_/A1 _10775_/C _10779_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__07653__A2 _07609_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11282__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08850__A1 _08863_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08602__A1 _08602_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07405__A2 _08825_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11327_ _11327_/D _11686_/RN _06705_/Z _11327_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__07169__A1 _05925_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11258_ _11258_/D input162/Z _11683_/CLK _11258_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_11189_ _11189_/D _11686_/RN _06705_/Z _11189_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10209_ _10209_/A1 _10209_/A2 _10209_/A3 _10209_/A4 _10209_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_05750_ input33/Z _06396_/A1 input28/Z _06398_/A2 _05750_/C _05775_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__08669__A1 _08355_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05681_ _05681_/I _09800_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XANTENNA__10476__A1 _10895_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07420_ _07424_/A2 _11250_/Q _07421_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07351_ _07076_/Z _07354_/A2 _07351_/B _07352_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11625__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06302_ _06302_/A1 _06302_/A2 _06302_/A3 _06302_/A4 _06303_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_07282_ _07282_/I _11201_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07644__A2 _07609_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08841__A1 _07426_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05655__A1 _08825_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09021_ _07431_/Z _09039_/A2 _09021_/B _09022_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06233_ _06217_/Z _11033_/A2 _11138_/Q _06234_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__09397__A2 _09397_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06164_ _11453_/Q _09299_/A1 _11445_/Q _09274_/A1 _06164_/C _06165_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_144_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10951__A2 _11672_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06095_ _06394_/A1 input6/Z _06096_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09923_ _10426_/A2 _10394_/A2 _10440_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__09149__A2 _09169_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09854_ _09950_/A1 _09938_/A1 _09939_/I _09855_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11196__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08805_ _06855_/Z _08820_/A2 _08805_/B _08806_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06907__A1 _06837_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09785_ _09798_/A2 _11606_/Q _09786_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06383__A2 _06238_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06997_ _10957_/A1 _06974_/I _06997_/B _06998_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11155__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08736_ _08740_/A2 _11276_/Q _08737_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05948_ _08890_/A1 _11328_/Q _05949_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_66_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05879_ _05879_/A1 _05879_/A2 _05880_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08667_ _08667_/A1 _08667_/A2 _08536_/I _08667_/A4 _08672_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_53_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07332__A1 _07310_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07618_ _07618_/I _07619_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_53_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10219__A1 _10378_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08598_ _08598_/I _08601_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05894__A1 _05894_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07549_ input97/Z _07733_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09085__A1 _09089_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output297_I _11071_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10560_ _10560_/A1 _06556_/I _10880_/C _10560_/C _10562_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_139_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10491_ _10914_/A1 _11595_/Q _10914_/B1 _11603_/Q _10492_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11120__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09219_ _09220_/A2 _11426_/Q _09220_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09388__A2 _09397_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10942__A2 _10934_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06071__A1 _11534_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05949__A2 _08742_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06071__B2 _05693_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11112_ _11112_/D _11672_/CLK _11112_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06610__A3 _06610_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11043_ _11050_/I _11690_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09560__A2 _09572_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11187__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07571__A1 _08339_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06374__A2 _11499_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11648__CLK _11658_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07323__A1 _10947_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05885__A1 _09197_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09076__A1 _09089_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10827_ _10922_/A1 _11362_/Q _10831_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10758_ _10758_/A1 _10758_/A2 _10759_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05637__A1 _07419_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09379__A2 _09397_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10689_ _10689_/I _10690_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput317 _11116_/Q wb_dat_o[13] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput306 _06696_/ZN serial_resetn VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput328 _11128_/Q wb_dat_o[23] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_113_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput339 _11212_/Q wb_dat_o[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__06062__A1 _08846_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10933__A2 input162/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11178__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06920_ _06924_/A2 _11105_/Q _06921_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09000__A1 _09013_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11178__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10146__B1 _10146_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10697__A1 _10924_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06851_ _09154_/I _06851_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__09551__A2 _09572_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09570_ _09570_/I _11537_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06782_ _06782_/A1 _06782_/A2 _06783_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05802_ _05717_/I _05802_/A2 _05624_/I _06217_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_48_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08521_ _08521_/A1 _11016_/A1 _08522_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05733_ _05753_/A2 _05741_/A2 _06192_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__09303__A2 _11452_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08452_ _08648_/A3 _08650_/A2 _08648_/A2 _08455_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__07314__A1 _10938_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07403_ _07081_/Z _07403_/A2 _07403_/B _07404_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05664_ _09724_/A1 _05668_/I _06872_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_08383_ _08383_/A1 _08649_/B _08454_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05595_ _11256_/Q _08523_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11350__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09067__A1 _09089_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07617__A2 _07593_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08814__A1 _06859_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07334_ _07334_/I _11215_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07265_ _06867_/Z _07265_/A2 _07265_/B _07266_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10621__A1 _10892_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11102__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08290__A2 _08395_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09004_ _06855_/Z _09013_/A2 _09004_/B _09005_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06216_ _09248_/A1 _11436_/Q _06219_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07196_ _07197_/A1 _11180_/Q _07197_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08042__A2 _08358_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06147_ _06147_/A1 _06147_/A2 _06148_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input56_I mgmt_gpio_in[28] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06078_ _11382_/Q _09066_/A1 _11358_/Q _08990_/A1 _06078_/C _06098_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__06053__B2 _09171_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06053__A1 _11422_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09906_ _09906_/I _11636_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_76_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11169__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09837_ _09837_/I _11622_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06356__A2 _11451_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_391 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_09768_ _09768_/I _11600_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_18_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08719_ _08799_/A1 _08719_/A2 _06838_/Z _08724_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_09699_ _09699_/A1 _09015_/I _09722_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XPHY_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07856__A2 split16/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05867__B2 _11561_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10860__A1 _10906_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11661_ _11661_/D input76/Z _11663_/CLK _11661_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XPHY_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09058__A1 _06859_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_11592_ _11592_/D _11686_/RN _06705_/Z _11592_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10612_ _10612_/A1 _10612_/A2 _11658_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08805__A1 _06855_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_10543_ _10920_/A1 _11340_/Q _10921_/A1 _11332_/Q _10547_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07748__I _07748_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08281__A2 _08519_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_74 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10474_ _10896_/A1 _11435_/Q _10477_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09230__A1 _09125_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06044__A1 _06044_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06044__B2 _10144_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11320__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07792__A1 _08328_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07483__I _08495_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11470__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10679__A1 _10679_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11026_ _11026_/I _11032_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06347__A2 _08795_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09297__A1 _09270_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09049__A1 _06847_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11332__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07050_ _06837_/Z _07053_/A2 _07050_/B _07051_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06283__A1 _09091_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06001_ _09549_/A1 _11535_/Q _06002_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11399__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput169 _06744_/Z debug_in VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_07952_ _08355_/I _08692_/A1 _07955_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06903_ _06903_/I _11100_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07883_ _07883_/A1 _08357_/B _07883_/A3 _07887_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__09524__A2 _09015_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09622_ _09270_/Z _09622_/A2 _09622_/B _09623_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06834_ _06835_/A1 _11078_/Q _06835_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09553_ _09572_/A2 _11532_/Q _09554_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08504_ _07508_/I _07572_/I _08504_/B _08504_/C _08690_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__09288__A1 _09158_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input110_I wb_adr_i[21] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06765_ _07110_/I _11056_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09484_ _09497_/A2 _11510_/Q _09485_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05716_ _05716_/A1 _05716_/A2 _05717_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06696_ _06696_/A1 _06696_/A2 _06696_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08435_ _08435_/A1 _08435_/A2 _08435_/A3 _08435_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_05647_ _05647_/I _05753_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10842__A1 _10884_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08366_ _08366_/I _08368_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05578_ _06510_/A2 _06786_/A1 _05507_/I _05578_/B1 _05578_/B2 _11688_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_07317_ _07310_/I _11210_/Q _07318_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09460__A1 _09154_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08297_ _08204_/I _07748_/I _08297_/B _08676_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06274__A1 _08839_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07248_ _07248_/I _11190_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11343__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07179_ _05925_/Z _09158_/I _07180_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06026__B2 input56/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10190_ _10190_/A1 _10382_/A2 _10190_/B _10190_/C _10192_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__11493__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07774__A1 _08328_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06577__A2 _06556_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09515__A2 _11520_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07526__A1 _07575_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06329__A2 _06329_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10125__A3 _10265_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11562__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09279__A1 _09121_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07829__A2 _08632_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11314__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10833__A1 _10833_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11644_ _11644_/D input76/Z _11665_/CLK _11644_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__09451__A1 _09116_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11575_ _11575_/D _11686_/RN _06705_/Z _11575_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__08254__A2 _08519_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput16 mask_rev_in[20] input16/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput27 mask_rev_in[30] input27/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput49 mgmt_gpio_in[21] input49/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10526_ _10894_/B2 _11484_/Q _10527_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput38 mgmt_gpio_in[11] input38/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10457_ _10457_/I _10922_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XANTENNA__11010__A1 _08493_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10388_ _10493_/A2 _10426_/A2 _10389_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06568__A2 _10433_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09506__A2 _11517_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11009_ _11016_/A1 input158/Z _11012_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10788__B _10788_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11553__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11216__CLK _11666_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06550_ _06550_/I _11089_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10824__A1 _10914_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06481_ _06481_/I _11065_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05501_ _06610_/A3 _11070_/Q _11069_/Q _05501_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__11305__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09690__A1 _09697_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06099__A4 _06099_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08220_ split7/I _08232_/A2 _08220_/B _08472_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11366__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08151_ _08481_/B _08567_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07048__A3 _06871_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08082_ split12/I _08519_/A1 split8/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__06256__A1 _07419_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07102_ _07102_/I _11157_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_161_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07033_ _07033_/I _11138_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09745__A2 _09725_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input158_I wb_dat_i[6] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08984_ _08988_/A2 _11353_/Q _08985_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07935_ split21/I _08364_/B _08441_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07866_ input105/Z _06591_/I input106/Z split16/I _07867_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__08181__A1 _08490_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09605_ _09605_/I _11548_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11544__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07797_ _07722_/I _08639_/B _07800_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input19_I mask_rev_in[23] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06817_ _06835_/A1 _11075_/Q _06818_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09536_ _09536_/I _11526_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06748_ _06748_/I _06748_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09467_ _09467_/I _11504_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09681__A1 _09697_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08418_ _08418_/A1 _08418_/A2 _08627_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06679_ input1/Z input2/Z _06680_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10291__A2 _10369_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09398_ _09398_/I _11482_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08349_ _08349_/A1 _07297_/I _08349_/A3 _08349_/A4 _08398_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__06247__A1 _09424_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09984__A2 _10030_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11360_ _11360_/D _11686_/RN _06705_/Z _11360_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__06798__A2 _11072_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10311_ _10350_/A1 _10311_/A2 _10312_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_152_336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10880__C _10880_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11291_ _11291_/D input76/Z _06705_/Z _11291_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__09736__A2 _09725_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10242_ _11401_/Q _10359_/A2 _11393_/Q _10359_/B2 _10242_/C _10247_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_10173_ _10173_/A1 _10173_/A2 _10173_/A3 _10173_/A4 _10190_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__11239__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07761__I _07761_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08172__A1 _08490_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11535__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11269__CLKN input68/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11389__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10806__A1 _10806_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09672__A1 _09270_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10282__A2 _11434_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09424__A1 _09424_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11627_ _11627_/D input76/Z _11665_/CLK _11627_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_11558_ _11558_/D _11686_/RN _06705_/Z _11558_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__10034__A2 _10265_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07986__A1 split14/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10509_ _10509_/A1 _10509_/A2 _10509_/A3 _10509_/A4 _10510_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_11489_ _11489_/D _11686_/RN _06705_/Z _11489_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__10990__B1 _08460_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09727__A2 _09725_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_935 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_924 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_913 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_902 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_946 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06410__A1 _08786_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_979 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_07720_ _07720_/I _08580_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__06961__A2 _06941_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05981_ _06785_/A1 _11075_/Q _05984_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11526__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07651_ _07651_/A1 _07651_/A2 _07656_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_0_wb_clk_i wb_clk_i clkbuf_0_wb_clk_i/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07582_ _07582_/I _07583_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06602_ _11222_/Q _10930_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06533_ _06533_/I _11224_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09321_ _09322_/A2 _11458_/Q _09322_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09663__A1 _09158_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06464_ _06488_/A1 _06490_/B1 _06484_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10273__A2 _10351_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09252_ _09272_/A2 _11436_/Q _09253_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09415__A1 _09422_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08218__A2 _07722_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08203_ _08203_/I _08206_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06395_ _08799_/A1 _11271_/Q _08719_/A2 _06397_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_21_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09183_ _09183_/I _11414_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08134_ _08134_/I _08222_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07977__A1 _08355_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08065_ _08202_/A1 _08043_/I _08571_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05988__B1 _11383_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09718__A2 _11585_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07016_ _07016_/I _11133_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06952__A2 _06941_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08967_ _07426_/Z _08988_/A2 _08967_/B _08968_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_75_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07918_ _07918_/I _08015_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08154__A1 _08434_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11531__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08898_ _06847_/Z _08913_/A2 _08898_/B _08899_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07849_ input128/Z input98/Z _07851_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10860_ _10906_/A1 _11685_/Q _10861_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07901__A1 _07685_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09519_ _09241_/Z _09522_/A2 _09519_/B _09520_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_17_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11085__SETN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11681__CLK _06687_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08457__A2 _08545_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09654__A1 _09121_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_10791_ _10887_/A2 _11426_/Q _10793_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06468__A1 _06491_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_289 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_130_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09406__A1 _09422_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_172_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11412_ _11412_/D _11686_/RN _06705_/Z _11412_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__07968__A1 _08355_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05979__B1 _06518_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11343_ _11343_/D _11686_/RN _06705_/Z _11343_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__09709__A2 _11582_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11061__CLK input68/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11274_ _11274_/D _11686_/RN _06705_/Z _11274_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10225_ _10225_/A1 _10225_/A2 _10225_/A3 _10226_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08393__A1 _08395_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10724__B1 _10897_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10156_ _10191_/A1 _10880_/C _10156_/B _10157_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08145__A1 _08161_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10087_ _10087_/A1 _06556_/I _10880_/C _10087_/C _10090_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08696__A2 _08696_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10989_ _08493_/B input149/Z _10991_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07120__A2 _09121_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10007__A2 _10265_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06180_ _09750_/A1 _11596_/Q _06181_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11404__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06631__A1 input77/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06570__I _08460_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09870_ _11631_/Q _09958_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__10092__I _10092_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_710 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11554__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_08821_ _08821_/I _11301_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_754 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08136__A1 _08161_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_08752_ _08759_/A2 _11281_/Q _08753_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05964_ _11352_/Q _05723_/Z _08990_/A1 _11360_/Q _05966_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08683_ _08683_/A1 _07297_/I _08684_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07703_ _08426_/A1 _08290_/C _07704_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07634_ _07634_/A1 _08534_/C _07639_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09884__B2 _09902_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06698__A1 _06266_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05895_ _10954_/A1 _05969_/I _05896_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07565_ _08677_/A2 _08339_/A1 _07566_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_07496_ _07496_/I _07675_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_3
X_09304_ _09121_/Z _09322_/A2 _09304_/B _09305_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06516_ _11643_/Q _09942_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09121__I _09121_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09235_ _09246_/A2 _11431_/Q _09236_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06447_ _06456_/A1 _06456_/A2 _06458_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input86_I spimemio_flash_io0_do VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06378_ _06238_/Z _11240_/Q _11033_/A2 _06380_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09166_ _06863_/Z _09169_/A2 _09166_/B _09167_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11084__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08117_ _08117_/A1 _08117_/A2 _08122_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09097_ _09097_/I _11388_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08048_ _08048_/A1 split16/Z _08067_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10010_ _10135_/A1 _09970_/I _10363_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__10182__A1 _10373_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09999_ _10369_/B1 _11499_/Q _10006_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08127__A1 _08434_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06138__B1 _07201_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10912_ _10912_/A1 _10912_/A2 _10913_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xsplit21 split21/I split21/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_32_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_10843_ _10886_/B2 _11131_/Q _10886_/A2 _11133_/Q _10844_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_10774_ _10774_/A1 _10774_/A2 _10775_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06655__I _06655_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11427__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06861__A1 _06859_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08602__A2 _11016_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07405__A3 _06838_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11577__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11326_ _11326_/D input76/Z _06705_/Z _11326_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_4_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05967__A3 _05967_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11257_ _11257_/D input162/Z _11683_/CLK _11257_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__07169__A2 _09125_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11188_ _11188_/D input76/Z _06705_/Z _11188_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10208_ _11448_/Q _10363_/A2 _11440_/Q _10363_/B2 _10208_/C _10209_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_10139_ _10360_/A1 _11430_/Q _10141_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06392__A3 _06392_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05680_ _08825_/A2 _05803_/A2 _05681_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09618__A1 _09622_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07350_ _07354_/A2 _11230_/Q _07351_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10228__A2 _10092_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06301_ _06301_/A1 _06301_/A2 _06301_/A3 _06302_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_07281_ _06855_/Z _07290_/A2 _07281_/B _07282_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09876__I _09876_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09020_ _09039_/A2 _11364_/Q _09021_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05655__A2 _08799_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06852__A1 _06869_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06232_ _07370_/A1 _11136_/Q _06217_/I _06234_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06163_ _06163_/A1 _06163_/A2 _06164_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06514__B _06514_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06094_ _06393_/A1 input14/Z _06096_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09922_ _10642_/A1 _09935_/B _09922_/B _09936_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09853_ _09853_/A1 _10047_/B _09866_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10164__A1 _11383_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09784_ _09784_/I _11605_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input140_I wb_dat_i[19] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08804_ _08820_/A2 _11296_/Q _08805_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10164__B2 _10355_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_573 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_06996_ _06974_/I _11128_/Q _06997_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09116__I _09116_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07580__A2 _08204_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08735_ _08735_/I _11275_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05947_ _05947_/I _05947_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_45_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05878_ _09374_/A1 _11481_/Q _05879_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08666_ _08666_/A1 _08666_/A2 _08666_/A3 _08667_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__09609__A1 _09622_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08597_ _08594_/Z _08642_/A3 _08642_/A1 _08675_/A1 _08601_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_07617_ _08264_/B _07593_/I _07618_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07548_ _07548_/I _08589_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
X_07479_ _07479_/A1 _07479_/A2 _07690_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_14_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10490_ _10910_/A1 _11563_/Q _10492_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output192_I _10634_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09218_ _09218_/I _11425_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09149_ _09121_/Z _09169_/A2 _09149_/B _09150_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_497 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11111_ _11111_/D _11672_/CLK _11111_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06071__A2 _09549_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10155__A1 _10155_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11042_ _11050_/I _11042_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07020__A1 _07370_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09848__A1 _09270_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10458__A2 _10406_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10826_ _10826_/A1 _10826_/A2 _10826_/A3 _10826_/A4 _10833_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_32_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05885__A2 _11425_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09076__A2 _11382_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07087__A1 _07076_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08823__A2 _08827_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10757_ _10887_/B1 _11433_/Q _10758_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10688_ _10688_/A1 _10688_/A2 _10689_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05637__A2 _08825_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06834__A1 _06835_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08587__A1 _07609_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput307 _06742_/Z spi_sdi VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput329 _11667_/Q wb_dat_o[24] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput318 _11117_/Q wb_dat_o[14] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__06062__A2 input64/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08339__A1 _08339_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11309_ _11309_/D _11686_/RN _06705_/Z _11309_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__10146__A1 _09972_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05892__C _05892_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09000__A2 _11358_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06850_ _06850_/I _11081_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07011__A1 _06843_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05801_ _11522_/Q _09499_/A1 _11514_/Q _09474_/A1 _05801_/C _05827_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__09839__A1 _09158_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06781_ _11684_/Q _05633_/B _06782_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08520_ _08520_/A1 _08344_/I _08601_/A3 _08520_/A4 _08521_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__10449__A2 _10449_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05732_ _05732_/I _05741_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08451_ _08448_/Z _08553_/A2 _08455_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05663_ _05590_/I _05598_/I _05668_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__11484__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07402_ _07403_/A2 _11245_/Q _07403_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08382_ _08382_/A1 _08650_/A3 _08648_/A3 _08648_/A4 _08392_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_05594_ _11205_/Q _05633_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__09067__A2 _11379_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08814__A2 _08820_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07333_ _10957_/A1 _07310_/I _07333_/B _07334_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07264_ _07265_/A2 _11196_/Q _07265_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11499__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05628__A2 _06466_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09003_ _09013_/A2 _11359_/Q _09004_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06215_ _09222_/A1 _11428_/Q _06219_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07195_ _11204_/Q _05925_/Z _07195_/B _07197_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06146_ _06146_/A1 _06146_/A2 _06146_/A3 _06146_/A4 _06147_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_144_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11122__CLK _11672_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07250__A1 _06847_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06053__A2 _09197_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06077_ _10613_/B1 _05764_/I _05768_/I _10137_/B2 _06078_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA_input49_I mgmt_gpio_in[21] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09905_ _09922_/B _11636_/Q _09905_/B _09906_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10137__B2 _10137_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09836_ _09154_/I _09848_/A2 _09836_/B _09837_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08750__A1 _06847_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11437__SETN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09767_ _09187_/I _09773_/A2 _09767_/B _09768_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05564__A1 _05519_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06979_ _06974_/I _11122_/Q _06980_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11272__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09698_ _09698_/I _11578_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08718_ _11050_/I _11270_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08649_ _08649_/A1 _08692_/A2 _08649_/B _08650_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05867__A2 _09649_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11660_ _11660_/D input76/Z _11663_/CLK _11660_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XPHY_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09058__A2 _09064_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_11591_ _11591_/D _11686_/RN _06705_/Z _11591_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__07069__A1 _07419_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10611_ _10881_/A1 _11658_/Q _10612_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08805__A2 _08820_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10542_ _10542_/A1 _10542_/A2 _10542_/A3 _10542_/A4 _10548_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__05619__A2 _05515_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10473_ _10406_/I _06563_/I _09920_/I _10896_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__09230__A2 _09246_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11615__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11025_ _11221_/Q _11025_/A2 _11025_/B _11222_/Q _11026_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_92_502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10143__A4 _10143_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10300__A1 _10378_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10851__A2 _10897_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09049__A2 _09064_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10809_ _10809_/A1 _10809_/A2 _10810_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06843__I _09121_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11096__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06000_ _05693_/Z _11527_/Q _06002_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11145__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07480__A1 _07513_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10367__A1 _10367_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07232__A1 _05924_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07951_ _08444_/B _08692_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06902_ _06867_/Z _06902_/A2 _06902_/B _06903_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05794__A1 _06238_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11295__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07882_ _08386_/A1 _07593_/I _07883_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09621_ _09622_/A2 _11554_/Q _09622_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06833_ _05616_/C _11682_/Q _06833_/B _09270_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_09552_ _09552_/I _11531_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06764_ _11055_/I _07110_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_08503_ _08497_/Z _08588_/A1 _08636_/I _08586_/A1 _08508_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_05715_ _05715_/I _05716_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09483_ _09483_/I _11509_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06695_ _06266_/I _11298_/Q _06696_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08434_ _08434_/A1 _08361_/B _08435_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05646_ _05646_/A1 _05610_/I _05647_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input103_I wb_adr_i[15] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08365_ split8/I _08607_/B _08365_/B _08366_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05577_ _11688_/Q _05578_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08799__A1 _08799_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07316_ _07316_/A1 _07316_/A2 _11209_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09460__A2 _09472_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08296_ _08296_/A1 _08431_/B _08349_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07247_ _07081_/Z _07265_/A2 _07247_/B _07248_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06274__A2 _07419_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07178_ _07178_/I _11176_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06026__A2 _05927_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06129_ _09649_/A1 _11565_/Q _06131_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11638__CLK _11666_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05785__A1 _06238_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09819_ _09823_/A2 _11617_/Q _09820_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10530__A1 _10897_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10833__A2 _10092_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11643_ _11643_/D input76/Z _11665_/CLK _11643_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__11168__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09451__A2 _09472_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10597__A1 _10900_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11574_ _11574_/D _11686_/RN _06705_/Z _11574_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xinput17 mask_rev_in[21] input17/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput28 mask_rev_in[31] input28/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10525_ _10891_/A1 _11476_/Q _10527_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput39 mgmt_gpio_in[12] input39/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10456_ _10456_/A1 _10506_/A2 _10457_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07214__A1 _07240_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07765__A2 _07761_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_253 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10387_ _10387_/I _10493_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__06568__A3 _09934_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08962__A1 _08963_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11250__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11008_ _11008_/I _11680_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07517__A2 _07522_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09911__B1 _09922_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05528__A1 _06446_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08190__A2 _07535_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10521__A1 _10913_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10788__C _10880_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06838__I _09015_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06480_ _06480_/A1 _06479_/C _06480_/B _06481_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05500_ _11159_/Q _06610_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
X_08150_ _08150_/A1 _08567_/C _08155_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10588__A1 _10911_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07101_ _07076_/Z _07104_/A2 _07101_/B _07102_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08081_ _08081_/A1 _08081_/A2 _08464_/A2 _08081_/A4 _08090_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__06256__A2 _06238_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07032_ _06843_/Z _07032_/A2 _07032_/B _07033_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06008__A2 _11463_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07205__A1 _07240_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08953__A1 _08963_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11241__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10760__A1 _10884_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08983_ _08983_/I _11352_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05767__A1 _07006_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07934_ split15/I _08364_/B _08369_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07865_ _07865_/A1 _07865_/A2 _07463_/Z _07867_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__10107__A4 _10107_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08181__A2 _08614_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09604_ _09121_/Z _09622_/A2 _09604_/B _09605_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07796_ _07796_/A1 _08507_/C _08325_/B _07796_/A4 _07800_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_06816_ _11694_/Q _05633_/B _06816_/B _09158_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_09535_ _09154_/Z _09547_/A2 _09535_/B _09536_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06747_ _11308_/Q input39/Z _06748_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09466_ _09187_/Z _09472_/A2 _09466_/B _09467_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06678_ _06678_/I _06678_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11310__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09130__A1 _06851_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08417_ split15/Z _08417_/A2 _08417_/B _08418_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05629_ _06480_/A1 _05515_/I _05630_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09397_ _09270_/Z _09397_/A2 _09397_/B _09398_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10579__A1 _10892_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08348_ _08348_/A1 _08348_/A2 _08348_/A3 _08348_/B _08349_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_164_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11460__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08279_ _08279_/A1 _08538_/A2 _08279_/A3 _08628_/B _08284_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_22_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11290_ _11290_/D input76/Z _06705_/Z _11290_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_10310_ _11101_/Q _10311_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11480__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10241_ _10241_/A1 _10241_/A2 _10242_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09197__A1 _09197_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08944__A1 _08963_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10751__A1 _11625_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11232__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05758__A1 _08791_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10172_ _11447_/Q _10363_/A2 _11439_/Q _10363_/B2 _10172_/C _10173_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_154_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10751__B2 _10915_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08172__A2 _08614_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10503__A1 _10506_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06183__A1 _09800_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_74 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09672__A2 _09672_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11299__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_11626_ _11626_/D _11686_/RN _06705_/Z _11626_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__09424__A2 _09015_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11557_ _11557_/D _11686_/RN _06705_/Z _11557_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_155_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10508_ _10889_/A1 _11403_/Q _10509_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11471__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11488_ _11488_/D _11686_/RN _06705_/Z _11488_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__10990__A1 _08431_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09188__A1 _09195_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10439_ _10913_/A2 _11587_/Q _10442_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_914 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_903 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08935__A1 _06863_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_958 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_947 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_936 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11223__RN input162/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05980_ _11277_/Q _08726_/A1 _11282_/Q _08742_/A1 _05980_/C _05984_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__06410__A2 _08799_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_969 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09360__A1 _09154_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06174__A1 _07201_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07650_ _08537_/B _08686_/A2 _07651_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11333__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06601_ _06616_/A1 _11216_/Q _10931_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07581_ _08669_/A2 _07593_/I _07582_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09320_ _09320_/I _11457_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06532_ _06749_/I _08672_/B _06532_/B _06533_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09663__A2 _09672_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09251_ _09251_/I _11435_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11483__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08202_ _08202_/A1 _08202_/A2 _08202_/B _08203_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06463_ _11062_/Q _11061_/Q _11060_/Q _06488_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_21_446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09415__A2 _11488_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06394_ _06394_/A1 input34/Z _06397_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09182_ _09154_/Z _09195_/A2 _09182_/B _09183_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08133_ _08133_/A1 _08565_/C _08138_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07977__A2 _08380_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08064_ split12/I _08202_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_161_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11462__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10981__A1 _11016_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09179__A1 _09125_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05988__B2 _09066_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07015_ _06837_/Z _07018_/A2 _07015_/B _07016_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08926__A1 _06851_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10733__A1 _10906_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input31_I mask_rev_in[5] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08966_ _08988_/A2 _11347_/Q _08967_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07917_ _07917_/A1 _08095_/A2 _07918_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09351__A1 _09116_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08897_ _08913_/A2 _11325_/Q _08898_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07848_ _07875_/A1 _08006_/A2 _07874_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05912__A1 _09424_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09518_ _09522_/A2 _11521_/Q _09519_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07779_ _08328_/B1 _08315_/B _08317_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08457__A3 _08656_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09654__A2 _09672_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_10790_ _10790_/A1 _10790_/A2 _11662_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_09449_ _09449_/A1 _09015_/Z _09472_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XPHY_257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09406__A2 _11485_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07417__A1 _07081_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11411_ _11411_/D _11686_/RN _06705_/Z _11411_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_149_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11342_ _11342_/D _11686_/RN _06705_/Z _11342_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_180_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10972__A1 _10972_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06941__I _06941_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05979__A1 _05833_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11206__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11273_ _11273_/D _11686_/RN _06705_/Z _11273_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10224_ _10375_/A1 _11544_/Q _10225_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08917__A1 _07426_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09590__A1 _09597_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08393__A2 _08545_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10724__B2 _11464_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11205__RN input162/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10155_ _10155_/A1 _06556_/I _10926_/C _10155_/C _10156_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__11356__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10086_ _10086_/A1 _06556_/I _10087_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06156__A1 _11517_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06156__B2 _09474_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05903__A1 _09624_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10988_ _11016_/A1 input155/Z _10991_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_175_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11609_ _11609_/D _11686_/RN _06705_/Z _11609_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__06851__I _09154_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06631__A2 input90/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09581__A1 _09597_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_08820_ _07431_/Z _08820_/A2 _08820_/B _08821_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10715__A1 _10884_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_711 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07682__I _07682_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_766 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10191__A2 _06556_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06395__A1 _08799_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08751_ _08751_/I _11280_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05963_ _11336_/Q _10195_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_57_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05894_ _05894_/A1 _05894_/A2 _05894_/A3 _05894_/A4 _10954_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_08682_ _08682_/A1 _08682_/A2 _08683_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07702_ _07702_/I _08426_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07633_ _07635_/I _08686_/A2 _08534_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07564_ _07564_/I _08677_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_07495_ _07690_/A2 _07495_/A2 _08423_/A2 _07689_/B _07539_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_09303_ _09322_/A2 _11452_/Q _09304_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06515_ _06515_/I _11056_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09234_ _09234_/I _11430_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06446_ _06446_/I _06456_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_119_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11683__RN input162/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11229__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09165_ _09169_/A2 _11409_/Q _09166_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08116_ split8/I _08575_/B _08117_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06377_ _09349_/A1 _11467_/Q _06380_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_174_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10954__A1 _10954_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input79_I spi_csb VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09096_ _07431_/Z _09114_/A2 _09096_/B _09097_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11268__CLKN input68/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08047_ _08048_/A1 _08047_/A2 _08114_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11379__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09572__A1 _09270_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08375__A2 _08355_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10706__A1 _10910_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10182__A2 _11519_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06386__A1 _09499_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09998_ _09998_/I _10369_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_130_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08949_ _08949_/I _11341_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10911_ _10911_/A1 _11146_/Q _10912_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08637__B _08637_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10842_ _10884_/A1 _11129_/Q _10844_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10773_ _10903_/A1 _11561_/Q _10774_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10642__B1 _10642_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06310__A1 _05925_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06861__A2 _06869_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10945__A1 _10945_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11426__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07810__A1 _08592_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11325_ _11325_/D _11686_/RN _06705_/Z _11325_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_11256_ _11256_/D input162/Z _11666_/CLK _11256_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_69_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09563__A1 _09158_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11187_ _11187_/D _11686_/RN _06705_/Z _11187_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10207_ _10207_/A1 _10207_/A2 _10208_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_395 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10138_ _11366_/Q _10353_/A1 _11358_/Q _10352_/A1 _10138_/C _10143_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__06129__A1 _09649_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10069_ _10366_/A1 _11468_/Q _10071_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06392__A4 _06392_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10228__A3 _10228_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07280_ _07290_/A2 _11201_/Q _07281_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06300_ _05723_/Z _11348_/Q _06301_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11665__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06231_ _09117_/A1 _11396_/Q _06234_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11521__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06162_ _09248_/A1 _11437_/Q _06163_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06065__B1 _09775_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10936__A1 _10934_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06093_ _06093_/A1 _06093_/A2 _06093_/A3 _06098_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__11417__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09921_ _10394_/A2 _10427_/A1 _10642_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__11084__SETN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09554__A1 _09121_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11671__CLK _11683_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09852_ _10092_/I _09935_/B _10047_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_541 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10164__A2 _10355_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_3_1__f_wb_clk_i_I clkbuf_0_wb_clk_i/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06368__A1 _07370_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09783_ _09125_/I _09798_/A2 _09783_/B _09784_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05925__I _05925_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08803_ _08803_/A1 _06904_/Z _08820_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_06995_ _06995_/I _11127_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input133_I wb_dat_i[12] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08734_ _06847_/Z _08740_/A2 _08734_/B _08735_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_05946_ _06266_/I _10385_/A1 _05946_/B _05947_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_38_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05877_ _09399_/A1 _11489_/Q _05879_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08665_ _08665_/A1 _08665_/A2 _08667_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_324 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08596_ _08596_/A1 _08596_/A2 _08596_/A3 _08596_/A4 _08675_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_07616_ _07616_/I _08264_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_14_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07547_ _07747_/A1 _08045_/A3 _07548_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07478_ _07478_/A1 _08006_/A2 _07875_/A3 _07479_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11656__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09217_ _06863_/Z _09220_/A2 _09217_/B _09218_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06429_ _08990_/A1 _11355_/Q _06432_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09148_ _09169_/A2 _11404_/Q _09149_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11408__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09079_ _09089_/A2 _11383_/Q _09080_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11110_ _11110_/D _11686_/RN _06705_/Z _11110_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__06359__A1 _08825_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11041_ _11050_/I _11688_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10155__A2 _06556_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07020__A2 _06217_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11605__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10825_ _10825_/A1 _10825_/A2 _10825_/A3 _10825_/A4 _10826_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__11544__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11647__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10756_ _10887_/A2 _11425_/Q _10758_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10687_ _10906_/A1 _11543_/Q _10688_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06834__A2 _11078_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08587__A2 _08592_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput308 _06723_/Z spimemio_flash_io0_di VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__11694__CLK input68/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10918__A1 _10918_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput319 _11118_/Q wb_dat_o[15] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_11308_ _11308_/D _11686_/RN _06705_/Z _11308_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_11239_ _11239_/D _11686_/RN _06705_/Z _11239_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__10146__A2 _10146_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05800_ _05800_/A1 _05800_/A2 _05801_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06780_ _05616_/C _11687_/Q _06782_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05731_ _11362_/Q _08990_/A1 _11354_/Q _05723_/Z _05731_/C _05775_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__11074__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05662_ _05662_/A1 _05662_/A2 _05662_/A3 _05662_/A4 _05683_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_08450_ _08450_/A1 _08450_/A2 _08553_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06576__I _09935_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08381_ _08656_/A1 _08649_/B _08648_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07401_ _07401_/I _11244_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05876__A3 _05876_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05593_ _06498_/A2 _06466_/B _05593_/B _05597_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_16_390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10606__B1 _10919_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07332_ _07310_/I _11215_/Q _07333_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08275__A1 _08400_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11638__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07263_ _07263_/I _11195_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10082__A1 _10378_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07194_ _05925_/Z _09270_/I _07195_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06214_ _06213_/Z _11227_/Q _06219_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09002_ _09002_/I _11358_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06145_ _09750_/A1 _11597_/Q _06146_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09775__A1 _09775_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10385__A2 _10880_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06076_ _11374_/Q _10137_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07250__A2 _07265_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09904_ _09927_/A2 _11636_/Q _09905_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09835_ _09848_/A2 _11622_/Q _09836_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11417__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_393 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_09766_ _09773_/A2 _11600_/Q _09767_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06978_ _10938_/A1 _06990_/A2 _06980_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08750__A2 _08759_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05929_ _05660_/Z _11624_/Q _05933_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09697_ _09270_/Z _09697_/A2 _09697_/B _09698_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08717_ _11050_/I _11269_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_66_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08648_ _08648_/A1 _08648_/A2 _08648_/A3 _08648_/A4 _08651_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__11567__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_08579_ _08579_/A1 _08622_/A1 _08582_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_25_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_11590_ _11590_/D _11686_/RN _06705_/Z _11590_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__07069__A2 _06238_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10610_ _10092_/Z _11657_/Q _10610_/B _10880_/C _10612_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__11629__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06816__A2 _05633_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10073__A1 _10371_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10541_ _10905_/A1 _11532_/Q _10542_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09766__A1 _09773_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10472_ _10887_/A2 _11419_/Q _10477_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07110__I _07110_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09518__A1 _09522_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11024_ _11024_/I _11683_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10128__A2 _10880_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11097__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10808_ _10900_/A1 _11514_/Q _10809_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08257__A1 _08449_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10739_ _10920_/A1 _11344_/Q _10920_/B1 _11352_/Q _10742_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08009__A1 split12/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09757__A1 _09773_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06064__C _06064_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07480__A2 split16/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06035__A3 _06035_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07232__A2 _09241_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07950_ _07950_/A1 _08692_/C _07955_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09509__A1 _09522_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06901_ _06902_/A2 _11100_/Q _06902_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05794__A2 _08719_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06991__A1 _06974_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07881_ _07988_/A1 _08013_/A2 _07885_/I _08357_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09620_ _09620_/I _11553_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06832_ _11697_/Q _05633_/B _06833_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__06743__A1 input36/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09551_ _09116_/Z _09572_/A2 _09551_/B _09552_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06763_ _06763_/I _11055_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05714_ _05714_/A1 _05714_/A2 _05714_/A3 _05828_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_08502_ _08502_/A1 _08502_/A2 _08586_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09482_ _09125_/Z _09497_/A2 _09482_/B _09483_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06694_ _06694_/A1 _11642_/Q _06696_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08433_ _08433_/A1 _08433_/A2 _08693_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05645_ _05645_/I _05930_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08364_ _08383_/A1 _08355_/I _08364_/B _08441_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_149_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08248__A1 split21/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05576_ _11690_/Q _11068_/Q _05576_/B _05576_/C _05578_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_23_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08799__A2 _08799_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10055__A1 _10353_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07315_ _07310_/I _11209_/Q _07316_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08295_ _08295_/A1 _08430_/A1 _08430_/A3 _08295_/A4 _08296_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_07246_ _07265_/A2 _11190_/Q _07247_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09748__A1 _09270_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07177_ _07197_/A1 _07177_/A2 _07177_/B _07178_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11004__B1 _08460_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input61_I mgmt_gpio_in[32] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07223__A2 _05924_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06128_ _06128_/A1 _06128_/A2 _06128_/A3 _06128_/A4 _06166_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_06059_ _05660_/Z _11622_/Q _06063_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05785__A2 _05995_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06982__A1 _10942_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_319 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09818_ _09818_/I _11616_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_19_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08723__A2 _11272_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09749_ _09749_/I _11594_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10530__A2 _11452_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11642_ _11642_/D input76/Z _11663_/CLK _11642_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__09987__A1 _09896_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10046__A1 _10046_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11573_ _11573_/D _11686_/RN _06705_/Z _11573_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_155_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput18 mask_rev_in[22] input18/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10524_ _10894_/A2 _11492_/Q _10527_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput29 mask_rev_in[3] input29/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08380__B _08380_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09739__A1 _09158_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10455_ _10920_/A1 _11339_/Q _10920_/B1 _11347_/Q _10468_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11483__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10386_ _10386_/I _11655_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_287 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11007_ _11007_/A1 _10966_/Z _11007_/B _11008_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_92_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07150__A1 _05927_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11421__SETN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10285__A1 _11450_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11112__CLK _11672_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09978__A1 _10378_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07100_ _07104_/A2 _11157_/Q _07101_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_158_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08080_ split7/I _08200_/B _08081_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11436__SETN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11262__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07031_ _07032_/A2 _11138_/Q _07032_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_161_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07685__I _07685_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08402__A1 split15/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06964__A1 _10957_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08982_ _06859_/Z _08988_/A2 _08982_/B _08983_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05767__A2 _08799_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07933_ _08607_/B _08364_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07864_ _07465_/I _07864_/A2 _07865_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_110_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08705__A2 _11261_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06815_ _11000_/A1 _05633_/B _06816_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09603_ _09622_/A2 _11548_/Q _09604_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06716__A1 _06753_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07795_ _08592_/A2 _08509_/A2 _07796_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09534_ _09547_/A2 _11526_/Q _09535_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06746_ _06746_/I _06746_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09465_ _09472_/A2 _11504_/Q _09466_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06677_ _11326_/Q _06701_/I _06677_/B _06678_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09130__A2 _09142_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08416_ _08535_/A2 _08535_/A3 _08420_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05628_ _06474_/B _06466_/B _11205_/Q _05630_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09396_ _09397_/A2 _11482_/Q _09397_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07692__A2 split5/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11605__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05559_ _11692_/Q _05561_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08347_ _08347_/A1 _08600_/A1 _11025_/B _08348_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_11_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08278_ _08400_/A1 _07643_/I _08278_/B _08628_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07229_ _07240_/A1 _11186_/Q _07230_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10240_ _10357_/A1 _11417_/Q _10241_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09197__A2 _09015_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output265_I _11274_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06955__A1 _06941_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10200__B2 _10355_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05758__A2 _08799_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10171_ _10171_/A1 _10171_/A2 _10172_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10751__A2 _10916_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08172__A3 _08656_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11135__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10267__A1 _10092_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05694__A1 _05693_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11285__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11625_ _11625_/D _11686_/RN _06705_/Z _11625_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_11556_ _11556_/D _11686_/RN _06705_/Z _11556_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_116_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10507_ _10507_/I _10889_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_11487_ _11487_/D _11686_/RN _06705_/Z _11487_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10438_ _10478_/A1 _09934_/I _10913_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XTAP_926 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_915 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_904 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_10369_ _11148_/Q _10369_/A2 _10369_/B1 _11253_/Q _10372_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_88_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06946__A1 _06941_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08935__A2 _08938_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_959 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_948 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_937 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06410__A3 _11292_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08699__A1 _08699_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09360__A2 _09372_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06600_ _06600_/A1 _06600_/A2 _06616_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07580_ _07530_/I _08204_/I _07593_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__10258__A1 _10377_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06531_ _11219_/Q _06532_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11628__CLK _11665_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09250_ _09116_/Z _09272_/A2 _09250_/B _09251_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08201_ _08205_/C _08242_/A1 _08202_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06462_ _06479_/C _06497_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06393_ _06393_/A1 input11/Z _06397_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09181_ _09195_/A2 _11414_/Q _09182_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08132_ split8/I _08134_/I _08565_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08063_ _08573_/A3 _08063_/A2 _08063_/A3 _08066_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__10430__A1 _10408_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09179__A2 _09195_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05988__A2 _09091_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07014_ _07018_/A2 _11133_/Q _07015_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input163_I wb_sel_i[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08926__A2 _08938_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10733__A2 _11544_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08965_ _05723_/Z _06838_/Z _08988_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__06401__A3 _05833_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07916_ _07916_/A1 _07916_/A2 _08435_/A2 _07916_/A4 _07923_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__11158__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input24_I mask_rev_in[28] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08896_ _08896_/I _11324_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07847_ _07847_/I _07875_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__09351__A2 _09372_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06165__A2 _06165_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07778_ _08696_/A2 _08315_/B _08504_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09517_ _09517_/I _11520_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10249__A1 _10366_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06729_ _11414_/Q _10615_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_169_213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_214 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08862__A1 _08863_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09448_ _09448_/I _11498_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05676__A1 _08825_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09379_ _09121_/Z _09397_/A2 _09379_/B _09380_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11150__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_149_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11410_ _11410_/D input76/Z _06705_/Z _11410_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_20_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11341_ _11341_/D _11686_/RN _06705_/Z _11341_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__10972__A2 _10966_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05979__A2 _05700_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11272_ _11272_/D input76/Z _06705_/Z _11272_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_165_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10223_ _10374_/A1 _11536_/Q _10225_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06928__A1 _06837_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08917__A2 _08938_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09590__A2 _11544_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10724__A2 _10897_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10154_ _10154_/A1 _06556_/I _10155_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10085_ _10558_/A1 _10382_/A2 _10085_/B _10085_/C _10087_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_66_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06156__A2 _09499_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10488__A1 _10916_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_355 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05903__A2 _11560_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10987_ _10987_/I _11677_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08853__A1 _08863_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10660__A1 _10910_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05667__A1 _06324_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11141__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11608_ _11608_/D _11686_/RN _06705_/Z _11608_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_30_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11539_ _11539_/D _11686_/RN _06705_/Z _11539_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__09030__A1 _06855_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09581__A2 _11541_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11300__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06919__A1 _07006_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_745 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06395__A2 _11271_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_789 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_05962_ _05962_/A1 _05962_/A2 _05962_/A3 _05962_/A4 _05967_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_08750_ _06847_/Z _08759_/A2 _08750_/B _08751_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10479__A1 _10897_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05893_ _05893_/A1 _05893_/A2 _05893_/A3 _05893_/A4 _05894_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_08681_ _08681_/A1 _11016_/A1 _08682_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07701_ _08294_/B _08394_/A1 _07702_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11450__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07344__A1 _07076_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07632_ _07640_/A1 _07694_/A2 _07635_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09884__A3 _09927_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07563_ _07836_/A1 _07579_/A1 _07564_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06528__B _06701_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09302_ _09302_/I _11451_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07494_ _07494_/I _08423_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08844__A1 _07431_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06514_ _06446_/I _06610_/B _06514_/B _06515_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06445_ _06445_/I _11172_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10651__A1 _10924_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09233_ _09154_/Z _09246_/A2 _09233_/B _09234_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11132__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09164_ _09164_/I _11408_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08115_ _08142_/A2 _08148_/A2 _08575_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06376_ _09324_/A1 _11459_/Q _06380_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09095_ _09114_/A2 _11388_/Q _09096_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08046_ _07995_/I _07506_/I _08046_/B _08047_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10954__A2 _10934_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06083__A1 _08742_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09021__A1 _07431_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09572__A2 _09572_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11199__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06386__A2 _11515_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09997_ _10000_/A1 _10042_/A2 _09998_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08948_ _06847_/Z _08963_/A2 _08948_/B _08949_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09324__A2 _09015_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08879_ _06855_/Z _08888_/A2 _08879_/B _08880_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06138__A2 _05927_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10910_ _10910_/A1 _11262_/Q _10912_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05897__A1 _05584_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xsplit12 split12/I split12/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09088__A1 _09089_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10841_ _10883_/A1 _11119_/Q _10844_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10772_ _10904_/A1 _11553_/Q _10774_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07638__A2 _08509_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10642__A1 _10642_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06310__A2 input72/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10945__A2 _10934_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11323__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11324_ _11324_/D _11686_/RN _06705_/Z _11324_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_11255_ _11255_/D input162/Z _06687_/A2 _11255_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_4_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09012__A1 _09013_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10206_ _10361_/A1 _11424_/Q _10207_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09563__A2 _09572_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11473__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11186_ _11186_/D input76/Z _06705_/Z _11186_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10137_ _10137_/A1 _10041_/I _10043_/I _10137_/B2 _10138_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_125_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10068_ _11452_/Q _10365_/A2 _10365_/B1 _11460_/Q _10071_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_35_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07326__A1 _10950_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07877__A2 _08358_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10330__B1 _10369_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05888__A1 _11409_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11362__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09079__A1 _09089_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07629__A2 _08417_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10633__A1 _10904_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06230_ _09144_/A1 _11404_/Q _06234_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06161_ _09222_/A1 _11429_/Q _06163_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06065__B2 _11606_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06065__A1 _11614_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06092_ _06092_/A1 _06092_/A2 _06092_/A3 _06092_/A4 _06093_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_09920_ _09920_/I _10427_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__09003__A1 _09013_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10149__B1 _11486_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07565__A1 _08677_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09554__A2 _09572_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09851_ _09950_/A1 _09939_/I _09853_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06368__A2 _11135_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09782_ _09798_/A2 _11605_/Q _09783_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06994_ _10954_/A1 _06974_/I _06994_/B _06995_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_08802_ _08802_/I _11295_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08733_ _08740_/A2 _11275_/Q _08734_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05945_ _06266_/I _11299_/Q _05946_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07317__A1 _07310_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05876_ _05876_/A1 _05876_/A2 _05876_/A3 _05876_/A4 _05894_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_08664_ _08664_/A1 _08664_/A2 _08664_/A3 _08664_/A4 _08667_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA_input126_I wb_adr_i[7] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08595_ _07609_/Z _08329_/B _08596_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07615_ _07640_/A1 _07649_/A2 _07616_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11353__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07546_ _07530_/I _07601_/I _07747_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08817__A1 _06863_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10624__A1 _10895_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11105__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07477_ _07477_/I _07875_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09490__A1 _09497_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08293__A2 _08358_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input91_I spimemio_flash_io2_oeb VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11346__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09216_ _09220_/A2 _11425_/Q _09217_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06772__I _07110_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06428_ _05723_/Z _11347_/Q _06432_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06359_ _08825_/A1 _11232_/Q _06217_/Z _06360_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08045__A2 _07513_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09147_ _09147_/I _11403_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09242__A1 _09246_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06056__A1 _06056_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06056__B2 _06056_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10927__A2 _10880_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09078_ _09078_/I _11382_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11496__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output178_I _06056_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08029_ _08562_/A1 _07885_/I _08563_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05803__A1 _06217_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07556__A1 _08589_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11040_ _11050_/I _11687_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07020__A3 _06871_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07108__I _07110_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11592__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11344__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10824_ _10914_/A1 _11602_/Q _10825_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08808__A1 _06851_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09481__A1 _09497_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10755_ _10755_/A1 _10755_/A2 _10755_/A3 _10755_/A4 _10780_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__10615__B2 _10615_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06295__A1 _08940_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10686_ _10905_/A1 _11535_/Q _10688_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09233__A1 _09154_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07795__A1 _08592_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput309 _06725_/Z spimemio_flash_io1_di VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_11307_ _11307_/D _11686_/RN _06705_/Z _11307_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_99_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11238_ _11238_/D _11686_/RN _06705_/Z _11238_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_11169_ _11169_/D _11686_/RN _06705_/Z _11169_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__10146__A3 _09876_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11583__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11219__CLK _11666_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05730_ _10272_/A2 _05991_/I _05730_/B _05731_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05661_ _05660_/Z _11626_/Q _05662_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10854__A1 _10900_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11335__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11267__CLKN input68/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08380_ _08383_/A1 _08355_/I _08380_/B _08648_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07400_ _07076_/Z _07403_/A2 _07400_/B _07401_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_90_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11369__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05876__A4 _05876_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05592_ _06466_/B _11062_/Q _05593_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10606__A1 _10922_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07331_ _07331_/I _11214_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09472__A1 _09270_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07262_ _06863_/Z _07265_/A2 _07262_/B _07263_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07193_ _07193_/I _11179_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06213_ _08795_/A1 _06217_/I _06213_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09001_ _06851_/Z _09013_/A2 _09001_/B _09002_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09224__A1 _09116_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06144_ _06324_/A1 _11589_/Q _06146_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09775__A2 _09015_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07786__A1 _08696_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06075_ _11390_/Q _10613_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09903_ _09903_/A1 _09935_/B _10265_/A3 _09922_/B _11635_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09834_ _09834_/I _11621_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06210__A1 _05703_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11574__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09765_ _09765_/I _11599_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06977_ _06977_/A1 _06977_/A2 _11121_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05928_ input49/Z _05927_/Z _07201_/A1 input57/Z _05933_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09696_ _09697_/A2 _11578_/Q _09697_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08716_ _11050_/I _11268_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06767__I _07110_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08647_ _08647_/I _08648_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10845__A1 _10891_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_05859_ _11393_/Q _09091_/A1 _11385_/Q _09066_/A1 _05859_/C _05860_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XPHY_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_08578_ _08486_/Z _08578_/A2 _08622_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09463__A1 _09158_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07529_ _06587_/I _07999_/A2 _07471_/B _07530_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XANTENNA__07069__A3 _06871_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10540_ _10902_/B2 _11516_/Q _10542_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06277__A1 _06785_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08018__A2 _08632_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10471_ _10471_/A1 _10406_/I _10887_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__06029__A1 _06029_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09518__A2 _11521_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11023_ _07300_/B _11023_/A2 _11023_/B _11024_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06201__A1 _09674_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11511__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11317__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11083__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09454__A1 _09121_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10807_ _10899_/A1 _11506_/Q _10809_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08257__A2 _07566_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11661__CLK _11663_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10738_ _10921_/A1 _11336_/Q _10742_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_158_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08009__A2 _08632_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11013__A1 _10966_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10669_ _10883_/A1 _11375_/Q _10671_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07768__A1 _08328_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09509__A2 _11518_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06440__A1 _10935_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06900_ _06900_/I _11099_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07880_ _07880_/A1 _07872_/I _07988_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08193__A1 _07297_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06743__A2 input1/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06831_ _06831_/I _11077_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09550_ _09572_/A2 _11531_/Q _09551_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06762_ _06701_/I _11686_/RN _06763_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11191__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05491__I input58/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05713_ _11586_/Q _09699_/A1 _11578_/Q _09674_/A1 _05713_/C _05714_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_09481_ _09497_/A2 _11509_/Q _09482_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08501_ _07572_/I _07727_/I _08637_/B _08502_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10827__A1 _10922_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11308__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08432_ _08449_/A1 _08442_/A1 _08557_/B _08433_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09693__A1 _09697_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_464 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06693_ _06693_/I _06693_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05644_ _05644_/A1 _05598_/I _05645_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08363_ _08548_/A3 _08363_/A2 _08435_/A1 _08653_/A2 _08363_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__08248__A2 _07609_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05575_ _05575_/A1 _11069_/Q _06456_/A2 _06510_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_08294_ _08395_/A2 _08345_/A2 _08294_/B _08294_/C _08295_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_07314_ _10938_/A1 _07326_/A2 _07316_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07245_ _07245_/I _11189_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11604__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11004__A1 _08431_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09748__A2 _09725_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07176_ _07197_/A1 _11176_/Q _07177_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06127_ _11389_/Q _09091_/A1 _11381_/Q _09066_/A1 _06127_/C _06128_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__11619__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_391 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06058_ _06058_/A1 _06058_/A2 _06058_/A3 _06058_/A4 _06099_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA_input54_I mgmt_gpio_in[26] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06982__A2 _06974_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11534__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08184__A1 _08490_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09817_ _09187_/I _09823_/A2 _09817_/B _09818_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_143_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09748_ _09270_/Z _09725_/Z _09748_/B _09749_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10818__A1 _10910_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output210_I _10613_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09684__A1 _09697_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09679_ _09121_/I _09697_/A2 _09679_/B _09680_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11684__CLK _06687_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output308_I _06723_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_464 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_146_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11641_ _11641_/D _11686_/RN _11666_/CLK _11641_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_14_147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11572_ _11572_/D _11686_/RN _06705_/Z _11572_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__10046__A2 _10046_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10523_ _10899_/A1 _11500_/Q _10527_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput19 mask_rev_in[23] input19/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09739__A2 _09725_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10454_ _10484_/A1 _10406_/I _10920_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__11064__CLK input68/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08411__A2 _08411_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10385_ _10385_/A1 _10880_/C _10385_/B _10386_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10754__B1 _10913_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06422__A1 _09066_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06973__A2 input162/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11538__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11006_ _10966_/Z _11006_/A2 _11007_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09911__A2 _09935_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09675__A1 _09697_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07150__A2 _09270_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_253 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10037__A2 _09973_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11407__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06661__A1 _11059_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07030_ _07030_/I _11137_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11557__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06964__A2 _06941_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08981_ _08988_/A2 _11352_/Q _08982_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07932_ _07932_/A1 _07932_/A2 _07937_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07863_ _07863_/I _07864_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11529__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06814_ _11679_/Q _11000_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09602_ _09602_/I _11547_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07913__A1 split15/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06716__A2 input87/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09533_ _09533_/I _11525_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07794_ _08639_/B _08509_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09666__A1 _09187_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06745_ _11307_/Q input71/Z _06746_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09464_ _09464_/I _11503_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06676_ _06701_/I _11689_/Q _06677_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07141__A2 _05927_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09418__A1 _09422_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09395_ _09395_/I _11481_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08415_ split15/Z _08417_/A2 _08415_/B _08535_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05627_ _11066_/Q _06474_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_24_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_08346_ _08346_/I _08348_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_11_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10028__A2 _09878_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05558_ _05558_/I _11694_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11087__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08277_ _08419_/B _08279_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07228_ _11320_/Q _05924_/Z _07228_/B _07230_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_152_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07159_ _05925_/Z _09116_/I _07160_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10200__A2 _10355_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10170_ _10361_/A1 _11423_/Q _10171_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08157__A1 split8/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09657__A1 _09125_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08656__B _08656_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09409__A1 _09422_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07132__A2 _07151_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_11624_ _11624_/D _11686_/RN _06705_/Z _11624_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_1176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05694__A2 _11530_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11555_ _11555_/D _11686_/RN _06705_/Z _11555_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__08632__A2 _08632_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11486_ _11486_/D _11686_/RN _06705_/Z _11486_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10506_ _10506_/A1 _10506_/A2 _10507_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10437_ _10460_/A1 _10460_/A3 _10478_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__07199__A2 _06701_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_916 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_10368_ _10368_/A1 _10368_/A2 _10368_/A3 _10381_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_69_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10299_ _10377_/A1 _11578_/Q _10377_/B1 _11570_/Q _10302_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_949 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_938 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_927 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08699__A2 _08036_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06530_ _08431_/B _08672_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__10387__I _10387_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06461_ _06461_/A1 _06610_/A3 _06479_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__09241__I _09241_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08320__A1 _08686_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08200_ split7/I _08232_/A2 _08200_/B _08464_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06392_ _06392_/A1 _06392_/A2 _06392_/A3 _06392_/A4 _06392_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_09180_ _09180_/I _11413_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08131_ _08142_/A2 _08169_/A2 _08134_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08623__A2 _08623_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09820__A1 _09241_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06634__A1 input77/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08062_ _08205_/C _08332_/A1 _08063_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10430__A2 _09912_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07013_ _07013_/A1 _06904_/Z _07018_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input156_I wb_dat_i[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08964_ _08964_/I _11346_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07915_ _07926_/I _08361_/B _07916_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08139__A1 _08656_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08895_ _07431_/Z _08913_/A2 _08895_/B _08896_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07846_ _07846_/A1 _07870_/A3 split16/I _07847_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__06165__A3 _06165_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_356 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07777_ _07777_/A1 _07777_/A2 _07783_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input17_I mask_rev_in[21] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09516_ _09187_/Z _09522_/A2 _09516_/B _09517_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06775__I _07110_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06728_ _11382_/Q _10137_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09447_ _09270_/Z _09447_/A2 _09447_/B _09448_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_06659_ _11173_/Q _06661_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05676__A2 _05805_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09378_ _09397_/A2 _11476_/Q _09379_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09811__A1 _09154_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08614__A2 _08614_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08329_ _08332_/A1 _08417_/A2 _08329_/B _08511_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10421__A2 _10427_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11340_ _11340_/D _11686_/RN _06705_/Z _11340_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__08378__A1 split8/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11271_ _11271_/D input76/Z _06705_/Z _11271_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10222_ _10373_/A1 _11520_/Q _10373_/B1 _11528_/Q _10225_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07050__A1 _06837_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10153_ _10153_/A1 _10382_/A2 _10153_/B _10153_/C _10155_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__11420__SETN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11102__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10084_ _10084_/A1 _10084_/A2 _10084_/A3 _10084_/A4 _10085_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_47_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10488__A2 _11619_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11435__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11252__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06685__I _06685_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10986_ _10986_/A1 _10966_/Z _10986_/B _10987_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09996__I _09996_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06864__A1 _06869_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11607_ _11607_/D _11686_/RN _06705_/Z _11607_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__09802__A1 _09116_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08605__A2 _07844_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06616__A1 _06616_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11538_ _11538_/D _11686_/RN _06705_/Z _11538_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_116_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11469_ _11469_/D _11686_/RN _06705_/Z _11469_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_143_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08369__A1 split8/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10176__A1 _10366_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09030__A2 _09039_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06919__A2 _11033_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07041__A1 _07412_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_713 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_746 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input9_I mask_rev_in[14] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06395__A3 _08719_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07700_ _07700_/I _08394_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_05961_ _08799_/A1 _11033_/A2 _05962_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09869__A1 _09927_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08680_ _08680_/A1 _08680_/A2 _08691_/A2 _08681_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05892_ _11457_/Q _09299_/A1 _11449_/Q _09274_/A1 _05892_/C _05893_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_07631_ _07631_/A1 _07631_/A2 _07631_/A3 _08271_/B _07634_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_26_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_07562_ _07562_/I _08248_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09301_ _09116_/Z _09322_/A2 _09301_/B _09302_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06513_ _11056_/Q _06514_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07493_ _08519_/A2 _08358_/A2 _07494_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10100__A1 _10357_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06444_ _06444_/A1 _06446_/I _06444_/B _06445_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10651__A2 _11326_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09232_ _09246_/A2 _11430_/Q _09233_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06375_ _06375_/A1 _06375_/A2 _06375_/A3 _06391_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09163_ _06859_/Z _09169_/A2 _09163_/B _09164_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08114_ _08114_/A1 split16/Z _08142_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10403__A2 _10406_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09094_ _09094_/I _11387_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08045_ _08054_/A1 _07513_/I _08045_/A3 _08048_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__07280__A1 _07290_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11125__CLK _11672_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09021__A2 _09039_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05830__A2 _05969_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07032__A1 _06843_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09996_ _09996_/I _10000_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08780__A1 _08784_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11275__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08947_ _08963_/A2 _11341_/Q _08948_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08878_ _08888_/A2 _11319_/Q _08879_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07829_ _08341_/B _08632_/A2 _07831_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07335__A2 _06904_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10840_ _11137_/Q _10888_/A1 _11135_/Q _10889_/A1 _10840_/C _10844_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
Xsplit13 split13/I split13/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10771_ _10771_/A1 _10771_/A2 _10771_/A3 _10771_/A4 _10780_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__07099__A1 _07099_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10642__A2 _10642_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07271__A1 _07290_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11323_ _11323_/D _11686_/RN _06705_/Z _11323_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_11254_ _11254_/D input162/Z _06687_/A2 _11254_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__05821__A2 _11434_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11618__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10205_ _10360_/A1 _11432_/Q _10207_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08771__A1 _08784_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11185_ _11185_/D input76/Z _06705_/Z _11185_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__05584__I _05584_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10173__A4 _10173_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10136_ _11398_/Q _10359_/A2 _11390_/Q _10359_/B2 _10136_/C _10143_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_10067_ _10067_/A1 _10067_/A2 _10067_/A3 _10067_/A4 _10085_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__08523__A1 _07844_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10330__B2 _11252_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09079__A2 _11383_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05888__A2 _09144_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11389__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10969_ _08431_/B input160/Z _08460_/B input137/Z _10970_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08826__A2 _07114_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11148__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10397__A1 _10433_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06160_ _11421_/Q _09197_/A1 _11413_/Q _09171_/A1 _06160_/C _06165_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__07262__A1 _06863_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06065__A2 _09800_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06091_ _08915_/A1 _11334_/Q _06092_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10149__B2 _10371_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11298__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07565__A2 _08339_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09850_ _09945_/A2 _10092_/I _09939_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08762__A1 _08784_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_532 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06368__A3 _06217_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09781_ _09781_/I _11604_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06993_ _06974_/I _11127_/Q _06994_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_08801_ _08801_/A1 _08827_/A2 _08801_/B _08802_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08732_ _08732_/I _11274_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05944_ _11655_/Q _10385_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_08663_ _08355_/I _08280_/B _08663_/B _08664_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05875_ input70/Z _05924_/I _05925_/I input41/Z _05876_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07614_ _07614_/A1 split16/Z _07640_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08594_ _08690_/A1 _08638_/A1 _08679_/A2 _08640_/A1 _08594_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_121_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input119_I wb_adr_i[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07545_ _08046_/B split16/Z _07601_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08817__A2 _08820_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07476_ input112/Z input111/Z _07477_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10624__A2 _11446_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08293__A3 _08677_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09215_ _09215_/I _11424_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06427_ _06427_/A1 _06427_/A2 _06427_/A3 _06438_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_input84_I spimemio_flash_clk VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06358_ _07419_/A2 _11228_/Q _06217_/Z _06360_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09146_ _09116_/Z _09169_/A2 _09146_/B _09147_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09242__A2 _11433_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07253__A1 _06851_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09077_ _06851_/Z _09089_/A2 _09077_/B _09078_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06289_ _09041_/A1 _11372_/Q _06291_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08028_ _08395_/B _08677_/A2 _08459_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05803__A2 _05803_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05567__A1 _05519_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09979_ _09979_/A1 _10040_/A2 _09980_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06359__A3 _06217_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08753__A1 _06851_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10560__A1 _10560_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08505__A1 _08696_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10312__B2 _10351_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10823_ _10914_/B1 _11610_/Q _10825_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08808__A2 _08820_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10076__B1 _10373_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10615__A2 _10615_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10754_ _11585_/Q _10913_/B2 _10913_/A2 _11593_/Q _10755_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_10685_ _10903_/A1 _11559_/Q _10690_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10379__A1 _10379_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09233__A2 _09246_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07244__A1 _07076_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11440__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07794__I _08639_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11306_ _11306_/D _11686_/RN _06705_/Z _11306_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__08992__A1 _07426_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11280__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11237_ _11237_/D _11686_/RN _06705_/Z _11237_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_11168_ _11168_/D _11686_/RN _06705_/Z _11168_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__11590__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08744__A1 _07426_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10153__C _10153_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10119_ _10119_/A1 _10119_/A2 _10119_/A3 _10124_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_121_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11099_ _11099_/D _11686_/RN _06705_/Z _11099_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__10303__A1 _10303_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05660_ _05660_/I _05660_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_05591_ _11061_/Q _06498_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07330_ _10954_/A1 _07310_/I _07330_/B _07331_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_91_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09472__A2 _09472_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11099__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07261_ _07265_/A2 _11195_/Q _07262_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09000_ _09013_/A2 _11358_/Q _09001_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07192_ _07197_/A1 _07192_/A2 _07192_/B _07193_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06212_ _06212_/A1 _06212_/A2 _06212_/A3 _06212_/A4 _06259_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__09224__A2 _09246_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06143_ _09800_/A1 _11613_/Q _06146_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07235__A1 _07240_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05797__A1 _06238_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06074_ _06074_/A1 _06074_/A2 _06074_/A3 _06099_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11271__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09902_ _09902_/I _09922_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
X_09833_ _09125_/I _09848_/A2 _09833_/B _09834_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07538__A2 _08592_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_09764_ _09158_/I _09773_/A2 _09764_/B _09765_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06976_ _06974_/I _11121_/Q _06977_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_395 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_05927_ _05927_/I _05927_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_09695_ _09695_/I _11577_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xrebuffer20 _08063_/A2 _08202_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlya_2
XANTENNA__06269__B _06269_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08715_ _11050_/I _11267_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11313__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08646_ _08646_/A1 _08646_/A2 _08646_/A3 _11258_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09160__A1 _09158_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05858_ _05858_/A1 _05858_/A2 _05859_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_05789_ _11490_/Q _09399_/A1 _11482_/Q _09374_/A1 _05789_/C _05827_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_08577_ _08662_/A1 _08577_/A2 _08697_/A3 _08579_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09463__A2 _09472_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07528_ _08400_/B _08400_/C _08294_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_07459_ _07996_/A2 _07445_/I split5/I _07471_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__11463__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06277__A2 _11072_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10470_ _10887_/B1 _11427_/Q _10477_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09129_ _09142_/A2 _11398_/Q _09130_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11262__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10781__A1 _10919_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11022_ _11022_/I _11682_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10533__A1 _10906_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09151__A1 _09169_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07701__A2 _08394_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_284 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09454__A2 _09472_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10806_ _10806_/A1 _10806_/A2 _10806_/A3 _10806_/A4 _10826_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_32_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06693__I _06693_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10737_ _10737_/A1 _10737_/A2 _10737_/A3 _10737_/A4 _10744_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__06268__A2 _11305_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07217__A1 _05924_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10668_ _10886_/B2 _11391_/Q _10886_/A2 _11399_/Q _10671_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_10599_ _10905_/A1 _11533_/Q _10603_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08965__A1 _05723_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10772__A1 _10904_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11253__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06440__A2 _05969_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08193__A2 _11254_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10524__A1 _10894_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09390__A1 _09397_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11336__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06830_ _06835_/A1 _09241_/I _06830_/B _06831_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06761_ _06761_/I _11218_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05951__A1 _08761_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05712_ _05712_/A1 _05712_/A2 _05713_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09480_ _09480_/I _11508_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08500_ _08509_/A1 _08587_/B _08500_/B _08500_/C _08636_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__09142__A1 _06867_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06692_ _11306_/Q _06692_/A2 _06692_/B _06693_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05643_ input71/Z _05924_/I _05925_/I input42/Z _05662_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08431_ _08431_/A1 _08431_/A2 _08431_/B _08522_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11486__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08362_ _08656_/A1 _08361_/B split15/I _08549_/A1 _08653_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05574_ _05574_/I _11690_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08293_ _08294_/B _08358_/A2 _08677_/A2 _08430_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_07313_ _07313_/A1 _07313_/A2 _11208_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07244_ _07076_/Z _07265_/A2 _07244_/B _07245_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07175_ _11200_/Q _05925_/Z _07175_/B _07177_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_253 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11244__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08956__A1 _08963_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06126_ _06126_/A1 _06126_/A2 _06127_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06057_ _11454_/Q _09299_/A1 _11446_/Q _09274_/A1 _06057_/C _06058_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA_input47_I mgmt_gpio_in[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_289 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10515__A1 _10914_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09381__A1 _09397_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09816_ _09823_/A2 _11616_/Q _09817_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06195__A1 _09624_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09154__I _09154_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06778__I _07110_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09747_ _09725_/Z _11594_/Q _09748_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06959_ _06959_/A1 _06959_/A2 _11116_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05942__A1 _08839_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09133__A1 _06855_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09678_ _09697_/A2 _11572_/Q _09679_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07695__A1 _07691_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08629_ _08688_/A2 _08665_/A2 _08629_/A3 _08664_/A1 _08631_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_42_435 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11640_ _11640_/D _11686_/RN _11666_/CLK _11640_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_11571_ _11571_/D _11686_/RN _06705_/Z _11571_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_52_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10522_ _10522_/A1 _10522_/A2 _10522_/A3 _10522_/A4 _10548_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_10_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11209__CLK _11656_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10453_ _10453_/I _10920_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XANTENNA__10754__A1 _11585_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10384_ _10384_/A1 _06556_/I _10926_/C _10384_/C _10385_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08947__A1 _08963_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11266__CLKN input68/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11235__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06422__A2 _11379_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05630__B1 _05633_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11359__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09372__A1 _09270_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08175__A2 _07492_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10506__A1 _10506_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11005_ _11005_/A1 _11005_/A2 _11005_/A3 _11006_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__05933__A1 _05933_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05528__A4 _06491_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06489__A2 _06491_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10993__A1 _10993_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11474__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06110__A1 _08839_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06661__A2 _06661_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08938__A1 _06867_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11226__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10745__A1 _10092_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08980_ _08980_/I _11351_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07931_ split6/I _08607_/B _07932_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07862_ _07874_/A1 _07862_/A2 _07880_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09363__A1 _09158_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08166__A2 _07535_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06177__A1 _08825_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09601_ _09116_/Z _09622_/A2 _09601_/B _09602_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06813_ _06813_/I _11074_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09532_ _09125_/Z _09547_/A2 _09532_/B _09533_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07793_ _07793_/A1 _07793_/A2 _08639_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__09666__A2 _09672_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06744_ _06744_/I _06744_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09463_ _09158_/Z _09472_/A2 _09463_/B _09464_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06675_ _06675_/I _06675_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_435 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09394_ _09241_/Z _09397_/A2 _09394_/B _09395_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08414_ _08414_/A1 _08687_/A3 _08414_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_05626_ _05626_/I _05718_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA_input101_I wb_adr_i[13] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09418__A2 _11489_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08345_ _08490_/A3 _08345_/A2 _08519_/B _08346_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05557_ _05557_/A1 _05519_/I _05557_/B _05558_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07429__A1 _07426_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11465__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08276_ split14/Z _07609_/Z _08276_/B _08419_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07227_ _05924_/Z _09187_/I _07228_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06652__A2 _06652_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11501__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07158_ _07201_/A1 _05925_/Z _07158_/B _09015_/I _07197_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XANTENNA__08929__A1 _06855_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11217__RN input162/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06109_ _11275_/Q _08726_/A1 _08742_/A1 _11280_/Q _06114_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06404__A2 _11273_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07089_ _07090_/A2 _11154_/Q _07090_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11082__SETN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09354__A1 _09121_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11651__CLK _11665_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05915__A1 _09144_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09657__A2 _09672_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_11623_ _11623_/D _11686_/RN _06705_/Z _11623_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__06340__A1 _05703_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09409__A2 _11486_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08672__B _08672_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11554_ _11554_/D _11686_/RN _06705_/Z _11554_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__11456__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10975__A1 _08493_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11485_ _11485_/D _11686_/RN _06705_/Z _11485_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_10505_ _10905_/A1 _11531_/Q _10509_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10436_ _10913_/B2 _11579_/Q _10442_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11181__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09593__A1 _09597_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10727__A1 _10900_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_917 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_906 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_10367_ _10367_/A1 _11241_/Q _10368_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10298_ _10298_/A1 _10298_/A2 _10298_/A3 _10303_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_939 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_928 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11603__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06460_ _06460_/A1 _06619_/A1 _06466_/B _06461_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06331__A1 _09549_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08130_ _08130_/A1 _08224_/B _08475_/A2 _08130_/A4 _08133_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_06391_ _06391_/A1 _06391_/A2 _06391_/A3 _06391_/A4 _06392_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__11524__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11447__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06634__A2 input93/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09820__A2 _09823_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08061_ _08467_/B _08205_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_07012_ _07012_/I _11132_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09584__A1 _09597_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10718__A1 _10891_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11674__CLK _11683_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08963_ _06867_/Z _08963_/A2 _08963_/B _08964_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input149_I wb_dat_i[27] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07914_ split21/I _08361_/B _08435_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08894_ _08913_/A2 _11324_/Q _08895_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07898__A1 _07685_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07845_ _07845_/A1 _07845_/A2 _08037_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07776_ _07722_/I _07508_/I _07777_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09515_ _09522_/A2 _11520_/Q _09516_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06727_ _11358_/Q _06727_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08311__A2 _08411_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09446_ _09447_/A2 _11498_/Q _09447_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_249 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11686__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06322__A1 _07398_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06658_ _06658_/A1 _06658_/A2 _06658_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06589_ _06589_/A1 _08006_/A2 _08005_/A2 _06588_/Z _06600_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_09377_ _09377_/I _11475_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05609_ _05609_/A1 _06497_/A3 _05633_/B _05609_/B2 _05610_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06873__A2 _11087_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_165_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08075__A1 split12/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08328_ _07593_/I _08329_/B _08328_/B1 _08509_/A2 _08596_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10957__A1 _10957_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09811__A2 _09823_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08259_ _08259_/A1 _08530_/I _08406_/A1 _08668_/I _08263_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__11438__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output270_I _11278_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09575__A1 _09597_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11270_ _11270_/D _11270_/RN input68/Z _11270_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
X_10221_ _10221_/A1 _10221_/A2 _10221_/A3 _10226_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__06389__A1 _08825_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10152_ _10152_/A1 _10152_/A2 _10152_/A3 _10152_/A4 _10153_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__11610__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10083_ _10083_/A1 _10083_/A2 _10083_/A3 _10084_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xoutput290 _11088_/Q pll_trim[25] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_47_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10985_ _10966_/Z _10985_/A2 _10986_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11677__RN input162/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11547__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11606_ _11606_/D _11686_/RN _06705_/Z _11606_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_11537_ _11537_/D _11686_/RN _06705_/Z _11537_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__09802__A2 _09823_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11697__CLK input68/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10948__A1 _10934_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11468_ _11468_/D _11686_/RN _06705_/Z _11468_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__09566__A1 _09187_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10419_ _10463_/A1 _09934_/I _10916_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_11399_ _11399_/D _11686_/RN _06705_/Z _11399_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__06919__A3 _06871_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07041__A2 _06217_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_714 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11601__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_05960_ _06398_/A2 input25/Z _05962_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05891_ _05891_/A1 _05891_/A2 _05892_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11077__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07630_ _08415_/B _08509_/A1 _08271_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07561_ _07607_/A1 _07649_/A2 _07562_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11557__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09300_ _09322_/A2 _11451_/Q _09301_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06512_ _11163_/Q _06610_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07492_ _07492_/I _08519_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__10100__A2 _11413_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06304__A1 _10938_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06443_ _06446_/I _11701_/Q _11172_/Q _06444_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09231_ _09231_/I _11429_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06374_ _09449_/A1 _11499_/Q _06375_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09162_ _09169_/A2 _11408_/Q _09163_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07804__A1 _08592_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08113_ _08113_/A1 _08212_/B _08470_/A2 _08113_/A4 _08117_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__10939__A1 _10934_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06607__A2 _11302_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09093_ _07426_/Z _09114_/A2 _09093_/B _09094_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08044_ _08162_/A1 _08167_/A1 _08251_/A2 _08063_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__09557__A1 _09125_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09995_ _10034_/A1 _09899_/I _09996_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__06791__A1 _06835_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08946_ _08946_/I _11340_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08877_ _08877_/I _11318_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07828_ _07828_/I _08632_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_17_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07759_ _07759_/A1 _08305_/B _07766_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xsplit14 split21/Z split14/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_10770_ _11457_/Q _10897_/A2 _10897_/B1 _11465_/Q _10771_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07099__A2 _06904_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11659__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09429_ _09121_/Z _09447_/A2 _09429_/B _09430_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10642__A3 _10427_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11322_ _11322_/D input76/Z _06705_/Z _11322_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_11253_ _11253_/D _11686_/RN _06705_/Z _11253_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_106_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10204_ _11400_/Q _10359_/A2 _11392_/Q _10359_/B2 _10204_/C _10209_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_11184_ _11184_/D input76/Z _06705_/Z _11184_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10135_ _10135_/A1 _10615_/A2 _09887_/I _10615_/B2 _10019_/I _10136_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_85_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10066_ _11444_/Q _10363_/A2 _11436_/Q _10363_/B2 _10066_/C _10067_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__10330__A2 _10369_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10968_ _08493_/B input146/Z _10970_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10094__A1 _11349_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10094__B2 _10351_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10899_ _10899_/A1 _11253_/Q _10901_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10397__A2 _10406_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07262__A2 _07265_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06090_ _08890_/A1 _11326_/Q _06092_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10149__A2 _10370_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_500 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_533 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_08800_ _08801_/A1 _11295_/Q _06904_/Z _08801_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__07990__I _07990_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09780_ _09121_/I _09798_/A2 _09780_/B _09781_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06992_ _06992_/A1 _06992_/A2 _11126_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08762__A2 _11284_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_08731_ _07431_/Z _08740_/A2 _08731_/B _08732_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05943_ _05943_/I _08742_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_577 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_08662_ _08662_/A1 _08662_/A2 _08662_/A3 _08673_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05874_ input50/Z _05927_/I _07201_/A1 input59/Z _05876_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07613_ _07613_/A1 _07613_/A2 _08411_/A2 _08265_/B _07619_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__06525__A1 input67/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08593_ _08593_/A1 _08593_/A2 _08593_/A3 _08593_/A4 _08640_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__10872__A3 _10872_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07544_ _07544_/A1 _07544_/A2 _07574_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08278__A1 _08400_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07475_ _07689_/A1 _06587_/I _07479_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06828__A2 _05633_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09214_ _09187_/Z _09220_/A2 _09214_/B _09215_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06426_ _08940_/A1 _11339_/Q _06427_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06357_ _09274_/A1 _11443_/Q _06360_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09145_ _09169_/A2 _11403_/Q _09146_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07253__A2 _07265_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09076_ _09089_/A2 _11382_/Q _09077_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input77_I qspi_enabled VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06288_ _09016_/A1 _11364_/Q _06966_/A1 _11120_/Q _06291_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08027_ _08033_/B _08395_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11242__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09978_ _10378_/A1 _11547_/Q _09983_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08753__A2 _08759_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11392__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10560__A2 _06556_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08929_ _06855_/Z _08938_/A2 _08929_/B _08930_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08505__A2 _08509_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10312__A2 _10351_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10822_ _10915_/A1 _11618_/Q _10916_/A1 _11626_/Q _10825_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_10753_ _10911_/A1 _11577_/Q _10755_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10076__B2 _11524_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10076__A1 _10373_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10684_ _10904_/A1 _11551_/Q _10690_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09769__A1 _09773_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07244__A2 _07265_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11305_ _11305_/D _11686_/RN _06705_/Z _11305_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__08992__A2 _09013_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11236_ _11236_/D _11686_/RN _06705_/Z _11236_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_11167_ _11167_/D _11686_/RN _06705_/Z _11167_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__08744__A2 _08759_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10118_ _10374_/A1 _11533_/Q _10119_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11098_ _11098_/D _11686_/RN _06705_/Z _11098_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10049_ _10086_/A1 _10880_/C _10049_/B _10050_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05590_ _05590_/I _05644_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11115__CLK _11672_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07260_ _07260_/I _11194_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07191_ _07197_/A1 _11179_/Q _07192_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06211_ _06211_/A1 _06211_/A2 _06211_/A3 _06211_/A4 _06212_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_06142_ _09775_/A1 _11605_/Q _06146_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08432__A1 _08449_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06073_ _11582_/Q _09699_/A1 _09674_/A1 _11574_/Q _06074_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__05797__A2 _08799_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06994__A1 _10954_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09901_ _09986_/I _09901_/A2 _09903_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09832_ _09848_/A2 _11621_/Q _09833_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05549__A2 _05519_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09763_ _09773_/A2 _11599_/Q _09764_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06210__A3 _07370_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_06975_ _10935_/A1 _06990_/A2 _06977_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input131_I wb_dat_i[10] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_08714_ _11050_/I _11266_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09694_ _09241_/Z _09697_/A2 _09694_/B _09695_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xrebuffer10 _08478_/A1 _08481_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlya_1
X_05926_ input69/Z _05924_/Z _05925_/Z input40/Z _05933_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08645_ _08645_/A1 _11221_/Q _11016_/A1 _08646_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__07171__A1 _07197_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09160__A2 _09169_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05857_ _09041_/A1 _11377_/Q _05858_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08576_ _08576_/A1 _08576_/A2 _08576_/A3 _08697_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XPHY_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_05788_ _05788_/A1 _05788_/A2 _05789_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09999__A1 _10369_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07527_ _07527_/I _08400_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10058__B2 _10355_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11608__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07458_ _07472_/A2 _07999_/A2 _07689_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07389_ _07081_/Z _07389_/A2 _07389_/B _07390_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11373__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06409_ _08795_/A1 _08799_/A1 _06408_/Z _06413_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09128_ _09128_/I _11397_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06985__A1 _10945_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09059_ _09059_/I _11376_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11388__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11021_ _11019_/Z _11021_/A2 _11022_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07844__B _07844_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08726__A2 _06904_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11138__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10297__A1 _10374_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07162__A1 _07197_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09151__A2 _11405_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06974__I _06974_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11326__SETN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10805_ _11458_/Q _10897_/A2 _10897_/B1 _11466_/Q _10806_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11288__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10736_ _10736_/A1 _10736_/A2 _10736_/A3 _10736_/A4 _10737_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_13_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10667_ _11415_/Q _10888_/A1 _11407_/Q _10889_/A1 _10667_/C _10671_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__07217__A2 _09154_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10598_ _10598_/A1 _10598_/A2 _10598_/A3 _10598_/A4 _10604_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__06976__A1 _06974_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08965__A2 _06838_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11219_ _11219_/D input162/Z _11666_/CLK _11219_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__09390__A2 _11480_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06760_ _06760_/A1 _08672_/B _06761_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10288__A1 _10366_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05711_ _09624_/A1 _11562_/Q _05712_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09142__A2 _09142_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06691_ _11306_/Q input94/Z _06692_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08430_ _08430_/A1 _08430_/A2 _08430_/A3 _08430_/A4 _08431_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_05642_ _05642_/I _05925_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
X_08361_ _08383_/A1 _08355_/I _08361_/B _08435_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05573_ _06610_/A2 _05572_/B _05573_/B _05574_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06259__A3 _06259_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08292_ _08292_/A1 _08292_/A2 _08541_/A3 _08292_/A4 _08295_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_07312_ _07310_/I _11208_/Q _07313_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_176_143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07243_ _07265_/A2 _11189_/Q _07244_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07208__A2 _05924_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10212__A1 _10366_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07174_ _05925_/Z _09154_/I _07175_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06125_ _09016_/A1 _11365_/Q _06126_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06056_ _06056_/A1 _05823_/I _05820_/I _06056_/B2 _06057_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__08708__A2 _11262_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09905__A1 _09922_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09815_ _09815_/I _11615_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06719__A1 _06753_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_355 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09381__A2 _11477_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09746_ _09746_/I _11593_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06958_ _06941_/I _11116_/Q _06959_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05909_ _05909_/A1 _05909_/A2 _05910_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09677_ _09677_/I _11571_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09133__A2 _09142_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05942__A2 _07370_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10279__A1 _10357_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06889_ _06902_/A2 _11096_/Q _06890_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08495__B _08495_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08628_ _08355_/I _08276_/B _08628_/B _08628_/C _08664_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_42_403 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11430__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08892__A1 _07426_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_285 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08559_ _08559_/A1 _08559_/A2 _08693_/A3 _08561_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11180__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11570_ _11570_/D _11686_/RN _06705_/Z _11570_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__11580__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10521_ _10913_/B2 _11580_/Q _10522_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10451__A1 _10514_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10452_ _10452_/A1 _10506_/A2 _10453_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06958__A1 _06941_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10383_ _10383_/A1 _06556_/I _10384_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10754__A2 _10913_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11004_ _08431_/B input134/Z _08460_/B input143/Z _11005_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10506__A2 _10506_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09372__A2 _09372_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07135__A1 _05927_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07686__A2 _07455_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11171__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08635__A1 _07844_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10719_ _10892_/A1 _11472_/Q _10720_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10993__A2 _10966_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11699_ _11699_/D _11699_/RN input68/Z _11699_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__06110__A2 _08795_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer1 _07870_/A3 _07669_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06949__A1 _10942_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09060__A1 _09064_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08938__A2 _08938_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07610__A2 _07609_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11303__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07930_ _07930_/A1 _07964_/A2 _08607_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_322 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07861_ _07861_/A1 _07999_/A2 _07862_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09363__A2 _09372_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11453__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06177__A2 _11033_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07792_ _08328_/B1 _08592_/B _08325_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09600_ _09622_/A2 _11547_/Q _09601_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06812_ _06835_/A1 _09154_/I _06812_/B _06813_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09531_ _09547_/A2 _11525_/Q _09532_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06743_ input36/Z input1/Z _06744_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09462_ _09472_/A2 _11503_/Q _09463_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07503__I split16/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06674_ _06674_/A1 input1/Z _06674_/B _06675_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09393_ _09397_/A2 _11481_/Q _09394_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10681__A1 _10900_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05688__A1 _05703_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08413_ _07616_/I _08419_/A1 _08413_/B _08413_/C _08687_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05625_ _05802_/A2 _05684_/A2 _05626_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08344_ _08344_/I _08348_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05556_ _05519_/I _11694_/Q _05557_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_177_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10433__A1 _10433_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08275_ _08400_/A1 _08537_/B _08275_/B _08538_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06101__A2 _05969_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07226_ _07226_/I _11185_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07157_ _07114_/B _07267_/A1 _07158_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05860__A1 _05860_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08929__A2 _08938_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09051__A1 _09064_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06108_ input22/Z _06398_/A2 _08799_/A1 _06108_/B2 _06108_/C _06128_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_07088_ _07088_/I _11153_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06039_ _10947_/A1 _06304_/A2 _06619_/B _06039_/C _06040_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__09354__A2 _09372_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07365__A1 _07076_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06168__A2 _05969_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09729_ _09725_/Z _11588_/Q _09730_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05915__A2 _11408_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08865__A1 _08865_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1145 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10672__A1 _10891_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11153__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_11622_ _11622_/D _11686_/RN _06705_/Z _11622_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__06340__A2 _08825_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11553_ _11553_/D _11686_/RN _06705_/Z _11553_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_11484_ _11484_/D _11686_/RN _06705_/Z _11484_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_10504_ _10504_/I _10905_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__11326__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10435_ _10480_/A1 _09934_/I _10913_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__09042__A1 _09064_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09593__A2 _11545_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11476__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_907 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_10366_ _10366_/A1 _11237_/Q _10368_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10297_ _10374_/A1 _11538_/Q _10298_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_929 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_918 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07356__A1 _08825_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11392__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10112__B1 _10369_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_285 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08856__A1 _08863_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11144__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06390_ _06390_/A1 _06390_/A2 _06390_/A3 _06390_/A4 _06391_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_14_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08060_ _08169_/A1 _08142_/A1 _08467_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_119_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07011_ _06843_/Z _07011_/A2 _07011_/B _07012_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05842__A1 _06839_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09033__A1 _06859_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10718__A2 _11480_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08962_ _08963_/A2 _11346_/Q _08963_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07913_ split15/I _08361_/B _07916_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08893_ _08893_/I _11323_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07844_ _07844_/A1 _11016_/A1 _07844_/B _07845_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07347__A1 _07081_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07775_ _07775_/A1 _08586_/A3 _08313_/B _07777_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11383__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09514_ _09514_/I _11519_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06726_ _11350_/Q _06726_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08847__A1 _08863_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09445_ _09445_/I _11497_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_06657_ _11058_/Q input68/Z _06658_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11135__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11265__CLKN input68/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05608_ _11255_/Q _05609_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06322__A2 _08825_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11349__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06588_ input128/Z input127/Z _06588_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_09376_ _09116_/Z _09397_/A2 _09376_/B _09377_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08075__A2 _08395_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08327_ _08327_/A1 _08327_/A2 _08640_/A3 _08509_/B _08330_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_05539_ _05539_/A1 _05539_/A2 _05540_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09272__A1 _09270_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08064__I split12/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08258_ _08400_/A1 _08405_/B _08258_/B _08668_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10957__A2 _10934_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06086__A1 _08761_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11499__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09024__A1 _06847_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07209_ _07240_/A1 _11182_/Q _07210_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10220_ _10377_/B1 _11568_/Q _10221_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08189_ _08189_/A1 _08492_/C _08189_/A3 _08245_/B _08192_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__06389__A2 _06238_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output263_I _11272_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10151_ _11526_/Q _10373_/B1 _11518_/Q _10373_/A1 _10151_/C _10152_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
Xoutput280 _11284_/Q pll_trim[16] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_10082_ _10378_/A1 _11548_/Q _10083_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput291 _11081_/Q pll_trim[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_58_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11374__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10984_ _10984_/A1 _10984_/A2 _10984_/A3 _10985_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__10645__A1 _10645_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11605_ _11605_/D _11686_/RN _06705_/Z _11605_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_11536_ _11536_/D _11686_/RN _06705_/Z _11536_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__10948__A2 _11671_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06077__A1 _10613_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06077__B2 _10137_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11467_ _11467_/D _11686_/RN _06705_/Z _11467_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__06092__A4 _06092_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09566__A2 _09572_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10418_ _10426_/A2 _10460_/A3 _10463_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_11398_ _11398_/D _11686_/RN _06705_/Z _11398_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10349_ _11102_/Q _10350_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07041__A3 _06871_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_715 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_748 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_726 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08526__B1 _07685_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07329__A1 _07310_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06001__A1 _09549_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05890_ _09222_/A1 _11433_/Q _05891_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10884__A1 _10884_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07560_ _07560_/I _07649_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06511_ _06511_/I _11057_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07491_ _07836_/A1 _07699_/A2 _07492_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_09230_ _09125_/Z _09246_/A2 _09230_/B _09231_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11081__SETN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06442_ _06442_/A1 _06442_/A2 _11263_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06373_ _08795_/A1 _06238_/Z _11147_/Q _06375_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11641__CLK _11666_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09161_ _09161_/I _11407_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08112_ split7/I _08213_/B _08113_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10939__A2 _11668_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09092_ _09114_/A2 _11387_/Q _09093_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08043_ _08043_/I _08251_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05815__A1 _08791_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09006__A1 _09013_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09557__A2 _09572_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_214 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input161_I wb_dat_i[9] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09994_ _09994_/I _10034_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06240__A1 _07370_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06791__A2 _11071_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08945_ _07431_/Z _08963_/A2 _08945_/B _08946_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input22_I mask_rev_in[26] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08876_ _06851_/Z _08888_/A2 _08876_/B _08877_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_29_336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07827_ _07827_/I _08341_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__10875__A1 _10919_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11171__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07758_ _08304_/B _08242_/A1 _08305_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11108__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06709_ _11057_/Q input67/Z _06710_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09493__A1 _09497_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07689_ _07689_/A1 _07689_/A2 _07689_/B _07690_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xsplit15 split15/I split15/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08296__A2 _08431_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09428_ _09447_/A2 _11492_/Q _09429_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08048__A2 split16/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09359_ _09372_/A2 _11470_/Q _09360_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09245__A1 _09246_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06059__A1 _05660_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11321_ _11321_/D _11686_/RN _06705_/Z _11321_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_180_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07559__A1 _07575_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11252_ _11252_/D _11686_/RN _06705_/Z _11252_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_4_468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11183_ _11183_/D input76/Z _06705_/Z _11183_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10203_ _10203_/A1 _10203_/A2 _10204_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10134_ _11350_/Q _10351_/A2 _11342_/Q _10351_/B2 _10134_/C _10143_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_69_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11514__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10065_ _10065_/A1 _10065_/A2 _10066_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10618__A1 _10887_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10967_ _11016_/A1 input130/Z _10970_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09484__A1 _09497_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11664__CLK _11665_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10898_ _10898_/A1 _10898_/A2 _10898_/A3 _10898_/A4 _10918_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__10094__A2 _10351_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06298__A1 _08990_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09236__A1 _09158_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07798__A1 _07727_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06217__I _06217_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11519_ _11519_/D _11686_/RN _06705_/Z _11519_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_152_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06222__A1 _07419_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_512 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11586__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07970__A1 split15/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06991_ _06974_/I _11126_/Q _06992_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11194__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08730_ _08740_/A2 _11274_/Q _08731_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05942_ _08839_/A1 _07370_/A1 _05943_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_05873_ _05660_/Z _11625_/Q _05876_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08661_ _08698_/A3 _08698_/A2 _08662_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10857__A1 _10903_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11338__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07612_ _08247_/B _08509_/A1 _08265_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08592_ _07609_/Z _08592_/A2 _08592_/B _08593_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10872__A4 _10872_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10609__A1 _10609_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09475__A1 _09497_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07543_ _07685_/I _07485_/I _07544_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_167_506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07474_ _07495_/A2 _07474_/A2 _07663_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06289__A1 _09041_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10085__A2 _10382_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11510__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07511__I _07511_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09213_ _09220_/A2 _11424_/Q _09214_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09227__A1 _09121_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06425_ _07006_/A2 _11105_/Q _11033_/A2 _06427_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09144_ _09144_/A1 _09015_/Z _09169_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_06356_ _09299_/A1 _11451_/Q _06360_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06287_ _06197_/I _05719_/I _06966_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09075_ _09075_/I _11381_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08026_ _08562_/A1 _08386_/A1 _08033_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11537__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06213__A1 _08795_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11577__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07961__A1 split14/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09977_ _09972_/I _09876_/I _10378_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_08928_ _08938_/A2 _11335_/Q _08929_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10848__B2 _10894_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11329__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08859_ _08863_/A2 _11313_/Q _08860_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09466__A1 _09187_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10821_ _11594_/Q _10913_/A2 _11586_/Q _10913_/B2 _10821_/C _10825_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_10752_ _10910_/A1 _11569_/Q _10755_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10683_ _11527_/Q _10902_/A2 _11519_/Q _10902_/B2 _10683_/C _10690_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__11541__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11067__CLK input68/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11304_ _11304_/D _11686_/RN _06705_/Z _11304_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__11556__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11235_ _11235_/D _11686_/RN _06705_/Z _11235_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_11166_ _11166_/D _11686_/RN _06705_/Z _11166_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__11568__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10000__A2 _10040_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11097_ _11097_/D _11686_/RN _06705_/Z _11097_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__07952__A1 _08355_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10117_ _10375_/A1 _11541_/Q _10119_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10048_ _11323_/Q _10382_/A2 _10048_/B _10049_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10450__C _10450_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07180__A2 _05925_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09457__A1 _09125_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06210_ _05703_/Z _11158_/Q _07370_/A1 _06211_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11016__A1 _11016_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11509__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07190_ _11203_/Q _05925_/Z _07190_/B _07192_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06691__A1 _11306_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06141_ _06141_/A1 _06141_/A2 _06141_/A3 _06141_/A4 _06147_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_06072_ _11566_/Q _09649_/A1 _09624_/A1 _11558_/Q _06074_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06443__A1 _06446_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06994__A2 _06974_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09900_ _09952_/I _10265_/A3 _09901_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09831_ _09831_/I _11620_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11559__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09762_ _09762_/I _11598_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06974_ _06974_/I _06990_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_05925_ _05925_/I _05925_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05954__B1 _09066_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08713_ _11050_/I _11265_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xrebuffer11 _08010_/I _08442_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlya_2
X_09693_ _09697_/A2 _11577_/Q _09694_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09696__A1 _09697_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08644_ _08691_/A1 _08680_/A2 _08644_/A3 _08644_/A4 _08645_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA_input124_I wb_adr_i[5] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05856_ _09016_/A1 _11369_/Q _05858_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05787_ _09349_/A1 _11474_/Q _05788_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08575_ split8/Z _07727_/I _08575_/B _08576_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09999__A2 _11499_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07526_ _07575_/A1 _07590_/A1 _07527_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10058__A2 _10355_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08120__A1 _08161_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07457_ _07457_/I _07999_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_167_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11007__A1 _11007_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07388_ _07389_/A2 _11241_/Q _07389_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06408_ _06408_/I _06408_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06339_ _09699_/A1 _11579_/Q _06341_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09127_ _09125_/Z _09142_/A2 _09127_/B _09128_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09058_ _06859_/Z _09064_/A2 _09058_/B _09059_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06434__A1 _09041_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08009_ split12/I _08632_/A2 _08010_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__06985__A2 _06974_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08187__A1 _08490_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11020_ _10966_/Z _11682_/Q _11021_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07934__A1 split15/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09687__A1 _09697_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10804_ _10896_/A1 _11442_/Q _10806_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10049__A2 _10880_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08111__A1 _08161_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10735_ _10735_/I _10736_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11702__CLK input68/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10666_ _10666_/A1 _10666_/A2 _10667_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10597_ _10900_/A1 _11509_/Q _10598_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06425__A1 _07006_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11218_ _11218_/D input162/Z _11666_/CLK _11218_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_11149_ _11149_/D _11686_/RN _06705_/Z _11149_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__07925__A1 split21/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09678__A1 _09697_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06690_ _11178_/Q _06692_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05710_ _05710_/I _09624_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
X_05641_ _08825_/A2 _08839_/A2 _05642_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11232__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08360_ _08437_/A1 _08439_/A2 _08549_/B _08363_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_23_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08102__A1 _08434_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05572_ input58/Z _05576_/C _05572_/B _05573_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07311_ _10935_/A1 _07326_/A2 _07313_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08291_ _08291_/I _08292_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07456__A3 _07455_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07242_ _05927_/Z _07242_/A2 _09015_/I _07265_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XANTENNA__10460__A2 _10506_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11382__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07173_ _07173_/I _11175_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08405__A2 _07586_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06416__A1 _08839_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06124_ _09041_/A1 _11373_/Q _06126_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06967__A2 _11119_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06055_ _11430_/Q _06056_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09814_ _09158_/I _09823_/A2 _09814_/B _09815_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06719__A2 input86/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10920__B1 _10920_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09669__A1 _09241_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09745_ _09241_/I _09725_/Z _09745_/B _09746_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06957_ _10950_/A1 _06957_/A2 _06959_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06888_ _06888_/I _11095_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05908_ _09349_/A1 _11472_/Q _05909_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09676_ _09116_/I _09697_/A2 _09676_/B _09677_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10279__A2 _11418_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08341__A1 _08677_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08627_ _08627_/I _08665_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05839_ _06266_/I _11300_/Q _05840_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07695__A3 _07492_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08892__A2 _08913_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08558_ _08558_/A1 _08558_/A2 _08558_/A3 _08693_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_07509_ _08315_/B split5/Z _07510_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08489_ _08480_/Z _08657_/A1 _08486_/Z _08582_/A2 _08493_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_168_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10520_ _10913_/A2 _11588_/Q _10522_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10451__A2 _10451_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10451_ _10514_/I _10451_/A2 _10451_/A3 _10510_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__10739__B1 _10920_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10382_ _10382_/A1 _10382_/A2 _10382_/B _10382_/C _10384_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__11105__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11003_ _08493_/B input151/Z _11005_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11255__CLK _06687_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08686__B _08686_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07135__A2 _09158_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08332__A1 _08332_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08635__A2 _11258_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10718_ _10891_/A1 _11480_/Q _10720_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11698_ _11698_/D _11698_/RN input68/Z _11698_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xrebuffer2 _08002_/A1 _08000_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10649_ _10922_/A1 _11358_/Q _10650_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07071__A1 _06837_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06949__A2 _06941_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07860_ _07860_/A1 _07859_/Z _07861_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07791_ _08696_/A2 _08592_/B _08507_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06811_ _06835_/A1 _11074_/Q _06812_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11372__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09530_ _09530_/I _11524_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06742_ _06742_/I _06742_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08323__A1 _08332_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09461_ _09461_/I _11502_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07126__A2 _05927_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06334__B1 _11523_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06673_ input3/Z input1/Z _06674_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09392_ _09392_/I _11480_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05688__A2 _05803_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08412_ _08412_/A1 _08411_/Z _08414_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05624_ _05624_/I _05684_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11387__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09823__A1 _09270_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05555_ _11693_/Q _05557_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08343_ _08580_/A2 _08677_/A2 _08519_/B _08344_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_11_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06637__A1 input77/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10433__A2 _10427_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08274_ _08274_/A1 _08418_/A1 _08274_/A3 _08535_/A2 _08279_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__10969__B1 _08460_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07225_ _07240_/A1 _07225_/A2 _07225_/B _07226_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11128__CLK _11683_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11041__I _11050_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10085__C _10085_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07156_ _05642_/I _06701_/I _07267_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__10197__A1 _10353_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07062__A1 _08795_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07087_ _07076_/Z _07090_/A2 _07087_/B _07088_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06107_ _06107_/A1 _06107_/A2 _06108_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input52_I mgmt_gpio_in[24] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06038_ _06304_/A2 _06102_/A1 _06039_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11278__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07989_ _07989_/A1 _07989_/A2 _07990_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09728_ _09728_/I _11587_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07117__A2 _07151_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10121__A1 _10379_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09659_ _09672_/A2 _11566_/Q _09660_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output306_I _06696_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08865__A2 _06838_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10672__A2 _11479_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_11621_ _11621_/D _11686_/RN _06705_/Z _11621_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_144_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09814__A1 _09158_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11552_ _11552_/D _11686_/RN _06705_/Z _11552_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__09290__A2 _11448_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11483_ _11483_/D _11686_/RN _06705_/Z _11483_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_10503_ _10506_/A1 _10503_/A2 _10504_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10434_ _10493_/A2 _10460_/A1 _10480_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_10365_ _11229_/Q _10365_/A2 _10365_/B1 _11233_/Q _10368_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07053__A1 _06843_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_908 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05603__A2 _05515_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10296_ _10375_/A1 _11546_/Q _10298_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_919 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07356__A2 _06217_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08305__A1 _08686_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10112__B2 _11501_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09805__A1 _09121_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06619__A1 _06619_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09281__A2 _11445_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10179__A1 _10371_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07010_ _07011_/A2 _11132_/Q _07011_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09033__A2 _09039_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11420__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08961_ _08961_/I _11345_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07912_ _07912_/A1 _07912_/A2 _07916_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08892_ _07426_/Z _08913_/A2 _08892_/B _08893_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11570__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07843_ _07843_/A1 _07843_/A2 _07843_/A3 _07843_/A4 _07844_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__10351__B2 _10351_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07774_ _08328_/B1 _07774_/A2 _08313_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09513_ _09158_/Z _09522_/A2 _09513_/B _09514_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06725_ _06725_/I _06725_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09444_ _09241_/Z _09447_/A2 _09444_/B _09445_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_06656_ _06668_/C _11174_/Q _06658_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_05607_ _06466_/B _11061_/Q _06497_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06587_ _06587_/I _08005_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09375_ _09397_/A2 _11475_/Q _09376_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05969__I _05969_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08326_ _07722_/I _07586_/I _08639_/B _08509_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05538_ _05536_/Z _05538_/A2 _11699_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09272__A2 _09272_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07283__A1 _07290_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08257_ _08449_/A1 _07566_/I _08405_/B _08406_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08188_ _08490_/A1 _08205_/C _08242_/A1 _08245_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_07208_ _11316_/Q _05924_/Z _07208_/B _07210_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07139_ _11169_/Q _07142_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09024__A2 _09039_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08783__A1 _08784_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10590__A1 _10914_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10150_ _10634_/A2 _09961_/I _09965_/I _10634_/B2 _10151_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
Xoutput270 _11278_/Q pll_sel[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA_output256_I _11704_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10081_ _10379_/A1 _11556_/Q _10083_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11279__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput281 _11285_/Q pll_trim[17] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput292 _11082_/Q pll_trim[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_181_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10983_ _08431_/B input131/Z _08460_/B input139/Z _10984_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_74_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06849__A1 _06847_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11604_ _11604_/D _11686_/RN _06705_/Z _11604_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_11535_ _11535_/D _11686_/RN _06705_/Z _11535_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__07274__A1 _07290_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11443__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11466_ _11466_/D _11686_/RN _06705_/Z _11466_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10417_ _10417_/I _10460_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
X_11397_ _11397_/D _11686_/RN _06705_/Z _11397_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__10581__A1 _10894_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11593__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08774__A1 _08784_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10348_ _11207_/Q _10382_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_749 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_10279_ _10357_/A1 _11418_/Q _10280_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08526__B2 _07485_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08526__A1 _08686_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06001__A2 _11535_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05760__A1 _06785_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08829__A2 _06904_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07490_ _07490_/I _07699_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_80_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06510_ _06610_/A2 _06510_/A2 _06510_/B _06511_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06441_ _05584_/I _11263_/Q _06442_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06372_ _09424_/A1 _11491_/Q _07427_/A1 _11252_/Q _06375_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09160_ _09158_/Z _09169_/A2 _09160_/B _09161_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07265__A1 _06867_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08111_ _08161_/A1 _08213_/B _08470_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09091_ _09091_/A1 _09015_/Z _09114_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_08042_ _08614_/A2 _08358_/A2 _08043_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05815__A2 _06217_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09993_ _09993_/A1 _11633_/Q _09994_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08765__A1 _08784_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input154_I wb_dat_i[31] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06240__A2 _06238_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08944_ _08963_/A2 _11340_/Q _08945_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08875_ _08888_/A2 _11318_/Q _08876_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07826_ _07826_/A1 _07826_/A2 _07831_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11316__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07740__A2 _08339_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07757_ _07757_/A1 _07757_/A2 _07759_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input15_I mask_rev_in[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06708_ _06753_/A1 input85/Z _06710_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xsplit16 split16/I split16/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07688_ _07688_/A1 _07688_/A2 _07704_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06639_ _06639_/I _06639_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11466__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09427_ _09427_/I _11491_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09358_ _09358_/I _11469_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09245__A2 _11434_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06059__A2 _11622_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07256__A1 _06855_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08309_ _08309_/I _08500_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10260__B1 _10373_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09289_ _09289_/I _11447_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11320_ _11320_/D input76/Z _06705_/Z _11320_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_176_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07008__A1 _06837_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11251_ _11251_/D _11686_/RN _06705_/Z _11251_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_109_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08756__A1 _06855_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10202_ _10357_/A1 _11416_/Q _10203_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11182_ _11182_/D _11686_/RN _06705_/Z _11182_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_69_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10133_ _10350_/A1 _10133_/A2 _10134_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10563__A1 _10886_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05990__A1 _08990_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10064_ _10361_/A1 _11420_/Q _10065_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09181__A1 _09195_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09484__A2 _11510_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10966_ _10966_/I _10966_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__10618__A2 _11430_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10897_ _11229_/Q _10897_/A2 _10897_/B1 _11233_/Q _10898_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07247__A1 _07081_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09236__A2 _09246_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07798__A2 _08639_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08995__A1 _07431_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11518_ _11518_/D _11686_/RN _06705_/Z _11518_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__11283__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08713__I _11050_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11449_ _11449_/D _11686_/RN _06705_/Z _11449_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_131_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08747__A1 _07431_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11264__CLKN input68/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10554__A1 _10887_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06990_ _10950_/A1 _06990_/A2 _06992_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_535 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11339__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05941_ _05941_/I _07370_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__05981__A1 _06785_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10306__A1 _10306_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input7_I mask_rev_in[12] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_568 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_05872_ _11617_/Q _09800_/A1 _11609_/Q _09775_/A1 _05872_/C _05876_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_08660_ _08464_/Z _08089_/I _08660_/A3 _08660_/A4 _08698_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__09172__A1 _09195_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11489__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07611_ _08417_/A2 _07774_/A2 _08411_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_08591_ _08591_/I _08679_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07542_ _07542_/A1 _07690_/A2 _07685_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__10609__A2 _10092_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07473_ _07689_/B _07474_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09212_ _09212_/I _11423_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06424_ _08915_/A1 _11331_/Q _06912_/A1 _11103_/Q _06427_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06355_ _06355_/A1 _06355_/A2 _06355_/A3 _06355_/A4 _06371_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_09143_ _09143_/I _11402_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07238__A1 _11322_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09227__A2 _09246_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11274__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09074_ _06847_/Z _09089_/A2 _09074_/B _09075_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06286_ _06286_/A1 _06286_/A2 _06286_/A3 _06302_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_08025_ _08393_/B _08545_/A2 _08032_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06461__A2 _06610_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07410__A1 _07081_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10545__A1 _10883_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06213__A2 _06217_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09976_ _10379_/A1 _11555_/Q _09983_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08927_ _08927_/I _11334_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05972__A1 _10950_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10848__A2 _10894_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09163__A1 _06859_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08858_ _08858_/I _11312_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07809_ _08674_/B _08332_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08910__A1 _06863_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08789_ _08789_/A1 _08827_/A2 _08789_/B _08790_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09466__A2 _09472_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10820_ _10820_/A1 _10820_/A2 _10821_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10751_ _11625_/Q _10916_/A1 _11617_/Q _10915_/A1 _10751_/C _10755_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_10682_ _10682_/A1 _10682_/A2 _10683_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07229__A1 _07240_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11025__A2 _11025_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10784__A1 _10921_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11303_ _11303_/D _11686_/RN _06705_/Z _11303_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_113_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11234_ _11234_/D _11686_/RN _06705_/Z _11234_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__08689__B _08689_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_470 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10536__A1 _10903_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11165_ _11165_/D _11686_/RN _06705_/Z _11165_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_136_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11096_ _11096_/D _11686_/RN _06705_/Z _11096_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10116_ _10373_/A1 _11517_/Q _10373_/B1 _11525_/Q _10119_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_96_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11080__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11631__CLK _11666_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10047_ _10047_/A1 _10382_/A2 _10047_/B _10048_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08901__A1 _06851_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09457__A2 _09472_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10949_ _10949_/A1 _10949_/A2 _11671_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06140__A1 _05660_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06691__A2 input94/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10775__A1 _11545_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06140_ _05660_/Z _11621_/Q _06141_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10775__B2 _10905_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06071_ _11534_/Q _09549_/A1 _11526_/Q _05693_/Z _06071_/C _06074_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__07640__A1 _07640_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11256__RN input162/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11161__CLK input68/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09393__A1 _09397_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08196__A2 _07722_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_470 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09830_ _09121_/I _09848_/A2 _09830_/B _09831_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09761_ _09154_/I _09773_/A2 _09761_/B _09762_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06973_ _11220_/Q input162/Z _06974_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_05924_ _05924_/I _05924_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09145__A1 _09169_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08712_ _11050_/I _11264_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09692_ _09692_/I _11576_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08643_ _08341_/B split5/Z _08644_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05706__A1 _05703_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05855_ input27/Z _06398_/A2 _05995_/A2 _08799_/A1 _05855_/C _05860_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_05786_ _05786_/I _09349_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
X_08574_ _08617_/A1 _08698_/A2 _08577_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input117_I wb_adr_i[28] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07525_ _07525_/I _07590_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07522__I _07522_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11044__I _11050_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07456_ _07846_/A1 _07470_/I _07455_/Z _07472_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11495__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11007__A2 _10966_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07387_ _07387_/I _11240_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06407_ _11690_/Q _11057_/Q _11294_/Q _06408_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__11504__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06338_ _06338_/A1 _06338_/A2 _06338_/A3 _06338_/A4 _06350_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA_input82_I spi_sdo VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08959__A1 _08963_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09126_ _09142_/A2 _11397_/Q _09127_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11247__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06269_ _06694_/A1 _05836_/I _06269_/B _06269_/C _06281_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09057_ _09064_/A2 _11376_/Q _09058_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08008_ _08008_/A1 _08041_/I split12/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__10518__B2 _10911_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08187__A2 _08395_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06198__A1 _05703_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09384__A1 _09397_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11654__CLK _11665_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09959_ _09959_/I _10042_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05945__A1 _06266_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09136__A1 _06859_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09912__I _09912_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10803_ _10895_/A1 _11450_/Q _10806_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10734_ _10734_/A1 _10734_/A2 _10735_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11486__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06673__A2 input1/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10665_ _10887_/B1 _11431_/Q _10666_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11184__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10596_ _10902_/B2 _11517_/Q _10598_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10757__A1 _10887_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11238__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09375__A1 _09397_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06189__A1 _09574_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11217_ _11217_/D input162/Z _11672_/CLK _11222_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_11148_ _11148_/D _11686_/RN _06705_/Z _11148_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__05936__A1 _06324_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11410__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09127__A1 _09125_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11079_ _11079_/D _11686_/RN _06705_/Z _11079_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_05640_ _05600_/I _09724_/A1 _08839_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__08350__A2 _08395_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10693__B1 _10920_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06361__A1 _09197_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05571_ _05575_/A1 _11068_/Q _05572_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07310_ _07310_/I _07326_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11527__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08290_ _08394_/A1 _08395_/A2 _08294_/B _08290_/C _08291_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__10996__A1 _08493_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09850__A2 _10092_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06113__A1 _08803_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06664__A2 _11187_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07241_ _07241_/I _11188_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_176_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07172_ _07197_/A1 _07172_/A2 _07172_/B _07173_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11677__CLK _06687_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10748__A1 _10914_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11229__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06416__A2 _11087_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06123_ _11349_/Q _05723_/Z _11357_/Q _08990_/A1 _06123_/C _06128_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_06054_ _11438_/Q _06056_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09366__A1 _09187_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09813_ _09823_/A2 _11615_/Q _09814_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11401__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09118__A1 _09142_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10920__A1 _10920_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09669__A2 _09672_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09744_ _09725_/Z _11593_/Q _09745_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11540__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06956_ _06956_/A1 _06956_/A2 _11115_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06887_ _06847_/Z _06902_/A2 _06887_/B _06888_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05907_ _09324_/A1 _11464_/Q _05909_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09675_ _09697_/A2 _11571_/Q _09676_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11057__CLK input68/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08626_ _08626_/A1 _08626_/A2 _08261_/I _08626_/A4 _08688_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_05838_ _11665_/Q _10927_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08557_ split6/Z _08546_/I _08557_/B _08558_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__11555__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05769_ _09041_/A1 _11378_/Q _05773_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09841__A2 _11624_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07508_ _07508_/I _08315_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_08488_ _08488_/A1 _08488_/A2 _08582_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_22_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07439_ input99/Z input98/Z _07440_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_167_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08083__I split8/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10450_ _11411_/Q _10888_/A1 _11371_/Q _10883_/A1 _10450_/C _10451_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__10739__A1 _10920_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09109_ _09109_/I _11392_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07604__A1 _07593_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10381_ _10381_/A1 _10381_/A2 _10381_/A3 _10381_/A4 _10382_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__06407__A2 _11057_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09357__A1 _09125_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11002_ _11016_/A1 input157/Z _11005_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10911__A1 _10911_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05918__B2 _09171_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05918__A1 _11424_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11508__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08332__A2 _08417_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10675__B1 _11487_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06343__A1 _05703_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10978__A1 _10966_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09832__A2 _11621_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10717_ _10717_/A1 _10717_/A2 _10717_/A3 _10717_/A4 _10737_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__06646__A2 _06646_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11697_ _11697_/D _11697_/RN input68/Z _11697_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__09596__A1 _09597_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer3 _07998_/A1 _08006_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10648_ _10921_/A1 _11334_/Q _10650_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10579_ _10892_/A1 _11469_/Q _10583_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_3_6__f_wb_clk_i_I clkbuf_0_wb_clk_i/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11631__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10902__B2 _10902_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08571__A2 _08696_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07790_ _08332_/A1 _08592_/B _07790_/B _07796_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06810_ _11693_/Q _05633_/B _06810_/B _09154_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_06741_ input63/Z input80/Z _06742_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__08323__A2 _08417_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09460_ _09154_/Z _09472_/A2 _09460_/B _09461_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06334__B2 _05693_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08411_ _08411_/A1 _08411_/A2 _08411_/A3 _08411_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_06672_ _11181_/Q _06674_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09391_ _09187_/Z _09397_/A2 _09391_/B _09392_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05623_ _05623_/A1 _11205_/Q _05623_/B _05624_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_08342_ _08342_/A1 _08641_/A1 _08515_/B _08599_/I _08348_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_05554_ _05554_/I _11695_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06637__A2 input91/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09823__A2 _09823_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08273_ split14/Z _07609_/Z _08415_/B _08535_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10969__A1 _08431_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07224_ _07240_/A1 _11185_/Q _07225_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09587__A1 _09597_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07155_ _11050_/I _11172_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05860__A3 _05860_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07062__A2 _06238_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07086_ _07090_/A2 _11153_/Q _07087_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06106_ _06396_/A1 input26/Z _06107_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06037_ _11266_/Q _06102_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input45_I mgmt_gpio_in[18] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08011__A1 _08434_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07988_ _07988_/A1 _08013_/A2 _08385_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08562__A2 _08562_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09727_ _09116_/I _09725_/Z _09727_/B _09728_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_498 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06939_ _06939_/I _11110_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10121__A2 _11557_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09658_ _09658_/I _11565_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06325__A1 _08825_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_09589_ _09589_/I _11543_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08609_ _08649_/A1 _08692_/A2 _08609_/B _08610_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06876__A2 _11088_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_11620_ _11620_/D _11686_/RN _06705_/Z _11620_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__08078__A1 split12/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07825__A1 _08204_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11551_ _11551_/D _11686_/RN _06705_/Z _11551_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__09814__A2 _09823_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06628__A2 input77/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10502_ _10502_/I _10506_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_10_143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_11482_ _11482_/D _11686_/RN _06705_/Z _11482_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_6_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09578__A1 _09597_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10433_ _10433_/A1 _10427_/B _10899_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_12_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_10364_ _10364_/A1 _10364_/A2 _10364_/A3 _10364_/A4 _10382_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__11613__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11222__CLK _11666_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10295_ _10373_/A1 _11522_/Q _10373_/B1 _11530_/Q _10298_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_909 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09750__A1 _09750_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07356__A3 _06871_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11372__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08305__A2 _07761_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06316__A1 _07201_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10112__A2 _10369_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08716__I _11050_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09805__A2 _09823_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09569__A1 _09241_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10179__A2 _11487_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06680__B _06680_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08792__A2 _11293_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08960_ _06863_/Z _08963_/A2 _08960_/B _08961_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07911_ _07911_/I _07912_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08891_ _08913_/A2 _11323_/Q _08892_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09741__A1 _09725_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07842_ _08519_/B _08345_/A2 _07843_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10887__B1 _10887_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10351__A2 _10351_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09512_ _09522_/A2 _11519_/Q _09513_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07773_ _08592_/A2 _08315_/B _08586_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10639__B1 _11614_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06724_ _06724_/A1 _11056_/Q _06725_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09443_ _09447_/A2 _11497_/Q _09444_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06655_ _06655_/I _06655_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09374_ _09374_/A1 _09015_/Z _09397_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XPHY_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_05606_ _11060_/Q _05515_/I _11205_/Q _05609_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06586_ input112/Z input111/Z _06587_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_08325_ _08686_/A2 _08639_/B _08325_/B _08640_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07807__A1 _08328_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05537_ _05537_/A1 _05539_/A2 _05538_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08256_ split21/I _08449_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__11245__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08187_ _08490_/A3 _08395_/A2 _08243_/B _08189_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07207_ _05924_/Z _09121_/I _07208_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07138_ _07138_/I _11168_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08232__A1 split7/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07069_ _07419_/A2 _06238_/Z _06871_/Z _07074_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__05597__A2 _05633_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput260 _11282_/Q pll90_sel[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput271 _11279_/Q pll_sel[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__11395__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10080_ _10377_/A1 _11572_/Q _10377_/B1 _11564_/Q _10083_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xoutput282 _11286_/Q pll_trim[18] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA_output249_I _06713_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput293 _11083_/Q pll_trim[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__09732__A1 _09725_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10982_ _08493_/B input148/Z _10984_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10131__I _11326_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09920__I _09920_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06849__A2 _06869_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11603_ _11603_/D _11686_/RN _06705_/Z _11603_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_11_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10802__B1 _11490_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11534_ _11534_/D _11686_/RN _06705_/Z _11534_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_11465_ _11465_/D _11686_/RN _06705_/Z _11465_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__11371__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10416_ _10416_/I _10914_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_11396_ _11396_/D _11686_/RN _06705_/Z _11396_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__05588__A2 _05515_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08774__A2 _11288_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10347_ _10347_/I _11654_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06785__A1 _06785_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10581__A2 _11485_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_10278_ _10356_/A1 _11410_/Q _10280_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11118__CLK _11672_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05760__A2 _11078_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_393 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06440_ _10935_/A1 _05969_/I _06619_/B _06442_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_73_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06371_ _06371_/A1 _06371_/A2 _06371_/A3 _06371_/A4 _06392_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__07265__A2 _07265_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08110_ _08434_/A1 _08213_/B _08212_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09090_ _09090_/I _11386_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08041_ _08041_/I _08167_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11339__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09962__A1 _10374_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09992_ _11459_/Q _10365_/B1 _11451_/Q _10365_/A2 _09992_/C _10006_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__05579__A2 _11687_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08943_ _08943_/I _11339_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08517__A2 _07564_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06528__A1 _11687_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07525__I _07525_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input147_I wb_dat_i[25] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08874_ _08874_/I _11317_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07825_ _08204_/I _07827_/I _07825_/B _07826_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11047__I _11050_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07756_ _08498_/C _07757_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06707_ _11057_/Q _06753_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
X_09426_ _09116_/Z _09447_/A2 _09426_/B _09427_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07687_ _08630_/C _07688_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06638_ _11614_/Q input77/Z _06638_/B _06639_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09357_ _09125_/Z _09372_/A2 _09357_/B _09358_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06569_ _11223_/Q _08460_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__07256__A2 _07265_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08308_ _08332_/A1 _08417_/A2 _08587_/B _08309_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09288_ _09158_/Z _09297_/A2 _09288_/B _09289_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10260__A1 _10373_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08239_ _08578_/A2 _08621_/A3 _08621_/A2 _08241_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_output199_I _06738_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09187__I _09187_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08205__A1 _08519_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11250_ _11250_/D _11686_/RN _06705_/Z _11250_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__08756__A2 _08759_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11181_ _11181_/D _11686_/RN _06705_/Z _11181_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10201_ _10356_/A1 _11408_/Q _10203_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10132_ _11334_/Q _10133_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10063_ _10360_/A1 _11428_/Q _10065_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07192__A1 _07197_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09181__A2 _11414_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10965_ _10965_/A1 _10965_/A2 _07297_/I _10966_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__11410__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10896_ _10896_/A1 _11144_/Q _10898_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11560__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08444__A1 _08449_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07247__A2 _07265_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11517_ _11517_/D _11686_/RN _06705_/Z _11517_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__10251__A1 _10251_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10745__B _10745_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08995__A2 _09013_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11448_ _11448_/D _11686_/RN _06705_/Z _11448_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__10003__A1 _09996_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08747__A2 _08759_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11379_ _11379_/D _11686_/RN _06705_/Z _11379_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XTAP_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06222__A3 _06217_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_05940_ _05940_/A1 _05940_/A2 _05941_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__05981__A2 _11075_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10306__A2 _06556_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_569 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_05871_ _05871_/A1 _05871_/A2 _05872_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09172__A2 _11411_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08590_ _08590_/A1 _08590_/A2 _08590_/A3 _08590_/A4 _08591_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
X_07610_ _08247_/B _07609_/Z _07613_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07541_ _07541_/I _07542_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11090__CLK _11665_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07472_ _07472_/A1 _07472_/A2 _07689_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10490__A1 _10910_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09211_ _09158_/Z _09220_/A2 _09211_/B _09212_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06423_ _06423_/A1 _06423_/A2 _06423_/A3 _06438_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06354_ _08786_/A1 _11143_/Q _06217_/Z _06355_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09142_ _06867_/Z _09142_/A2 _09142_/B _09143_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07238__A2 _05924_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06997__A1 _10957_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09073_ _09089_/A2 _11381_/Q _09074_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10242__B2 _10359_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06285_ _09066_/A1 _11380_/Q _06286_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08024_ _08391_/B _08393_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09935__A1 _10911_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09975_ _09975_/I _10379_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__11216__SETN input162/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08926_ _06851_/Z _08938_/A2 _08926_/B _08927_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07174__A1 _05925_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09163__A2 _09169_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08857_ _06851_/Z _08863_/A2 _08857_/B _08858_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07808_ _07808_/A1 _07808_/A2 _08674_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08910__A2 _08913_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11433__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06921__A1 _06837_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08788_ _08789_/A1 _07114_/C _11292_/Q _08789_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07739_ _08589_/A1 _08580_/A2 _08302_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08674__A1 _07566_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11583__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10750_ _10750_/A1 _10750_/A2 _10751_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09409_ _09422_/A2 _11486_/Q _09410_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10681_ _10900_/A1 _11511_/Q _10682_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10481__A1 _10897_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07229__A2 _11186_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10233__A1 _10350_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06988__A1 _06974_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11302_ _11302_/D _11686_/RN _06705_/Z _11302_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_11233_ _11233_/D _11686_/RN _06705_/Z _11233_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_20_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_11164_ _11164_/D _11686_/RN _06705_/Z _11164_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__09941__A4 _09922_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11095_ _11095_/D _11686_/RN _06705_/Z _11095_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10115_ _10115_/A1 _10115_/A2 _10115_/A3 _10124_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_10046_ _10046_/A1 _10046_/A2 _10046_/A3 _10046_/A4 _10047_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__08362__B1 split15/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08901__A2 _08913_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10948_ _10934_/I _11671_/Q _10949_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_176_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10472__A1 _10887_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06140__A2 _11621_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10879_ _10879_/A1 _10092_/Z _10877_/Z _10879_/A4 _10880_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__10224__A1 _10375_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08417__A1 split15/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06979__A1 _06974_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10775__A2 _10906_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06070_ _10146_/A2 _05689_/I _05691_/I _10634_/B2 _06071_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__11306__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09917__B2 _09902_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11456__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09760_ _09773_/A2 _11598_/Q _09761_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06972_ _06972_/I _11120_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_09691_ _09187_/I _09697_/A2 _09691_/B _09692_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05923_ _05923_/A1 _05923_/A2 _05923_/A3 _05923_/A4 _05939_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_399 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09145__A2 _11403_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05954__A2 _09091_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08711_ _11050_/I _11263_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08642_ _08642_/A1 _08642_/A2 _08642_/A3 _08644_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__05706__A2 _08799_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05854_ _05854_/A1 _05854_/A2 _05854_/A3 _05855_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_66_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08573_ _08573_/A1 _08573_/A2 _08573_/A3 _08573_/A4 _08698_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_05785_ _06238_/I _05995_/A2 _05786_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11192__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_07524_ _07524_/A1 _07524_/A2 _07525_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08656__A1 _08656_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_167_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07455_ _07996_/A2 split5/I _07455_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_06406_ _06406_/A1 _06406_/A2 _06406_/A3 _06406_/A4 _06419_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_07386_ _07076_/Z _07389_/A2 _07386_/B _07387_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09125_ _09125_/I _09125_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__10215__A1 _10371_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06337_ _09574_/A1 _11539_/Q _07092_/A1 _11155_/Q _06338_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input75_I pad_flash_io1_di VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09056_ _09056_/I _11375_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06268_ _08829_/A1 _11305_/Q _06269_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08007_ _08007_/A1 _08007_/A2 _08041_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_135_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10518__A2 _10915_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06199_ _05703_/Z _08795_/A1 _11146_/Q _06200_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__06198__A2 _08786_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09384__A2 _11478_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09958_ _09958_/A1 _11632_/Q _09959_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_08909_ _08913_/A2 _11329_/Q _08910_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09136__A2 _09142_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09889_ _09889_/I _10023_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_66_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10151__B1 _11518_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07698__A2 _08614_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08895__A1 _07431_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11183__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10802_ _11498_/Q _10894_/A2 _11490_/Q _10894_/B2 _10802_/C _10806_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_13_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10733_ _10906_/A1 _11544_/Q _10734_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11263__CLKN input68/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11329__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10664_ _10887_/A2 _11423_/Q _10666_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05881__A1 _09499_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10595_ _10902_/A2 _11525_/Q _10598_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10757__A2 _11433_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11479__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07622__A2 _08509_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06425__A3 _11033_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10509__A2 _10509_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11216_ _11216_/D input162/Z _11666_/CLK _11216_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__07386__A1 _07076_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11147_ _11147_/D _11686_/RN _06705_/Z _11147_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__05936__A2 _11592_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09127__A2 _09142_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput160 wb_dat_i[8] input160/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11078_ _11078_/D _11686_/RN _06705_/Z _11078_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__10142__B1 _11438_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10029_ _10135_/A1 _09893_/I _10351_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__11174__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10693__A1 _10920_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06361__A2 _11419_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05570_ _11690_/Q _06610_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_44_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07240_ _07240_/A1 _07240_/A2 _07240_/B _07241_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05872__B2 _09775_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07171_ _07197_/A1 _11175_/Q _07172_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09063__A1 _09064_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06122_ _10607_/A1 _05991_/I _06122_/B _06123_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08810__A1 _08820_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06416__A3 _06872_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06053_ _11422_/Q _09197_/A1 _11414_/Q _09171_/A1 _06053_/C _06058_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__09366__A2 _09372_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07377__A1 _08825_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09812_ _09812_/I _11614_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09743_ _09743_/I _11592_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06955_ _06941_/I _11115_/Q _06956_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06886_ _06902_/A2 _11095_/Q _06887_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05906_ _05906_/A1 _05906_/A2 _05906_/A3 _05906_/A4 _05939_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_09674_ _09674_/A1 _09015_/I _09697_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__10684__A1 _10904_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08625_ _08686_/A1 _08686_/A2 _08625_/B _08626_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__11165__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05837_ _11301_/Q _06266_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08556_ _08647_/I _08651_/A2 _08559_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_14_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07507_ _07793_/A1 _08045_/A3 _07508_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__10436__A1 _10913_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05768_ _05768_/I _09041_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
X_08487_ _08487_/I _08488_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05699_ _05753_/A1 _05699_/A2 _05700_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_07438_ input128/Z input127/Z _07440_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11621__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07201__C _09015_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07369_ _07369_/I _11235_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09054__A1 _09064_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09108_ _06859_/Z _09114_/A2 _09108_/B _09109_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10380_ _10380_/A1 _10380_/A2 _10380_/A3 _10381_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__05615__A1 _06466_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output181_I _10144_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output279_I _11078_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09039_ _06867_/Z _09039_/A2 _09039_/B _09040_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09357__A2 _09372_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11001_ _11001_/I _11679_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07368__A1 _07081_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_293 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05918__A2 _09197_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10675__B2 _10894_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11156__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06343__A2 _07419_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11151__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11696_ _11696_/D _11696_/RN input68/Z _11696_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10716_ _10886_/B2 _11392_/Q _10886_/A2 _11400_/Q _10717_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_10647_ _10920_/A1 _11342_/Q _10920_/B1 _11350_/Q _10650_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09045__A1 _09064_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer4 _07998_/A1 _08002_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09596__A2 _11546_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10578_ _10578_/A1 _10578_/A2 _10578_/A3 _10578_/A4 _10578_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__06031__A1 _09775_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10902__A2 _10902_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08859__A1 _08863_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06740_ _06740_/I _06740_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11147__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06671_ _06671_/A1 _06671_/A2 _11056_/Q _06724_/A1 _06671_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06334__A2 _07099_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05622_ _08684_/A1 _11205_/Q _05623_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08410_ split15/Z _08247_/B _08411_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09390_ _09397_/A2 _11480_/Q _09391_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08341_ _08677_/A2 _08345_/A2 _08341_/B _08599_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05553_ _05553_/A1 _05519_/I _05553_/B _05554_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11644__CLK _11665_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07834__A2 _08358_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08272_ _08534_/B _08274_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06098__A1 _06098_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09036__A1 _06863_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07223_ _11319_/Q _05924_/Z _07223_/B _07225_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09587__A2 _11543_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07154_ _11055_/I _11050_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__07062__A3 _06871_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07085_ _08825_/A1 _06238_/Z _06871_/Z _07090_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_06105_ input13/Z _06393_/A1 _06394_/A1 input5/Z _06107_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06036_ _06036_/A1 _06036_/A2 _10947_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06270__A1 _08890_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10382__C _10382_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07987_ _07987_/A1 _08454_/A2 _08454_/A3 _07993_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_input38_I mgmt_gpio_in[11] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11386__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07770__A1 _08332_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09726_ _09725_/Z _11587_/Q _09727_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11174__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06938_ _06843_/Z _06938_/A2 _06938_/B _06939_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10106__B1 _11437_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10657__A1 _10914_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11138__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_09657_ _09125_/I _09672_/A2 _09657_/B _09658_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06325__A2 _11238_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06869_ _06867_/Z _06869_/A2 _06869_/B _06870_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08608_ _08608_/A1 _08366_/I _08608_/A3 _08608_/A4 _08693_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XTAP_1137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_09588_ _09158_/Z _09597_/A2 _09588_/B _09589_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_63_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08078__A2 _08545_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10409__A1 _10506_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08539_ _08539_/A1 _08629_/A3 _08665_/A1 _08541_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_11550_ _11550_/D _11686_/RN _06705_/Z _11550_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10501_ _10501_/A1 _10501_/A2 _10502_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11481_ _11481_/D _11686_/RN _06705_/Z _11481_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_6_115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09027__A1 _06851_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11310__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10432_ _10432_/I _10906_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_10363_ _11227_/Q _10363_/A2 _11144_/Q _10363_/B2 _10363_/C _10364_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__06261__A1 _08799_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10294_ _10294_/A1 _10294_/A2 _10294_/A3 _10303_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__06013__A1 _09424_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11517__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09750__A2 _09015_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10896__A1 _10896_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11377__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11129__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10648__A1 _10921_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11667__CLK _11683_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07816__A2 _08513_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05827__A1 _05827_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11679_ _11679_/D input162/Z _06687_/A2 _11679_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__11301__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09018__A1 _07426_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09569__A2 _09572_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07910_ _07921_/A1 _08361_/B _07911_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__11197__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08890_ _08890_/A1 _06838_/Z _08913_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_68_111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09741__A2 _11592_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06004__A1 _09649_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07841_ _08545_/A2 _08677_/A2 _08519_/B _07843_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11368__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07772_ _07774_/A2 _08696_/A2 _07772_/B _07775_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09511_ _09511_/I _11518_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10639__A1 _11622_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06723_ _06723_/I _06723_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10639__B2 _10915_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09442_ _09442_/I _11496_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06654_ _06786_/A1 _11059_/Q _06654_/B _06655_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06585_ _06585_/I _08006_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
X_09373_ _09373_/I _11474_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_05605_ _05605_/I _05646_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08324_ _08507_/B _08327_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05536_ _05537_/A1 _05539_/A2 _05536_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__10811__A1 _10904_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08255_ _08400_/A1 _07596_/I _08255_/B _08530_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09009__A1 _09013_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11507__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08186_ _08243_/B _08394_/A1 _08492_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07206_ _07206_/I _11181_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07137_ _07137_/A1 _07151_/B _07137_/B _07138_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_145_182 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06243__A1 _09374_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07068_ _07068_/I _11148_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xoutput261 _11283_/Q pll90_sel[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput250 _06754_/ZN pad_flash_clk_oe VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput283 _11287_/Q pll_trim[19] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput272 _11280_/Q pll_sel[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput294 _11084_/Q pll_trim[5] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_06019_ _11423_/Q _09197_/A1 _11415_/Q _09171_/A1 _06019_/C _06024_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_59_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11359__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10878__A1 _10924_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10981_ _11016_/A1 input152/Z _10984_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09709_ _09722_/A2 _11582_/Q _09710_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09496__A1 _09497_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11602_ _11602_/D _11686_/RN _06705_/Z _11602_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__05809__A1 _09144_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10802__B2 _10894_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11533_ _11533_/D _11686_/RN _06705_/Z _11533_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_90_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11464_ _11464_/D _11686_/RN _06705_/Z _11464_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10415_ _10452_/A1 _10415_/A2 _10416_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11395_ _11395_/D _11686_/RN _06705_/Z _11395_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__11598__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10346_ _10383_/A1 _10880_/C _10346_/B _10347_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06785__A2 _09015_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10030__A2 _10030_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_10277_ _11386_/Q _10355_/A2 _11378_/Q _10355_/B2 _10277_/C _10286_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08501__B _08637_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10869__A1 _10914_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09487__A1 _09497_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11522__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09239__A1 _09187_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06370_ _06370_/A1 _06370_/A2 _06370_/A3 _06370_/A4 _06371_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_9_74 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_174_255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08040_ _08167_/A2 _08167_/A3 _08162_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06225__A1 _09197_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11493__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09991_ _09991_/A1 _09991_/A2 _09992_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08942_ _07426_/Z _08963_/A2 _08942_/B _08943_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08873_ _06847_/Z _08888_/A2 _08873_/B _08874_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07824_ _08600_/A1 _08494_/A2 _08332_/B _07825_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__09478__A1 _09497_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07755_ _08304_/B _08490_/A3 _08498_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06706_ _11486_/Q _06706_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07686_ _08281_/A1 _07455_/Z _08630_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06637_ input77/Z input91/Z _06638_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11513__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09425_ _09447_/A2 _11491_/Q _09426_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11212__CLK _11656_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09356_ _09372_/A2 _11469_/Q _09357_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06568_ _06557_/Z _10433_/A1 _09934_/I _09945_/A2 _06568_/B2 _11092_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__08453__A2 _08562_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09650__A1 _09672_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08307_ _08307_/A1 _08498_/B _08588_/A2 _08312_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06499_ _06499_/I _11061_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09287_ _09297_/A2 _11447_/Q _09288_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05519_ _05519_/I _05529_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10260__A2 _11521_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08238_ _08490_/A1 _08656_/B _08242_/A1 _08621_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11362__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08205__A2 _08623_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08169_ _08169_/A1 _08169_/A2 _08170_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10200_ _11384_/Q _10355_/A2 _11376_/Q _10355_/B2 _10200_/C _10209_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_11180_ _11180_/D _11686_/RN _06705_/Z _11180_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA_output261_I _11283_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09953__A2 _10265_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10131_ _11326_/Q _10153_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10062_ _11396_/Q _10359_/A2 _11388_/Q _10359_/B2 _10062_/C _10067_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_94_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09469__A1 _09241_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_10964_ _08431_/B _11029_/A1 _11027_/A1 _08460_/B _10965_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_43_320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11504__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08692__A2 _08692_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06152__B1 _11477_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10895_ _10895_/A1 _11227_/Q _10898_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11028__A1 _11028_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09641__A1 _09187_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11516_ _11516_/D _11686_/RN _06705_/Z _11516_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_129_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10745__C _10880_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11447_ _11447_/D _11686_/RN _06705_/Z _11447_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__06207__A1 _05693_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10003__A2 _09973_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11378_ _11378_/D _11686_/RN _06705_/Z _11378_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10329_ _10329_/A1 _10329_/A2 _10329_/A3 _10342_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06530__I _08431_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_537 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_05870_ _09750_/A1 _11601_/Q _05871_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11235__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07540_ _07540_/A1 _07689_/B _07541_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08132__A1 split8/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07471_ _07471_/A1 _07471_/A2 _07471_/B _07472_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08683__A2 _07297_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11019__A1 _10966_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06694__A1 _06694_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11385__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09210_ _09220_/A2 _11423_/Q _09211_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06422_ _09066_/A1 _11379_/Q _06423_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06353_ _09222_/A1 _11427_/Q _06355_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09141_ _09142_/A2 _11402_/Q _09142_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09632__A1 _09125_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10778__B1 _10902_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10242__A2 _10359_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09072_ _09072_/I _11380_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08023_ _08023_/A1 _08023_/A2 _08032_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06997__A2 _06974_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06284_ _07419_/A2 _07006_/A2 _11132_/Q _06286_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_128_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07946__A1 split15/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09974_ _09979_/A1 _10030_/A2 _09975_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09699__A1 _09699_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08925_ _08938_/A2 _11334_/Q _08926_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input20_I mask_rev_in[24] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08856_ _08863_/A2 _11312_/Q _08857_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07174__A2 _09154_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07807_ _08328_/B1 _08329_/B _08331_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08787_ _06904_/Z _08787_/A2 _08787_/A3 _08827_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_05999_ _05999_/A1 _05999_/A2 _05999_/A3 _06036_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_07738_ _07738_/A1 _08298_/B _07738_/A3 _07738_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_25_320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07669_ _07669_/I _07938_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_13_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09408_ _09408_/I _11485_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10680_ _10899_/A1 _11503_/Q _10682_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10481__A2 _11451_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09339_ _09339_/I _11463_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11108__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11301_ _11301_/D input76/Z _06705_/Z _11301_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_11232_ _11232_/D _11686_/RN _06705_/Z _11232_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_11163_ _11163_/D _11163_/RN input68/Z _11163_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10114_ _10371_/A1 _11485_/Q _10115_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11323__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11094_ _11094_/D _11686_/RN _06705_/Z _11094_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xsplit5 split5/I split5/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11258__CLK _11683_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10045_ _10045_/A1 _10045_/A2 _10045_/A3 _10045_/A4 _10046_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__07165__A2 _05925_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08362__A1 _08656_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06912__A2 _06904_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07114__C _07114_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10947_ _10947_/A1 _10950_/A2 _10949_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06676__A1 _06701_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10472__A2 _11419_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10878_ _10924_/A1 _11206_/Q _10879_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08417__A2 _08417_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06428__A1 _05723_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10224__A2 _11544_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09917__A2 _09927_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06971_ _06843_/Z _06971_/A2 _06971_/B _06972_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_09690_ _09697_/A2 _11576_/Q _09691_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05922_ _11456_/Q _09299_/A1 _11448_/Q _09274_/A1 _05922_/C _05923_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_08710_ _08710_/I _11262_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_08641_ _08641_/A1 _07825_/B _08642_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07156__A2 _06701_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05853_ _06396_/A1 input32/Z _05854_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10160__B2 _10351_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08572_ split12/Z _08572_/A2 _08573_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05784_ _09324_/A1 _11466_/Q _05788_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_07523_ _07888_/A2 _07675_/B _07524_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08656__A2 _08696_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07454_ _07533_/I _07490_/I split5/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__10463__A2 _10427_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06667__A1 _06701_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_06405_ _11306_/Q _08829_/A1 _08803_/A1 _11645_/Q _06406_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07385_ _07389_/A2 _11240_/Q _07386_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10215__A2 _11488_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06336_ _05703_/Z _07412_/A1 _11151_/Q _06338_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09124_ _09124_/I _11396_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05890__A2 _11433_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07092__A1 _07092_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06267_ _11279_/Q _08742_/A1 _08726_/A1 _11274_/Q _06269_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09055_ _06855_/Z _09064_/A2 _09055_/B _09056_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08006_ _08006_/A1 _08006_/A2 _07477_/I _08007_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_input68_I mgmt_gpio_in[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06198_ _05703_/Z _08786_/A1 _11262_/Q _06200_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11400__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08592__A1 _07609_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06198__A3 _11262_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09957_ _09957_/I _10373_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
X_08908_ _08908_/I _11328_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07147__A2 _07151_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11550__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_890 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_09888_ _09898_/A1 _09960_/A2 _09889_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10151__A1 _11526_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10151__B2 _10373_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08895__A2 _08913_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08839_ _08839_/A1 _08839_/A2 _06838_/Z _08844_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_10801_ _10801_/A1 _10801_/A2 _10802_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10732_ _10905_/A1 _11536_/Q _10734_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10454__A2 _10406_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_10663_ _10663_/A1 _10663_/A2 _10663_/A3 _10663_/A4 _10691_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__05881__A2 _11521_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10594_ _10899_/A1 _11501_/Q _10598_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10206__A2 _11424_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07083__A1 _07081_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_500 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06830__A1 _06835_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10509__A3 _10509_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11080__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10914__B1 _10914_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11215_ _11215_/D _11672_/CLK _11215_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11146_ _11146_/D _11686_/RN _06705_/Z _11146_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_11077_ _11077_/D _11686_/RN _06705_/Z _11077_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
Xinput150 wb_dat_i[28] input150/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput161 wb_dat_i[9] input161/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10028_ _09893_/I _09878_/I _09899_/I _10351_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__10142__A1 _11446_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05872__A2 _09800_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07170_ _11199_/Q _05925_/Z _07170_/B _07172_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07074__A1 _06843_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11423__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06121_ _08940_/A1 _11341_/Q _06122_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06821__A1 _11007_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07613__A3 _08411_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06052_ _10615_/A2 _05808_/I _05811_/I _10613_/A2 _06053_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_172_364 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09811_ _09154_/I _09823_/A2 _09811_/B _09812_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11573__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07377__A2 _11033_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09742_ _09187_/I _09725_/Z _09742_/B _09743_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08326__A1 _07722_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06954_ _10947_/A1 _06957_/A2 _06956_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06885_ _06885_/I _11094_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09673_ _09673_/I _11570_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05905_ _11584_/Q _09699_/A1 _09674_/A1 _11576_/Q _05906_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06337__B1 _07092_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10133__A1 _10350_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08624_ _08697_/A1 _08624_/A2 _08624_/A3 _08624_/A4 _08634_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA_input122_I wb_adr_i[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05836_ _05836_/I _08803_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_08555_ _08555_/A1 _08555_/A2 _08651_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05767_ _07006_/A2 _08799_/A2 _05768_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07506_ _07506_/I _08045_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__05560__A1 _05519_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05698_ _11554_/Q _09599_/A1 _11546_/Q _09574_/A1 _05698_/C _05714_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_08486_ _08486_/A1 _08486_/A2 _08486_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_07437_ _07437_/A1 _07437_/A2 _07441_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07368_ _07081_/Z _07368_/A2 _07368_/B _07369_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06319_ _09800_/A1 _11611_/Q _06323_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09107_ _09114_/A2 _11392_/Q _09108_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07299_ _11023_/B _07300_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06812__A1 _06835_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08801__A2 _08827_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output174_I _10615_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09038_ _09039_/A2 _11370_/Q _09039_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11000_ _11000_/A1 _10966_/Z _11000_/B _11001_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08317__A1 _08686_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10675__A2 _10894_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06879__A1 _07201_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09817__A1 _09187_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10427__A2 _09912_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09293__A2 _11449_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11695_ _11695_/D _11695_/RN input68/Z _11695_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__11446__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10715_ _10884_/A1 _11384_/Q _10717_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10646_ _10919_/A1 _11366_/Q _10650_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11596__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10577_ _10895_/A1 _11445_/Q _10578_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05606__A2 _05515_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11092__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10363__A1 _11227_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08308__A1 _08332_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11129_ _11129_/D _11686_/RN _06705_/Z _11129_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__05790__A1 _08791_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06670_ input75/Z _06724_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05621_ _11259_/Q _08684_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09808__A1 _09125_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08340_ _08632_/A2 _08614_/A2 _08341_/B _08515_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05552_ _05519_/I _11695_/Q _05553_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09284__A2 _11446_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08271_ _08400_/A1 _07635_/I _08271_/B _08534_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07222_ _05924_/Z _09158_/I _07223_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07153_ _07153_/I _11171_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09036__A2 _09039_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07598__A2 _08417_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06104_ _05941_/I _05726_/I _06108_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08795__A1 _08795_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09992__B1 _11451_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07084_ _07084_/I _11152_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06035_ _06035_/A1 _06035_/A2 _06035_/A3 _06035_/A4 _06036_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__06270__A2 _11324_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08547__A1 _08692_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07986_ split14/Z _08649_/B _08454_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11319__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09725_ _09725_/I _09725_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_86_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06937_ _06938_/A2 _11110_/Q _06938_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10106__A1 _11445_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09656_ _09672_/A2 _11565_/Q _09657_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08607_ split6/Z _08546_/I _08607_/B _08608_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_1105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06325__A3 _11033_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06868_ _06869_/A2 _11086_/Q _06869_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_09587_ _09597_/A2 _11543_/Q _09588_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11469__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_05819_ _06217_/I _08719_/A2 _05820_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06799_ _06835_/A1 _09121_/I _06799_/B _06800_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08538_ _08538_/A1 _08538_/A2 _08538_/A3 _08665_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__07286__A1 _07290_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08469_ _08464_/Z _08570_/A1 _08573_/A1 _08473_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__06089__A2 _11276_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10500_ _11523_/Q _10902_/A2 _10902_/B2 _11515_/Q _10509_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_11480_ _11480_/D _11686_/RN _06705_/Z _11480_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_10_145 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09027__A2 _09039_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10431_ _10444_/A1 _10503_/A2 _10432_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10362_ _10362_/A1 _10362_/A2 _10363_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08786__A1 _08786_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10293_ _10370_/A1 _11498_/Q _10294_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06261__A2 _11272_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09934__I _09934_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10345__A1 _10345_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07210__A1 _07240_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05772__A1 _09016_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07277__A1 _07290_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05827__A2 _05827_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11678_ _11678_/D input162/Z _06687_/A2 _11678_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__07292__A4 _11219_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07029__A1 _06837_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09018__A2 _09039_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10629_ _10900_/A1 _11510_/Q _10630_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08777__A1 _08784_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10584__A1 _10584_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10336__A1 _10375_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07840_ _07840_/I _08545_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__07201__A1 _07201_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10887__A2 _10887_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07771_ _07771_/A1 _08310_/A2 _07771_/A3 _08311_/A1 _07772_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_09510_ _09154_/Z _09522_/A2 _09510_/B _09511_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11611__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06722_ _06753_/A1 input74/Z _06723_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__05763__A1 _08791_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10639__A2 _10916_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08701__A1 _07844_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07504__A2 _07513_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09441_ _09187_/Z _09447_/A2 _09441_/B _09442_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06653_ _11059_/Q _11175_/Q _06654_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06584_ _07457_/I _07470_/I _06585_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09372_ _09270_/Z _09372_/A2 _09372_/B _09373_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05604_ _05616_/C _11254_/Q _05604_/B _05605_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08323_ _08332_/A1 _08417_/A2 _08592_/B _08507_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07268__A1 _07290_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05535_ _05541_/A2 _05541_/A1 _05539_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08254_ _08281_/A1 _08519_/A2 _08400_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_08185_ _08185_/I _08243_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07205_ _07240_/A1 _07205_/A2 _07205_/B _07206_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07136_ _11193_/Q _05927_/Z _07151_/B _07136_/C _07137_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08768__A1 _08784_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10575__A1 _10897_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07067_ _06843_/Z _07067_/A2 _07067_/B _07068_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input50_I mgmt_gpio_in[22] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput240 _06633_/Z mgmt_gpio_out[36] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput251 _06710_/ZN pad_flash_csb VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput262 _11292_/Q pll_bypass VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_06018_ _06018_/A1 _06018_/A2 _06019_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11141__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10327__A1 _10367_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07991__A2 _08395_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput273 _11079_/Q pll_trim[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput284 _11080_/Q pll_trim[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput295 _11085_/Q pll_trim[6] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__08940__A1 _08940_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09708_ _09708_/I _11581_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07969_ split14/Z _08609_/B _07971_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11291__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05754__A1 _06204_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_10980_ _10980_/I _11676_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09639_ _09639_/I _11559_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_output304_I _05841_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07259__A1 _06859_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11601_ _11601_/D _11686_/RN _06705_/Z _11601_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__09248__A2 _09015_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11614__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10802__A2 _10894_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11532_ _11532_/D _11686_/RN _06705_/Z _11532_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__05809__A2 _11410_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11295__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11463_ _11463_/D _11686_/RN _06705_/Z _11463_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10414_ _10414_/I _10452_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08759__A1 _06859_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11394_ _11394_/D _11686_/RN _06705_/Z _11394_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__10566__A1 _10886_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10345_ _10345_/A1 _06556_/I _10926_/C _10345_/C _10346_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__10030__A3 _10265_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_719 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_10276_ _10276_/A1 _10276_/A2 _10277_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10318__A1 _10357_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09184__A1 _09195_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11634__CLK _11658_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08931__A1 _08938_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09239__A2 _09246_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08998__A1 _06847_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11164__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10557__A1 _10548_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09990_ _10367_/A1 _11475_/Q _09991_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_08941_ _08963_/A2 _11339_/Q _08942_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08872_ _08888_/A2 _11317_/Q _08873_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09175__A1 _09195_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07823_ _08600_/A1 _07823_/A2 _07827_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08922__A1 _08938_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09478__A2 _11508_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07754_ _07754_/A1 _07754_/A2 _08678_/A2 _08297_/B _07757_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_07685_ _07685_/I _08281_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
X_06705_ _06705_/I _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
XFILLER_44_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06636_ _06636_/I _06636_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09424_ _09424_/A1 _09015_/Z _09447_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_09355_ _09355_/I _11468_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06567_ _06567_/I _06568_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11507__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08306_ _08306_/I _08588_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06498_ _06500_/A1 _06498_/A2 _06498_/B _06499_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05518_ _05523_/A1 _11161_/Q _05519_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_09286_ _09286_/I _11446_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input98_I wb_adr_i[10] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10796__A1 _10884_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08237_ split12/Z _08614_/A2 _08205_/C _08621_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11277__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08168_ _08168_/I _08490_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_118_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11657__CLK _11658_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07119_ _11165_/Q _07122_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08099_ _08656_/A1 _08209_/B _08100_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05975__A1 _08839_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10130_ _11649_/Q _10191_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09166__A1 _06863_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10061_ _10061_/A1 _10061_/A2 _10062_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08913__A1 _06867_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11201__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05727__A1 _07006_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09469__A2 _09472_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10963_ input168/Z input165/Z _11027_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06152__A1 _11485_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06152__B2 _09374_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10894_ _11249_/Q _10894_/A2 _11245_/Q _10894_/B2 _10894_/C _10898_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_70_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11187__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09641__A2 _09647_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11515_ _11515_/D _11686_/RN _06705_/Z _11515_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_11_251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10787__A1 _10787_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_429 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10539__A1 _10902_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11446_ _11446_/D _11686_/RN _06705_/Z _11446_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__06207__A2 _11524_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11377_ _11377_/D _11686_/RN _06705_/Z _11377_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10328_ _10366_/A1 _11236_/Q _10329_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11440__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10259_ _10259_/A1 _10259_/A2 _10259_/A3 _10264_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08904__A1 _06855_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10711__A1 _10887_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08380__A2 _08355_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_287 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07470_ _07470_/I _07471_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__06143__A1 _09800_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06421_ _07419_/A2 _07006_/A2 _11131_/Q _06423_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06352_ _09248_/A1 _11435_/Q _06355_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09140_ _09140_/I _11401_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09632__A2 _09647_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10778__B2 _11521_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11259__RN input162/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09071_ _07431_/Z _09089_/A2 _09071_/B _09072_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06283_ _09091_/A1 _11388_/Q _07013_/A1 _11134_/Q _06286_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08022_ _08391_/B _08204_/I _08023_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09396__A1 _09397_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09973_ _09973_/I _10030_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__06721__I _06721_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10950__A1 _10950_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input152_I wb_dat_i[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09148__A1 _09169_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11431__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08924_ _08924_/I _11333_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_split8_I split8/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09699__A2 _09015_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08855_ _08855_/I _11311_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10702__A1 _10914_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05709__A1 _05703_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07806_ _08696_/A2 _08329_/B _08511_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06382__A1 _09399_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08786_ _08786_/A1 _08799_/A1 _08789_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07737_ _07885_/I _08339_/A1 _07738_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05998_ _05998_/A1 _06265_/A2 _05998_/A3 _05998_/A4 _05999_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA_input13_I mask_rev_in[18] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07668_ _07890_/A1 _07890_/A2 _07672_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11498__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06134__A1 _09549_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09871__A2 _09935_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09407_ _09125_/Z _09422_/A2 _09407_/B _09408_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07599_ _08262_/B _08509_/A1 _08260_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06619_ _06619_/A1 _06619_/A2 _06619_/B _06620_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10218__B1 _10379_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09338_ _09158_/Z _09347_/A2 _09338_/B _09339_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_111_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10769__A1 _10895_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09269_ _09269_/I _11441_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11300_ _11300_/D input76/Z _06705_/Z _11300_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__09387__A1 _09397_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11231_ _11231_/D _11686_/RN _06705_/Z _11231_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_20_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07727__I _07727_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11162_ _11162_/D _11162_/RN input68/Z _11162_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__10941__A1 _10934_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10113_ _10370_/A1 _11493_/Q _10115_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05948__A1 _08890_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09139__A1 _06863_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11422__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11093_ _11093_/D _11686_/RN _06705_/Z _11093_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xsplit6 split6/I split6/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10044_ _11379_/Q _10355_/A2 _10355_/B2 _11371_/Q _10045_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06373__A1 _08795_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08114__A2 split16/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11489__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11492__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10946_ _10946_/I _11670_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_16_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06125__A1 _09016_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10877_ _10877_/A1 _10877_/A2 _10877_/A3 _10877_/A4 _10877_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_1
XPHY_360 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07625__A1 _08686_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09378__A1 _09397_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11661__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11429_ _11429_/D input76/Z _06705_/Z _11429_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_6_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11202__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06970_ _06971_/A2 _11120_/Q _06971_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05921_ _05921_/A1 _05921_/A2 _05922_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input5_I mask_rev_in[10] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09550__A1 _09572_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08640_ _08640_/A1 _08640_/A2 _08640_/A3 _08640_/A4 _08680_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__11445__SETN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05852_ _06394_/A1 input9/Z _05854_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10160__A2 _10351_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11352__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_287 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06364__A1 _07412_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08571_ _08200_/B _08696_/A2 _08571_/B _08573_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05783_ _05783_/I _09324_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XPHY_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10999__A1 _10966_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07522_ _07522_/I _07675_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_81_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06116__A1 _06785_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07453_ _07496_/I input97/Z _07490_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_34_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05875__B1 _05925_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06404_ _08726_/A1 _11273_/Q _06406_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07384_ _06238_/Z _11033_/A2 _06838_/Z _07389_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_09123_ _09121_/Z _09142_/A2 _09123_/B _09124_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06335_ _09599_/A1 _11547_/Q _06338_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07092__A2 _06904_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06266_ _06266_/I _06694_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09054_ _09064_/A2 _11375_/Q _09055_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08005_ _08005_/A1 _08005_/A2 _08007_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09369__A1 _09241_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11652__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06197_ _06197_/I _08786_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__08592__A2 _08592_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09956_ _10023_/A1 _09899_/I _09957_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_880 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_09887_ _09887_/I _09960_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08907_ _06859_/Z _08913_/A2 _08907_/B _08908_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09541__A1 _09187_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_08838_ _08838_/I _11306_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10151__A2 _10373_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08769_ _06847_/Z _08784_/A2 _08769_/B _08770_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10800_ _10892_/A1 _11474_/Q _10801_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09844__A2 _11625_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10731_ _10903_/A1 _11560_/Q _10736_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10662_ _11583_/Q _10913_/B2 _10913_/A2 _11591_/Q _10663_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_10593_ _10589_/Z _10593_/A2 _10593_/A3 _10593_/A4 _10604_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__08280__A1 split14/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11225__CLK _06687_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11643__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06830__A2 _09241_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11214_ _11214_/D _11672_/CLK _11214_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10914__B2 _11239_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10914__A1 _10914_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09780__A1 _09121_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08583__A2 _08493_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11145_ _11145_/D _11686_/RN _06705_/Z _11145_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__11375__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11076_ _11076_/D _11686_/RN _06705_/Z _11076_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
Xinput151 wb_dat_i[29] input151/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput140 wb_dat_i[19] input140/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09532__A1 _09125_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10678__B1 _10897_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput162 wb_rstn_i input162/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_48_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10027_ _10027_/A1 _10027_/A2 _10027_/A3 _10027_/A4 _10046_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__06346__A1 _09649_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08099__A1 _08656_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09835__A2 _11622_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10929_ _11666_/Q _10931_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06649__A2 _06649_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07141__B _07151_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09599__A1 _09599_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05609__B1 _05633_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08271__A1 _08400_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06120_ _11333_/Q _10607_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06051_ _11398_/Q _10613_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11634__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06821__A2 _05633_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10905__A1 _10905_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09810_ _09823_/A2 _11614_/Q _09811_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07377__A3 _06838_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09741_ _09725_/Z _11592_/Q _09742_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06953_ _06953_/I _11114_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08326__A2 _07586_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05904_ _09649_/A1 _11568_/Q _05906_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06884_ _06843_/Z _06902_/A2 _06884_/B _06885_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09672_ _09270_/Z _09672_/A2 _09672_/B _09673_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06337__A1 _09574_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08623_ _08242_/B _08623_/A2 _08624_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05835_ _08839_/A1 _11033_/A2 _05836_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_08554_ _08375_/B _08692_/A2 _08554_/B _08554_/C _08555_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA_input115_I wb_adr_i[26] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05766_ _05766_/I _09066_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XANTENNA__09826__A2 _11619_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07505_ _07505_/I _07793_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
X_05697_ _05697_/A1 _05697_/A2 _05698_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08485_ _08485_/I _08486_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07436_ input103/Z input102/Z _07437_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06446__I _06446_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07367_ _07368_/A2 _11235_/Q _07368_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11248__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06318_ _06318_/A1 _06318_/A2 _06318_/A3 _06318_/A4 _06329_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__08262__A1 split21/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09106_ _09106_/I _11391_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input80_I spi_enabled VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11625__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07298_ _07844_/B _10930_/B _11023_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09037_ _09037_/I _11369_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06249_ _08795_/A1 _06238_/Z _11148_/Q _06252_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__06812__A2 _09154_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11398__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08565__A2 _08696_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06025__B1 _05925_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output334_I _11672_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08317__A2 _08689_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09939_ _09939_/I _09940_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_172_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06879__A2 _06838_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09817__A2 _09823_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_split16_I split16/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11694_ _11694_/D _11694_/RN input68/Z _11694_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_9_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10714_ _10883_/A1 _11376_/Q _10717_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10645_ _10645_/A1 _10645_/A2 _10645_/A3 _10645_/A4 _10652_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_42_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11616__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10576_ _10896_/A1 _11437_/Q _10578_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10060__A1 _10357_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06803__A2 _05633_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11128_ _11128_/D _11683_/CLK _11128_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08308__A2 _08417_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07136__B _07151_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05790__A2 _06238_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06319__A1 _09800_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11059_ _11059_/D _11059_/RN input68/Z _11059_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_05620_ _06480_/A1 _05515_/I _05620_/B _05623_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09808__A2 _09823_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05551_ _11694_/Q _05553_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08270_ split14/Z _07609_/Z _08417_/B _08418_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06098__A3 _06098_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06266__I _06266_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07221_ _07221_/I _11184_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07152_ _07152_/A1 _07151_/B _07152_/B _07153_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11540__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11607__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06103_ _06103_/I _11266_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_172_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07083_ _07081_/Z _07083_/A2 _07083_/B _07084_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08795__A2 _08799_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06034_ _06034_/A1 _06034_/A2 _06034_/A3 _06034_/A4 _06035_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_99_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09744__A1 _09725_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11690__CLK input68/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07985_ _08355_/I _08649_/B _08454_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_435 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09724_ _09724_/A1 _05636_/I _05668_/I _07114_/C _09725_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_1
X_06936_ _06936_/I _11109_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06867_ _09270_/I _06867_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_09655_ _09655_/I _11564_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08606_ _08606_/I _11257_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05818_ _05818_/I _09274_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_09586_ _09586_/I _11542_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_06798_ _06835_/A1 _11072_/Q _06799_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_08537_ _08686_/A1 _08686_/A2 _08537_/B _08538_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05749_ _05749_/A1 _05749_/A2 _05750_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11070__CLK input68/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08468_ _08468_/A1 _08203_/I _08573_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06176__I _11239_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10290__A1 _10290_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07419_ _05703_/Z _07419_/A2 _06838_/Z _07424_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_23_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08399_ _08399_/I _11255_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10430_ _10408_/I _09912_/I _10444_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_10_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output284_I _11080_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06904__I _09015_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10361_ _10361_/A1 _11140_/Q _10362_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08786__A2 _08799_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10292_ _10371_/A1 _11490_/Q _10294_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06261__A3 _08719_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09735__A1 _09725_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10345__A2 _06556_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06549__B2 _11302_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05772__A2 _11370_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11413__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11563__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10805__B1 _10897_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_474 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10281__B2 _10359_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11677_ _11677_/D input162/Z _06687_/A2 _11677_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_146_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05827__A3 _05827_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10628_ _10899_/A1 _11502_/Q _10630_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06788__A1 _10972_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10559_ _10559_/A1 _06556_/I _10560_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10033__B2 _10351_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10584__A2 _10578_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09726__A1 _09725_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08529__A2 _08529_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07201__A2 _05924_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07770_ _08332_/A1 _07774_/A2 _08311_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11093__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06960__A1 _06941_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06721_ _06721_/I _06721_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05763__A2 _07006_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09440_ _09447_/A2 _11496_/Q _09441_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06652_ _06652_/A1 _06652_/A2 _06652_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06712__A1 _11056_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06583_ _06583_/A1 _06583_/A2 _06583_/A3 _06583_/A4 _06589_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_09371_ _09372_/A2 _11474_/Q _09372_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05603_ _06500_/B1 _05515_/I _05603_/B _05616_/C _05604_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08322_ _08322_/A1 _08593_/A1 _08593_/A2 _08327_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05534_ _11698_/Q _05541_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08253_ _08403_/A1 _08253_/A2 _08528_/A2 _08528_/A3 _08259_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__10272__A1 _10350_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07204_ _07240_/A1 _11181_/Q _07205_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08217__A1 split7/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08184_ _08490_/A1 _08205_/C _08185_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07135_ _05927_/Z _09158_/I _07136_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10575__A2 _11461_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07066_ _07067_/A2 _11148_/Q _07067_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput230 _11096_/Q mgmt_gpio_out[27] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput241 _06629_/Z mgmt_gpio_out[37] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput252 _06753_/ZN pad_flash_csb_oe VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_06017_ _09117_/A1 _11399_/Q _06018_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input43_I mgmt_gpio_in[16] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput274 _11073_/Q pll_trim[10] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput285 _11288_/Q pll_trim[20] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput263 _11272_/Q pll_dco_ena VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput296 _11086_/Q pll_trim[7] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__11436__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07968_ _08355_/I _08609_/B _07971_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08940__A2 _06838_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09707_ _09125_/I _09722_/A2 _09707_/B _09708_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06951__A1 _06941_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06919_ _07006_/A2 _11033_/A2 _06871_/Z _06924_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__05754__A2 _05738_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07899_ _07899_/I split21/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__11586__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09638_ _09158_/Z _09647_/A2 _09638_/B _09639_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09569_ _09241_/Z _09572_/A2 _09569_/B _09570_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07259__A2 _07265_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11600_ _11600_/D _11686_/RN _06705_/Z _11600_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_11531_ _11531_/D _11686_/RN _06705_/Z _11531_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_135_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11462_ _11462_/D _11686_/RN _06705_/Z _11462_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_7_426 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05690__A1 _05703_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10413_ _10460_/A1 _10501_/A1 _10414_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09956__A1 _10023_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08759__A2 _08759_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11393_ _11393_/D _11686_/RN _06705_/Z _11393_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10344_ _10344_/A1 _06556_/I _10345_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_151_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10275_ _10352_/A1 _11362_/Q _10276_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06942__A1 _10935_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07498__A2 _07522_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10254__A1 _10370_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08998__A2 _09013_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05588__C _05616_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11309__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10557__A2 _10924_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11459__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08940_ _08940_/A1 _06838_/Z _08963_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__09175__A2 _11412_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08871_ _08871_/I _11316_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07822_ _07822_/I _07823_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07186__A1 _07197_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07753_ _08589_/A1 _08242_/A1 _08297_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06704_ _07242_/A2 _06704_/A2 _05616_/C _11023_/A2 _06705_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_4
X_07684_ _07684_/A1 _07684_/A2 _08540_/A2 _07684_/A4 _07688_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__08686__A1 _08686_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06635_ _11622_/Q input77/Z _06635_/B _06636_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09423_ _09423_/I _11490_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09354_ _09121_/Z _09372_/A2 _09354_/B _09355_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08305_ _08686_/A2 _07761_/I _08305_/B _08306_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06566_ _10425_/A2 _11641_/Q _09934_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_06497_ _06497_/A1 _11060_/Q _06497_/A3 _06498_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05517_ _05517_/I _05523_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
X_09285_ _09154_/Z _09297_/A2 _09285_/B _09286_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_60_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08236_ _08236_/I _08578_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07661__A2 _07609_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08167_ _08167_/A1 _08167_/A2 _08167_/A3 _08168_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__05672__A1 _09750_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07118_ _07118_/I _11164_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08098_ _08098_/I _08209_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
X_07049_ _07053_/A2 _11143_/Q _07050_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05975__A2 _05995_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09166__A2 _09169_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10060_ _10357_/A1 _11412_/Q _10061_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07177__A1 _07197_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08913__A2 _08913_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05727__A2 _05995_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06924__A1 _06843_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10962_ input168/Z input164/Z _11029_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06629__I _06629_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06152__A2 _09399_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10893_ _10893_/A1 _10893_/A2 _10894_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07101__A1 _07076_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10236__A1 _10352_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11514_ _11514_/D _11686_/RN _06705_/Z _11514_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__10787__A2 _10092_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11445_ _11445_/D _11686_/RN _06705_/Z _11445_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_50_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11601__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10539__A2 _11524_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11376_ _11376_/D _11686_/RN _06705_/Z _11376_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10327_ _10367_/A1 _11240_/Q _10329_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06612__B1 _06466_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_462 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_10258_ _10377_/B1 _11569_/Q _10259_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08904__A2 _08913_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10189_ _10189_/A1 _10189_/A2 _10189_/A3 _10189_/A4 _10190_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__10711__A2 _11432_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10172__B1 _11439_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10475__A1 _10642_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07340__A1 _07081_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06420_ _09091_/A1 _11387_/Q _07013_/A1 _11133_/Q _06423_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11131__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06351_ _06213_/Z _11226_/Q _06355_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09093__A1 _07426_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10778__A2 _10902_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06282_ _06204_/I _05719_/I _07013_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09070_ _09089_/A2 _11380_/Q _09071_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08021_ _08021_/A1 _08390_/A2 _08021_/A3 _08023_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11281__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09396__A2 _11482_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09972_ _09972_/I _09979_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08923_ _06847_/Z _08938_/A2 _08923_/B _08924_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07159__A1 _05925_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08854_ _06847_/Z _08863_/A2 _08854_/B _08855_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05709__A2 _08719_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input145_I wb_dat_i[23] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11195__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07805_ _07805_/A1 _08226_/A2 _08596_/A2 _07805_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
X_08785_ _08785_/I _11291_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05997_ _06398_/A2 input24/Z _05998_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07736_ _07828_/I _08495_/B _07885_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_44_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10466__A1 _10894_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07667_ _07674_/A2 _07505_/I _07890_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09406_ _09422_/A2 _11485_/Q _09407_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07598_ _08262_/B _08417_/A2 _08408_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07882__A2 _07593_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06618_ _06604_/B _06610_/B _06619_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11624__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10218__B2 _11560_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09337_ _09347_/A2 _11463_/Q _09338_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06549_ _06567_/I _09945_/A2 _09946_/A1 _11302_/Q _06550_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__10769__A2 _11449_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09268_ _09241_/Z _09272_/A2 _09268_/B _09269_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08219_ _08696_/B _08221_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_output197_I _10642_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08831__A1 _06847_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09199_ _09116_/Z _09220_/A2 _09199_/B _09200_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09387__A2 _11479_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07398__A1 _07398_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11230_ _11230_/D _11686_/RN _06705_/Z _11230_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_11161_ _11161_/D _11161_/RN input68/Z _11161_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__06070__B2 _10634_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10112_ _11509_/Q _10369_/A2 _10369_/B1 _11501_/Q _10115_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06070__A1 _10146_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05948__A2 _11328_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09139__A2 _09142_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xsplit7 split7/I split7/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_136_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11092_ _11092_/D input76/Z _11663_/CLK _11092_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08898__A1 _06847_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10043_ _10043_/I _10355_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__11186__RN input76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11154__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06373__A2 _06238_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10945_ _10945_/A1 _10934_/I _10945_/B _10946_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10876_ _10922_/A1 _11107_/Q _10877_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05884__B2 _09424_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05884__A1 _11505_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07625__A2 _08686_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11110__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11428_ _11428_/D input76/Z _06705_/Z _11428_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__07389__A1 _07081_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11359_ _11359_/D _11686_/RN _06705_/Z _11359_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__06061__A1 _07201_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05939__A2 _05939_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_05920_ _09222_/A1 _11432_/Q _05921_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11177__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05851_ _06393_/A1 input18/Z _05854_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08570_ _08570_/A1 _08570_/A2 _08100_/I _07763_/I _08617_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_81_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07521_ _07521_/A1 _07521_/A2 _07575_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05782_ _06238_/I _06872_/A2 _05783_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10448__A1 _10903_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11647__CLK _11663_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06116__A2 _11073_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07452_ _07487_/I input119/Z _07533_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__05875__A1 input70/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_07383_ _07383_/I _11239_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06403_ _08742_/A1 _11278_/Q _06406_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09066__A1 _09066_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06334_ _11157_/Q _07099_/A1 _11523_/Q _05693_/Z _06334_/C _06338_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_09122_ _09142_/A2 _11396_/Q _09123_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08813__A1 _08820_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10620__A1 _10891_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09053_ _09053_/I _11374_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06265_ _06265_/A1 _06265_/A2 _06265_/A3 _06265_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__11101__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_08004_ _08167_/A3 _08039_/I _08008_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__09369__A2 _09372_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_06196_ _09649_/A1 _11564_/Q _06200_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06052__A1 _10615_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09955_ _09973_/I _09887_/I _10265_/A3 _10373_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__06052__B2 _10613_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11177__CLK _06705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09886_ _09892_/A2 _11634_/Q _09887_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_08906_ _08913_/A2 _11328_/Q _08907_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11168__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09541__A2 _09547_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10687__A1 _10906_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_892 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_881 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_08837_ _07426_/Z _08837_/A2 _08837_/B _08838_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_122_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08768_ _08784_/A2 _11286_/Q _08769_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10439__A1 _10913_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07719_ _07719_/A1 _08431_/B _07845_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08699_ _08699_/A1 _08036_/B _11028_/A2 _08699_/B2 _08700_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_25_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07304__A1 _07076_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10730_ _10904_/A1 _11552_/Q _10736_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05866__A1 _09674_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10661_ _10911_/A1 _11575_/Q _10663_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09057__A1 _09064_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10592_ _10915_/A1 _11613_/Q _10916_/A1 _11621_/Q _10593_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08804__A1 _08820_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08280__A2 _07609_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11213_ _11213_/D _11656_/CLK _11213_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09780__A2 _09798_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11144_ _11144_/D _11686_/RN _06705_/Z _11144_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__07791__A1 _08696_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06594__A2 input129/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_11075_ _11075_/D _11686_/RN _06705_/Z _11075_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xinput163 wb_sel_i[0] input163/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput152 wb_dat_i[2] input152/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput130 wb_dat_i[0] input130/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput141 wb_dat_i[1] input141/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09532__A2 _09547_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10678__B2 _11463_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10026_ _10359_/B2 _11387_/Q _10359_/A2 _11395_/Q _10027_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07543__A1 _07685_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10928_ _10928_/I _11665_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10850__A1 _10896_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05857__A1 _09041_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_10859_ _10905_/A1 _11157_/Q _10861_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09048__A1 _09064_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09599__A2 _09015_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_180 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10602__A1 _10906_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05609__B2 _05609_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08271__A2 _07635_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06050_ _11406_/Q _10615_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06282__A1 _06204_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09220__A1 _06867_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11398__RN _11686_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07782__A1 _08592_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_09740_ _09740_/I _11591_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06952_ _10945_/A1 _06941_/I _06952_/B _06953_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
.ends

