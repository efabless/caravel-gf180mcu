VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO digital_pll
  CLASS BLOCK ;
  FOREIGN digital_pll ;
  ORIGIN 0.000 0.000 ;
  SIZE 170.000 BY 100.000 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 24.650 3.620 26.250 94.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 64.350 3.620 65.950 94.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 104.050 3.620 105.650 94.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 143.750 3.620 145.350 94.380 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 5.300 14.640 164.380 16.240 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 5.300 37.680 164.380 39.280 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 5.300 60.720 164.380 62.320 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 5.300 83.760 164.380 85.360 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 44.500 3.620 46.100 94.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 84.200 3.620 85.800 94.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 123.900 3.620 125.500 94.380 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 5.300 26.160 164.380 27.760 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 5.300 49.200 164.380 50.800 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 5.300 72.240 164.380 73.840 ;
    END
  END VSS
  PIN clockp[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3.080 4.000 3.640 ;
    END
  END clockp[0]
  PIN clockp[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 9.240 4.000 9.800 ;
    END
  END clockp[1]
  PIN dco
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 52.920 4.000 53.480 ;
    END
  END dco
  PIN div[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 15.400 4.000 15.960 ;
    END
  END div[0]
  PIN div[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 21.560 4.000 22.120 ;
    END
  END div[1]
  PIN div[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 27.720 4.000 28.280 ;
    END
  END div[2]
  PIN div[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 33.880 4.000 34.440 ;
    END
  END div[3]
  PIN div[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 40.040 4.000 40.600 ;
    END
  END div[4]
  PIN enable
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 46.200 4.000 46.760 ;
    END
  END enable
  PIN ext_trim[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 59.080 4.000 59.640 ;
    END
  END ext_trim[0]
  PIN ext_trim[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 45.080 96.000 45.640 100.000 ;
    END
  END ext_trim[10]
  PIN ext_trim[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 57.960 96.000 58.520 100.000 ;
    END
  END ext_trim[11]
  PIN ext_trim[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 70.840 96.000 71.400 100.000 ;
    END
  END ext_trim[12]
  PIN ext_trim[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 84.280 96.000 84.840 100.000 ;
    END
  END ext_trim[13]
  PIN ext_trim[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 97.160 96.000 97.720 100.000 ;
    END
  END ext_trim[14]
  PIN ext_trim[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 110.600 96.000 111.160 100.000 ;
    END
  END ext_trim[15]
  PIN ext_trim[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 123.480 96.000 124.040 100.000 ;
    END
  END ext_trim[16]
  PIN ext_trim[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 136.360 96.000 136.920 100.000 ;
    END
  END ext_trim[17]
  PIN ext_trim[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 149.800 96.000 150.360 100.000 ;
    END
  END ext_trim[18]
  PIN ext_trim[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 162.680 96.000 163.240 100.000 ;
    END
  END ext_trim[19]
  PIN ext_trim[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 65.240 4.000 65.800 ;
    END
  END ext_trim[1]
  PIN ext_trim[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 166.000 91.000 170.000 91.560 ;
    END
  END ext_trim[20]
  PIN ext_trim[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 166.000 74.200 170.000 74.760 ;
    END
  END ext_trim[21]
  PIN ext_trim[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 166.000 57.960 170.000 58.520 ;
    END
  END ext_trim[22]
  PIN ext_trim[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 166.000 41.160 170.000 41.720 ;
    END
  END ext_trim[23]
  PIN ext_trim[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 166.000 24.360 170.000 24.920 ;
    END
  END ext_trim[24]
  PIN ext_trim[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 166.000 8.120 170.000 8.680 ;
    END
  END ext_trim[25]
  PIN ext_trim[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 71.400 4.000 71.960 ;
    END
  END ext_trim[2]
  PIN ext_trim[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 77.560 4.000 78.120 ;
    END
  END ext_trim[3]
  PIN ext_trim[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 83.720 4.000 84.280 ;
    END
  END ext_trim[4]
  PIN ext_trim[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 89.880 4.000 90.440 ;
    END
  END ext_trim[5]
  PIN ext_trim[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 96.040 4.000 96.600 ;
    END
  END ext_trim[6]
  PIN ext_trim[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 5.880 96.000 6.440 100.000 ;
    END
  END ext_trim[7]
  PIN ext_trim[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 18.760 96.000 19.320 100.000 ;
    END
  END ext_trim[8]
  PIN ext_trim[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 31.640 96.000 32.200 100.000 ;
    END
  END ext_trim[9]
  PIN osc
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 127.400 0.000 127.960 4.000 ;
    END
  END osc
  PIN resetb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 42.280 0.000 42.840 4.000 ;
    END
  END resetb
  OBS
      LAYER Metal1 ;
        RECT 5.600 2.670 164.080 94.380 ;
      LAYER Metal2 ;
        RECT 4.340 95.700 5.580 96.000 ;
        RECT 6.740 95.700 18.460 96.000 ;
        RECT 19.620 95.700 31.340 96.000 ;
        RECT 32.500 95.700 44.780 96.000 ;
        RECT 45.940 95.700 57.660 96.000 ;
        RECT 58.820 95.700 70.540 96.000 ;
        RECT 71.700 95.700 83.980 96.000 ;
        RECT 85.140 95.700 96.860 96.000 ;
        RECT 98.020 95.700 110.300 96.000 ;
        RECT 111.460 95.700 123.180 96.000 ;
        RECT 124.340 95.700 136.060 96.000 ;
        RECT 137.220 95.700 149.500 96.000 ;
        RECT 150.660 95.700 162.380 96.000 ;
        RECT 4.340 4.300 163.100 95.700 ;
        RECT 4.340 2.610 41.980 4.300 ;
        RECT 43.140 2.610 127.100 4.300 ;
        RECT 128.260 2.610 163.100 4.300 ;
      LAYER Metal3 ;
        RECT 4.300 95.740 166.000 96.460 ;
        RECT 4.000 91.860 166.000 95.740 ;
        RECT 4.000 90.740 165.700 91.860 ;
        RECT 4.300 90.700 165.700 90.740 ;
        RECT 4.300 89.580 166.000 90.700 ;
        RECT 4.000 84.580 166.000 89.580 ;
        RECT 4.300 83.420 166.000 84.580 ;
        RECT 4.000 78.420 166.000 83.420 ;
        RECT 4.300 77.260 166.000 78.420 ;
        RECT 4.000 75.060 166.000 77.260 ;
        RECT 4.000 73.900 165.700 75.060 ;
        RECT 4.000 72.260 166.000 73.900 ;
        RECT 4.300 71.100 166.000 72.260 ;
        RECT 4.000 66.100 166.000 71.100 ;
        RECT 4.300 64.940 166.000 66.100 ;
        RECT 4.000 59.940 166.000 64.940 ;
        RECT 4.300 58.820 166.000 59.940 ;
        RECT 4.300 58.780 165.700 58.820 ;
        RECT 4.000 57.660 165.700 58.780 ;
        RECT 4.000 53.780 166.000 57.660 ;
        RECT 4.300 52.620 166.000 53.780 ;
        RECT 4.000 47.060 166.000 52.620 ;
        RECT 4.300 45.900 166.000 47.060 ;
        RECT 4.000 42.020 166.000 45.900 ;
        RECT 4.000 40.900 165.700 42.020 ;
        RECT 4.300 40.860 165.700 40.900 ;
        RECT 4.300 39.740 166.000 40.860 ;
        RECT 4.000 34.740 166.000 39.740 ;
        RECT 4.300 33.580 166.000 34.740 ;
        RECT 4.000 28.580 166.000 33.580 ;
        RECT 4.300 27.420 166.000 28.580 ;
        RECT 4.000 25.220 166.000 27.420 ;
        RECT 4.000 24.060 165.700 25.220 ;
        RECT 4.000 22.420 166.000 24.060 ;
        RECT 4.300 21.260 166.000 22.420 ;
        RECT 4.000 16.260 166.000 21.260 ;
        RECT 4.300 15.100 166.000 16.260 ;
        RECT 4.000 10.100 166.000 15.100 ;
        RECT 4.300 8.980 166.000 10.100 ;
        RECT 4.300 8.940 165.700 8.980 ;
        RECT 4.000 7.820 165.700 8.940 ;
        RECT 4.000 3.940 166.000 7.820 ;
        RECT 4.300 3.220 166.000 3.940 ;
      LAYER Metal4 ;
        RECT 6.020 4.850 24.350 92.030 ;
        RECT 26.550 4.850 44.200 92.030 ;
        RECT 46.400 4.850 64.050 92.030 ;
        RECT 66.250 4.850 83.900 92.030 ;
        RECT 86.100 4.850 103.750 92.030 ;
        RECT 105.950 4.850 123.600 92.030 ;
        RECT 125.800 4.850 138.460 92.030 ;
      LAYER Metal5 ;
        RECT 7.620 85.860 138.540 92.020 ;
        RECT 7.620 74.340 138.540 83.260 ;
        RECT 7.620 62.820 138.540 71.740 ;
        RECT 7.620 51.300 138.540 60.220 ;
        RECT 7.620 39.780 138.540 48.700 ;
        RECT 7.620 28.260 138.540 37.180 ;
        RECT 7.620 16.880 138.540 25.660 ;
  END
END digital_pll
END LIBRARY

